module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84, po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96, po97);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71, po72, po73, po74, po75, po76, po77, po78, po79, po80, po81, po82, po83, po84, po85, po86, po87, po88, po89, po90, po91, po92, po93, po94, po95, po96, po97;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396;
assign w0 = pi026 & ~w179;
assign w1 = pi045 & ~w371;
assign w2 = (pi088 & ~w371) | (pi088 & w8) | (~w371 & w8);
assign w3 = ~w177 & ~w258;
assign w4 = pi015 & pi010;
assign w5 = w95 & w337;
assign w6 = (pi088 & ~w371) | (pi088 & w348) | (~w371 & w348);
assign w7 = pi018 & ~w179;
assign w8 = pi085 & pi088;
assign w9 = ~w210 & w35;
assign w10 = pi015 & w95;
assign w11 = pi021 & ~pi092;
assign w12 = ~w216 & w291;
assign w13 = ~w39 & w228;
assign w14 = pi033 & w95;
assign w15 = ~w164 & ~w310;
assign w16 = pi069 & w333;
assign w17 = ~pi041 & pi088;
assign w18 = ~w234 & ~w393;
assign w19 = ~pi015 & pi011;
assign w20 = ~w270 & ~w207;
assign w21 = ~w0 & w238;
assign w22 = pi044 & ~w371;
assign w23 = ~w189 & w332;
assign w24 = (pi088 & ~w179) | (pi088 & w348) | (~w179 & w348);
assign w25 = ~w328 & ~w11;
assign w26 = ~w120 & w362;
assign w27 = ~w10 & ~w53;
assign w28 = w184 & ~w285;
assign w29 = ~w87 & ~w305;
assign w30 = pi079 & ~pi104;
assign w31 = pi075 & w333;
assign w32 = pi063 & ~w93;
assign w33 = w184 & ~w342;
assign w34 = ~w80 & ~w274;
assign w35 = w184 & ~w75;
assign w36 = pi051 & ~w371;
assign w37 = w95 & w380;
assign w38 = ~w52 & ~w255;
assign w39 = pi022 & ~w179;
assign w40 = (pi088 & ~w371) | (pi088 & w239) | (~w371 & w239);
assign w41 = ~w77 & ~w73;
assign w42 = w184 & ~w344;
assign w43 = pi074 & w333;
assign w44 = pi046 & ~w371;
assign w45 = ~pi094 & ~w187;
assign w46 = pi038 & ~w371;
assign w47 = ~w227 & w6;
assign w48 = ~w60 & ~w292;
assign w49 = ~pi090 & w93;
assign w50 = pi040 & ~w371;
assign w51 = ~w193 & w257;
assign w52 = pi032 & pi092;
assign w53 = pi053 & ~w95;
assign w54 = w184 & ~w173;
assign w55 = (pi001 & ~w95) | (pi001 & w302) | (~w95 & w302);
assign w56 = ~w31 & ~w51;
assign w57 = ~w195 & w79;
assign w58 = pi015 & pi013;
assign w59 = pi029 & ~w179;
assign w60 = pi083 & w333;
assign w61 = ~pi059 & ~pi093;
assign w62 = pi100 & pi104;
assign w63 = pi064 & ~w93;
assign w64 = ~w272 & w54;
assign w65 = ~w209 & w91;
assign w66 = ~w163 & ~w340;
assign w67 = pi097 & pi105;
assign w68 = pi078 & ~pi104;
assign w69 = ~pi047 & pi088;
assign w70 = w82 & w14;
assign w71 = ~w101 & w236;
assign w72 = pi015 & pi006;
assign w73 = pi083 & ~pi104;
assign w74 = (pi010 & ~w95) | (pi010 & w229) | (~w95 & w229);
assign w75 = w95 & w99;
assign w76 = pi095 & ~w138;
assign w77 = pi096 & pi104;
assign w78 = pi060 & ~w95;
assign w79 = (pi088 & ~w179) | (pi088 & w125) | (~w179 & w125);
assign w80 = pi103 & pi105;
assign w81 = pi021 & ~w179;
assign w82 = pi036 & w299;
assign w83 = pi015 & pi009;
assign w84 = pi037 & ~w371;
assign w85 = w95 & w277;
assign w86 = ~pi015 & pi007;
assign w87 = pi068 & w333;
assign w88 = pi082 & ~pi104;
assign w89 = (~pi034 & ~w37) | (~pi034 & w359) | (~w37 & w359);
assign w90 = (pi088 & ~w179) | (pi088 & w320) | (~w179 & w320);
assign w91 = w184 & ~w268;
assign w92 = pi015 & ~pi014;
assign w93 = pi067 & ~pi084;
assign w94 = ~pi060 & pi093;
assign w95 = ~pi067 & pi084;
assign w96 = pi019 & pi092;
assign w97 = (pi088 & ~w371) | (pi088 & w320) | (~w371 & w320);
assign w98 = (pi088 & ~w179) | (pi088 & w383) | (~w179 & w383);
assign w99 = pi015 & pi001;
assign w100 = pi094 & ~w200;
assign w101 = pi043 & ~w371;
assign w102 = ~w145 & w183;
assign w103 = (pi088 & ~w371) | (pi088 & w69) | (~w371 & w69);
assign w104 = ~pi037 & pi088;
assign w105 = ~w160 & ~w106;
assign w106 = pi071 & ~pi105;
assign w107 = pi018 & pi092;
assign w108 = ~pi015 & pi005;
assign w109 = (~pi035 & ~w95) | (~pi035 & w226) | (~w95 & w226);
assign w110 = pi080 & ~pi105;
assign w111 = pi026 & ~pi092;
assign w112 = ~w32 & ~w49;
assign w113 = ~w346 & ~w364;
assign w114 = pi074 & ~pi105;
assign w115 = w95 & w341;
assign w116 = ~pi043 & pi088;
assign w117 = pi025 & ~pi092;
assign w118 = ~w186 & w347;
assign w119 = (pi088 & ~w179) | (pi088 & w288) | (~w179 & w288);
assign w120 = ~pi061 & ~pi093;
assign w121 = ~pi015 & pi012;
assign w122 = pi041 & ~w371;
assign w123 = ~w353 & ~w190;
assign w124 = w10 & w82;
assign w125 = ~pi038 & pi088;
assign w126 = pi072 & w333;
assign w127 = ~w254 & ~w271;
assign w128 = ~w339 & ~w335;
assign w129 = pi057 & ~w95;
assign w130 = pi052 & ~w371;
assign w131 = ~w55 & w28;
assign w132 = ~w43 & ~w167;
assign w133 = ~w304 & w252;
assign w134 = ~pi015 & pi004;
assign w135 = ~w202 & ~w208;
assign w136 = pi049 & ~w371;
assign w137 = ~w70 & w378;
assign w138 = ~w263 & ~w26;
assign w139 = pi024 & ~w179;
assign w140 = pi054 & ~w95;
assign w141 = ~w46 & w97;
assign w142 = ~pi015 & pi006;
assign w143 = pi023 & ~pi092;
assign w144 = ~w223 & w369;
assign w145 = pi030 & ~w179;
assign w146 = (pi088 & ~w179) | (pi088 & w116) | (~w179 & w116);
assign w147 = ~w67 & ~w249;
assign w148 = ~pi015 & pi003;
assign w149 = (pi088 & ~w179) | (pi088 & w354) | (~w179 & w354);
assign w150 = pi098 & pi104;
assign w151 = ~w316 & ~w143;
assign w152 = ~w324 & w357;
assign w153 = ~w205 & ~w375;
assign w154 = ~w333 & ~w137;
assign w155 = ~w232 & ~w30;
assign w156 = ~pi095 & ~w222;
assign w157 = pi094 & ~w269;
assign w158 = ~pi046 & pi088;
assign w159 = pi099 & pi104;
assign w160 = pi102 & pi105;
assign w161 = w184 & ~w185;
assign w162 = pi015 & pi005;
assign w163 = pi078 & w333;
assign w164 = pi102 & pi104;
assign w165 = ~pi015 & pi009;
assign w166 = pi055 & ~w95;
assign w167 = ~w74 & w33;
assign w168 = (~pi000 & ~w95) | (~pi000 & w211) | (~w95 & w211);
assign w169 = ~pi015 & ~pi053;
assign w170 = (pi088 & ~w371) | (pi088 & w17) | (~w371 & w17);
assign w171 = (pi004 & ~w95) | (pi004 & w134) | (~w95 & w134);
assign w172 = ~pi015 & pi002;
assign w173 = w95 & w162;
assign w174 = pi101 & pi104;
assign w175 = ~w130 & w181;
assign w176 = ~w7 & w149;
assign w177 = pi079 & w333;
assign w178 = (pi088 & ~w371) | (pi088 & w368) | (~w371 & w368);
assign w179 = w95 & w313;
assign w180 = ~w122 & w225;
assign w181 = (pi088 & ~w371) | (pi088 & w383) | (~w371 & w383);
assign w182 = pi054 & w95;
assign w183 = (pi088 & ~w179) | (pi088 & w17) | (~w179 & w17);
assign w184 = ~pi062 & pi088;
assign w185 = w95 & w323;
assign w186 = pi025 & ~w179;
assign w187 = ~pi056 & pi093;
assign w188 = ~pi015 & ~pi016;
assign w189 = ~pi036 & ~w37;
assign w190 = pi076 & ~pi104;
assign w191 = ~w373 & w301;
assign w192 = ~w16 & ~w191;
assign w193 = (pi012 & ~w95) | (pi012 & w121) | (~w95 & w121);
assign w194 = (pi088 & ~w371) | (pi088 & w315) | (~w371 & w315);
assign w195 = pi031 & ~w179;
assign w196 = ~w321 & ~w273;
assign w197 = ~w338 & ~w199;
assign w198 = w184 & ~w240;
assign w199 = pi029 & ~pi092;
assign w200 = ~pi054 & ~pi093;
assign w201 = w95 & w83;
assign w202 = pi058 & ~w95;
assign w203 = pi015 & pi008;
assign w204 = ~w336 & w24;
assign w205 = pi101 & pi105;
assign w206 = pi099 & pi105;
assign w207 = ~w201 & w352;
assign w208 = pi055 & w95;
assign w209 = (pi011 & ~w95) | (pi011 & w19) | (~w95 & w19);
assign w210 = (pi002 & ~w95) | (pi002 & w172) | (~w95 & w172);
assign w211 = ~pi015 & ~pi000;
assign w212 = ~w129 & ~w261;
assign w213 = ~w126 & ~w267;
assign w214 = ~w94 & w100;
assign w215 = pi023 & ~w179;
assign w216 = (pi008 & ~w95) | (pi008 & w217) | (~w95 & w217);
assign w217 = ~pi015 & pi008;
assign w218 = ~pi063 & w95;
assign w219 = ~w44 & w367;
assign w220 = ~w382 & w327;
assign w221 = w95 & w298;
assign w222 = ~w214 & ~w286;
assign w223 = pi020 & ~w179;
assign w224 = ~w78 & ~w182;
assign w225 = (pi088 & ~w371) | (pi088 & w325) | (~w371 & w325);
assign w226 = ~pi015 & ~pi035;
assign w227 = pi042 & ~w371;
assign w228 = (pi088 & ~w179) | (pi088 & w368) | (~w179 & w368);
assign w229 = ~pi015 & pi010;
assign w230 = w184 & ~w296;
assign w231 = pi056 & w95;
assign w232 = pi103 & pi104;
assign w233 = pi015 & ~pi016;
assign w234 = pi056 & ~w95;
assign w235 = pi071 & w333;
assign w236 = (pi088 & ~w371) | (pi088 & w354) | (~w371 & w354);
assign w237 = pi059 & ~w95;
assign w238 = (pi088 & ~w179) | (pi088 & w315) | (~w179 & w315);
assign w239 = ~pi039 & pi088;
assign w240 = w95 & w203;
assign w241 = w184 & ~w5;
assign w242 = ~pi091 & w93;
assign w243 = ~w59 & w303;
assign w244 = ~pi055 & pi093;
assign w245 = pi070 & w333;
assign w246 = ~w379 & ~w64;
assign w247 = ~w174 & ~w396;
assign w248 = pi060 & w95;
assign w249 = pi072 & ~pi105;
assign w250 = ~w350 & ~w9;
assign w251 = (pi013 & ~w95) | (pi013 & w360) | (~w95 & w360);
assign w252 = (pi088 & ~w179) | (pi088 & w325) | (~w179 & w325);
assign w253 = ~w1 & w178;
assign w254 = pi017 & pi092;
assign w255 = pi022 & ~pi092;
assign w256 = ~w96 & ~w111;
assign w257 = w184 & ~w85;
assign w258 = ~w295 & w42;
assign w259 = ~pi044 & pi088;
assign w260 = (pi088 & ~w371) | (pi088 & w104) | (~w371 & w104);
assign w261 = pi058 & w95;
assign w262 = (pi088 & ~w371) | (pi088 & w259) | (~w371 & w259);
assign w263 = ~w266 & w157;
assign w264 = ~pi033 & ~w124;
assign w265 = ~w150 & ~w281;
assign w266 = ~pi057 & pi093;
assign w267 = ~w343 & w198;
assign w268 = w95 & w4;
assign w269 = ~pi058 & ~pi093;
assign w270 = pi073 & w333;
assign w271 = pi024 & ~pi092;
assign w272 = (pi006 & ~w95) | (pi006 & w142) | (~w95 & w142);
assign w273 = pi073 & ~pi105;
assign w274 = pi069 & ~pi105;
assign w275 = pi039 & ~w371;
assign w276 = ~pi036 & pi088;
assign w277 = pi015 & pi011;
assign w278 = ~w308 & w146;
assign w279 = ~w140 & ~w231;
assign w280 = pi088 & ~w37;
assign w281 = pi077 & ~pi104;
assign w282 = ~w50 & w388;
assign w283 = pi015 & pi012;
assign w284 = ~w139 & w330;
assign w285 = w95 & w92;
assign w286 = ~w61 & w45;
assign w287 = ~w136 & w262;
assign w288 = ~pi045 & pi088;
assign w289 = pi082 & w333;
assign w290 = ~w264 & ~w384;
assign w291 = w184 & ~w115;
assign w292 = ~w10 & w381;
assign w293 = ~w289 & ~w152;
assign w294 = pi076 & w333;
assign w295 = (pi007 & ~w95) | (pi007 & w86) | (~w95 & w86);
assign w296 = w95 & w283;
assign w297 = pi061 & ~w95;
assign w298 = pi015 & pi002;
assign w299 = pi034 & pi035;
assign w300 = ~w36 & w170;
assign w301 = w184 & ~w168;
assign w302 = ~pi015 & pi001;
assign w303 = (pi088 & ~w179) | (pi088 & w239) | (~w179 & w239);
assign w304 = pi032 & ~w179;
assign w305 = ~w311 & w161;
assign w306 = pi048 & ~w371;
assign w307 = ~w275 & w2;
assign w308 = pi019 & ~w179;
assign w309 = ~w366 & ~w12;
assign w310 = pi081 & ~pi104;
assign w311 = (pi005 & ~w95) | (pi005 & w108) | (~w95 & w108);
assign w312 = ~w76 & ~w156;
assign w313 = ~pi015 & pi053;
assign w314 = ~w329 & w103;
assign w315 = ~pi050 & pi088;
assign w316 = pi030 & pi092;
assign w317 = ~w63 & ~w242;
assign w318 = pi027 & ~w179;
assign w319 = ~w159 & ~w88;
assign w320 = ~pi048 & pi088;
assign w321 = pi098 & pi105;
assign w322 = ~w251 & w230;
assign w323 = pi015 & pi004;
assign w324 = (pi003 & ~w95) | (pi003 & w148) | (~w95 & w148);
assign w325 = ~pi040 & pi088;
assign w326 = ~w107 & ~w117;
assign w327 = (pi088 & ~w371) | (pi088 & w158) | (~w371 & w158);
assign w328 = pi031 & pi092;
assign w329 = pi050 & ~w371;
assign w330 = (pi088 & ~w179) | (pi088 & w158) | (~w179 & w158);
assign w331 = ~w166 & ~w345;
assign w332 = (pi088 & ~w37) | (pi088 & w276) | (~w37 & w276);
assign w333 = pi062 & pi088;
assign w334 = w390 & ~w89;
assign w335 = pi020 & ~pi092;
assign w336 = pi017 & ~w179;
assign w337 = pi015 & pi003;
assign w338 = pi027 & pi092;
assign w339 = pi028 & pi092;
assign w340 = ~w171 & w241;
assign w341 = pi015 & pi007;
assign w342 = w95 & w233;
assign w343 = (pi009 & ~w95) | (pi009 & w165) | (~w95 & w165);
assign w344 = w95 & w72;
assign w345 = pi061 & w95;
assign w346 = pi100 & pi105;
assign w347 = (pi088 & ~w179) | (pi088 & w69) | (~w179 & w69);
assign w348 = ~pi051 & pi088;
assign w349 = (~pi016 & ~w95) | (~pi016 & w188) | (~w95 & w188);
assign w350 = pi077 & w333;
assign w351 = ~w245 & ~w65;
assign w352 = w184 & ~w349;
assign w353 = pi097 & pi104;
assign w354 = ~pi042 & pi088;
assign w355 = pi096 & pi105;
assign w356 = ~w235 & ~w322;
assign w357 = w184 & ~w221;
assign w358 = ~w355 & ~w110;
assign w359 = ~pi036 & ~pi034;
assign w360 = ~pi015 & pi013;
assign w361 = ~w318 & w392;
assign w362 = ~pi094 & ~w244;
assign w363 = ~w81 & w98;
assign w364 = pi070 & ~pi105;
assign w365 = ~w297 & ~w248;
assign w366 = pi080 & w333;
assign w367 = (pi088 & ~w371) | (pi088 & w288) | (~w371 & w288);
assign w368 = ~pi052 & pi088;
assign w369 = (pi088 & ~w179) | (pi088 & w259) | (~w179 & w259);
assign w370 = ~w206 & ~w114;
assign w371 = w93 & ~w169;
assign w372 = ~w306 & w260;
assign w373 = w95 & w58;
assign w374 = ~w22 & w40;
assign w375 = pi075 & ~pi105;
assign w376 = ~pi065 & ~pi066;
assign w377 = pi028 & ~w179;
assign w378 = pi015 & pi088;
assign w379 = pi081 & w333;
assign w380 = pi015 & pi035;
assign w381 = pi014 & w184;
assign w382 = pi047 & ~w371;
assign w383 = ~pi049 & pi088;
assign w384 = ~w137 & ~w390;
assign w385 = ~w294 & ~w131;
assign w386 = ~w215 & w119;
assign w387 = ~w109 & w280;
assign w388 = (pi088 & ~w371) | (pi088 & w125) | (~w371 & w125);
assign w389 = ~w84 & w194;
assign w390 = pi088 & ~w124;
assign w391 = ~w237 & ~w218;
assign w392 = (pi088 & ~w179) | (pi088 & w104) | (~w179 & w104);
assign w393 = pi059 & w95;
assign w394 = ~w377 & w90;
assign w395 = ~w62 & ~w68;
assign w396 = pi068 & ~pi104;
assign one = 1;
assign po00 = pi000;// level 0
assign po01 = w197;// level 2
assign po02 = w128;// level 2
assign po03 = w25;// level 2
assign po04 = w38;// level 2
assign po05 = w151;// level 2
assign po06 = w127;// level 2
assign po07 = w326;// level 2
assign po08 = w256;// level 2
assign po09 = pi087;// level 0
assign po10 = ~w192;// level 5
assign po11 = ~w385;// level 5
assign po12 = ~w250;// level 5
assign po13 = ~w293;// level 5
assign po14 = ~w66;// level 5
assign po15 = ~w29;// level 5
assign po16 = ~w246;// level 5
assign po17 = ~w3;// level 5
assign po18 = ~w309;// level 5
assign po19 = ~w213;// level 5
assign po20 = ~w132;// level 5
assign po21 = ~w351;// level 5
assign po22 = ~w56;// level 5
assign po23 = ~w356;// level 5
assign po24 = ~w48;// level 4
assign po25 = one;// level 0
assign po26 = ~w154;// level 5
assign po27 = ~w20;// level 5
assign po28 = w204;// level 4
assign po29 = w176;// level 4
assign po30 = w278;// level 4
assign po31 = w144;// level 4
assign po32 = w363;// level 4
assign po33 = w13;// level 4
assign po34 = w386;// level 4
assign po35 = w284;// level 4
assign po36 = w118;// level 4
assign po37 = w21;// level 4
assign po38 = w361;// level 4
assign po39 = w394;// level 4
assign po40 = w243;// level 4
assign po41 = w102;// level 4
assign po42 = w57;// level 4
assign po43 = w133;// level 4
assign po44 = w290;// level 6
assign po45 = w334;// level 5
assign po46 = w387;// level 4
assign po47 = w23;// level 4
assign po48 = w389;// level 4
assign po49 = w141;// level 4
assign po50 = w307;// level 4
assign po51 = w282;// level 4
assign po52 = w180;// level 4
assign po53 = w47;// level 4
assign po54 = w71;// level 4
assign po55 = w374;// level 4
assign po56 = w253;// level 4
assign po57 = w219;// level 4
assign po58 = w220;// level 4
assign po59 = w372;// level 4
assign po60 = w287;// level 4
assign po61 = w314;// level 4
assign po62 = w300;// level 4
assign po63 = w175;// level 4
assign po64 = ~w27;// level 3
assign po65 = ~w279;// level 3
assign po66 = ~w331;// level 3
assign po67 = ~w18;// level 3
assign po68 = ~w212;// level 3
assign po69 = ~w135;// level 3
assign po70 = ~w391;// level 3
assign po71 = ~w224;// level 3
assign po72 = ~w365;// level 3
assign po73 = w376;// level 1
assign po74 = w112;// level 3
assign po75 = w317;// level 3
assign po76 = ~pi066;// level 0
assign po77 = ~w312;// level 6
assign po78 = pi084;// level 0
assign po79 = ~w247;// level 2
assign po80 = ~w34;// level 2
assign po81 = ~w113;// level 2
assign po82 = ~w105;// level 2
assign po83 = ~w147;// level 2
assign po84 = ~w196;// level 2
assign po85 = ~w370;// level 2
assign po86 = ~w153;// level 2
assign po87 = ~w123;// level 2
assign po88 = ~w265;// level 2
assign po89 = ~w395;// level 2
assign po90 = ~w155;// level 2
assign po91 = ~w358;// level 2
assign po92 = ~w15;// level 2
assign po93 = ~w319;// level 2
assign po94 = ~w41;// level 2
assign po95 = pi086;// level 0
assign po96 = ~pi064;// level 0
assign po97 = pi089;// level 0
endmodule
