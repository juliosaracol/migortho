module top (
            pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, 
            po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24);
input pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19;
output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23, po24;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515;
assign w0 = pi01 & ~pi02;
assign w1 = (~pi04 & w0) | (~pi04 & w6577) | (w0 & w6577);
assign w2 = ~pi07 & ~pi08;
assign w3 = ~pi06 & w2;
assign w4 = ~pi17 & ~pi18;
assign w5 = ~pi13 & ~pi19;
assign w6 = w4 & w5;
assign w7 = ~pi15 & ~pi16;
assign w8 = ~pi12 & ~pi14;
assign w9 = w7 & w8;
assign w10 = w6 & w9;
assign w11 = ~pi11 & ~pi12;
assign w12 = ~pi09 & ~pi10;
assign w13 = w11 & w12;
assign w14 = w10 & w13;
assign w15 = w2 & w6578;
assign w16 = w10 & w6579;
assign w17 = ~w1 & w16;
assign w18 = ~pi10 & ~pi11;
assign w19 = ~pi08 & ~pi09;
assign w20 = w18 & w19;
assign w21 = pi06 & w2;
assign w22 = w10 & w6580;
assign w23 = pi13 & ~pi14;
assign w24 = ~pi19 & w4;
assign w25 = w7 & w24;
assign w26 = w24 & w6047;
assign w27 = pi16 & ~pi19;
assign w28 = pi15 & ~pi18;
assign w29 = ~pi19 & ~w28;
assign w30 = pi17 & ~pi18;
assign w31 = pi11 & ~pi12;
assign w32 = pi09 & ~pi12;
assign w33 = w18 & w32;
assign w34 = ~w31 & ~w33;
assign w35 = ~pi16 & ~pi19;
assign w36 = w4 & w35;
assign w37 = ~pi13 & ~pi14;
assign w38 = ~pi15 & w37;
assign w39 = w36 & w38;
assign w40 = ~w34 & w39;
assign w41 = (~w30 & w29) | (~w30 & w6581) | (w29 & w6581);
assign w42 = ~w26 & w41;
assign w43 = ~w40 & w42;
assign w44 = ~w22 & w43;
assign w45 = ~w17 & ~w44;
assign w46 = ~pi03 & ~pi04;
assign w47 = w16 & w46;
assign w48 = ~pi01 & ~pi02;
assign w49 = ~pi00 & w48;
assign w50 = w16 & w6582;
assign w51 = ~w45 & ~w50;
assign w52 = w16 & w6583;
assign w53 = ~pi19 & ~w4;
assign w54 = ~w11 & w37;
assign w55 = (~w53 & ~w25) | (~w53 & w6584) | (~w25 & w6584);
assign w56 = ~w2 & w14;
assign w57 = ~w16 & ~w55;
assign w58 = ~w56 & w57;
assign w59 = ~w52 & ~w58;
assign w60 = w11 & w37;
assign w61 = w10 & w6585;
assign w62 = (~pi19 & ~w25) | (~pi19 & w6586) | (~w25 & w6586);
assign w63 = ~w61 & w62;
assign w64 = ~w47 & ~w63;
assign w65 = w25 & ~w61;
assign w66 = ~pi14 & ~pi15;
assign w67 = pi04 & ~pi13;
assign w68 = w66 & w67;
assign w69 = pi07 & pi15;
assign w70 = pi05 & ~pi15;
assign w71 = w23 & w70;
assign w72 = pi06 & ~pi15;
assign w73 = pi14 & w72;
assign w74 = ~w68 & ~w69;
assign w75 = ~w71 & ~w73;
assign w76 = w74 & w75;
assign w77 = w36 & ~w76;
assign w78 = w30 & w6048;
assign w79 = pi11 & pi19;
assign w80 = pi18 & ~pi19;
assign w81 = pi10 & w80;
assign w82 = w4 & w27;
assign w83 = pi08 & w82;
assign w84 = ~w79 & ~w81;
assign w85 = ~w78 & w84;
assign w86 = ~w83 & w85;
assign w87 = ~w77 & w86;
assign w88 = ~w10 & ~w87;
assign w89 = pi03 & ~pi15;
assign w90 = w37 & w89;
assign w91 = w36 & w90;
assign w92 = w31 & w91;
assign w93 = pi00 & pi08;
assign w94 = w10 & w6049;
assign w95 = pi10 & w11;
assign w96 = pi02 & w39;
assign w97 = w39 & w6050;
assign w98 = pi01 & w39;
assign w99 = w39 & w6051;
assign w100 = ~w92 & ~w94;
assign w101 = ~w97 & ~w99;
assign w102 = w100 & w101;
assign w103 = ~w88 & w102;
assign w104 = w37 & w70;
assign w105 = w36 & w104;
assign w106 = pi12 & pi19;
assign w107 = pi11 & w80;
assign w108 = w30 & w6052;
assign w109 = pi09 & w82;
assign w110 = pi15 & w36;
assign w111 = w36 & w6053;
assign w112 = pi14 & w36;
assign w113 = pi07 & ~pi15;
assign w114 = w36 & w6054;
assign w115 = ~w106 & ~w107;
assign w116 = ~w105 & w115;
assign w117 = ~w108 & ~w109;
assign w118 = w116 & w117;
assign w119 = ~w111 & ~w114;
assign w120 = (~w10 & ~w118) | (~w10 & w6055) | (~w118 & w6055);
assign w121 = pi07 & w19;
assign w122 = w19 & w6056;
assign w123 = pi04 & pi11;
assign w124 = pi02 & pi09;
assign w125 = ~w123 & ~w124;
assign w126 = ~w122 & w125;
assign w127 = ~w18 & ~w123;
assign w128 = w10 & ~w127;
assign w129 = ~w126 & w128;
assign w130 = pi01 & ~pi09;
assign w131 = pi08 & ~pi16;
assign w132 = w66 & w131;
assign w133 = w6 & w132;
assign w134 = ~pi12 & w18;
assign w135 = w133 & w6587;
assign w136 = w91 & w95;
assign w137 = w36 & w6057;
assign w138 = ~w136 & ~w137;
assign w139 = ~w129 & w138;
assign w140 = ~w135 & w139;
assign w141 = ~w120 & w140;
assign w142 = w103 & w141;
assign w143 = w24 & w6058;
assign w144 = w10 & w6588;
assign w145 = (pi08 & w144) | (pi08 & w6589) | (w144 & w6589);
assign w146 = pi06 & ~pi13;
assign w147 = w66 & w146;
assign w148 = w36 & w147;
assign w149 = pi10 & w82;
assign w150 = pi13 & pi19;
assign w151 = w30 & w6059;
assign w152 = ~w148 & ~w150;
assign w153 = ~w149 & ~w151;
assign w154 = w152 & w153;
assign w155 = ~w10 & ~w154;
assign w156 = w36 & w6060;
assign w157 = w36 & w68;
assign w158 = w95 & w157;
assign w159 = w36 & w6061;
assign w160 = w13 & w21;
assign w161 = pi00 & w39;
assign w162 = w160 & w161;
assign w163 = w10 & w18;
assign w164 = pi03 & pi09;
assign w165 = w19 & w6590;
assign w166 = ~w164 & ~w165;
assign w167 = w163 & ~w166;
assign w168 = w31 & w105;
assign w169 = pi12 & w80;
assign w170 = ~w156 & ~w169;
assign w171 = ~w158 & ~w159;
assign w172 = ~w168 & w171;
assign w173 = ~w162 & w170;
assign w174 = ~w167 & w173;
assign w175 = ~w155 & w172;
assign w176 = w174 & w175;
assign w177 = ~w145 & w176;
assign w178 = ~w142 & w177;
assign w179 = w142 & ~w177;
assign w180 = ~w178 & ~w179;
assign w181 = w36 & w6062;
assign w182 = ~w110 & ~w181;
assign w183 = ~pi11 & pi15;
assign w184 = pi10 & w143;
assign w185 = pi15 & pi19;
assign w186 = pi14 & w80;
assign w187 = pi12 & w82;
assign w188 = w30 & w6063;
assign w189 = ~w185 & ~w186;
assign w190 = ~w133 & w189;
assign w191 = ~w187 & ~w188;
assign w192 = w190 & w191;
assign w193 = ~w184 & w192;
assign w194 = (~w10 & ~w193) | (~w10 & w6064) | (~w193 & w6064);
assign w195 = pi04 & ~pi05;
assign w196 = pi00 & w195;
assign w197 = w16 & ~w196;
assign w198 = w95 & w148;
assign w199 = w13 & w24;
assign w200 = w68 & w131;
assign w201 = w199 & w200;
assign w202 = w33 & w105;
assign w203 = w121 & w134;
assign w204 = w91 & w203;
assign w205 = pi07 & w39;
assign w206 = w39 & w6065;
assign w207 = w3 & w196;
assign w208 = ~pi01 & ~pi06;
assign w209 = ~pi02 & pi06;
assign w210 = w2 & ~w208;
assign w211 = ~w209 & w210;
assign w212 = ~w207 & ~w211;
assign w213 = w14 & ~w212;
assign w214 = ~w198 & ~w201;
assign w215 = ~w202 & ~w204;
assign w216 = w214 & w215;
assign w217 = ~w206 & ~w213;
assign w218 = w216 & w217;
assign w219 = ~w197 & ~w218;
assign w220 = ~w194 & ~w219;
assign w221 = pi03 & pi08;
assign w222 = w2 & w6066;
assign w223 = ~w221 & ~w222;
assign w224 = w14 & ~w223;
assign w225 = w33 & w157;
assign w226 = w95 & w105;
assign w227 = w2 & w130;
assign w228 = w134 & w227;
assign w229 = ~w31 & ~w228;
assign w230 = w148 & ~w229;
assign w231 = pi02 & pi07;
assign w232 = w10 & w6067;
assign w233 = ~w225 & ~w226;
assign w234 = ~w224 & w233;
assign w235 = ~w230 & ~w232;
assign w236 = w234 & w235;
assign w237 = ~w16 & ~w236;
assign w238 = w36 & w6068;
assign w239 = pi14 & pi19;
assign w240 = pi13 & w80;
assign w241 = pi11 & w82;
assign w242 = ~pi09 & pi14;
assign w243 = ~pi08 & ~pi14;
assign w244 = ~w37 & ~w242;
assign w245 = ~w243 & w244;
assign w246 = w25 & w245;
assign w247 = w30 & w6591;
assign w248 = ~w239 & ~w240;
assign w249 = ~w241 & w248;
assign w250 = ~w205 & ~w238;
assign w251 = ~w246 & w250;
assign w252 = (~w10 & ~w251) | (~w10 & w6069) | (~w251 & w6069);
assign w253 = ~w237 & ~w252;
assign w254 = w177 & ~w253;
assign w255 = w142 & w254;
assign w256 = w177 & w253;
assign w257 = w142 & w256;
assign w258 = (w253 & ~w256) | (w253 & w6592) | (~w256 & w6592);
assign w259 = ~w255 & ~w258;
assign w260 = ~w220 & ~w259;
assign w261 = pi03 & w160;
assign w262 = (~w31 & ~w13) | (~w31 & w6328) | (~w13 & w6328);
assign w263 = pi08 & ~w262;
assign w264 = pi06 & w33;
assign w265 = w11 & w6329;
assign w266 = ~w264 & ~w265;
assign w267 = ~w261 & w266;
assign w268 = (w39 & ~w267) | (w39 & w6330) | (~w267 & w6330);
assign w269 = pi09 & w39;
assign w270 = (pi12 & w269) | (pi12 & w6070) | (w269 & w6070);
assign w271 = w157 & w203;
assign w272 = w30 & w6071;
assign w273 = pi15 & w80;
assign w274 = pi16 & ~w5;
assign w275 = ~w53 & w274;
assign w276 = pi10 & w26;
assign w277 = pi11 & w143;
assign w278 = pi01 & w195;
assign w279 = (~pi02 & ~w195) | (~pi02 & w48) | (~w195 & w48);
assign w280 = w3 & ~w279;
assign w281 = w14 & w280;
assign w282 = ~pi04 & pi05;
assign w283 = ~pi06 & ~pi07;
assign w284 = ~w282 & w283;
assign w285 = pi00 & ~pi04;
assign w286 = ~pi12 & w285;
assign w287 = w20 & w286;
assign w288 = w284 & w287;
assign w289 = w91 & w288;
assign w290 = ~w272 & ~w273;
assign w291 = ~w275 & w290;
assign w292 = ~w271 & w291;
assign w293 = ~w276 & ~w277;
assign w294 = ~w281 & ~w289;
assign w295 = w293 & w294;
assign w296 = ~w270 & w292;
assign w297 = w295 & w296;
assign w298 = w14 & w6331;
assign w299 = ~w289 & w298;
assign w300 = (~w299 & ~w295) | (~w299 & w6332) | (~w295 & w6332);
assign w301 = (~w268 & w297) | (~w268 & w6072) | (w297 & w6072);
assign w302 = w142 & w220;
assign w303 = w256 & w302;
assign w304 = w301 & ~w303;
assign w305 = ~w301 & w303;
assign w306 = ~w304 & ~w305;
assign w307 = ~w141 & ~w306;
assign w308 = ~w103 & w301;
assign w309 = w301 & w303;
assign w310 = (pi17 & w28) | (pi17 & w6333) | (w28 & w6333);
assign w311 = w146 & w199;
assign w312 = (~w95 & ~w199) | (~w95 & w6334) | (~w199 & w6334);
assign w313 = w133 & ~w312;
assign w314 = pi05 & ~pi08;
assign w315 = (pi07 & w314) | (pi07 & w6335) | (w314 & w6335);
assign w316 = ~pi03 & pi05;
assign w317 = ~pi09 & ~w316;
assign w318 = w3 & w317;
assign w319 = ~w315 & ~w318;
assign w320 = w163 & ~w319;
assign w321 = pi14 & ~pi17;
assign w322 = ~pi18 & ~w321;
assign w323 = w27 & ~w322;
assign w324 = w36 & w6336;
assign w325 = pi10 & w39;
assign w326 = (pi12 & w325) | (pi12 & w6337) | (w325 & w6337);
assign w327 = (pi11 & w32) | (pi11 & w6593) | (w32 & w6593);
assign w328 = w67 & w160;
assign w329 = w36 & w66;
assign w330 = (w329 & w328) | (w329 & w6338) | (w328 & w6338);
assign w331 = ~w310 & ~w323;
assign w332 = ~w324 & w331;
assign w333 = ~w320 & w332;
assign w334 = ~w313 & w333;
assign w335 = ~w326 & ~w330;
assign w336 = pi00 & ~pi03;
assign w337 = (pi02 & w336) | (pi02 & w6594) | (w336 & w6594);
assign w338 = pi01 & ~pi04;
assign w339 = pi03 & w338;
assign w340 = ~w337 & ~w339;
assign w341 = w16 & w340;
assign w342 = (~w341 & ~w334) | (~w341 & w6339) | (~w334 & w6339);
assign w343 = pi10 & pi19;
assign w344 = pi09 & w80;
assign w345 = w30 & w6073;
assign w346 = pi07 & w82;
assign w347 = w36 & w6074;
assign w348 = w36 & w6075;
assign w349 = ~w343 & ~w344;
assign w350 = ~w91 & w349;
assign w351 = ~w345 & ~w346;
assign w352 = w350 & w351;
assign w353 = ~w347 & ~w348;
assign w354 = (~w10 & ~w352) | (~w10 & w6076) | (~w352 & w6076);
assign w355 = pi04 & w26;
assign w356 = pi02 & pi11;
assign w357 = pi00 & pi09;
assign w358 = w18 & w357;
assign w359 = ~w356 & ~w358;
assign w360 = w10 & ~w359;
assign w361 = w39 & w6595;
assign w362 = ~w355 & ~w360;
assign w363 = ~w361 & w362;
assign w364 = ~w354 & w363;
assign w365 = ~w342 & ~w364;
assign w366 = (w365 & ~w303) | (w365 & w6077) | (~w303 & w6077);
assign w367 = ~w268 & ~w364;
assign w368 = ~w300 & w367;
assign w369 = w342 & w368;
assign w370 = w303 & w369;
assign w371 = ~w366 & ~w370;
assign w372 = w308 & ~w371;
assign w373 = ~w307 & ~w372;
assign w374 = ~w141 & ~w342;
assign w375 = ~w103 & ~w364;
assign w376 = w374 & w375;
assign w377 = ~w303 & w6596;
assign w378 = ~w373 & ~w377;
assign w379 = ~w336 & w6597;
assign w380 = ~pi03 & ~w338;
assign w381 = ~w379 & ~w380;
assign w382 = w16 & ~w381;
assign w383 = w10 & w6340;
assign w384 = ~w31 & ~w32;
assign w385 = w39 & w6341;
assign w386 = ~pi07 & ~pi09;
assign w387 = w133 & w6342;
assign w388 = ~pi05 & ~pi07;
assign w389 = w7 & w243;
assign w390 = ~w388 & w389;
assign w391 = w311 & w390;
assign w392 = ~w383 & ~w385;
assign w393 = ~w387 & ~w391;
assign w394 = w392 & w393;
assign w395 = ~w28 & w6598;
assign w396 = ~pi18 & ~w27;
assign w397 = (~w395 & w112) | (~w395 & w6599) | (w112 & w6599);
assign w398 = pi11 & ~pi14;
assign w399 = ~pi13 & ~w398;
assign w400 = ~w8 & ~w399;
assign w401 = w25 & w400;
assign w402 = ~w397 & ~w401;
assign w403 = (w402 & w394) | (w402 & w6343) | (w394 & w6343);
assign w404 = ~w268 & ~w342;
assign w405 = w256 & w6344;
assign w406 = w220 & ~w300;
assign w407 = w257 & w6078;
assign w408 = ~w403 & ~w407;
assign w409 = w220 & w6600;
assign w410 = w405 & w409;
assign w411 = (~w364 & ~w405) | (~w364 & w6079) | (~w405 & w6079);
assign w412 = ~w408 & w411;
assign w413 = ~w103 & ~w342;
assign w414 = ~w408 & w6345;
assign w415 = (~w413 & w408) | (~w413 & w6346) | (w408 & w6346);
assign w416 = ~w414 & ~w415;
assign w417 = w378 & ~w416;
assign w418 = ~w378 & w416;
assign w419 = ~w417 & ~w418;
assign w420 = ~w103 & w220;
assign w421 = ~w219 & w6347;
assign w422 = w256 & w6348;
assign w423 = ~w368 & ~w420;
assign w424 = ~w422 & w423;
assign w425 = w308 & w421;
assign w426 = ~w309 & ~w425;
assign w427 = ~w424 & w426;
assign w428 = ~w103 & w253;
assign w429 = w421 & w428;
assign w430 = ~w141 & w253;
assign w431 = ~w429 & ~w430;
assign w432 = w428 & w6349;
assign w433 = ~w431 & ~w432;
assign w434 = w427 & w433;
assign w435 = ~w177 & w253;
assign w436 = ~w432 & ~w435;
assign w437 = (w436 & ~w427) | (w436 & w6080) | (~w427 & w6080);
assign w438 = ~w141 & w220;
assign w439 = w308 & ~w421;
assign w440 = w438 & ~w439;
assign w441 = ~w438 & w439;
assign w442 = ~w440 & ~w441;
assign w443 = w371 & ~w442;
assign w444 = ~w371 & w442;
assign w445 = ~w443 & ~w444;
assign w446 = ~w437 & ~w445;
assign w447 = w425 & ~w432;
assign w448 = (w435 & w429) | (w435 & w6350) | (w429 & w6350);
assign w449 = ~w424 & w448;
assign w450 = ~w447 & w449;
assign w451 = (~w255 & ~w449) | (~w255 & w6601) | (~w449 & w6601);
assign w452 = ~w446 & w451;
assign w453 = w220 & w6351;
assign w454 = w308 & ~w453;
assign w455 = ~w371 & w454;
assign w456 = (~w308 & ~w303) | (~w308 & w6352) | (~w303 & w6352);
assign w457 = ~w425 & ~w438;
assign w458 = (~w457 & ~w456) | (~w457 & w6081) | (~w456 & w6081);
assign w459 = ~w455 & w458;
assign w460 = ~w177 & w459;
assign w461 = ~w177 & w220;
assign w462 = ~w459 & ~w461;
assign w463 = ~w460 & ~w462;
assign w464 = w452 & ~w463;
assign w465 = ~w452 & w463;
assign w466 = ~w464 & ~w465;
assign w467 = w419 & w466;
assign w468 = (~w452 & w419) | (~w452 & w6353) | (w419 & w6353);
assign w469 = ~w467 & w6354;
assign w470 = (~w260 & w467) | (~w260 & w6355) | (w467 & w6355);
assign w471 = ~w469 & ~w470;
assign w472 = ~w194 & w218;
assign w473 = ~w253 & w472;
assign w474 = w463 & w473;
assign w475 = ~w419 & w474;
assign w476 = w459 & w6602;
assign w477 = (~w473 & ~w459) | (~w473 & w6603) | (~w459 & w6603);
assign w478 = ~w476 & ~w477;
assign w479 = (~w478 & w419) | (~w478 & w6604) | (w419 & w6604);
assign w480 = ~w475 & ~w479;
assign w481 = ~w177 & w301;
assign w482 = w373 & ~w481;
assign w483 = ~w413 & ~w481;
assign w484 = (w483 & w408) | (w483 & w6356) | (w408 & w6356);
assign w485 = (w413 & ~w304) | (w413 & w6082) | (~w304 & w6082);
assign w486 = ~w481 & w485;
assign w487 = w412 & w486;
assign w488 = ~w484 & ~w487;
assign w489 = ~w482 & w488;
assign w490 = w412 & w485;
assign w491 = ~w177 & ~w373;
assign w492 = ~w415 & ~w490;
assign w493 = w491 & w492;
assign w494 = w489 & ~w493;
assign w495 = ~w103 & w403;
assign w496 = w364 & ~w495;
assign w497 = w374 & ~w496;
assign w498 = w364 & w495;
assign w499 = ~w374 & ~w498;
assign w500 = (w499 & ~w411) | (w499 & w6605) | (~w411 & w6605);
assign w501 = (~w497 & w414) | (~w497 & w6606) | (w414 & w6606);
assign w502 = ~w494 & w501;
assign w503 = w494 & ~w501;
assign w504 = ~w502 & ~w503;
assign w505 = ~w480 & w504;
assign w506 = w480 & ~w504;
assign w507 = ~w505 & ~w506;
assign w508 = w471 & w507;
assign w509 = ~w471 & ~w507;
assign w510 = ~w508 & ~w509;
assign w511 = ~w180 & ~w301;
assign w512 = ~w180 & ~w253;
assign w513 = w426 & w6357;
assign w514 = ~w427 & ~w433;
assign w515 = ~w434 & ~w514;
assign w516 = ~w141 & w177;
assign w517 = ~w103 & ~w141;
assign w518 = ~w420 & ~w517;
assign w519 = ~w516 & ~w518;
assign w520 = ~w375 & ~w517;
assign w521 = w256 & ~w520;
assign w522 = w177 & w453;
assign w523 = ~w179 & ~w521;
assign w524 = ~w522 & w523;
assign w525 = ~w519 & ~w524;
assign w526 = w426 & w6358;
assign w527 = w178 & ~w253;
assign w528 = ~w453 & w527;
assign w529 = (~w528 & w526) | (~w528 & w6607) | (w526 & w6607);
assign w530 = (w529 & ~w515) | (w529 & w7431) | (~w515 & w7431);
assign w531 = ~w437 & ~w450;
assign w532 = w445 & ~w531;
assign w533 = ~w445 & w531;
assign w534 = ~w532 & ~w533;
assign w535 = ~w530 & w534;
assign w536 = w513 & w525;
assign w537 = ~w180 & ~w220;
assign w538 = ~w536 & ~w537;
assign w539 = (w538 & ~w534) | (w538 & w7432) | (~w534 & w7432);
assign w540 = ~w220 & w536;
assign w541 = (w515 & w6608) | (w515 & w6609) | (w6608 & w6609);
assign w542 = (w541 & w534) | (w541 & w7433) | (w534 & w7433);
assign w543 = ~w539 & ~w542;
assign w544 = ~w419 & ~w466;
assign w545 = ~w467 & ~w544;
assign w546 = w543 & w545;
assign w547 = (w545 & w7434) | (w545 & w7435) | (w7434 & w7435);
assign w548 = (w6361 & ~w545) | (w6361 & w7436) | (~w545 & w7436);
assign w549 = ~w547 & ~w548;
assign w550 = w510 & w549;
assign w551 = ~w510 & ~w549;
assign w552 = ~w550 & ~w551;
assign w553 = ~w142 & ~w517;
assign w554 = w342 & w553;
assign w555 = ~w220 & w553;
assign w556 = ~w524 & w6362;
assign w557 = ~w515 & ~w556;
assign w558 = ~w253 & w553;
assign w559 = (~w220 & ~w256) | (~w220 & w6084) | (~w256 & w6084);
assign w560 = ~w303 & ~w364;
assign w561 = ~w559 & w560;
assign w562 = w428 & ~w516;
assign w563 = ~w428 & w516;
assign w564 = ~w562 & ~w563;
assign w565 = w561 & w564;
assign w566 = w561 & w6363;
assign w567 = w515 & w556;
assign w568 = ~w177 & w553;
assign w569 = w103 & ~w364;
assign w570 = w430 & w569;
assign w571 = ~w568 & ~w570;
assign w572 = ~w561 & ~w564;
assign w573 = ~w565 & ~w572;
assign w574 = w430 & w6610;
assign w575 = ~w558 & ~w574;
assign w576 = (w575 & w573) | (w575 & w6086) | (w573 & w6086);
assign w577 = ~w567 & ~w576;
assign w578 = w577 & w6087;
assign w579 = (~w555 & ~w577) | (~w555 & w6088) | (~w577 & w6088);
assign w580 = ~w578 & ~w579;
assign w581 = w530 & ~w534;
assign w582 = ~w535 & ~w581;
assign w583 = w580 & w582;
assign w584 = w577 & w6516;
assign w585 = ~w301 & w553;
assign w586 = (~w585 & ~w577) | (~w585 & w6517) | (~w577 & w6517);
assign w587 = ~w584 & ~w586;
assign w588 = ~w583 & w587;
assign w589 = w583 & ~w587;
assign w590 = ~w588 & ~w589;
assign w591 = ~w543 & ~w545;
assign w592 = ~w546 & ~w591;
assign w593 = ~w590 & ~w592;
assign w594 = (w585 & w583) | (w585 & w6611) | (w583 & w6611);
assign w595 = (w554 & w593) | (w554 & w6364) | (w593 & w6364);
assign w596 = ~w593 & w6365;
assign w597 = (~w403 & w593) | (~w403 & w6612) | (w593 & w6612);
assign w598 = (w597 & w552) | (w597 & w6366) | (w552 & w6366);
assign w599 = ~w595 & ~w596;
assign w600 = w552 & w599;
assign w601 = ~w403 & w553;
assign w602 = ~w601 & ~w595;
assign w603 = (w602 & ~w552) | (w602 & w6367) | (~w552 & w6367);
assign w604 = ~w598 & ~w603;
assign w605 = ~w180 & w342;
assign w606 = w605 & w7474;
assign w607 = w510 & w606;
assign w608 = ~w546 & w6613;
assign w609 = (~w608 & ~w510) | (~w608 & w6368) | (~w510 & w6368);
assign w610 = (~w605 & w546) | (~w605 & w6614) | (w546 & w6614);
assign w611 = (w610 & ~w510) | (w610 & w6369) | (~w510 & w6369);
assign w612 = w609 & ~w611;
assign w613 = ~w259 & ~w301;
assign w614 = ~w469 & ~w613;
assign w615 = (w614 & ~w507) | (w614 & w6370) | (~w507 & w6370);
assign w616 = ~w301 & ~w470;
assign w617 = (w616 & w507) | (w616 & w6371) | (w507 & w6371);
assign w618 = ~w615 & ~w617;
assign w619 = ~w493 & ~w501;
assign w620 = w489 & ~w619;
assign w621 = ~w141 & w403;
assign w622 = w403 & ~w520;
assign w623 = (~w621 & w520) | (~w621 & w6615) | (w520 & w6615);
assign w624 = ~w498 & w621;
assign w625 = ~w623 & ~w624;
assign w626 = w405 & w6089;
assign w627 = w103 & ~w621;
assign w628 = ~w626 & w627;
assign w629 = ~w625 & ~w628;
assign w630 = ~w496 & w6616;
assign w631 = (~w342 & ~w303) | (~w342 & w948) | (~w303 & w948);
assign w632 = w303 & w6090;
assign w633 = ~w631 & ~w632;
assign w634 = (~w177 & w496) | (~w177 & w6617) | (w496 & w6617);
assign w635 = (~w630 & w633) | (~w630 & w6372) | (w633 & w6372);
assign w636 = w629 & ~w635;
assign w637 = ~w629 & w635;
assign w638 = ~w636 & ~w637;
assign w639 = w295 & w6618;
assign w640 = ~w253 & w639;
assign w641 = ~w638 & ~w640;
assign w642 = w638 & w640;
assign w643 = ~w641 & ~w642;
assign w644 = ~w620 & w643;
assign w645 = w620 & ~w643;
assign w646 = ~w644 & ~w645;
assign w647 = ~w479 & ~w504;
assign w648 = w256 & w6619;
assign w649 = (~w648 & ~w459) | (~w648 & w6620) | (~w459 & w6620);
assign w650 = ~w475 & w649;
assign w651 = ~w647 & w650;
assign w652 = w646 & ~w651;
assign w653 = ~w646 & w651;
assign w654 = ~w652 & ~w653;
assign w655 = w618 & w654;
assign w656 = ~w618 & ~w654;
assign w657 = ~w655 & ~w656;
assign w658 = w612 & ~w657;
assign w659 = ~w612 & w657;
assign w660 = ~w658 & ~w659;
assign w661 = w604 & w660;
assign w662 = ~w604 & ~w660;
assign w663 = ~w661 & ~w662;
assign w664 = (~w364 & ~w176) | (~w364 & w6621) | (~w176 & w6621);
assign w665 = w253 & ~w664;
assign w666 = w141 & ~w177;
assign w667 = ~w516 & ~w666;
assign w668 = (~w364 & w237) | (~w364 & w6622) | (w237 & w6622);
assign w669 = ~w667 & w668;
assign w670 = w553 & w6623;
assign w671 = w571 & ~w670;
assign w672 = ~w573 & w671;
assign w673 = (~w669 & ~w573) | (~w669 & w6091) | (~w573 & w6091);
assign w674 = ~w672 & w673;
assign w675 = ~w674 & w6624;
assign w676 = (w220 & w674) | (w220 & w6625) | (w674 & w6625);
assign w677 = ~w557 & ~w567;
assign w678 = ~w566 & ~w576;
assign w679 = ~w677 & ~w678;
assign w680 = w677 & w678;
assign w681 = ~w679 & ~w680;
assign w682 = (w301 & w674) | (w301 & w6626) | (w674 & w6626);
assign w683 = (w682 & ~w681) | (w682 & w6627) | (~w681 & w6627);
assign w684 = ~w580 & ~w582;
assign w685 = ~w103 & ~w583;
assign w686 = ~w683 & ~w684;
assign w687 = w685 & w686;
assign w688 = ~w103 & ~w301;
assign w689 = ~w687 & w6092;
assign w690 = w590 & w592;
assign w691 = ~w593 & ~w690;
assign w692 = (w342 & w687) | (w342 & w6093) | (w687 & w6093);
assign w693 = ~w103 & ~w403;
assign w694 = (~w687 & w6373) | (~w687 & w6374) | (w6373 & w6374);
assign w695 = (w694 & ~w691) | (w694 & w6629) | (~w691 & w6629);
assign w696 = ~w495 & ~w695;
assign w697 = ~w552 & ~w599;
assign w698 = ~w600 & ~w697;
assign w699 = ~w103 & w342;
assign w700 = ~w687 & w6094;
assign w701 = (~w693 & w687) | (~w693 & w6375) | (w687 & w6375);
assign w702 = (w701 & w691) | (w701 & w6630) | (w691 & w6630);
assign w703 = ~w695 & ~w702;
assign w704 = ~w692 & ~w700;
assign w705 = w691 & ~w704;
assign w706 = ~w691 & w704;
assign w707 = ~w705 & ~w706;
assign w708 = w703 & w707;
assign w709 = ~w698 & w708;
assign w710 = ~w696 & w709;
assign w711 = w663 & ~w710;
assign w712 = w698 & ~w703;
assign w713 = (~w696 & ~w698) | (~w696 & w6095) | (~w698 & w6095);
assign w714 = ~w703 & w707;
assign w715 = w698 & w714;
assign w716 = ~w709 & ~w715;
assign w717 = ~w713 & ~w716;
assign w718 = ~w663 & ~w717;
assign w719 = ~w711 & ~w718;
assign w720 = ~w713 & w716;
assign w721 = w663 & w720;
assign w722 = ~w709 & w713;
assign w723 = ~w663 & w722;
assign w724 = ~w721 & ~w723;
assign w725 = ~w719 & w724;
assign w726 = ~w180 & w725;
assign w727 = ~w698 & w703;
assign w728 = ~w712 & ~w727;
assign w729 = ~w707 & ~w728;
assign w730 = (~w180 & w707) | (~w180 & w6631) | (w707 & w6631);
assign w731 = w729 & w730;
assign w732 = ~w707 & w728;
assign w733 = w728 & w6632;
assign w734 = ~w303 & ~w559;
assign w735 = w259 & w734;
assign w736 = ~w260 & ~w735;
assign w737 = ~w707 & ~w736;
assign w738 = ~w707 & w734;
assign w739 = (w259 & w707) | (w259 & w6633) | (w707 & w6633);
assign w740 = (~w737 & ~w728) | (~w737 & w6634) | (~w728 & w6634);
assign w741 = ~w733 & ~w740;
assign w742 = ~w731 & ~w741;
assign w743 = w725 & w6635;
assign w744 = w729 & w6636;
assign w745 = (~w744 & ~w726) | (~w744 & w6096) | (~w726 & w6096);
assign w746 = ~w180 & ~w403;
assign w747 = ~w607 & w6097;
assign w748 = (~w403 & w607) | (~w403 & w6098) | (w607 & w6098);
assign w749 = ~w747 & ~w748;
assign w750 = w658 & ~w749;
assign w751 = ~w658 & w749;
assign w752 = ~w750 & ~w751;
assign w753 = ~w259 & w342;
assign w754 = ~w301 & w734;
assign w755 = ~w646 & w754;
assign w756 = ~w651 & w755;
assign w757 = w646 & ~w754;
assign w758 = ~w475 & w6099;
assign w759 = ~w647 & w758;
assign w760 = ~w757 & ~w759;
assign w761 = ~w756 & w760;
assign w762 = (~w641 & w620) | (~w641 & w6376) | (w620 & w6376);
assign w763 = ~w220 & w301;
assign w764 = ~w496 & w6637;
assign w765 = ~w636 & ~w764;
assign w766 = ~w253 & ~w342;
assign w767 = ~w177 & ~w403;
assign w768 = ~w622 & ~w767;
assign w769 = w667 & ~w768;
assign w770 = ~w667 & w768;
assign w771 = ~w769 & ~w770;
assign w772 = w766 & ~w771;
assign w773 = ~w766 & w771;
assign w774 = ~w772 & ~w773;
assign w775 = w765 & ~w774;
assign w776 = ~w765 & w774;
assign w777 = ~w775 & ~w776;
assign w778 = ~w763 & ~w777;
assign w779 = w763 & w777;
assign w780 = ~w778 & ~w779;
assign w781 = w762 & ~w780;
assign w782 = ~w762 & w780;
assign w783 = ~w781 & ~w782;
assign w784 = w761 & ~w783;
assign w785 = ~w761 & w783;
assign w786 = ~w784 & ~w785;
assign w787 = ~w753 & ~w786;
assign w788 = w753 & w786;
assign w789 = ~w787 & ~w788;
assign w790 = (~w615 & ~w618) | (~w615 & w6100) | (~w618 & w6100);
assign w791 = w789 & w790;
assign w792 = ~w789 & ~w790;
assign w793 = ~w791 & ~w792;
assign w794 = ~w752 & w793;
assign w795 = w752 & ~w793;
assign w796 = ~w794 & ~w795;
assign w797 = ~w598 & ~w661;
assign w798 = ~w661 & w6101;
assign w799 = w796 & w798;
assign w800 = ~w796 & ~w798;
assign w801 = ~w799 & ~w800;
assign w802 = ~w663 & w713;
assign w803 = (~w103 & w663) | (~w103 & w6102) | (w663 & w6102);
assign w804 = ~w718 & w6377;
assign w805 = (w803 & w718) | (w803 & w6378) | (w718 & w6378);
assign w806 = ~w804 & ~w805;
assign w807 = w801 & w806;
assign w808 = ~w801 & ~w806;
assign w809 = ~w807 & ~w808;
assign w810 = ~w301 & ~w707;
assign w811 = (w734 & w728) | (w734 & w6103) | (w728 & w6103);
assign w812 = ~w306 & ~w734;
assign w813 = ~w707 & w812;
assign w814 = ~w813 & ~w811;
assign w815 = ~w707 & w6638;
assign w816 = ~w728 & w815;
assign w817 = ~w814 & w816;
assign w818 = w728 & w810;
assign w819 = w811 & ~w818;
assign w820 = (~w813 & w728) | (~w813 & w6639) | (w728 & w6639);
assign w821 = ~w819 & w820;
assign w822 = ~w817 & ~w821;
assign w823 = ~w259 & w725;
assign w824 = w822 & w823;
assign w825 = ~w822 & ~w823;
assign w826 = ~w824 & ~w825;
assign w827 = (~w745 & w826) | (~w745 & w6379) | (w826 & w6379);
assign w828 = w809 & w826;
assign w829 = w827 & ~w828;
assign w830 = ~w180 & w809;
assign w831 = w745 & w826;
assign w832 = w830 & w831;
assign w833 = w745 & ~w826;
assign w834 = ~w830 & w833;
assign w835 = ~w832 & ~w834;
assign w836 = ~w829 & w835;
assign w837 = ~w731 & w741;
assign w838 = (~w837 & ~w725) | (~w837 & w6640) | (~w725 & w6640);
assign w839 = ~w743 & ~w838;
assign w840 = w663 & ~w713;
assign w841 = ~w802 & ~w840;
assign w842 = w725 & ~w737;
assign w843 = (w731 & w841) | (w731 & w6641) | (w841 & w6641);
assign w844 = ~w842 & w843;
assign w845 = ~w839 & ~w844;
assign w846 = w553 & w809;
assign w847 = ~w845 & w846;
assign w848 = ~w728 & w6104;
assign w849 = w728 & ~w730;
assign w850 = ~w848 & ~w849;
assign w851 = ~w707 & w6642;
assign w852 = ~w850 & ~w851;
assign w853 = w841 & w852;
assign w854 = ~w841 & ~w852;
assign w855 = ~w853 & ~w854;
assign w856 = ~w553 & w716;
assign w857 = w178 & ~w517;
assign w858 = ~w728 & w6643;
assign w859 = ~w553 & ~w716;
assign w860 = ~w841 & w859;
assign w861 = (~w858 & ~w841) | (~w858 & w6105) | (~w841 & w6105);
assign w862 = ~w860 & w861;
assign w863 = ~w855 & w862;
assign w864 = (w553 & ~w855) | (w553 & w6644) | (~w855 & w6644);
assign w865 = ~w863 & w864;
assign w866 = (~w865 & ~w846) | (~w865 & w6645) | (~w846 & w6645);
assign w867 = w845 & ~w846;
assign w868 = ~w180 & w403;
assign w869 = (~w868 & w658) | (~w868 & w6646) | (w658 & w6646);
assign w870 = ~w794 & ~w869;
assign w871 = ~w259 & ~w403;
assign w872 = (~w871 & ~w786) | (~w871 & w6647) | (~w786 & w6647);
assign w873 = (w872 & ~w789) | (w872 & w6648) | (~w789 & w6648);
assign w874 = ~w788 & ~w790;
assign w875 = (~w403 & w786) | (~w403 & w6380) | (w786 & w6380);
assign w876 = ~w874 & w875;
assign w877 = w342 & w734;
assign w878 = (~w756 & ~w761) | (~w756 & w6106) | (~w761 & w6106);
assign w879 = w877 & ~w878;
assign w880 = ~w877 & w878;
assign w881 = ~w879 & ~w880;
assign w882 = ~w220 & ~w342;
assign w883 = (w882 & w776) | (w882 & w6649) | (w776 & w6649);
assign w884 = ~w776 & w6650;
assign w885 = ~w883 & ~w884;
assign w886 = ~w408 & ~w410;
assign w887 = ~w408 & w6381;
assign w888 = w177 & ~w887;
assign w889 = ~w177 & w887;
assign w890 = ~w888 & ~w889;
assign w891 = ~w623 & ~w857;
assign w892 = w890 & w891;
assign w893 = ~w890 & ~w891;
assign w894 = ~w892 & ~w893;
assign w895 = w885 & w894;
assign w896 = ~w885 & ~w894;
assign w897 = ~w895 & ~w896;
assign w898 = (~w305 & w782) | (~w305 & w6651) | (w782 & w6651);
assign w899 = w897 & ~w898;
assign w900 = ~w897 & w898;
assign w901 = ~w899 & ~w900;
assign w902 = w881 & ~w901;
assign w903 = ~w881 & w901;
assign w904 = ~w902 & ~w903;
assign w905 = ~w873 & w6107;
assign w906 = (w904 & w873) | (w904 & w6108) | (w873 & w6108);
assign w907 = ~w905 & ~w906;
assign w908 = w870 & ~w907;
assign w909 = ~w870 & w907;
assign w910 = ~w908 & ~w909;
assign w911 = (w797 & ~w796) | (w797 & w6109) | (~w796 & w6109);
assign w912 = ~w910 & ~w911;
assign w913 = w910 & w911;
assign w914 = ~w912 & ~w913;
assign w915 = ~w801 & w804;
assign w916 = w801 & w805;
assign w917 = ~w915 & ~w916;
assign w918 = w914 & w917;
assign w919 = ~w914 & ~w917;
assign w920 = ~w918 & ~w919;
assign w921 = w553 & w920;
assign w922 = ~w867 & w921;
assign w923 = ~w866 & w922;
assign w924 = (w865 & w846) | (w865 & w6652) | (w846 & w6652);
assign w925 = ~w847 & ~w921;
assign w926 = ~w924 & w925;
assign w927 = ~w923 & ~w926;
assign w928 = w836 & ~w927;
assign w929 = ~w836 & w927;
assign w930 = ~w928 & ~w929;
assign w931 = ~w728 & w6653;
assign w932 = w716 & ~w732;
assign w933 = ~w732 & w6654;
assign w934 = ~w180 & ~w707;
assign w935 = ~w933 & ~w934;
assign w936 = (~w931 & ~w725) | (~w931 & w6655) | (~w725 & w6655);
assign w937 = ~w809 & w936;
assign w938 = w809 & ~w936;
assign w939 = w855 & ~w862;
assign w940 = ~w863 & ~w939;
assign w941 = ~w938 & w940;
assign w942 = (~w920 & w941) | (~w920 & w6110) | (w941 & w6110);
assign w943 = ~w103 & ~w942;
assign w944 = (~w180 & ~w870) | (~w180 & w6111) | (~w870 & w6111);
assign w945 = ~w876 & w904;
assign w946 = ~w873 & ~w945;
assign w947 = (~w259 & w945) | (~w259 & w6656) | (w945 & w6656);
assign w948 = ~w301 & ~w342;
assign w949 = ~w220 & w403;
assign w950 = (w253 & ~w890) | (w253 & w6657) | (~w890 & w6657);
assign w951 = (~w889 & ~w890) | (~w889 & w6659) | (~w890 & w6659);
assign w952 = ~w950 & w951;
assign w953 = w949 & ~w952;
assign w954 = ~w949 & w952;
assign w955 = ~w953 & ~w954;
assign w956 = w948 & ~w955;
assign w957 = ~w948 & w955;
assign w958 = ~w956 & ~w957;
assign w959 = (~w883 & ~w885) | (~w883 & w6660) | (~w885 & w6660);
assign w960 = w958 & w959;
assign w961 = ~w958 & ~w959;
assign w962 = ~w960 & ~w961;
assign w963 = ~w306 & w342;
assign w964 = ~w898 & w6661;
assign w965 = (~w963 & w898) | (~w963 & w6662) | (w898 & w6662);
assign w966 = ~w964 & ~w965;
assign w967 = ~w962 & w966;
assign w968 = w962 & ~w966;
assign w969 = ~w967 & ~w968;
assign w970 = (w901 & ~w878) | (w901 & w6663) | (~w878 & w6663);
assign w971 = (~w403 & w970) | (~w403 & w6382) | (w970 & w6382);
assign w972 = ~w403 & w734;
assign w973 = ~w970 & w6383;
assign w974 = ~w971 & ~w973;
assign w975 = w969 & w974;
assign w976 = ~w969 & ~w974;
assign w977 = ~w975 & ~w976;
assign w978 = w947 & ~w977;
assign w979 = ~w947 & w977;
assign w980 = ~w978 & ~w979;
assign w981 = ~w944 & w980;
assign w982 = w944 & ~w980;
assign w983 = ~w981 & ~w982;
assign w984 = w801 & w803;
assign w985 = ~w913 & w984;
assign w986 = ~w985 & w6112;
assign w987 = (~w983 & w985) | (~w983 & w6113) | (w985 & w6113);
assign w988 = ~w986 & ~w987;
assign w989 = ~w914 & w915;
assign w990 = (w719 & w910) | (w719 & w6114) | (w910 & w6114);
assign w991 = w985 & w990;
assign w992 = ~w989 & ~w991;
assign w993 = ~w103 & w992;
assign w994 = ~w983 & w991;
assign w995 = (~w994 & ~w993) | (~w994 & w6115) | (~w993 & w6115);
assign w996 = ~w943 & w995;
assign w997 = ~w847 & ~w867;
assign w998 = w865 & ~w997;
assign w999 = ~w941 & w6116;
assign w1000 = (~w999 & ~w997) | (~w999 & w6384) | (~w997 & w6384);
assign w1001 = w995 & ~w998;
assign w1002 = (~w996 & ~w1001) | (~w996 & w6385) | (~w1001 & w6385);
assign w1003 = ~w998 & w1000;
assign w1004 = w988 & ~w992;
assign w1005 = ~w988 & w992;
assign w1006 = ~w1004 & ~w1005;
assign w1007 = w943 & w1006;
assign w1008 = ~w1003 & w1007;
assign w1009 = w1002 & ~w1008;
assign w1010 = w930 & ~w1009;
assign w1011 = ~w930 & w1009;
assign w1012 = ~w1010 & ~w1011;
assign w1013 = (~w971 & ~w974) | (~w971 & w6664) | (~w974 & w6664);
assign w1014 = ~w306 & ~w403;
assign w1015 = (w1014 & w967) | (w1014 & w6665) | (w967 & w6665);
assign w1016 = ~w967 & w6666;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = (~w957 & ~w958) | (~w957 & w6667) | (~w958 & w6667);
assign w1019 = ~w301 & w403;
assign w1020 = w220 & w951;
assign w1021 = (w890 & w6668) | (w890 & w6669) | (w6668 & w6669);
assign w1022 = ~w1020 & w6670;
assign w1023 = (w1019 & w1020) | (w1019 & w6671) | (w1020 & w6671);
assign w1024 = ~w1022 & ~w1023;
assign w1025 = w1018 & ~w1024;
assign w1026 = ~w632 & w1024;
assign w1027 = ~w1018 & w1026;
assign w1028 = ~w1025 & ~w1027;
assign w1029 = w1017 & ~w1028;
assign w1030 = ~w1017 & w1028;
assign w1031 = ~w1029 & ~w1030;
assign w1032 = w1013 & w6672;
assign w1033 = (w1031 & ~w1013) | (w1031 & w6673) | (~w1013 & w6673);
assign w1034 = ~w1032 & ~w1033;
assign w1035 = ~w259 & w977;
assign w1036 = ~w946 & ~w1035;
assign w1037 = w1034 & ~w1036;
assign w1038 = ~w1034 & w1036;
assign w1039 = ~w1037 & ~w1038;
assign w1040 = ~w912 & ~w982;
assign w1041 = ~w985 & w1040;
assign w1042 = (w1039 & w1041) | (w1039 & w6117) | (w1041 & w6117);
assign w1043 = ~w1041 & w6118;
assign w1044 = ~w1042 & ~w1043;
assign w1045 = w1004 & w1044;
assign w1046 = ~w403 & ~w633;
assign w1047 = (~w1046 & ~w1018) | (~w1046 & w6674) | (~w1018 & w6674);
assign w1048 = w1018 & w6675;
assign w1049 = ~w1047 & ~w1048;
assign w1050 = w342 & w403;
assign w1051 = w301 & ~w1021;
assign w1052 = (w1019 & ~w951) | (w1019 & w6678) | (~w951 & w6678);
assign w1053 = (w1050 & w1052) | (w1050 & w6679) | (w1052 & w6679);
assign w1054 = ~w1052 & w6680;
assign w1055 = ~w1053 & ~w1054;
assign w1056 = ~w1049 & w1055;
assign w1057 = w1049 & ~w1055;
assign w1058 = ~w1056 & ~w1057;
assign w1059 = (~w1016 & ~w1017) | (~w1016 & w6681) | (~w1017 & w6681);
assign w1060 = ~w1059 & w6682;
assign w1061 = (~w1058 & w1059) | (~w1058 & w6683) | (w1059 & w6683);
assign w1062 = ~w1060 & ~w1061;
assign w1063 = ~w1032 & w6684;
assign w1064 = (w1062 & w1032) | (w1062 & w6685) | (w1032 & w6685);
assign w1065 = ~w1063 & ~w1064;
assign w1066 = ~w1038 & ~w1042;
assign w1067 = w1065 & w1066;
assign w1068 = ~w1065 & ~w1066;
assign w1069 = ~w1067 & ~w1068;
assign w1070 = w1045 & ~w1069;
assign w1071 = (w890 & w6686) | (w890 & w6687) | (w6686 & w6687);
assign w1072 = ~w410 & ~w631;
assign w1073 = (w951 & w6688) | (w951 & w6689) | (w6688 & w6689);
assign w1074 = ~w1071 & ~w1073;
assign w1075 = (~w1074 & ~w1018) | (~w1074 & w6690) | (~w1018 & w6690);
assign w1076 = (w1075 & ~w1049) | (w1075 & w6691) | (~w1049 & w6691);
assign w1077 = ~w633 & ~w1076;
assign w1078 = (w633 & w1073) | (w633 & w6692) | (w1073 & w6692);
assign w1079 = ~w1059 & w6693;
assign w1080 = ~w1060 & w1079;
assign w1081 = ~w1064 & w1080;
assign w1082 = (~w1081 & ~w1066) | (~w1081 & w6694) | (~w1066 & w6694);
assign w1083 = ~w1063 & w1080;
assign w1084 = w1066 & w1083;
assign w1085 = ~w1082 & ~w1084;
assign w1086 = w1045 & w6695;
assign w1087 = (w1085 & ~w1045) | (w1085 & w6696) | (~w1045 & w6696);
assign w1088 = ~w1086 & ~w1087;
assign w1089 = ~w1045 & w1069;
assign w1090 = ~w1070 & ~w1089;
assign w1091 = ~w1004 & ~w1044;
assign w1092 = ~w1045 & ~w1091;
assign w1093 = w886 & w1006;
assign w1094 = (w886 & w841) | (w886 & w1211) | (w841 & w1211);
assign w1095 = (w841 & w6697) | (w841 & w6698) | (w6697 & w6698);
assign w1096 = ~w801 & ~w803;
assign w1097 = ~w984 & ~w1096;
assign w1098 = (~w732 & w841) | (~w732 & w6699) | (w841 & w6699);
assign w1099 = ~w719 & w1097;
assign w1100 = (w886 & w1097) | (w886 & w6119) | (w1097 & w6119);
assign w1101 = ~w1099 & w1100;
assign w1102 = ~w1095 & ~w1101;
assign w1103 = ~w410 & w725;
assign w1104 = (~w1103 & w1097) | (~w1103 & w6700) | (w1097 & w6700);
assign w1105 = w809 & ~w1104;
assign w1106 = ~w1102 & w1105;
assign w1107 = (~w920 & w1102) | (~w920 & w6701) | (w1102 & w6701);
assign w1108 = w1006 & w6702;
assign w1109 = ~w1092 & ~w1108;
assign w1110 = w1088 & ~w1109;
assign w1111 = (w1090 & w1110) | (w1090 & w6703) | (w1110 & w6703);
assign w1112 = ~w633 & w1092;
assign w1113 = w886 & w920;
assign w1114 = w1095 & ~w1104;
assign w1115 = ~w809 & ~w1114;
assign w1116 = w1113 & ~w1115;
assign w1117 = ~w1107 & ~w1116;
assign w1118 = w1093 & ~w1117;
assign w1119 = ~w1093 & w1117;
assign w1120 = ~w1118 & ~w1119;
assign w1121 = ~w1112 & w1120;
assign w1122 = w1112 & ~w1120;
assign w1123 = ~w1121 & ~w1122;
assign w1124 = ~w633 & w1006;
assign w1125 = ~w633 & w920;
assign w1126 = ~w707 & w841;
assign w1127 = w1094 & ~w1126;
assign w1128 = (~w886 & w732) | (~w886 & w6704) | (w732 & w6704);
assign w1129 = ~w1127 & ~w1128;
assign w1130 = w633 & w886;
assign w1131 = ~w707 & ~w1130;
assign w1132 = (~w1131 & ~w728) | (~w1131 & w6120) | (~w728 & w6120);
assign w1133 = (w728 & w6705) | (w728 & w6706) | (w6705 & w6706);
assign w1134 = w841 & w1133;
assign w1135 = (~w633 & w1134) | (~w633 & w6121) | (w1134 & w6121);
assign w1136 = w1097 & w1135;
assign w1137 = ~w1134 & w6122;
assign w1138 = ~w1097 & w1137;
assign w1139 = ~w1136 & ~w1138;
assign w1140 = ~w1129 & ~w1139;
assign w1141 = ~w1134 & w1139;
assign w1142 = ~w1140 & ~w1141;
assign w1143 = w1125 & w1142;
assign w1144 = ~w1125 & ~w1142;
assign w1145 = ~w1143 & ~w1144;
assign w1146 = w1095 & w1097;
assign w1147 = (w1103 & w1101) | (w1103 & w6707) | (w1101 & w6707);
assign w1148 = ~w1101 & w6708;
assign w1149 = ~w1147 & ~w1148;
assign w1150 = w1145 & w1149;
assign w1151 = (~w1143 & ~w1145) | (~w1143 & w6123) | (~w1145 & w6123);
assign w1152 = ~w1124 & w1151;
assign w1153 = w1124 & ~w1151;
assign w1154 = ~w1106 & w6709;
assign w1155 = (w1113 & w1106) | (w1113 & w6710) | (w1106 & w6710);
assign w1156 = ~w1154 & ~w1155;
assign w1157 = (w1156 & w1151) | (w1156 & w6711) | (w1151 & w6711);
assign w1158 = ~w1152 & ~w1157;
assign w1159 = w1123 & ~w1158;
assign w1160 = (~w1121 & ~w1123) | (~w1121 & w6712) | (~w1123 & w6712);
assign w1161 = w1090 & w1160;
assign w1162 = ~w633 & w1090;
assign w1163 = ~w1160 & ~w1162;
assign w1164 = ~w1161 & ~w1163;
assign w1165 = w886 & w1092;
assign w1166 = ~w1006 & ~w1116;
assign w1167 = ~w1108 & ~w1166;
assign w1168 = w1165 & ~w1167;
assign w1169 = ~w1165 & w1167;
assign w1170 = ~w1168 & ~w1169;
assign w1171 = w1164 & ~w1170;
assign w1172 = (~w1161 & ~w1164) | (~w1161 & w6713) | (~w1164 & w6713);
assign w1173 = w886 & w1090;
assign w1174 = w1165 & ~w1166;
assign w1175 = ~w1109 & ~w1174;
assign w1176 = ~w1173 & w1175;
assign w1177 = w1173 & ~w1175;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = (w1172 & w6715) | (w1172 & w6716) | (w6715 & w6716);
assign w1180 = w1110 & w1174;
assign w1181 = w886 & ~w1090;
assign w1182 = ~w1180 & w1181;
assign w1183 = ~w1111 & ~w1182;
assign w1184 = w1183 & ~w1179;
assign w1185 = (w1172 & w6719) | (w1172 & w6720) | (w6719 & w6720);
assign w1186 = w1088 & ~w1185;
assign w1187 = ~w1185 & w1188;
assign w1188 = ~w306 & w1088;
assign w1189 = (w1188 & w1180) | (w1188 & w6722) | (w1180 & w6722);
assign w1190 = w633 & ~w1086;
assign w1191 = ~w1189 & w1190;
assign w1192 = (~w1191 & w1185) | (~w1191 & w6723) | (w1185 & w6723);
assign w1193 = w306 & ~w1186;
assign w1194 = ~w1187 & ~w1193;
assign w1195 = ~w1164 & w1170;
assign w1196 = ~w1171 & ~w1195;
assign w1197 = ~w1088 & ~w1172;
assign w1198 = ~w1123 & w1158;
assign w1199 = ~w1159 & ~w1198;
assign w1200 = ~w306 & w1090;
assign w1201 = ~w1199 & w1200;
assign w1202 = ~w306 & w1092;
assign w1203 = ~w306 & w1006;
assign w1204 = w1129 & w1139;
assign w1205 = ~w1140 & ~w1204;
assign w1206 = ~w306 & w920;
assign w1207 = w1205 & ~w1206;
assign w1208 = ~w1205 & w1206;
assign w1209 = ~w306 & w6724;
assign w1210 = ~w728 & w6725;
assign w1211 = ~w707 & w886;
assign w1212 = ~w732 & w6124;
assign w1213 = ~w1211 & ~w1212;
assign w1214 = w306 & ~w633;
assign w1215 = w403 & w1214;
assign w1216 = ~w728 & w6726;
assign w1217 = ~w1210 & ~w1216;
assign w1218 = ~w1213 & w1217;
assign w1219 = ~w306 & w725;
assign w1220 = w1218 & w1219;
assign w1221 = (~w1210 & ~w1219) | (~w1210 & w6727) | (~w1219 & w6727);
assign w1222 = (w1132 & ~w725) | (w1132 & w6386) | (~w725 & w6386);
assign w1223 = ~w1134 & ~w1222;
assign w1224 = ~w809 & ~w1223;
assign w1225 = (~w1221 & w809) | (~w1221 & w6728) | (w809 & w6728);
assign w1226 = w809 & w1223;
assign w1227 = w809 & w6729;
assign w1228 = ~w1225 & ~w1227;
assign w1229 = (w1228 & w1205) | (w1228 & w6730) | (w1205 & w6730);
assign w1230 = w1203 & w6731;
assign w1231 = (~w1203 & w1229) | (~w1203 & w6125) | (w1229 & w6125);
assign w1232 = ~w1145 & ~w1149;
assign w1233 = ~w1150 & ~w1232;
assign w1234 = w1202 & w7475;
assign w1235 = ~w1230 & w7476;
assign w1236 = ~w1234 & ~w1235;
assign w1237 = ~w1152 & ~w1153;
assign w1238 = w1156 & w1237;
assign w1239 = ~w1156 & ~w1237;
assign w1240 = ~w1238 & ~w1239;
assign w1241 = w1236 & ~w1240;
assign w1242 = ~w1234 & ~w1241;
assign w1243 = w1199 & ~w1200;
assign w1244 = ~w1201 & ~w1243;
assign w1245 = ~w1242 & w1244;
assign w1246 = (w1188 & w1199) | (w1188 & w6732) | (w1199 & w6732);
assign w1247 = (w1246 & ~w1244) | (w1246 & w6733) | (~w1244 & w6733);
assign w1248 = ~w1197 & ~w1247;
assign w1249 = ~w1196 & ~w1248;
assign w1250 = w1196 & w1248;
assign w1251 = ~w1249 & ~w1250;
assign w1252 = w1242 & ~w1244;
assign w1253 = ~w1245 & ~w1252;
assign w1254 = ~w1236 & w1240;
assign w1255 = ~w1241 & ~w1254;
assign w1256 = w734 & w1090;
assign w1257 = w734 & w1092;
assign w1258 = w734 & w1006;
assign w1259 = w734 & w920;
assign w1260 = ~w963 & ~w1214;
assign w1261 = ~w728 & w6127;
assign w1262 = w306 & w707;
assign w1263 = w633 & ~w707;
assign w1264 = ~w1262 & ~w1263;
assign w1265 = w728 & w1264;
assign w1266 = ~w1261 & ~w1265;
assign w1267 = ~w728 & w6734;
assign w1268 = ~w1266 & w1267;
assign w1269 = w1266 & ~w1267;
assign w1270 = ~w1268 & ~w1269;
assign w1271 = w716 & w734;
assign w1272 = w841 & w1271;
assign w1273 = ~w716 & w734;
assign w1274 = ~w841 & w1273;
assign w1275 = ~w1272 & ~w1274;
assign w1276 = w1270 & ~w1275;
assign w1277 = (~w1268 & w1275) | (~w1268 & w6128) | (w1275 & w6128);
assign w1278 = ~w1218 & ~w1219;
assign w1279 = ~w1220 & ~w1278;
assign w1280 = w1277 & ~w1279;
assign w1281 = ~w1277 & w1279;
assign w1282 = w734 & w809;
assign w1283 = ~w1281 & ~w1282;
assign w1284 = (~w1259 & w1283) | (~w1259 & w6388) | (w1283 & w6388);
assign w1285 = ~w1283 & w6389;
assign w1286 = ~w1284 & ~w1285;
assign w1287 = (w1221 & ~w809) | (w1221 & w6735) | (~w809 & w6735);
assign w1288 = ~w1224 & ~w1226;
assign w1289 = ~w1287 & w1288;
assign w1290 = w1287 & ~w1288;
assign w1291 = ~w1289 & ~w1290;
assign w1292 = w1286 & ~w1291;
assign w1293 = (~w1284 & ~w1286) | (~w1284 & w6129) | (~w1286 & w6129);
assign w1294 = ~w1258 & ~w1293;
assign w1295 = w1258 & w1293;
assign w1296 = ~w1207 & ~w1208;
assign w1297 = ~w1228 & ~w1296;
assign w1298 = w1228 & w1296;
assign w1299 = ~w1297 & ~w1298;
assign w1300 = ~w1295 & w1299;
assign w1301 = (~w1257 & w1300) | (~w1257 & w6736) | (w1300 & w6736);
assign w1302 = w1257 & ~w1294;
assign w1303 = ~w1300 & w1302;
assign w1304 = ~w1230 & ~w1231;
assign w1305 = w1233 & w1304;
assign w1306 = ~w1233 & ~w1304;
assign w1307 = ~w1305 & ~w1306;
assign w1308 = ~w1303 & ~w1307;
assign w1309 = ~w1308 & w6390;
assign w1310 = ~w1255 & ~w1309;
assign w1311 = (~w1256 & w1308) | (~w1256 & w6391) | (w1308 & w6391);
assign w1312 = w1088 & ~w1311;
assign w1313 = (w734 & w1310) | (w734 & w6737) | (w1310 & w6737);
assign w1314 = ~w1253 & w1313;
assign w1315 = w1251 & w1314;
assign w1316 = ~w1178 & w7477;
assign w1317 = ~w1179 & ~w1316;
assign w1318 = w1251 & w6738;
assign w1319 = w734 & ~w1318;
assign w1320 = (w1172 & w6739) | (w1172 & w6740) | (w6739 & w6740);
assign w1321 = ~w1184 & ~w1320;
assign w1322 = (w1321 & ~w1249) | (w1321 & w6741) | (~w1249 & w6741);
assign w1323 = w1319 & w1322;
assign w1324 = (~w1322 & w1318) | (~w1322 & w6742) | (w1318 & w6742);
assign w1325 = ~w1323 & ~w1324;
assign w1326 = ~w259 & w1092;
assign w1327 = ~w259 & w1006;
assign w1328 = ~w259 & w920;
assign w1329 = ~w1270 & w1275;
assign w1330 = ~w1276 & ~w1329;
assign w1331 = (~w817 & ~w823) | (~w817 & w6130) | (~w823 & w6130);
assign w1332 = w809 & ~w1331;
assign w1333 = ~w1330 & ~w1332;
assign w1334 = ~w259 & w809;
assign w1335 = (w1331 & ~w809) | (w1331 & w6131) | (~w809 & w6131);
assign w1336 = ~w1333 & ~w1335;
assign w1337 = w1328 & w1336;
assign w1338 = ~w1328 & ~w1336;
assign w1339 = ~w1280 & ~w1281;
assign w1340 = w1282 & ~w1339;
assign w1341 = ~w1282 & w1339;
assign w1342 = ~w1340 & ~w1341;
assign w1343 = ~w1338 & ~w1342;
assign w1344 = ~w1343 & w6132;
assign w1345 = (w1327 & w1343) | (w1327 & w6133) | (w1343 & w6133);
assign w1346 = ~w1286 & w1291;
assign w1347 = ~w1292 & ~w1346;
assign w1348 = (w6134 & w6392) | (w6134 & w6393) | (w6392 & w6393);
assign w1349 = (~w6134 & w6394) | (~w6134 & w6395) | (w6394 & w6395);
assign w1350 = ~w1348 & ~w1349;
assign w1351 = ~w1294 & ~w1295;
assign w1352 = w1299 & w1351;
assign w1353 = ~w1299 & ~w1351;
assign w1354 = ~w1352 & ~w1353;
assign w1355 = w1350 & ~w1354;
assign w1356 = ~w1085 & w1090;
assign w1357 = ~w1301 & ~w1303;
assign w1358 = ~w1307 & w1357;
assign w1359 = w1307 & ~w1357;
assign w1360 = ~w1358 & ~w1359;
assign w1361 = ~w1090 & w1348;
assign w1362 = ~w259 & w1090;
assign w1363 = ~w1348 & w1362;
assign w1364 = ~w1361 & ~w1363;
assign w1365 = w1355 & ~w1364;
assign w1366 = ~w1355 & w1364;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = ~w1360 & w1367;
assign w1369 = ~w259 & w7478;
assign w1370 = (w1369 & ~w1367) | (w1369 & w7437) | (~w1367 & w7437);
assign w1371 = ~w1309 & ~w1311;
assign w1372 = w1255 & ~w1371;
assign w1373 = ~w1255 & w1371;
assign w1374 = ~w1372 & ~w1373;
assign w1375 = w1370 & w1374;
assign w1376 = w1253 & ~w1313;
assign w1377 = ~w1314 & ~w1376;
assign w1378 = w1375 & w1377;
assign w1379 = (~w259 & ~w1378) | (~w259 & w6744) | (~w1378 & w6744);
assign w1380 = ~w1315 & w6745;
assign w1381 = (w1317 & w1315) | (w1317 & w6746) | (w1315 & w6746);
assign w1382 = ~w1380 & ~w1381;
assign w1383 = w1379 & ~w1382;
assign w1384 = ~w1370 & ~w1374;
assign w1385 = ~w1375 & ~w1384;
assign w1386 = ~w180 & w1090;
assign w1387 = ~w1344 & ~w1345;
assign w1388 = w1347 & w1387;
assign w1389 = ~w1347 & ~w1387;
assign w1390 = ~w1388 & ~w1389;
assign w1391 = ~w180 & w920;
assign w1392 = ~w832 & w6396;
assign w1393 = w1330 & w1331;
assign w1394 = ~w1330 & ~w1331;
assign w1395 = ~w1393 & ~w1394;
assign w1396 = w1334 & w1395;
assign w1397 = ~w1334 & ~w1395;
assign w1398 = ~w1396 & ~w1397;
assign w1399 = ~w1392 & ~w1398;
assign w1400 = ~w180 & w992;
assign w1401 = w988 & w1400;
assign w1402 = ~w180 & ~w992;
assign w1403 = ~w988 & w1402;
assign w1404 = ~w1401 & ~w1403;
assign w1405 = (w1391 & w832) | (w1391 & w6397) | (w832 & w6397);
assign w1406 = w1404 & ~w1405;
assign w1407 = ~w1399 & w1406;
assign w1408 = w1398 & ~w1405;
assign w1409 = ~w1392 & ~w1404;
assign w1410 = ~w1408 & w1409;
assign w1411 = ~w1407 & ~w1410;
assign w1412 = ~w1337 & ~w1338;
assign w1413 = ~w1342 & w1412;
assign w1414 = w1342 & ~w1412;
assign w1415 = ~w1413 & ~w1414;
assign w1416 = w1411 & ~w1415;
assign w1417 = ~w180 & w1092;
assign w1418 = ~w1407 & w1417;
assign w1419 = w1407 & ~w1417;
assign w1420 = ~w1418 & ~w1419;
assign w1421 = ~w1416 & w1420;
assign w1422 = w1416 & w1417;
assign w1423 = ~w1421 & ~w1422;
assign w1424 = ~w1390 & ~w1423;
assign w1425 = ~w1416 & w1418;
assign w1426 = (w6135 & w6398) | (w6135 & w6399) | (w6398 & w6399);
assign w1427 = ~w1350 & w1354;
assign w1428 = ~w1355 & ~w1427;
assign w1429 = (~w6135 & w6400) | (~w6135 & w6401) | (w6400 & w6401);
assign w1430 = ~w1426 & ~w1429;
assign w1431 = ~w1428 & w1430;
assign w1432 = (~w1426 & ~w1430) | (~w1426 & w6747) | (~w1430 & w6747);
assign w1433 = w1360 & ~w1367;
assign w1434 = ~w1368 & ~w1433;
assign w1435 = (w1088 & w1434) | (w1088 & w6748) | (w1434 & w6748);
assign w1436 = ~w1375 & ~w1377;
assign w1437 = ~w1378 & ~w1436;
assign w1438 = w1432 & w1434;
assign w1439 = w1385 & w6749;
assign w1440 = (~w180 & ~w1437) | (~w180 & w6750) | (~w1437 & w6750);
assign w1441 = (w1251 & w1378) | (w1251 & w1315) | (w1378 & w1315);
assign w1442 = ~w1378 & w6751;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = w1440 & ~w1443;
assign w1445 = ~w1440 & w1443;
assign w1446 = ~w1444 & ~w1445;
assign w1447 = w1428 & ~w1430;
assign w1448 = ~w1431 & ~w1447;
assign w1449 = w553 & w1090;
assign w1450 = ~w836 & ~w923;
assign w1451 = w553 & w992;
assign w1452 = w988 & w1451;
assign w1453 = w553 & ~w992;
assign w1454 = ~w988 & w1453;
assign w1455 = ~w1452 & ~w1454;
assign w1456 = ~w926 & ~w1455;
assign w1457 = ~w1450 & w1456;
assign w1458 = ~w1392 & ~w1405;
assign w1459 = ~w1398 & w1458;
assign w1460 = w1398 & ~w1458;
assign w1461 = ~w1459 & ~w1460;
assign w1462 = ~w1457 & ~w1461;
assign w1463 = (w1455 & w1450) | (w1455 & w6136) | (w1450 & w6136);
assign w1464 = w1092 & ~w1463;
assign w1465 = ~w1462 & w1464;
assign w1466 = w553 & w1092;
assign w1467 = w1463 & ~w1466;
assign w1468 = ~w1457 & ~w1466;
assign w1469 = ~w1461 & w1468;
assign w1470 = ~w1467 & ~w1469;
assign w1471 = ~w1411 & w1415;
assign w1472 = ~w1416 & ~w1471;
assign w1473 = w1470 & ~w1472;
assign w1474 = (w1449 & w1473) | (w1449 & w6137) | (w1473 & w6137);
assign w1475 = w1390 & w1423;
assign w1476 = ~w1424 & ~w1475;
assign w1477 = ~w1473 & w6138;
assign w1478 = (w1088 & w1473) | (w1088 & w6752) | (w1473 & w6752);
assign w1479 = (w1478 & w1476) | (w1478 & w6753) | (w1476 & w6753);
assign w1480 = w553 & ~w1479;
assign w1481 = w1448 & w1480;
assign w1482 = ~w180 & w1088;
assign w1483 = ~w1426 & ~w1482;
assign w1484 = w1426 & w1482;
assign w1485 = ~w1483 & ~w1484;
assign w1486 = ~w1431 & w1485;
assign w1487 = w1434 & w1486;
assign w1488 = w1481 & ~w1487;
assign w1489 = w1434 & ~w1486;
assign w1490 = ~w180 & ~w1489;
assign w1491 = ~w1435 & w1490;
assign w1492 = w1385 & w1488;
assign w1493 = ~w1491 & w1492;
assign w1494 = w553 & ~w1493;
assign w1495 = w1385 & w1491;
assign w1496 = w1491 & w6754;
assign w1497 = w1437 & ~w1495;
assign w1498 = ~w1496 & ~w1497;
assign w1499 = w1494 & w1498;
assign w1500 = ~w1448 & ~w1480;
assign w1501 = ~w1481 & ~w1500;
assign w1502 = ~w930 & w1002;
assign w1503 = ~w103 & w1092;
assign w1504 = (~w1503 & w1003) | (~w1503 & w6139) | (w1003 & w6139);
assign w1505 = ~w1502 & w1504;
assign w1506 = ~w1457 & ~w1463;
assign w1507 = w1461 & ~w1506;
assign w1508 = ~w1461 & w1506;
assign w1509 = ~w1507 & ~w1508;
assign w1510 = ~w1505 & ~w1509;
assign w1511 = ~w103 & w1090;
assign w1512 = (w1503 & w1502) | (w1503 & w6140) | (w1502 & w6140);
assign w1513 = ~w1511 & ~w1512;
assign w1514 = ~w1510 & w1513;
assign w1515 = (~w6404 & w6755) | (~w6404 & w6756) | (w6755 & w6756);
assign w1516 = (w1511 & w1502) | (w1511 & w6141) | (w1502 & w6141);
assign w1517 = ~w1509 & w1516;
assign w1518 = (w1502 & w6405) | (w1502 & w6406) | (w6405 & w6406);
assign w1519 = ~w1517 & ~w1518;
assign w1520 = ~w1514 & w1519;
assign w1521 = (w1472 & ~w1470) | (w1472 & w6407) | (~w1470 & w6407);
assign w1522 = w1470 & w6408;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = w1520 & ~w1523;
assign w1525 = w1520 & w6757;
assign w1526 = (~w1515 & ~w1520) | (~w1515 & w6758) | (~w1520 & w6758);
assign w1527 = ~w1474 & ~w1477;
assign w1528 = w1476 & ~w1527;
assign w1529 = ~w1476 & w1527;
assign w1530 = ~w1528 & ~w1529;
assign w1531 = ~w1526 & w1530;
assign w1532 = ~w1525 & ~w1531;
assign w1533 = ~w1487 & ~w1532;
assign w1534 = w1501 & w1533;
assign w1535 = ~w1491 & w1534;
assign w1536 = ~w103 & ~w1535;
assign w1537 = (w1385 & w1491) | (w1385 & w1492) | (w1491 & w1492);
assign w1538 = ~w1491 & w6759;
assign w1539 = ~w1537 & ~w1538;
assign w1540 = w1536 & ~w1539;
assign w1541 = ~w1494 & ~w1498;
assign w1542 = ~w1499 & ~w1541;
assign w1543 = w1540 & w1542;
assign w1544 = (~w1499 & ~w1542) | (~w1499 & w6760) | (~w1542 & w6760);
assign w1545 = w1446 & ~w1544;
assign w1546 = ~w1379 & w1382;
assign w1547 = ~w1383 & ~w1546;
assign w1548 = w1547 & w7479;
assign w1549 = (w1325 & w1548) | (w1325 & w6762) | (w1548 & w6762);
assign w1550 = (w1548 & w6763) | (w1548 & w6764) | (w6763 & w6764);
assign w1551 = w1319 & w6765;
assign w1552 = (w1548 & w6768) | (w1548 & w6769) | (w6768 & w6769);
assign w1553 = ~w1130 & w7480;
assign w1554 = w1552 & ~w1553;
assign w1555 = ~w1552 & w1553;
assign w1556 = ~w1554 & ~w1555;
assign w1557 = ~w220 & ~w1556;
assign w1558 = (~w1194 & ~w1319) | (~w1194 & w6771) | (~w1319 & w6771);
assign w1559 = ~w1551 & ~w1558;
assign w1560 = ~w1559 & ~w1549;
assign w1561 = ~w1550 & ~w1560;
assign w1562 = ~w1548 & w6772;
assign w1563 = ~w1549 & ~w1562;
assign w1564 = ~w301 & w1563;
assign w1565 = (w1544 & w6773) | (w1544 & w6774) | (w6773 & w6774);
assign w1566 = ~w1548 & ~w1565;
assign w1567 = ~w1446 & w1544;
assign w1568 = ~w1545 & ~w1567;
assign w1569 = ~w1540 & ~w1542;
assign w1570 = ~w1543 & ~w1569;
assign w1571 = ~w1536 & w1539;
assign w1572 = ~w1540 & ~w1571;
assign w1573 = ~w301 & w1572;
assign w1574 = ~w1501 & w1532;
assign w1575 = w1501 & ~w1532;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = w342 & ~w1576;
assign w1578 = ~w1520 & w1523;
assign w1579 = ~w1524 & ~w1578;
assign w1580 = w342 & ~w1579;
assign w1581 = ~w1505 & ~w1512;
assign w1582 = ~w1509 & ~w1581;
assign w1583 = w1509 & w1581;
assign w1584 = ~w1582 & ~w1583;
assign w1585 = (~w1012 & w1584) | (~w1012 & w6775) | (w1584 & w6775);
assign w1586 = w1580 & ~w1585;
assign w1587 = ~w1525 & ~w1526;
assign w1588 = ~w1530 & w1587;
assign w1589 = w1530 & ~w1587;
assign w1590 = ~w1588 & ~w1589;
assign w1591 = w1586 & w1590;
assign w1592 = w342 & w1590;
assign w1593 = ~w1586 & ~w1592;
assign w1594 = ~w403 & w1012;
assign w1595 = ~w1584 & ~w1594;
assign w1596 = ~w1579 & w6776;
assign w1597 = (w1595 & w1579) | (w1595 & w6777) | (w1579 & w6777);
assign w1598 = ~w1596 & ~w1597;
assign w1599 = ~w1593 & w6778;
assign w1600 = ~w1591 & ~w1599;
assign w1601 = w1577 & ~w1600;
assign w1602 = ~w1577 & w1600;
assign w1603 = ~w1601 & ~w1602;
assign w1604 = ~w403 & w1590;
assign w1605 = ~w1584 & w1594;
assign w1606 = w1579 & ~w1605;
assign w1607 = ~w1579 & w6779;
assign w1608 = ~w1606 & ~w1607;
assign w1609 = ~w1604 & w1608;
assign w1610 = w1604 & ~w1608;
assign w1611 = ~w1609 & ~w1610;
assign w1612 = w1603 & ~w1611;
assign w1613 = ~w1603 & w1611;
assign w1614 = ~w1612 & ~w1613;
assign w1615 = ~w301 & ~w1576;
assign w1616 = ~w301 & w1012;
assign w1617 = ~w1584 & w6780;
assign w1618 = ~w1579 & w1617;
assign w1619 = (~w1617 & w1579) | (~w1617 & w6781) | (w1579 & w6781);
assign w1620 = ~w1618 & ~w1619;
assign w1621 = (w1594 & w1584) | (w1594 & w6782) | (w1584 & w6782);
assign w1622 = ~w1584 & w6783;
assign w1623 = ~w1621 & ~w1622;
assign w1624 = ~w1619 & w6409;
assign w1625 = (~w1618 & ~w6409) | (~w1618 & w6784) | (~w6409 & w6784);
assign w1626 = ~w301 & w1590;
assign w1627 = w1625 & ~w1626;
assign w1628 = w1590 & ~w1625;
assign w1629 = ~w1627 & ~w1628;
assign w1630 = ~w1585 & ~w1605;
assign w1631 = w342 & w1012;
assign w1632 = (w1579 & w6786) | (w1579 & w6787) | (w6786 & w6787);
assign w1633 = ~w1586 & ~w1632;
assign w1634 = w1629 & ~w1633;
assign w1635 = (~w1627 & ~w1629) | (~w1627 & w6788) | (~w1629 & w6788);
assign w1636 = ~w1615 & ~w1635;
assign w1637 = (w1598 & w1593) | (w1598 & w6789) | (w1593 & w6789);
assign w1638 = ~w1599 & ~w1637;
assign w1639 = w1615 & w1635;
assign w1640 = ~w1636 & ~w1639;
assign w1641 = ~w1638 & w1640;
assign w1642 = (~w1636 & ~w1640) | (~w1636 & w6790) | (~w1640 & w6790);
assign w1643 = ~w1614 & ~w1642;
assign w1644 = (~w1487 & ~w1490) | (~w1487 & w6791) | (~w1490 & w6791);
assign w1645 = (~w1481 & w1532) | (~w1481 & w6410) | (w1532 & w6410);
assign w1646 = w1644 & ~w1645;
assign w1647 = ~w1644 & w1645;
assign w1648 = ~w1646 & ~w1647;
assign w1649 = ~w301 & ~w1648;
assign w1650 = w1614 & w1642;
assign w1651 = ~w1643 & ~w1650;
assign w1652 = ~w1649 & w1651;
assign w1653 = (~w1643 & ~w1651) | (~w1643 & w6792) | (~w1651 & w6792);
assign w1654 = ~w1573 & ~w1653;
assign w1655 = w342 & ~w1648;
assign w1656 = (~w1601 & ~w1603) | (~w1601 & w6793) | (~w1603 & w6793);
assign w1657 = ~w403 & ~w1576;
assign w1658 = w1590 & w6794;
assign w1659 = ~w1590 & ~w1607;
assign w1660 = ~w1658 & ~w1659;
assign w1661 = w1657 & ~w1660;
assign w1662 = ~w1657 & w1660;
assign w1663 = ~w1661 & ~w1662;
assign w1664 = ~w1656 & ~w1663;
assign w1665 = w1656 & w1663;
assign w1666 = ~w1664 & ~w1665;
assign w1667 = w1655 & w1666;
assign w1668 = ~w1655 & ~w1666;
assign w1669 = ~w1667 & ~w1668;
assign w1670 = w1573 & w1653;
assign w1671 = ~w1654 & ~w1670;
assign w1672 = ~w1669 & w1671;
assign w1673 = (~w1654 & ~w1671) | (~w1654 & w6795) | (~w1671 & w6795);
assign w1674 = w1570 & w1673;
assign w1675 = w342 & w1572;
assign w1676 = (~w1664 & ~w1666) | (~w1664 & w6796) | (~w1666 & w6796);
assign w1677 = ~w403 & ~w1648;
assign w1678 = w1576 & ~w1658;
assign w1679 = ~w1576 & w6797;
assign w1680 = ~w1678 & ~w1679;
assign w1681 = w1677 & ~w1680;
assign w1682 = ~w1677 & w1680;
assign w1683 = ~w1681 & ~w1682;
assign w1684 = w1676 & w1683;
assign w1685 = ~w1676 & ~w1683;
assign w1686 = ~w1684 & ~w1685;
assign w1687 = ~w1675 & w1686;
assign w1688 = w1675 & ~w1686;
assign w1689 = ~w1687 & ~w1688;
assign w1690 = ~w301 & w1570;
assign w1691 = ~w1673 & ~w1690;
assign w1692 = ~w1674 & ~w1691;
assign w1693 = ~w1689 & w1692;
assign w1694 = (~w1674 & ~w1692) | (~w1674 & w6798) | (~w1692 & w6798);
assign w1695 = w1568 & ~w1694;
assign w1696 = w342 & w1570;
assign w1697 = (~w1684 & ~w1686) | (~w1684 & w6799) | (~w1686 & w6799);
assign w1698 = ~w403 & w1572;
assign w1699 = w1677 & ~w1678;
assign w1700 = w1648 & ~w1679;
assign w1701 = ~w1699 & ~w1700;
assign w1702 = ~w1698 & w1701;
assign w1703 = w1698 & ~w1701;
assign w1704 = ~w1702 & ~w1703;
assign w1705 = w1697 & ~w1704;
assign w1706 = ~w1697 & w1704;
assign w1707 = ~w1705 & ~w1706;
assign w1708 = w1696 & w1707;
assign w1709 = ~w1696 & ~w1707;
assign w1710 = ~w1708 & ~w1709;
assign w1711 = ~w301 & w1568;
assign w1712 = w1694 & ~w1711;
assign w1713 = ~w1695 & ~w1712;
assign w1714 = w1710 & w1713;
assign w1715 = (~w1695 & ~w1713) | (~w1695 & w6800) | (~w1713 & w6800);
assign w1716 = w1566 & ~w1715;
assign w1717 = ~w301 & w1566;
assign w1718 = w1715 & ~w1717;
assign w1719 = w342 & w1568;
assign w1720 = ~w1572 & ~w1699;
assign w1721 = w1572 & w6801;
assign w1722 = ~w1720 & ~w1721;
assign w1723 = (w1722 & ~w1570) | (w1722 & w6802) | (~w1570 & w6802);
assign w1724 = w1570 & w6803;
assign w1725 = ~w1723 & ~w1724;
assign w1726 = (~w1705 & ~w1707) | (~w1705 & w6804) | (~w1707 & w6804);
assign w1727 = ~w1725 & ~w1726;
assign w1728 = w1725 & w1726;
assign w1729 = ~w1727 & ~w1728;
assign w1730 = w1719 & w1729;
assign w1731 = ~w1719 & ~w1729;
assign w1732 = ~w1730 & ~w1731;
assign w1733 = ~w1718 & w1732;
assign w1734 = ~w1733 & w6805;
assign w1735 = (w1563 & w1733) | (w1563 & w6806) | (w1733 & w6806);
assign w1736 = w342 & w1566;
assign w1737 = ~w403 & w1568;
assign w1738 = ~w1720 & ~w1723;
assign w1739 = ~w1737 & ~w1738;
assign w1740 = w1568 & w1738;
assign w1741 = ~w1739 & ~w1740;
assign w1742 = ~w1570 & w1741;
assign w1743 = w1570 & ~w1741;
assign w1744 = ~w1742 & ~w1743;
assign w1745 = (~w1727 & ~w1729) | (~w1727 & w6807) | (~w1729 & w6807);
assign w1746 = ~w1744 & ~w1745;
assign w1747 = w1744 & w1745;
assign w1748 = ~w1746 & ~w1747;
assign w1749 = w1736 & w1748;
assign w1750 = ~w1736 & ~w1748;
assign w1751 = ~w1749 & ~w1750;
assign w1752 = ~w1735 & ~w1751;
assign w1753 = ~w1752 & w6808;
assign w1754 = w342 & w1563;
assign w1755 = (~w1746 & ~w1748) | (~w1746 & w6809) | (~w1748 & w6809);
assign w1756 = ~w403 & w1566;
assign w1757 = ~w1723 & w6811;
assign w1758 = ~w1568 & ~w1757;
assign w1759 = (w1741 & w6812) | (w1741 & w6813) | (w6812 & w6813);
assign w1760 = ~w1756 & w1759;
assign w1761 = w1756 & ~w1759;
assign w1762 = ~w1760 & ~w1761;
assign w1763 = ~w1755 & ~w1762;
assign w1764 = w1755 & w1762;
assign w1765 = ~w1763 & ~w1764;
assign w1766 = w1754 & w1765;
assign w1767 = ~w1754 & ~w1765;
assign w1768 = ~w1766 & ~w1767;
assign w1769 = ~w301 & w1561;
assign w1770 = (~w1769 & w1752) | (~w1769 & w6814) | (w1752 & w6814);
assign w1771 = ~w1753 & ~w1770;
assign w1772 = w1768 & w1771;
assign w1773 = w1192 & w7481;
assign w1774 = ~w1552 & ~w1773;
assign w1775 = ~w301 & w1774;
assign w1776 = ~w1772 & w6815;
assign w1777 = (w1774 & w1772) | (w1774 & w6816) | (w1772 & w6816);
assign w1778 = ~w1776 & ~w1777;
assign w1779 = w342 & w1561;
assign w1780 = (~w1763 & ~w1765) | (~w1763 & w6817) | (~w1765 & w6817);
assign w1781 = ~w403 & w1563;
assign w1782 = (w1741 & w6818) | (w1741 & w6819) | (w6818 & w6819);
assign w1783 = w1756 & ~w1758;
assign w1784 = ~w1782 & w6820;
assign w1785 = (w1781 & w1782) | (w1781 & w6821) | (w1782 & w6821);
assign w1786 = ~w1784 & ~w1785;
assign w1787 = ~w1780 & ~w1786;
assign w1788 = w1780 & w1786;
assign w1789 = ~w1787 & ~w1788;
assign w1790 = w1779 & w1789;
assign w1791 = ~w1779 & ~w1789;
assign w1792 = ~w1790 & ~w1791;
assign w1793 = w1778 & ~w1792;
assign w1794 = ~w1778 & w1792;
assign w1795 = ~w1793 & ~w1794;
assign w1796 = ~w220 & w1561;
assign w1797 = ~w220 & w1563;
assign w1798 = ~w220 & w1566;
assign w1799 = ~w220 & w1568;
assign w1800 = ~w220 & w1570;
assign w1801 = ~w220 & w1572;
assign w1802 = ~w220 & ~w1576;
assign w1803 = ~w220 & ~w1579;
assign w1804 = ~w220 & w1012;
assign w1805 = (~w301 & ~w1012) | (~w301 & w6822) | (~w1012 & w6822);
assign w1806 = (~w1631 & w1584) | (~w1631 & w6823) | (w1584 & w6823);
assign w1807 = ~w1584 & w1804;
assign w1808 = ~w1584 & w6824;
assign w1809 = (~w1808 & ~w1803) | (~w1808 & w6825) | (~w1803 & w6825);
assign w1810 = ~w220 & w1590;
assign w1811 = w1809 & ~w1810;
assign w1812 = w1590 & ~w1809;
assign w1813 = ~w1811 & ~w1812;
assign w1814 = ~w1620 & w1623;
assign w1815 = ~w1624 & ~w1814;
assign w1816 = w1813 & ~w1815;
assign w1817 = (~w1811 & ~w1813) | (~w1811 & w6411) | (~w1813 & w6411);
assign w1818 = w1802 & w1817;
assign w1819 = ~w1629 & w1633;
assign w1820 = ~w1634 & ~w1819;
assign w1821 = ~w1802 & ~w1817;
assign w1822 = ~w1818 & ~w1821;
assign w1823 = ~w1820 & w1822;
assign w1824 = (~w1818 & ~w1822) | (~w1818 & w6826) | (~w1822 & w6826);
assign w1825 = ~w1648 & ~w1824;
assign w1826 = w1638 & ~w1640;
assign w1827 = ~w1641 & ~w1826;
assign w1828 = ~w220 & ~w1648;
assign w1829 = w1824 & ~w1828;
assign w1830 = ~w1825 & ~w1829;
assign w1831 = ~w1827 & w1830;
assign w1832 = (~w1825 & ~w1830) | (~w1825 & w6827) | (~w1830 & w6827);
assign w1833 = ~w1801 & w1832;
assign w1834 = w1801 & ~w1832;
assign w1835 = ~w1833 & ~w1834;
assign w1836 = w1649 & ~w1651;
assign w1837 = ~w1652 & ~w1836;
assign w1838 = w1835 & w1837;
assign w1839 = ~w1838 & w6828;
assign w1840 = (~w1800 & w1838) | (~w1800 & w6829) | (w1838 & w6829);
assign w1841 = w1669 & ~w1671;
assign w1842 = ~w1672 & ~w1841;
assign w1843 = (~w1839 & w1842) | (~w1839 & w6830) | (w1842 & w6830);
assign w1844 = ~w1799 & w1843;
assign w1845 = w1689 & ~w1692;
assign w1846 = ~w1693 & ~w1845;
assign w1847 = w1799 & ~w1843;
assign w1848 = ~w1844 & ~w1847;
assign w1849 = ~w1846 & w1848;
assign w1850 = ~w1849 & w6831;
assign w1851 = (~w1798 & w1849) | (~w1798 & w6832) | (w1849 & w6832);
assign w1852 = ~w1850 & ~w1851;
assign w1853 = ~w1710 & ~w1713;
assign w1854 = ~w1714 & ~w1853;
assign w1855 = w1852 & w1854;
assign w1856 = (w1797 & w1855) | (w1797 & w6833) | (w1855 & w6833);
assign w1857 = ~w1855 & w6834;
assign w1858 = ~w1856 & ~w1857;
assign w1859 = ~w1716 & ~w1718;
assign w1860 = ~w1732 & w1859;
assign w1861 = w1732 & ~w1859;
assign w1862 = ~w1860 & ~w1861;
assign w1863 = w1858 & ~w1862;
assign w1864 = (w1796 & w1863) | (w1796 & w6835) | (w1863 & w6835);
assign w1865 = ~w1863 & w6836;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = ~w1734 & ~w1735;
assign w1868 = w1751 & ~w1867;
assign w1869 = ~w1751 & w1867;
assign w1870 = ~w1868 & ~w1869;
assign w1871 = w1866 & ~w1870;
assign w1872 = (~w1864 & ~w1866) | (~w1864 & w6837) | (~w1866 & w6837);
assign w1873 = ~w1768 & ~w1771;
assign w1874 = ~w1772 & ~w1873;
assign w1875 = ~w1872 & w1874;
assign w1876 = ~w220 & w1774;
assign w1877 = w1872 & ~w1874;
assign w1878 = ~w1875 & ~w1877;
assign w1879 = w1876 & w1878;
assign w1880 = (~w1875 & ~w1878) | (~w1875 & w6838) | (~w1878 & w6838);
assign w1881 = ~w1795 & ~w1880;
assign w1882 = w1795 & w1880;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = w1557 & w1883;
assign w1885 = ~w1557 & ~w1883;
assign w1886 = ~w1884 & ~w1885;
assign w1887 = ~w1866 & w1870;
assign w1888 = ~w1871 & ~w1887;
assign w1889 = ~w253 & w1570;
assign w1890 = ~w253 & w1572;
assign w1891 = ~w253 & ~w1648;
assign w1892 = ~w253 & ~w1576;
assign w1893 = (~w253 & ~w1579) | (~w253 & w6412) | (~w1579 & w6412);
assign w1894 = ~w1584 & w6413;
assign w1895 = (w1616 & w1584) | (w1616 & w6414) | (w1584 & w6414);
assign w1896 = ~w1894 & ~w1895;
assign w1897 = (w1896 & w1579) | (w1896 & w6839) | (w1579 & w6839);
assign w1898 = w1893 & ~w1897;
assign w1899 = w1590 & w1898;
assign w1900 = w220 & w1617;
assign w1901 = (w1806 & w1579) | (w1806 & w6840) | (w1579 & w6840);
assign w1902 = (~w1900 & ~w1803) | (~w1900 & w6841) | (~w1803 & w6841);
assign w1903 = ~w1901 & w1902;
assign w1904 = ~w253 & w1530;
assign w1905 = w1587 & w1904;
assign w1906 = ~w253 & ~w1530;
assign w1907 = ~w1587 & w1906;
assign w1908 = ~w1905 & ~w1907;
assign w1909 = ~w1898 & w1908;
assign w1910 = w1903 & ~w1909;
assign w1911 = ~w1899 & ~w1910;
assign w1912 = w1892 & ~w1911;
assign w1913 = ~w1813 & w1815;
assign w1914 = ~w1816 & ~w1913;
assign w1915 = ~w1892 & w1911;
assign w1916 = ~w1912 & ~w1915;
assign w1917 = ~w1914 & w1916;
assign w1918 = (w1891 & w1917) | (w1891 & w6415) | (w1917 & w6415);
assign w1919 = w1820 & ~w1822;
assign w1920 = ~w1823 & ~w1919;
assign w1921 = ~w1917 & w6416;
assign w1922 = ~w1918 & ~w1921;
assign w1923 = w1920 & w1922;
assign w1924 = (w1890 & w1923) | (w1890 & w6842) | (w1923 & w6842);
assign w1925 = w1827 & ~w1830;
assign w1926 = ~w1831 & ~w1925;
assign w1927 = ~w1923 & w6843;
assign w1928 = ~w1924 & ~w1927;
assign w1929 = w1926 & w1928;
assign w1930 = (w1889 & w1929) | (w1889 & w6844) | (w1929 & w6844);
assign w1931 = ~w1835 & ~w1837;
assign w1932 = ~w1838 & ~w1931;
assign w1933 = ~w1929 & w6845;
assign w1934 = ~w1930 & ~w1933;
assign w1935 = ~w1932 & w1934;
assign w1936 = (w1568 & w1935) | (w1568 & w6846) | (w1935 & w6846);
assign w1937 = ~w253 & w1568;
assign w1938 = ~w1935 & w6847;
assign w1939 = ~w1936 & ~w1938;
assign w1940 = ~w1839 & ~w1840;
assign w1941 = w1842 & ~w1940;
assign w1942 = ~w1842 & w1940;
assign w1943 = ~w1941 & ~w1942;
assign w1944 = w1939 & w1943;
assign w1945 = ~w253 & w1566;
assign w1946 = ~w1944 & w6848;
assign w1947 = w1846 & ~w1848;
assign w1948 = ~w1849 & ~w1947;
assign w1949 = (w1566 & w1944) | (w1566 & w6849) | (w1944 & w6849);
assign w1950 = (~w1946 & ~w1948) | (~w1946 & w6850) | (~w1948 & w6850);
assign w1951 = w1563 & w1950;
assign w1952 = ~w1852 & ~w1854;
assign w1953 = ~w1855 & ~w1952;
assign w1954 = ~w253 & w1563;
assign w1955 = ~w1950 & ~w1954;
assign w1956 = ~w1951 & ~w1955;
assign w1957 = w1953 & w1956;
assign w1958 = (w1561 & w1957) | (w1561 & w6851) | (w1957 & w6851);
assign w1959 = ~w1858 & w1862;
assign w1960 = ~w1863 & ~w1959;
assign w1961 = ~w253 & w1561;
assign w1962 = ~w1957 & w6852;
assign w1963 = ~w1958 & ~w1962;
assign w1964 = w1960 & w1963;
assign w1965 = (w1774 & w1964) | (w1774 & w6853) | (w1964 & w6853);
assign w1966 = ~w253 & w1774;
assign w1967 = ~w1964 & w6854;
assign w1968 = ~w1965 & ~w1967;
assign w1969 = w1888 & w1968;
assign w1970 = (w1553 & w1964) | (w1553 & w6855) | (w1964 & w6855);
assign w1971 = w1965 & w1970;
assign w1972 = (~w1971 & ~w1969) | (~w1971 & w6856) | (~w1969 & w6856);
assign w1973 = ~w1876 & ~w1878;
assign w1974 = ~w1879 & ~w1973;
assign w1975 = ~w253 & ~w1556;
assign w1976 = ~w1975 & ~w1965;
assign w1977 = ~w1969 & w1976;
assign w1978 = w1972 & ~w1977;
assign w1979 = w1974 & w1978;
assign w1980 = ~w253 & w1972;
assign w1981 = ~w1979 & w1980;
assign w1982 = ~w1886 & w1981;
assign w1983 = (~w253 & w1886) | (~w253 & w6857) | (w1886 & w6857);
assign w1984 = w342 & w1774;
assign w1985 = (~w1984 & w1784) | (~w1984 & w6858) | (w1784 & w6858);
assign w1986 = ~w403 & w1561;
assign w1987 = ~w1563 & ~w1986;
assign w1988 = w1559 & w1563;
assign w1989 = w1563 & w6859;
assign w1990 = ~w1987 & ~w1989;
assign w1991 = w1985 & ~w1990;
assign w1992 = ~w1985 & w1990;
assign w1993 = ~w1991 & ~w1992;
assign w1994 = (~w1787 & ~w1789) | (~w1787 & w6860) | (~w1789 & w6860);
assign w1995 = ~w220 & ~w1881;
assign w1996 = (w1994 & w1884) | (w1994 & w6861) | (w1884 & w6861);
assign w1997 = ~w1884 & w6862;
assign w1998 = ~w1996 & ~w1997;
assign w1999 = (w1556 & w1793) | (w1556 & w6863) | (w1793 & w6863);
assign w2000 = (~w301 & w1793) | (~w301 & w6864) | (w1793 & w6864);
assign w2001 = ~w1556 & ~w2000;
assign w2002 = ~w1999 & ~w2001;
assign w2003 = w1998 & ~w2002;
assign w2004 = ~w1998 & w2002;
assign w2005 = ~w2003 & ~w2004;
assign w2006 = ~w1993 & ~w2005;
assign w2007 = (~w1983 & ~w2005) | (~w1983 & w6865) | (~w2005 & w6865);
assign w2008 = ~w2006 & w2007;
assign w2009 = ~w103 & ~w1556;
assign w2010 = ~w103 & w1774;
assign w2011 = ~w177 & w1566;
assign w2012 = ~w177 & w1568;
assign w2013 = ~w177 & w1570;
assign w2014 = ~w177 & w1572;
assign w2015 = (~w1804 & w1584) | (~w1804 & w6866) | (w1584 & w6866);
assign w2016 = ~w177 & w1012;
assign w2017 = (~w253 & ~w1012) | (~w253 & w254) | (~w1012 & w254);
assign w2018 = (~w1804 & w1584) | (~w1804 & w6867) | (w1584 & w6867);
assign w2019 = ~w177 & ~w1523;
assign w2020 = w1520 & w2019;
assign w2021 = ~w177 & w1523;
assign w2022 = ~w1520 & w2021;
assign w2023 = ~w2020 & ~w2022;
assign w2024 = (~w2015 & ~w2023) | (~w2015 & w6142) | (~w2023 & w6142);
assign w2025 = w1590 & w2024;
assign w2026 = ~w1579 & w6868;
assign w2027 = (w1579 & w6869) | (w1579 & w6870) | (w6869 & w6870);
assign w2028 = (~w2027 & ~w1898) | (~w2027 & w6871) | (~w1898 & w6871);
assign w2029 = ~w177 & ~w2024;
assign w2030 = w1590 & w2029;
assign w2031 = ~w1590 & w2024;
assign w2032 = ~w2030 & ~w2031;
assign w2033 = w2028 & ~w2032;
assign w2034 = (~w2025 & w2032) | (~w2025 & w6872) | (w2032 & w6872);
assign w2035 = ~w177 & ~w1576;
assign w2036 = ~w1899 & ~w1909;
assign w2037 = ~w1903 & w2036;
assign w2038 = w1903 & ~w2036;
assign w2039 = ~w2037 & ~w2038;
assign w2040 = ~w2035 & w2039;
assign w2041 = (~w2034 & ~w2039) | (~w2034 & w6873) | (~w2039 & w6873);
assign w2042 = w2035 & ~w2039;
assign w2043 = ~w177 & ~w1648;
assign w2044 = ~w2042 & ~w2043;
assign w2045 = ~w2041 & w2044;
assign w2046 = w1914 & ~w1916;
assign w2047 = ~w1917 & ~w2046;
assign w2048 = (w2034 & w2039) | (w2034 & w6874) | (w2039 & w6874);
assign w2049 = ~w2040 & w2043;
assign w2050 = ~w2048 & w2049;
assign w2051 = ~w2045 & ~w2050;
assign w2052 = ~w2047 & w2051;
assign w2053 = (~w2045 & ~w2051) | (~w2045 & w6417) | (~w2051 & w6417);
assign w2054 = w2014 & w2053;
assign w2055 = ~w2014 & ~w2053;
assign w2056 = ~w2054 & ~w2055;
assign w2057 = ~w1920 & ~w1922;
assign w2058 = ~w1923 & ~w2057;
assign w2059 = w2056 & w2058;
assign w2060 = (~w2054 & ~w2056) | (~w2054 & w6875) | (~w2056 & w6875);
assign w2061 = ~w2013 & w2060;
assign w2062 = w2013 & ~w2060;
assign w2063 = ~w2061 & ~w2062;
assign w2064 = ~w1926 & ~w1928;
assign w2065 = ~w1929 & ~w2064;
assign w2066 = w2063 & ~w2065;
assign w2067 = (~w2061 & ~w2063) | (~w2061 & w6876) | (~w2063 & w6876);
assign w2068 = w2012 & w2067;
assign w2069 = w1932 & ~w1934;
assign w2070 = ~w1935 & ~w2069;
assign w2071 = ~w2012 & ~w2067;
assign w2072 = ~w2068 & ~w2071;
assign w2073 = w2070 & w2072;
assign w2074 = (~w2068 & ~w2072) | (~w2068 & w6877) | (~w2072 & w6877);
assign w2075 = w2011 & ~w2074;
assign w2076 = ~w2011 & w2074;
assign w2077 = ~w2075 & ~w2076;
assign w2078 = ~w1939 & ~w1943;
assign w2079 = ~w1944 & ~w2078;
assign w2080 = w2077 & w2079;
assign w2081 = ~w2077 & ~w2079;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = ~w141 & w1566;
assign w2084 = ~w141 & w1568;
assign w2085 = ~w141 & w1570;
assign w2086 = ~w141 & ~w1648;
assign w2087 = ~w141 & ~w1576;
assign w2088 = ~w1584 & w6878;
assign w2089 = w2023 & w6879;
assign w2090 = w2018 & ~w2023;
assign w2091 = ~w2089 & ~w2090;
assign w2092 = ~w253 & w666;
assign w2093 = w930 & w2092;
assign w2094 = w1009 & w2093;
assign w2095 = ~w930 & w2092;
assign w2096 = ~w1009 & w2095;
assign w2097 = ~w2094 & ~w2096;
assign w2098 = w1582 & ~w2097;
assign w2099 = ~w253 & w1012;
assign w2100 = (w177 & ~w1012) | (w177 & w256) | (~w1012 & w256);
assign w2101 = w1509 & ~w2097;
assign w2102 = (~w2100 & ~w2101) | (~w2100 & w6418) | (~w2101 & w6418);
assign w2103 = ~w2098 & w2102;
assign w2104 = ~w141 & w930;
assign w2105 = w1009 & w2104;
assign w2106 = ~w141 & ~w930;
assign w2107 = ~w1009 & w2106;
assign w2108 = ~w2105 & ~w2107;
assign w2109 = w1583 & w2108;
assign w2110 = ~w1509 & w2108;
assign w2111 = (~w2099 & ~w2110) | (~w2099 & w6419) | (~w2110 & w6419);
assign w2112 = ~w2109 & w2111;
assign w2113 = w2103 & ~w2112;
assign w2114 = ~w141 & ~w1523;
assign w2115 = w1520 & w2114;
assign w2116 = ~w141 & w1523;
assign w2117 = ~w1520 & w2116;
assign w2118 = ~w2115 & ~w2117;
assign w2119 = w2113 & w2118;
assign w2120 = w1584 & ~w2099;
assign w2121 = w2103 & ~w2120;
assign w2122 = ~w2119 & w2121;
assign w2123 = w1590 & w2122;
assign w2124 = w2091 & ~w2123;
assign w2125 = (~w141 & w2119) | (~w141 & w6143) | (w2119 & w6143);
assign w2126 = w1590 & w2125;
assign w2127 = ~w2122 & ~w2126;
assign w2128 = ~w2124 & ~w2127;
assign w2129 = ~w2087 & ~w2128;
assign w2130 = w2087 & w2128;
assign w2131 = ~w2028 & w2032;
assign w2132 = ~w2033 & ~w2131;
assign w2133 = ~w2130 & ~w2132;
assign w2134 = ~w2133 & w6880;
assign w2135 = ~w2040 & ~w2042;
assign w2136 = ~w2034 & ~w2135;
assign w2137 = w2034 & w2135;
assign w2138 = ~w2136 & ~w2137;
assign w2139 = ~w141 & w1572;
assign w2140 = (~w2086 & w2133) | (~w2086 & w6881) | (w2133 & w6881);
assign w2141 = w2139 & ~w2140;
assign w2142 = (w2141 & ~w2138) | (w2141 & w6882) | (~w2138 & w6882);
assign w2143 = w2047 & ~w2051;
assign w2144 = ~w2052 & ~w2143;
assign w2145 = ~w2134 & ~w2139;
assign w2146 = (w2145 & w2138) | (w2145 & w6883) | (w2138 & w6883);
assign w2147 = ~w2144 & ~w2146;
assign w2148 = ~w2147 & w6420;
assign w2149 = (w2085 & w2147) | (w2085 & w6421) | (w2147 & w6421);
assign w2150 = ~w2148 & ~w2149;
assign w2151 = ~w2056 & ~w2058;
assign w2152 = ~w2059 & ~w2151;
assign w2153 = w2150 & ~w2152;
assign w2154 = ~w2153 & w6884;
assign w2155 = ~w2063 & w2065;
assign w2156 = ~w2066 & ~w2155;
assign w2157 = (~w2084 & w2153) | (~w2084 & w6885) | (w2153 & w6885);
assign w2158 = ~w2154 & ~w2157;
assign w2159 = ~w2156 & w2158;
assign w2160 = ~w2159 & w6886;
assign w2161 = (w2083 & w2159) | (w2083 & w6887) | (w2159 & w6887);
assign w2162 = ~w2160 & ~w2161;
assign w2163 = ~w2070 & ~w2072;
assign w2164 = ~w2073 & ~w2163;
assign w2165 = w2162 & ~w2164;
assign w2166 = ~w141 & w1563;
assign w2167 = (~w2166 & w2165) | (~w2166 & w6888) | (w2165 & w6888);
assign w2168 = ~w2165 & w6889;
assign w2169 = ~w2167 & ~w2168;
assign w2170 = ~w2082 & w2169;
assign w2171 = w2082 & ~w2169;
assign w2172 = ~w2170 & ~w2171;
assign w2173 = ~w103 & w1561;
assign w2174 = ~w2162 & w2164;
assign w2175 = ~w2165 & ~w2174;
assign w2176 = ~w103 & w1563;
assign w2177 = ~w103 & w1566;
assign w2178 = ~w2150 & w2152;
assign w2179 = ~w2153 & ~w2178;
assign w2180 = ~w2142 & ~w2146;
assign w2181 = w2144 & ~w2180;
assign w2182 = ~w2144 & w2180;
assign w2183 = ~w2181 & ~w2182;
assign w2184 = ~w103 & w1012;
assign w2185 = w1012 & w6890;
assign w2186 = ~w103 & w1523;
assign w2187 = ~w1520 & w2186;
assign w2188 = ~w1524 & ~w2187;
assign w2189 = ~w141 & w1461;
assign w2190 = ~w1506 & w2189;
assign w2191 = ~w141 & ~w1461;
assign w2192 = w1506 & w2191;
assign w2193 = ~w2190 & ~w2192;
assign w2194 = w2016 & w2193;
assign w2195 = w568 & ~w930;
assign w2196 = ~w2193 & ~w2195;
assign w2197 = ~w1581 & ~w2196;
assign w2198 = ~w2194 & w2197;
assign w2199 = ~w141 & w1509;
assign w2200 = ~w2016 & w6145;
assign w2201 = ~w2198 & ~w2200;
assign w2202 = (w2201 & ~w6144) | (w2201 & w6891) | (~w6144 & w6891);
assign w2203 = ~w2113 & ~w2118;
assign w2204 = ~w2119 & ~w2203;
assign w2205 = w2202 & ~w2204;
assign w2206 = ~w1590 & ~w2205;
assign w2207 = ~w2202 & w2204;
assign w2208 = (~w103 & ~w2204) | (~w103 & w6146) | (~w2204 & w6146);
assign w2209 = ~w2206 & w2208;
assign w2210 = ~w1531 & w6892;
assign w2211 = ~w1501 & w2210;
assign w2212 = ~w1575 & ~w2211;
assign w2213 = ~w2209 & w2212;
assign w2214 = ~w1590 & w2122;
assign w2215 = ~w2126 & ~w2214;
assign w2216 = ~w2091 & w2215;
assign w2217 = w2091 & ~w2215;
assign w2218 = ~w2216 & ~w2217;
assign w2219 = ~w2213 & ~w2218;
assign w2220 = ~w103 & w1646;
assign w2221 = ~w1576 & w2209;
assign w2222 = ~w1481 & w7482;
assign w2223 = ~w1644 & w2222;
assign w2224 = (~w2223 & ~w2209) | (~w2223 & w6894) | (~w2209 & w6894);
assign w2225 = ~w2220 & w2224;
assign w2226 = ~w2219 & w2225;
assign w2227 = ~w1535 & ~w1539;
assign w2228 = ~w1571 & ~w2227;
assign w2229 = w2226 & ~w2228;
assign w2230 = ~w2213 & ~w2221;
assign w2231 = w2218 & w2230;
assign w2232 = ~w1648 & ~w2213;
assign w2233 = ~w2231 & w2232;
assign w2234 = ~w2129 & ~w2130;
assign w2235 = ~w2132 & w2234;
assign w2236 = w2132 & ~w2234;
assign w2237 = ~w2235 & ~w2236;
assign w2238 = (~w2228 & w2231) | (~w2228 & w6895) | (w2231 & w6895);
assign w2239 = w2237 & w2238;
assign w2240 = ~w2229 & ~w2239;
assign w2241 = ~w2226 & ~w2233;
assign w2242 = w2237 & w2241;
assign w2243 = ~w2226 & w2228;
assign w2244 = (w2243 & ~w2241) | (w2243 & w6896) | (~w2241 & w6896);
assign w2245 = w2240 & ~w2244;
assign w2246 = ~w2134 & ~w2140;
assign w2247 = ~w2138 & w2246;
assign w2248 = w2138 & ~w2246;
assign w2249 = ~w2247 & ~w2248;
assign w2250 = w2245 & ~w2249;
assign w2251 = ~w103 & w1570;
assign w2252 = ~w2240 & ~w2251;
assign w2253 = w2240 & w2251;
assign w2254 = ~w2252 & ~w2253;
assign w2255 = ~w2250 & w2254;
assign w2256 = w2245 & w6147;
assign w2257 = ~w2255 & ~w2256;
assign w2258 = w2183 & ~w2257;
assign w2259 = ~w2250 & w6148;
assign w2260 = ~w103 & w1568;
assign w2261 = (w2260 & w2250) | (w2260 & w6149) | (w2250 & w6149);
assign w2262 = ~w2259 & ~w2261;
assign w2263 = w2258 & ~w2262;
assign w2264 = ~w2258 & w2262;
assign w2265 = ~w2263 & ~w2264;
assign w2266 = ~w2179 & w2265;
assign w2267 = w2260 & ~w2265;
assign w2268 = ~w2266 & ~w2267;
assign w2269 = w2177 & ~w2268;
assign w2270 = w2156 & ~w2158;
assign w2271 = ~w2159 & ~w2270;
assign w2272 = ~w2177 & w2268;
assign w2273 = ~w2269 & ~w2272;
assign w2274 = w2271 & w2273;
assign w2275 = (~w2269 & ~w2273) | (~w2269 & w6150) | (~w2273 & w6150);
assign w2276 = w2176 & ~w2275;
assign w2277 = ~w2176 & w2275;
assign w2278 = ~w2276 & ~w2277;
assign w2279 = ~w2175 & w2278;
assign w2280 = ~w2275 & w6897;
assign w2281 = (~w2280 & ~w2278) | (~w2280 & w6898) | (~w2278 & w6898);
assign w2282 = w2173 & ~w2281;
assign w2283 = (~w2173 & w2275) | (~w2173 & w6899) | (w2275 & w6899);
assign w2284 = (w2283 & ~w2278) | (w2283 & w6900) | (~w2278 & w6900);
assign w2285 = ~w2282 & ~w2284;
assign w2286 = ~w2282 & w6901;
assign w2287 = ~w2281 & w6902;
assign w2288 = (w2010 & w2286) | (w2010 & w6903) | (w2286 & w6903);
assign w2289 = ~w141 & w1561;
assign w2290 = (~w2289 & w2170) | (~w2289 & w6904) | (w2170 & w6904);
assign w2291 = ~w2170 & w6905;
assign w2292 = ~w2290 & ~w2291;
assign w2293 = ~w177 & w1563;
assign w2294 = (~w2075 & ~w2077) | (~w2075 & w6906) | (~w2077 & w6906);
assign w2295 = w2293 & ~w2294;
assign w2296 = ~w2293 & w2294;
assign w2297 = ~w2295 & ~w2296;
assign w2298 = ~w1946 & ~w1949;
assign w2299 = w1948 & w2298;
assign w2300 = ~w1948 & ~w2298;
assign w2301 = ~w2299 & ~w2300;
assign w2302 = w2297 & ~w2301;
assign w2303 = ~w2297 & w2301;
assign w2304 = ~w2302 & ~w2303;
assign w2305 = w2292 & ~w2304;
assign w2306 = ~w2292 & w2304;
assign w2307 = ~w2305 & ~w2306;
assign w2308 = (~w2010 & w2281) | (~w2010 & w6907) | (w2281 & w6907);
assign w2309 = ~w2286 & w2308;
assign w2310 = ~w2288 & ~w2309;
assign w2311 = ~w2307 & w2310;
assign w2312 = (~w2288 & ~w2310) | (~w2288 & w6908) | (~w2310 & w6908);
assign w2313 = ~w2009 & w2312;
assign w2314 = ~w177 & w1561;
assign w2315 = (~w2295 & ~w2297) | (~w2295 & w6909) | (~w2297 & w6909);
assign w2316 = ~w2314 & w2315;
assign w2317 = w2314 & ~w2315;
assign w2318 = ~w2316 & ~w2317;
assign w2319 = ~w1953 & ~w1956;
assign w2320 = ~w1957 & ~w2319;
assign w2321 = w2318 & ~w2320;
assign w2322 = ~w2318 & w2320;
assign w2323 = ~w2321 & ~w2322;
assign w2324 = ~w2305 & w6910;
assign w2325 = ~w141 & w1774;
assign w2326 = (~w2325 & w2305) | (~w2325 & w6911) | (w2305 & w6911);
assign w2327 = ~w2324 & ~w2326;
assign w2328 = ~w2323 & w2327;
assign w2329 = w2323 & ~w2327;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = w2009 & ~w2312;
assign w2332 = ~w2313 & ~w2331;
assign w2333 = ~w2330 & w2332;
assign w2334 = (~w2313 & ~w2332) | (~w2313 & w6912) | (~w2332 & w6912);
assign w2335 = ~w177 & w1774;
assign w2336 = ~w1960 & ~w1963;
assign w2337 = ~w1964 & ~w2336;
assign w2338 = (~w2316 & ~w2318) | (~w2316 & w6913) | (~w2318 & w6913);
assign w2339 = ~w2337 & ~w2338;
assign w2340 = w2337 & w2338;
assign w2341 = ~w2339 & ~w2340;
assign w2342 = ~w2335 & w2341;
assign w2343 = w2335 & ~w2341;
assign w2344 = ~w2342 & ~w2343;
assign w2345 = (~w1556 & w2328) | (~w1556 & w6914) | (w2328 & w6914);
assign w2346 = ~w141 & ~w1556;
assign w2347 = ~w2328 & w6915;
assign w2348 = ~w2345 & ~w2347;
assign w2349 = ~w2344 & w2348;
assign w2350 = w2344 & ~w2348;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = ~w2334 & ~w2351;
assign w2353 = w2334 & w2351;
assign w2354 = ~w2352 & ~w2353;
assign w2355 = w103 & w2354;
assign w2356 = (~w2352 & ~w2354) | (~w2352 & w6916) | (~w2354 & w6916);
assign w2357 = ~w177 & ~w1556;
assign w2358 = ~w1888 & ~w1968;
assign w2359 = ~w1969 & ~w2358;
assign w2360 = (~w2339 & ~w2341) | (~w2339 & w6917) | (~w2341 & w6917);
assign w2361 = w2359 & w2360;
assign w2362 = ~w2359 & ~w2360;
assign w2363 = ~w2361 & ~w2362;
assign w2364 = w2357 & w2363;
assign w2365 = ~w2357 & ~w2363;
assign w2366 = ~w2364 & ~w2365;
assign w2367 = (~w2345 & w2344) | (~w2345 & w6918) | (w2344 & w6918);
assign w2368 = ~w141 & w2367;
assign w2369 = w2366 & ~w2368;
assign w2370 = ~w2366 & w2368;
assign w2371 = ~w2369 & ~w2370;
assign w2372 = w2356 & ~w2371;
assign w2373 = ~w2356 & w2371;
assign w2374 = ~w2372 & ~w2373;
assign w2375 = w2330 & ~w2332;
assign w2376 = ~w2333 & ~w2375;
assign w2377 = ~w364 & w1774;
assign w2378 = ~w364 & w1561;
assign w2379 = ~w364 & w1563;
assign w2380 = ~w364 & w1566;
assign w2381 = ~w364 & w1568;
assign w2382 = ~w364 & w1570;
assign w2383 = ~w364 & w1572;
assign w2384 = ~w364 & ~w1648;
assign w2385 = ~w103 & ~w1461;
assign w2386 = ~w1506 & w2385;
assign w2387 = ~w103 & w1461;
assign w2388 = w1506 & w2387;
assign w2389 = ~w2386 & ~w2388;
assign w2390 = ~w2108 & w2389;
assign w2391 = w1581 & ~w2390;
assign w2392 = ~w141 & w364;
assign w2393 = w930 & w2392;
assign w2394 = w1009 & w2393;
assign w2395 = ~w930 & w2392;
assign w2396 = ~w1009 & w2395;
assign w2397 = ~w2394 & ~w2396;
assign w2398 = ~w1506 & ~w2387;
assign w2399 = w1506 & ~w2385;
assign w2400 = ~w2398 & ~w2399;
assign w2401 = w2397 & w2400;
assign w2402 = ~w1581 & ~w2401;
assign w2403 = ~w2391 & ~w2402;
assign w2404 = ~w2108 & ~w2400;
assign w2405 = ~w1581 & w2404;
assign w2406 = ~w2389 & w2397;
assign w2407 = w1581 & w2406;
assign w2408 = ~w2405 & ~w2407;
assign w2409 = ~w2403 & w2408;
assign w2410 = ~w364 & w930;
assign w2411 = w1009 & w2410;
assign w2412 = ~w364 & ~w930;
assign w2413 = ~w1009 & w2412;
assign w2414 = ~w2411 & ~w2413;
assign w2415 = ~w2389 & ~w2414;
assign w2416 = w1581 & ~w2415;
assign w2417 = w2400 & ~w2414;
assign w2418 = ~w1581 & ~w2417;
assign w2419 = ~w2416 & ~w2418;
assign w2420 = w141 & w2419;
assign w2421 = ~w364 & ~w1523;
assign w2422 = w1520 & w2421;
assign w2423 = ~w364 & w1523;
assign w2424 = ~w1520 & w2423;
assign w2425 = ~w2422 & ~w2424;
assign w2426 = (~w2409 & ~w2425) | (~w2409 & w6151) | (~w2425 & w6151);
assign w2427 = ~w2198 & w6919;
assign w2428 = ~w2188 & w2427;
assign w2429 = w2188 & ~w2427;
assign w2430 = ~w2428 & ~w2429;
assign w2431 = w2426 & w2430;
assign w2432 = ~w1590 & ~w2431;
assign w2433 = ~w2426 & ~w2430;
assign w2434 = (~w364 & w2430) | (~w364 & w6152) | (w2430 & w6152);
assign w2435 = ~w2432 & w2434;
assign w2436 = (~w364 & w1531) | (~w364 & w6920) | (w1531 & w6920);
assign w2437 = w1501 & ~w2436;
assign w2438 = ~w1531 & w6921;
assign w2439 = ~w1501 & ~w2438;
assign w2440 = ~w2437 & ~w2439;
assign w2441 = ~w2435 & ~w2440;
assign w2442 = ~w1576 & w2435;
assign w2443 = ~w103 & w1590;
assign w2444 = ~w2205 & ~w2207;
assign w2445 = ~w2443 & w2444;
assign w2446 = w2443 & ~w2444;
assign w2447 = ~w2445 & ~w2446;
assign w2448 = ~w2442 & w2447;
assign w2449 = (~w2384 & w2448) | (~w2384 & w6922) | (w2448 & w6922);
assign w2450 = ~w2448 & w6923;
assign w2451 = ~w2218 & ~w2230;
assign w2452 = ~w2231 & ~w2451;
assign w2453 = ~w2450 & w2452;
assign w2454 = (~w2449 & ~w2452) | (~w2449 & w6924) | (~w2452 & w6924);
assign w2455 = ~w2383 & ~w2454;
assign w2456 = ~w2453 & w6153;
assign w2457 = ~w2237 & ~w2241;
assign w2458 = ~w2242 & ~w2457;
assign w2459 = ~w2456 & w2458;
assign w2460 = ~w2459 & w6154;
assign w2461 = (~w2382 & w2459) | (~w2382 & w6155) | (w2459 & w6155);
assign w2462 = ~w2245 & w2249;
assign w2463 = ~w2250 & ~w2462;
assign w2464 = (w6156 & w6925) | (w6156 & w6926) | (w6925 & w6926);
assign w2465 = (~w6156 & w6927) | (~w6156 & w6928) | (w6927 & w6928);
assign w2466 = ~w2183 & w2257;
assign w2467 = ~w2258 & ~w2466;
assign w2468 = (~w2464 & w2467) | (~w2464 & w6157) | (w2467 & w6157);
assign w2469 = w2380 & w2468;
assign w2470 = ~w2380 & ~w2468;
assign w2471 = w2179 & ~w2265;
assign w2472 = ~w2266 & ~w2471;
assign w2473 = (~w2469 & ~w2472) | (~w2469 & w6158) | (~w2472 & w6158);
assign w2474 = ~w2379 & w2473;
assign w2475 = ~w2271 & ~w2273;
assign w2476 = ~w2274 & ~w2475;
assign w2477 = w2379 & ~w2473;
assign w2478 = ~w2474 & ~w2477;
assign w2479 = ~w2476 & w2478;
assign w2480 = (~w2474 & w2476) | (~w2474 & w6159) | (w2476 & w6159);
assign w2481 = ~w2378 & ~w2480;
assign w2482 = w2378 & w2480;
assign w2483 = ~w2481 & ~w2482;
assign w2484 = w2175 & ~w2278;
assign w2485 = ~w2279 & ~w2484;
assign w2486 = w2483 & ~w2485;
assign w2487 = (~w2377 & w2486) | (~w2377 & w6929) | (w2486 & w6929);
assign w2488 = w2172 & ~w2285;
assign w2489 = ~w2286 & ~w2488;
assign w2490 = w1561 & w6930;
assign w2491 = (~w2490 & ~w2480) | (~w2490 & w6931) | (~w2480 & w6931);
assign w2492 = ~w2486 & ~w2491;
assign w2493 = ~w2487 & ~w2492;
assign w2494 = ~w2489 & w2493;
assign w2495 = ~w364 & w1556;
assign w2496 = (w2495 & w2494) | (w2495 & w6932) | (w2494 & w6932);
assign w2497 = w2307 & ~w2310;
assign w2498 = ~w2311 & ~w2497;
assign w2499 = ~w2494 & w6933;
assign w2500 = ~w364 & ~w2496;
assign w2501 = w2500 & w6934;
assign w2502 = ~w2496 & ~w2501;
assign w2503 = w2376 & ~w2502;
assign w2504 = ~w364 & ~w2503;
assign w2505 = ~w103 & ~w2354;
assign w2506 = ~w2355 & ~w2505;
assign w2507 = w2504 & ~w2506;
assign w2508 = ~w2376 & w2502;
assign w2509 = ~w2503 & ~w2508;
assign w2510 = ~w50 & ~w342;
assign w2511 = w303 & w6935;
assign w2512 = ~w1071 & ~w2511;
assign w2513 = w1086 & ~w2512;
assign w2514 = w39 & w6936;
assign w2515 = w39 & w6937;
assign w2516 = pi08 & w80;
assign w2517 = pi06 & w82;
assign w2518 = w36 & w6938;
assign w2519 = pi05 & w110;
assign w2520 = pi04 & w143;
assign w2521 = w30 & w6939;
assign w2522 = pi09 & pi19;
assign w2523 = ~w2516 & ~w2522;
assign w2524 = ~w2517 & w2523;
assign w2525 = ~w2521 & w2524;
assign w2526 = ~w96 & ~w2518;
assign w2527 = ~w2519 & w2526;
assign w2528 = ~w2520 & w2525;
assign w2529 = w2527 & w2528;
assign w2530 = ~w2514 & ~w2515;
assign w2531 = (w2530 & w2529) | (w2530 & w6940) | (w2529 & w6940);
assign w2532 = w2513 & ~w2531;
assign w2533 = ~w1556 & ~w2531;
assign w2534 = w1774 & ~w2531;
assign w2535 = w1563 & ~w2531;
assign w2536 = w1566 & ~w2531;
assign w2537 = w1570 & ~w2531;
assign w2538 = w1572 & ~w2531;
assign w2539 = ~w1648 & ~w2531;
assign w2540 = ~w1531 & w6941;
assign w2541 = ~w1501 & w2540;
assign w2542 = (~w2531 & w1531) | (~w2531 & w6942) | (w1531 & w6942);
assign w2543 = w1501 & w2542;
assign w2544 = ~w2541 & ~w2543;
assign w2545 = ~w2414 & ~w2531;
assign w2546 = ~w1584 & w2545;
assign w2547 = w1581 & w6422;
assign w2548 = ~w364 & ~w1509;
assign w2549 = ~w1581 & w2548;
assign w2550 = ~w2184 & ~w2549;
assign w2551 = ~w2547 & w2550;
assign w2552 = ~w2419 & ~w2551;
assign w2553 = ~w2546 & ~w2552;
assign w2554 = ~w1584 & w6943;
assign w2555 = ~w1523 & ~w2531;
assign w2556 = w1520 & w2555;
assign w2557 = w1523 & ~w2531;
assign w2558 = ~w1520 & w2557;
assign w2559 = ~w2556 & ~w2558;
assign w2560 = ~w2554 & w2559;
assign w2561 = ~w2553 & ~w2560;
assign w2562 = ~w2409 & ~w2420;
assign w2563 = w2425 & ~w2562;
assign w2564 = ~w2425 & w2562;
assign w2565 = ~w2563 & ~w2564;
assign w2566 = w2561 & w2565;
assign w2567 = ~w1590 & ~w2566;
assign w2568 = ~w2561 & ~w2565;
assign w2569 = (~w2531 & w2565) | (~w2531 & w6423) | (w2565 & w6423);
assign w2570 = ~w2567 & w2569;
assign w2571 = ~w2544 & w2570;
assign w2572 = w2544 & ~w2570;
assign w2573 = ~w364 & w1590;
assign w2574 = ~w2431 & ~w2433;
assign w2575 = ~w2573 & w2574;
assign w2576 = w2573 & ~w2574;
assign w2577 = ~w2575 & ~w2576;
assign w2578 = ~w2572 & ~w2577;
assign w2579 = (w2539 & w2578) | (w2539 & w6424) | (w2578 & w6424);
assign w2580 = ~w2578 & w6425;
assign w2581 = ~w2441 & ~w2442;
assign w2582 = w2447 & w2581;
assign w2583 = ~w2447 & ~w2581;
assign w2584 = ~w2582 & ~w2583;
assign w2585 = ~w2580 & ~w2584;
assign w2586 = (w2538 & w2585) | (w2538 & w6160) | (w2585 & w6160);
assign w2587 = ~w2585 & w6161;
assign w2588 = ~w2449 & ~w2450;
assign w2589 = w2452 & w2588;
assign w2590 = ~w2452 & ~w2588;
assign w2591 = ~w2589 & ~w2590;
assign w2592 = w2537 & w7483;
assign w2593 = ~w2586 & w7484;
assign w2594 = ~w2592 & ~w2593;
assign w2595 = ~w2455 & ~w2456;
assign w2596 = ~w2458 & w2595;
assign w2597 = w2458 & ~w2595;
assign w2598 = ~w2596 & ~w2597;
assign w2599 = w2594 & w2598;
assign w2600 = w1568 & ~w2531;
assign w2601 = ~w2592 & ~w2600;
assign w2602 = ~w2599 & w2601;
assign w2603 = w1568 & w2592;
assign w2604 = ~w2593 & w2600;
assign w2605 = w2598 & w2604;
assign w2606 = ~w2603 & ~w2605;
assign w2607 = ~w2460 & ~w2461;
assign w2608 = ~w2463 & w2607;
assign w2609 = w2463 & ~w2607;
assign w2610 = ~w2608 & ~w2609;
assign w2611 = (~w2602 & w2610) | (~w2602 & w6945) | (w2610 & w6945);
assign w2612 = w2536 & w2611;
assign w2613 = ~w2464 & ~w2465;
assign w2614 = ~w2467 & w2613;
assign w2615 = w2467 & ~w2613;
assign w2616 = ~w2614 & ~w2615;
assign w2617 = ~w2612 & w2616;
assign w2618 = ~w2536 & ~w2611;
assign w2619 = ~w2617 & w6946;
assign w2620 = (~w2535 & w2617) | (~w2535 & w2634) | (w2617 & w2634);
assign w2621 = ~w2469 & ~w2470;
assign w2622 = ~w2472 & w2621;
assign w2623 = w2472 & ~w2621;
assign w2624 = ~w2622 & ~w2623;
assign w2625 = ~w2620 & ~w2624;
assign w2626 = w1561 & ~w2531;
assign w2627 = ~w2619 & ~w2626;
assign w2628 = ~w2625 & w2627;
assign w2629 = w2476 & ~w2478;
assign w2630 = ~w2479 & ~w2629;
assign w2631 = ~w2619 & ~w2620;
assign w2632 = w2624 & w2631;
assign w2633 = (~w1988 & w2617) | (~w1988 & w6947) | (w2617 & w6947);
assign w2634 = ~w2535 & w2618;
assign w2635 = ~w2633 & ~w2634;
assign w2636 = ~w2632 & w2635;
assign w2637 = ~w2628 & ~w2636;
assign w2638 = w2630 & w2637;
assign w2639 = (~w2628 & ~w2630) | (~w2628 & w6948) | (~w2630 & w6948);
assign w2640 = w2534 & w2639;
assign w2641 = ~w2483 & w2485;
assign w2642 = ~w2486 & ~w2641;
assign w2643 = ~w2534 & ~w2639;
assign w2644 = ~w2640 & ~w2643;
assign w2645 = ~w2642 & w2644;
assign w2646 = (w2533 & w2645) | (w2533 & w6949) | (w2645 & w6949);
assign w2647 = w2489 & ~w2493;
assign w2648 = ~w2494 & ~w2647;
assign w2649 = ~w2645 & w6950;
assign w2650 = ~w2646 & ~w2649;
assign w2651 = ~w2648 & w2650;
assign w2652 = (w2498 & ~w2500) | (w2498 & w6951) | (~w2500 & w6951);
assign w2653 = ~w2501 & ~w2652;
assign w2654 = ~w1086 & ~w2531;
assign w2655 = ~w2651 & w6952;
assign w2656 = ~w2653 & w2655;
assign w2657 = ~w2651 & w6953;
assign w2658 = ~w2656 & w2657;
assign w2659 = w2509 & w2658;
assign w2660 = ~w2509 & ~w2658;
assign w2661 = ~w2659 & ~w2660;
assign w2662 = w2653 & ~w2655;
assign w2663 = ~w2656 & ~w2662;
assign w2664 = w39 & w6954;
assign w2665 = w36 & w6955;
assign w2666 = pi07 & w80;
assign w2667 = w30 & w6956;
assign w2668 = pi08 & pi19;
assign w2669 = pi03 & w143;
assign w2670 = pi02 & w26;
assign w2671 = pi05 & w82;
assign w2672 = ~w2666 & ~w2668;
assign w2673 = ~w2667 & w2672;
assign w2674 = ~w2671 & w2673;
assign w2675 = ~w98 & ~w2665;
assign w2676 = w2674 & w2675;
assign w2677 = ~w2669 & ~w2670;
assign w2678 = (~w10 & ~w2676) | (~w10 & w6957) | (~w2676 & w6957);
assign w2679 = ~w2664 & ~w2678;
assign w2680 = w1086 & w6958;
assign w2681 = ~w1556 & ~w2679;
assign w2682 = ~w2624 & ~w2631;
assign w2683 = ~w2632 & ~w2682;
assign w2684 = w1774 & ~w2679;
assign w2685 = w1566 & ~w2679;
assign w2686 = ~w1576 & ~w2679;
assign w2687 = w1509 & ~w2679;
assign w2688 = w1581 & w2687;
assign w2689 = ~w1509 & ~w2679;
assign w2690 = ~w1581 & w2689;
assign w2691 = ~w2688 & ~w2690;
assign w2692 = w1012 & ~w2531;
assign w2693 = w1012 & w6959;
assign w2694 = ~w2691 & w2693;
assign w2695 = ~w1581 & w6960;
assign w2696 = w1509 & ~w2531;
assign w2697 = w1581 & w2696;
assign w2698 = w2414 & ~w2697;
assign w2699 = ~w2695 & w2698;
assign w2700 = ~w2694 & ~w2699;
assign w2701 = ~w1523 & ~w2679;
assign w2702 = w1520 & w2701;
assign w2703 = w1523 & ~w2679;
assign w2704 = ~w1520 & w2703;
assign w2705 = ~w2702 & ~w2704;
assign w2706 = w2700 & ~w2705;
assign w2707 = (~w2694 & w2705) | (~w2694 & w6163) | (w2705 & w6163);
assign w2708 = w1590 & ~w2707;
assign w2709 = ~w1590 & w2707;
assign w2710 = (~w2554 & w2552) | (~w2554 & w6961) | (w2552 & w6961);
assign w2711 = ~w2531 & ~w2705;
assign w2712 = ~w2710 & w2711;
assign w2713 = ~w2553 & w2560;
assign w2714 = w2560 & w6164;
assign w2715 = ~w2712 & ~w2714;
assign w2716 = ~w2709 & ~w2715;
assign w2717 = ~w2708 & ~w2716;
assign w2718 = ~w2686 & w2717;
assign w2719 = w1590 & ~w2531;
assign w2720 = ~w2566 & ~w2568;
assign w2721 = w2719 & w2720;
assign w2722 = ~w2719 & ~w2720;
assign w2723 = ~w2721 & ~w2722;
assign w2724 = ~w2718 & w2723;
assign w2725 = w2686 & ~w2717;
assign w2726 = ~w2679 & ~w1645;
assign w2727 = w1644 & w2726;
assign w2728 = ~w1481 & w7485;
assign w2729 = ~w1644 & w2728;
assign w2730 = ~w2727 & ~w2729;
assign w2731 = ~w2725 & w2730;
assign w2732 = ~w2724 & w2731;
assign w2733 = ~w2571 & ~w2572;
assign w2734 = ~w2577 & w2733;
assign w2735 = w2577 & ~w2733;
assign w2736 = ~w2734 & ~w2735;
assign w2737 = ~w2732 & w2736;
assign w2738 = (~w2679 & w1535) | (~w2679 & w6963) | (w1535 & w6963);
assign w2739 = ~w1539 & w2738;
assign w2740 = ~w1535 & w6964;
assign w2741 = w1539 & w2740;
assign w2742 = ~w2739 & ~w2741;
assign w2743 = ~w2723 & ~w2725;
assign w2744 = ~w2718 & ~w2730;
assign w2745 = ~w2743 & w2744;
assign w2746 = w2742 & ~w2745;
assign w2747 = ~w2737 & w2746;
assign w2748 = ~w2579 & ~w2580;
assign w2749 = ~w2584 & w2748;
assign w2750 = w2584 & ~w2748;
assign w2751 = ~w2749 & ~w2750;
assign w2752 = ~w2747 & w2751;
assign w2753 = (~w2745 & ~w2736) | (~w2745 & w6165) | (~w2736 & w6165);
assign w2754 = ~w2742 & ~w2753;
assign w2755 = ~w1540 & ~w2679;
assign w2756 = w1542 & w2755;
assign w2757 = w1540 & ~w2679;
assign w2758 = ~w1542 & w2757;
assign w2759 = ~w2756 & ~w2758;
assign w2760 = ~w2754 & w2759;
assign w2761 = ~w2752 & w2760;
assign w2762 = w2754 & ~w2759;
assign w2763 = (~w2759 & w2737) | (~w2759 & w6426) | (w2737 & w6426);
assign w2764 = w2751 & w2763;
assign w2765 = ~w2762 & ~w2764;
assign w2766 = ~w2761 & w2765;
assign w2767 = ~w2586 & ~w2587;
assign w2768 = ~w2591 & w2767;
assign w2769 = w2591 & ~w2767;
assign w2770 = ~w2768 & ~w2769;
assign w2771 = w2766 & ~w2770;
assign w2772 = w1568 & ~w2679;
assign w2773 = ~w2761 & w2772;
assign w2774 = (w2773 & ~w2766) | (w2773 & w6965) | (~w2766 & w6965);
assign w2775 = w2685 & w2774;
assign w2776 = ~w2594 & ~w2598;
assign w2777 = ~w2599 & ~w2776;
assign w2778 = w2761 & ~w2772;
assign w2779 = ~w2764 & w6966;
assign w2780 = ~w2770 & w2779;
assign w2781 = ~w2778 & ~w2780;
assign w2782 = ~w2780 & w6166;
assign w2783 = w2777 & w2782;
assign w2784 = ~w2775 & ~w2783;
assign w2785 = ~w2602 & w2606;
assign w2786 = w2610 & ~w2785;
assign w2787 = ~w2610 & w2785;
assign w2788 = ~w2786 & ~w2787;
assign w2789 = w2784 & w2788;
assign w2790 = w1563 & ~w2679;
assign w2791 = ~w2774 & w2781;
assign w2792 = w2777 & w2791;
assign w2793 = ~w2685 & ~w2774;
assign w2794 = ~w2792 & w2793;
assign w2795 = (w2790 & w2792) | (w2790 & w6967) | (w2792 & w6967);
assign w2796 = ~w2789 & w2795;
assign w2797 = ~w2792 & w6968;
assign w2798 = w2784 & ~w2790;
assign w2799 = w2788 & w2798;
assign w2800 = ~w2797 & ~w2799;
assign w2801 = ~w2796 & w2800;
assign w2802 = ~w2612 & ~w2618;
assign w2803 = ~w2616 & w2802;
assign w2804 = w2616 & ~w2802;
assign w2805 = ~w2803 & ~w2804;
assign w2806 = w2801 & w2805;
assign w2807 = w1561 & ~w2679;
assign w2808 = (~w2807 & w2789) | (~w2807 & w6969) | (w2789 & w6969);
assign w2809 = ~w2806 & w2808;
assign w2810 = (w2684 & w2806) | (w2684 & w6970) | (w2806 & w6970);
assign w2811 = ~w2683 & w2810;
assign w2812 = ~w2799 & w6971;
assign w2813 = (w2812 & w2805) | (w2812 & w6972) | (w2805 & w6972);
assign w2814 = ~w1192 & w2813;
assign w2815 = ~w2811 & ~w2814;
assign w2816 = ~w2809 & ~w2813;
assign w2817 = ~w2683 & w2816;
assign w2818 = ~w2684 & ~w2813;
assign w2819 = (w2818 & ~w2816) | (w2818 & w6973) | (~w2816 & w6973);
assign w2820 = w2815 & ~w2819;
assign w2821 = ~w2630 & ~w2637;
assign w2822 = ~w2638 & ~w2821;
assign w2823 = w2820 & ~w2822;
assign w2824 = (w2815 & w2822) | (w2815 & w6974) | (w2822 & w6974);
assign w2825 = ~w2681 & w2824;
assign w2826 = w2642 & ~w2644;
assign w2827 = ~w2645 & ~w2826;
assign w2828 = w2681 & ~w2824;
assign w2829 = ~w2825 & ~w2828;
assign w2830 = ~w2827 & w2829;
assign w2831 = w2648 & ~w2650;
assign w2832 = ~w2651 & ~w2831;
assign w2833 = ~w1086 & ~w2679;
assign w2834 = (w2833 & w2830) | (w2833 & w6975) | (w2830 & w6975);
assign w2835 = w2832 & w2834;
assign w2836 = (~w2680 & w2830) | (~w2680 & w6976) | (w2830 & w6976);
assign w2837 = ~w2835 & w2836;
assign w2838 = w2663 & ~w2837;
assign w2839 = ~w2832 & ~w2834;
assign w2840 = ~w2835 & ~w2839;
assign w2841 = pi02 & w143;
assign w2842 = pi07 & pi19;
assign w2843 = w30 & w6977;
assign w2844 = pi06 & w80;
assign w2845 = pi04 & w82;
assign w2846 = w36 & w6978;
assign w2847 = pi01 & w26;
assign w2848 = ~w2842 & ~w2844;
assign w2849 = ~w2843 & w2848;
assign w2850 = ~w2845 & w2849;
assign w2851 = ~w161 & ~w2846;
assign w2852 = w2850 & w2851;
assign w2853 = ~w2841 & ~w2847;
assign w2854 = (~w10 & ~w2852) | (~w10 & w6979) | (~w2852 & w6979);
assign w2855 = w2513 & w2854;
assign w2856 = ~w2820 & w2822;
assign w2857 = ~w2823 & ~w2856;
assign w2858 = w1566 & w2854;
assign w2859 = w1570 & w2854;
assign w2860 = ~w2732 & ~w2745;
assign w2861 = ~w1535 & w6980;
assign w2862 = w1539 & w2861;
assign w2863 = (w2854 & w1535) | (w2854 & w6981) | (w1535 & w6981);
assign w2864 = ~w1539 & w2863;
assign w2865 = ~w2862 & ~w2864;
assign w2866 = ~w2736 & ~w2865;
assign w2867 = w2860 & w2866;
assign w2868 = w2736 & ~w2865;
assign w2869 = ~w2860 & w2868;
assign w2870 = ~w2867 & ~w2869;
assign w2871 = ~w1648 & w2854;
assign w2872 = w1012 & w2854;
assign w2873 = ~w2691 & w2872;
assign w2874 = ~w2691 & w6982;
assign w2875 = w2691 & ~w2692;
assign w2876 = ~w1523 & w2854;
assign w2877 = w1520 & w2876;
assign w2878 = w1523 & w2854;
assign w2879 = ~w1520 & w2878;
assign w2880 = ~w2877 & ~w2879;
assign w2881 = ~w2875 & ~w2880;
assign w2882 = (~w2874 & w2880) | (~w2874 & w6983) | (w2880 & w6983);
assign w2883 = ~w1584 & w6984;
assign w2884 = w2700 & ~w2883;
assign w2885 = w2705 & ~w2884;
assign w2886 = ~w2706 & ~w2885;
assign w2887 = ~w2882 & w2886;
assign w2888 = ~w1590 & ~w2887;
assign w2889 = w2882 & ~w2886;
assign w2890 = (w2854 & w2886) | (w2854 & w6985) | (w2886 & w6985);
assign w2891 = ~w2888 & w2890;
assign w2892 = ~w1576 & w2891;
assign w2893 = ~w1576 & w2854;
assign w2894 = ~w2891 & ~w2893;
assign w2895 = ~w2559 & ~w2710;
assign w2896 = ~w2713 & ~w2895;
assign w2897 = ~w2679 & w2707;
assign w2898 = w1590 & ~w2897;
assign w2899 = ~w2709 & ~w2898;
assign w2900 = ~w2896 & w2899;
assign w2901 = w2896 & ~w2899;
assign w2902 = ~w2900 & ~w2901;
assign w2903 = ~w2894 & w2902;
assign w2904 = (w2871 & w2903) | (w2871 & w6986) | (w2903 & w6986);
assign w2905 = ~w2903 & w6987;
assign w2906 = ~w2718 & ~w2725;
assign w2907 = ~w2723 & w2906;
assign w2908 = w2723 & ~w2906;
assign w2909 = ~w2907 & ~w2908;
assign w2910 = (~w2904 & w2909) | (~w2904 & w6988) | (w2909 & w6988);
assign w2911 = w2870 & w2910;
assign w2912 = ~w2736 & w2865;
assign w2913 = ~w2860 & w2912;
assign w2914 = ~w2745 & w2865;
assign w2915 = w2737 & w2914;
assign w2916 = ~w2913 & ~w2915;
assign w2917 = (~w2859 & w2911) | (~w2859 & w6167) | (w2911 & w6167);
assign w2918 = w2859 & w2916;
assign w2919 = ~w2911 & w2918;
assign w2920 = ~w2917 & ~w2919;
assign w2921 = ~w2747 & ~w2754;
assign w2922 = ~w2751 & w2921;
assign w2923 = w2751 & ~w2921;
assign w2924 = ~w2922 & ~w2923;
assign w2925 = w2920 & w2924;
assign w2926 = w1568 & w2854;
assign w2927 = ~w2917 & w2926;
assign w2928 = ~w2925 & w2927;
assign w2929 = w2917 & ~w2926;
assign w2930 = ~w2919 & ~w2926;
assign w2931 = w2924 & w2930;
assign w2932 = ~w2929 & ~w2931;
assign w2933 = ~w2766 & w2770;
assign w2934 = ~w2771 & ~w2933;
assign w2935 = w2932 & ~w2934;
assign w2936 = (w2858 & w2935) | (w2858 & w6168) | (w2935 & w6168);
assign w2937 = ~w2935 & w6169;
assign w2938 = ~w2936 & ~w2937;
assign w2939 = ~w2777 & ~w2791;
assign w2940 = ~w2792 & ~w2939;
assign w2941 = (~w2936 & ~w2938) | (~w2936 & w6989) | (~w2938 & w6989);
assign w2942 = w2784 & ~w2794;
assign w2943 = w1563 & w2854;
assign w2944 = ~w2610 & w2943;
assign w2945 = w2785 & ~w2944;
assign w2946 = w2610 & w2943;
assign w2947 = ~w2785 & ~w2946;
assign w2948 = ~w2945 & ~w2947;
assign w2949 = ~w2942 & w2948;
assign w2950 = w2785 & ~w2946;
assign w2951 = ~w2785 & ~w2944;
assign w2952 = ~w2950 & ~w2951;
assign w2953 = w2942 & w2952;
assign w2954 = ~w2949 & ~w2953;
assign w2955 = w2941 & w2954;
assign w2956 = w1561 & w2610;
assign w2957 = w2785 & ~w2956;
assign w2958 = w1561 & ~w2610;
assign w2959 = ~w2785 & ~w2958;
assign w2960 = ~w2957 & ~w2959;
assign w2961 = w1561 & ~w2788;
assign w2962 = ~w2942 & w2961;
assign w2963 = (~w1988 & ~w2942) | (~w1988 & w6170) | (~w2942 & w6170);
assign w2964 = ~w2962 & w2963;
assign w2965 = ~w2955 & ~w2964;
assign w2966 = w1774 & w2854;
assign w2967 = w2965 & w2966;
assign w2968 = ~w2801 & ~w2805;
assign w2969 = ~w2806 & ~w2968;
assign w2970 = w2610 & ~w2943;
assign w2971 = w2785 & ~w2970;
assign w2972 = ~w2610 & ~w2943;
assign w2973 = ~w2785 & ~w2972;
assign w2974 = ~w2971 & ~w2973;
assign w2975 = ~w2942 & w2974;
assign w2976 = w2785 & ~w2972;
assign w2977 = ~w2785 & ~w2970;
assign w2978 = ~w2976 & ~w2977;
assign w2979 = w2942 & w2978;
assign w2980 = ~w2975 & ~w2979;
assign w2981 = ~w2941 & w2980;
assign w2982 = w1561 & w2854;
assign w2983 = w2954 & ~w2982;
assign w2984 = ~w2981 & w2983;
assign w2985 = w2966 & ~w2984;
assign w2986 = w2969 & w2985;
assign w2987 = ~w2967 & ~w2986;
assign w2988 = ~w2965 & ~w2984;
assign w2989 = w2969 & w2988;
assign w2990 = ~w2965 & ~w2966;
assign w2991 = ~w2989 & w2990;
assign w2992 = w2987 & ~w2991;
assign w2993 = w2683 & ~w2816;
assign w2994 = ~w2817 & ~w2993;
assign w2995 = w2992 & w2994;
assign w2996 = ~w1556 & w2854;
assign w2997 = ~w2986 & w6171;
assign w2998 = (w2996 & w2986) | (w2996 & w6172) | (w2986 & w6172);
assign w2999 = ~w2997 & ~w2998;
assign w3000 = ~w2995 & w2999;
assign w3001 = w2992 & w6173;
assign w3002 = ~w3000 & ~w3001;
assign w3003 = w2857 & ~w3002;
assign w3004 = (w2996 & w2995) | (w2996 & w6990) | (w2995 & w6990);
assign w3005 = (~w3004 & w3002) | (~w3004 & w6991) | (w3002 & w6991);
assign w3006 = w2827 & ~w2829;
assign w3007 = ~w2830 & ~w3006;
assign w3008 = ~w1086 & w2854;
assign w3009 = w3005 & w3008;
assign w3010 = ~w3007 & w3009;
assign w3011 = ~w2855 & w3005;
assign w3012 = ~w3010 & w3011;
assign w3013 = w2840 & ~w3012;
assign w3014 = ~w2840 & w3012;
assign w3015 = ~w3013 & ~w3014;
assign w3016 = w3007 & ~w3009;
assign w3017 = ~w3010 & ~w3016;
assign w3018 = w30 & w6992;
assign w3019 = pi00 & w26;
assign w3020 = pi05 & w80;
assign w3021 = pi06 & pi19;
assign w3022 = pi03 & w82;
assign w3023 = w36 & w6993;
assign w3024 = pi01 & w143;
assign w3025 = ~w3020 & ~w3021;
assign w3026 = ~w3022 & w3025;
assign w3027 = ~w3023 & w3026;
assign w3028 = w3027 & w6994;
assign w3029 = ~w3018 & w3028;
assign w3030 = w1774 & ~w3029;
assign w3031 = w1566 & ~w3029;
assign w3032 = ~w2920 & ~w2924;
assign w3033 = ~w2925 & ~w3032;
assign w3034 = w2870 & w2916;
assign w3035 = ~w2910 & w3034;
assign w3036 = w2910 & ~w3034;
assign w3037 = ~w3035 & ~w3036;
assign w3038 = ~w2904 & ~w2905;
assign w3039 = ~w2909 & w3038;
assign w3040 = w2909 & ~w3038;
assign w3041 = ~w3039 & ~w3040;
assign w3042 = ~w1576 & ~w3029;
assign w3043 = ~w2692 & ~w2872;
assign w3044 = ~w2691 & ~w3043;
assign w3045 = ~w2875 & ~w3044;
assign w3046 = w2880 & ~w3045;
assign w3047 = ~w2881 & ~w3046;
assign w3048 = ~w2691 & w6995;
assign w3049 = w1579 & ~w3048;
assign w3050 = ~w1579 & ~w2874;
assign w3051 = ~w3049 & ~w3050;
assign w3052 = ~w3047 & ~w3051;
assign w3053 = w1590 & ~w3052;
assign w3054 = ~w3052 & w6174;
assign w3055 = ~w1590 & w3052;
assign w3056 = ~w1584 & w6996;
assign w3057 = w2679 & w3056;
assign w3058 = w1012 & ~w2679;
assign w3059 = (~w3058 & w1584) | (~w3058 & w6997) | (w1584 & w6997);
assign w3060 = ~w2873 & ~w3059;
assign w3061 = ~w3056 & ~w3060;
assign w3062 = ~w1579 & ~w3029;
assign w3063 = (~w3057 & ~w3062) | (~w3057 & w6998) | (~w3062 & w6998);
assign w3064 = (~w3063 & ~w3052) | (~w3063 & w7438) | (~w3052 & w7438);
assign w3065 = ~w3054 & ~w3064;
assign w3066 = ~w3042 & w3065;
assign w3067 = w1590 & w2854;
assign w3068 = ~w2887 & ~w2889;
assign w3069 = w3067 & ~w3068;
assign w3070 = ~w3067 & w3068;
assign w3071 = ~w3069 & ~w3070;
assign w3072 = ~w3066 & ~w3071;
assign w3073 = w3042 & ~w3065;
assign w3074 = ~w3029 & ~w1645;
assign w3075 = w1644 & w3074;
assign w3076 = ~w1481 & w7486;
assign w3077 = ~w1644 & w3076;
assign w3078 = ~w3075 & ~w3077;
assign w3079 = (w3078 & w3065) | (w3078 & w7000) | (w3065 & w7000);
assign w3080 = ~w3072 & w3079;
assign w3081 = w3071 & ~w3073;
assign w3082 = (~w3078 & ~w3065) | (~w3078 & w7001) | (~w3065 & w7001);
assign w3083 = ~w3081 & w3082;
assign w3084 = ~w3080 & ~w3083;
assign w3085 = ~w2892 & ~w2894;
assign w3086 = w2902 & w3085;
assign w3087 = ~w2902 & ~w3085;
assign w3088 = ~w3086 & ~w3087;
assign w3089 = w3084 & ~w3088;
assign w3090 = (~w3029 & w1535) | (~w3029 & w7002) | (w1535 & w7002);
assign w3091 = ~w1539 & w3090;
assign w3092 = ~w1535 & w7003;
assign w3093 = w1539 & w3092;
assign w3094 = ~w3091 & ~w3093;
assign w3095 = (~w3094 & w3072) | (~w3094 & w7004) | (w3072 & w7004);
assign w3096 = ~w3072 & w7005;
assign w3097 = ~w3095 & ~w3096;
assign w3098 = ~w3089 & ~w3097;
assign w3099 = w3084 & w6175;
assign w3100 = ~w3098 & w7006;
assign w3101 = (w3095 & ~w3084) | (w3095 & w7007) | (~w3084 & w7007);
assign w3102 = ~w3089 & w6176;
assign w3103 = w1570 & ~w3029;
assign w3104 = ~w3101 & w3103;
assign w3105 = ~w3102 & ~w3104;
assign w3106 = w3100 & ~w3105;
assign w3107 = ~w3100 & w3105;
assign w3108 = ~w3106 & ~w3107;
assign w3109 = w3037 & w3108;
assign w3110 = w3103 & ~w3108;
assign w3111 = ~w3109 & ~w3110;
assign w3112 = (w3031 & ~w3111) | (w3031 & w6177) | (~w3111 & w6177);
assign w3113 = ~w1568 & w3031;
assign w3114 = (w3113 & w3111) | (w3113 & w6178) | (w3111 & w6178);
assign w3115 = w3112 & ~w3114;
assign w3116 = (~w3031 & w3111) | (~w3031 & w6179) | (w3111 & w6179);
assign w3117 = ~w3112 & ~w3116;
assign w3118 = w1568 & ~w3029;
assign w3119 = ~w1566 & w3118;
assign w3120 = (w3119 & ~w3111) | (w3119 & w6180) | (~w3111 & w6180);
assign w3121 = ~w3114 & ~w3120;
assign w3122 = ~w3117 & w3121;
assign w3123 = ~w2928 & w2932;
assign w3124 = w2934 & ~w3123;
assign w3125 = ~w2934 & w3123;
assign w3126 = ~w3124 & ~w3125;
assign w3127 = ~w3122 & w3126;
assign w3128 = (~w3115 & w3122) | (~w3115 & w7008) | (w3122 & w7008);
assign w3129 = w1563 & ~w3029;
assign w3130 = w2940 & ~w3129;
assign w3131 = w2938 & w3130;
assign w3132 = ~w2940 & ~w3129;
assign w3133 = ~w2938 & w3132;
assign w3134 = ~w3131 & ~w3133;
assign w3135 = ~w3128 & w3134;
assign w3136 = w1561 & ~w3029;
assign w3137 = ~w2938 & ~w2940;
assign w3138 = (w3129 & ~w2938) | (w3129 & w6427) | (~w2938 & w6427);
assign w3139 = ~w3137 & w3138;
assign w3140 = ~w3136 & ~w3139;
assign w3141 = ~w3135 & w3140;
assign w3142 = w2954 & w2980;
assign w3143 = w2941 & ~w3142;
assign w3144 = ~w2941 & w3142;
assign w3145 = ~w3143 & ~w3144;
assign w3146 = ~w3141 & w3145;
assign w3147 = w3134 & w3136;
assign w3148 = ~w3128 & w3147;
assign w3149 = w1561 & w3139;
assign w3150 = ~w3148 & ~w3149;
assign w3151 = (w3030 & w3146) | (w3030 & w6181) | (w3146 & w6181);
assign w3152 = w1553 & w3151;
assign w3153 = ~w3148 & w6182;
assign w3154 = ~w3146 & w3153;
assign w3155 = ~w2969 & ~w2988;
assign w3156 = ~w2989 & ~w3155;
assign w3157 = ~w3154 & w3156;
assign w3158 = ~w1556 & ~w3029;
assign w3159 = w3157 & w3158;
assign w3160 = ~w3152 & ~w3159;
assign w3161 = w1086 & w7009;
assign w3162 = ~w1086 & ~w3029;
assign w3163 = ~w3151 & ~w3158;
assign w3164 = ~w3157 & w3163;
assign w3165 = w3162 & w3164;
assign w3166 = ~w2624 & w3162;
assign w3167 = ~w2631 & ~w3166;
assign w3168 = w2624 & w3162;
assign w3169 = w2631 & ~w3168;
assign w3170 = ~w3167 & ~w3169;
assign w3171 = w2816 & w3170;
assign w3172 = ~w2631 & w3168;
assign w3173 = w2631 & w3166;
assign w3174 = ~w3172 & ~w3173;
assign w3175 = ~w2816 & ~w3174;
assign w3176 = ~w3171 & ~w3175;
assign w3177 = ~w2992 & ~w3176;
assign w3178 = ~w2816 & ~w3170;
assign w3179 = w2816 & w3174;
assign w3180 = ~w3178 & ~w3179;
assign w3181 = w2992 & w3180;
assign w3182 = ~w3177 & ~w3181;
assign w3183 = w3160 & ~w3182;
assign w3184 = ~w3165 & ~w3183;
assign w3185 = ~w2857 & w3002;
assign w3186 = ~w3003 & ~w3185;
assign w3187 = ~w3184 & w3186;
assign w3188 = w3160 & ~w3164;
assign w3189 = ~w2992 & ~w2994;
assign w3190 = ~w2995 & ~w3189;
assign w3191 = w3188 & w3190;
assign w3192 = ~w3159 & w7010;
assign w3193 = (w3192 & ~w3188) | (w3192 & w7011) | (~w3188 & w7011);
assign w3194 = (w3193 & ~w3186) | (w3193 & w7012) | (~w3186 & w7012);
assign w3195 = w3017 & ~w3194;
assign w3196 = ~w3017 & w3194;
assign w3197 = ~w3195 & ~w3196;
assign w3198 = pi03 & w80;
assign w3199 = w36 & w7013;
assign w3200 = w30 & w7014;
assign w3201 = pi04 & pi19;
assign w3202 = pi01 & w82;
assign w3203 = ~w3198 & ~w3201;
assign w3204 = ~w3200 & w3203;
assign w3205 = w3204 & w7015;
assign w3206 = w2513 & ~w3205;
assign w3207 = ~w1086 & ~w3205;
assign w3208 = ~w3141 & w3150;
assign w3209 = w3145 & w3208;
assign w3210 = ~w3145 & ~w3208;
assign w3211 = ~w3209 & ~w3210;
assign w3212 = pi04 & w80;
assign w3213 = w30 & w7016;
assign w3214 = pi05 & pi19;
assign w3215 = pi02 & w82;
assign w3216 = w36 & w7017;
assign w3217 = pi00 & w143;
assign w3218 = ~w3213 & ~w3214;
assign w3219 = ~w3215 & w3218;
assign w3220 = ~w3216 & w3219;
assign w3221 = ~w3217 & w3220;
assign w3222 = w3220 & w7018;
assign w3223 = w1561 & ~w3222;
assign w3224 = w1563 & ~w3222;
assign w3225 = w1570 & ~w3222;
assign w3226 = w1572 & ~w3222;
assign w3227 = (~w2872 & w1584) | (~w2872 & w7019) | (w1584 & w7019);
assign w3228 = ~w3056 & ~w3227;
assign w3229 = ~w1584 & w7020;
assign w3230 = ~w1579 & w3229;
assign w3231 = (~w3228 & w1579) | (~w3228 & w7021) | (w1579 & w7021);
assign w3232 = (~w3222 & ~w1579) | (~w3222 & w7022) | (~w1579 & w7022);
assign w3233 = ~w3231 & w3232;
assign w3234 = w1530 & ~w3222;
assign w3235 = w1587 & ~w3234;
assign w3236 = ~w1530 & ~w3222;
assign w3237 = ~w1587 & ~w3236;
assign w3238 = ~w3235 & ~w3237;
assign w3239 = w3233 & w3238;
assign w3240 = ~w3233 & ~w3238;
assign w3241 = ~w3239 & ~w3240;
assign w3242 = ~w3057 & ~w3061;
assign w3243 = w3062 & ~w3242;
assign w3244 = ~w3062 & w3242;
assign w3245 = ~w3243 & ~w3244;
assign w3246 = w3241 & ~w3245;
assign w3247 = (~w3239 & ~w3241) | (~w3239 & w7023) | (~w3241 & w7023);
assign w3248 = ~w3053 & ~w3055;
assign w3249 = w1590 & w3029;
assign w3250 = w3063 & ~w3249;
assign w3251 = w3248 & ~w3250;
assign w3252 = ~w3248 & w3250;
assign w3253 = ~w3251 & ~w3252;
assign w3254 = ~w3247 & w3253;
assign w3255 = ~w1576 & ~w3222;
assign w3256 = (~w3255 & ~w3253) | (~w3255 & w6183) | (~w3253 & w6183);
assign w3257 = ~w1648 & ~w3222;
assign w3258 = w3247 & ~w3253;
assign w3259 = (w3257 & w3253) | (w3257 & w7024) | (w3253 & w7024);
assign w3260 = ~w3256 & w3259;
assign w3261 = ~w3066 & ~w3073;
assign w3262 = ~w3071 & w3261;
assign w3263 = w3071 & ~w3261;
assign w3264 = ~w3262 & ~w3263;
assign w3265 = ~w3260 & ~w3264;
assign w3266 = (w3255 & w3253) | (w3255 & w6184) | (w3253 & w6184);
assign w3267 = (~w3257 & ~w3253) | (~w3257 & w7025) | (~w3253 & w7025);
assign w3268 = ~w3266 & w3267;
assign w3269 = (~w3226 & w3265) | (~w3226 & w6185) | (w3265 & w6185);
assign w3270 = w1572 & ~w3268;
assign w3271 = ~w3265 & w3270;
assign w3272 = ~w3084 & w3088;
assign w3273 = ~w3089 & ~w3272;
assign w3274 = ~w3271 & w3273;
assign w3275 = ~w3274 & w6186;
assign w3276 = (~w3041 & w3098) | (~w3041 & w7026) | (w3098 & w7026);
assign w3277 = ~w3100 & ~w3276;
assign w3278 = ~w3275 & ~w3277;
assign w3279 = (~w3225 & w3274) | (~w3225 & w6187) | (w3274 & w6187);
assign w3280 = w1568 & ~w3279;
assign w3281 = ~w3278 & w3280;
assign w3282 = ~w3037 & ~w3108;
assign w3283 = ~w3109 & ~w3282;
assign w3284 = ~w3281 & ~w3283;
assign w3285 = w1566 & ~w3222;
assign w3286 = w1568 & ~w3222;
assign w3287 = ~w3286 & w7487;
assign w3288 = w3285 & ~w3287;
assign w3289 = ~w3284 & w3288;
assign w3290 = ~w3285 & w3287;
assign w3291 = (~w3285 & w3278) | (~w3285 & w6189) | (w3278 & w6189);
assign w3292 = ~w3283 & w3291;
assign w3293 = ~w3290 & ~w3292;
assign w3294 = ~w3289 & w3293;
assign w3295 = ~w2924 & w3118;
assign w3296 = w2924 & ~w3118;
assign w3297 = ~w3295 & ~w3296;
assign w3298 = w2920 & ~w3297;
assign w3299 = ~w2920 & w3297;
assign w3300 = ~w3298 & ~w3299;
assign w3301 = w3111 & w3300;
assign w3302 = ~w3111 & ~w3300;
assign w3303 = ~w3301 & ~w3302;
assign w3304 = w3294 & w3303;
assign w3305 = (~w3224 & w3284) | (~w3224 & w7027) | (w3284 & w7027);
assign w3306 = ~w3304 & w3305;
assign w3307 = ~w3304 & w7028;
assign w3308 = w3122 & ~w3126;
assign w3309 = ~w3127 & ~w3308;
assign w3310 = ~w3284 & w7029;
assign w3311 = ~w3292 & w6190;
assign w3312 = w3303 & w3311;
assign w3313 = (~w3310 & ~w3303) | (~w3310 & w7030) | (~w3303 & w7030);
assign w3314 = ~w3312 & w6428;
assign w3315 = ~w3309 & w3314;
assign w3316 = (~w3307 & w3309) | (~w3307 & w7031) | (w3309 & w7031);
assign w3317 = (w3223 & w3304) | (w3223 & w7032) | (w3304 & w7032);
assign w3318 = (w3317 & w3309) | (w3317 & w7033) | (w3309 & w7033);
assign w3319 = w3316 & ~w3318;
assign w3320 = w3134 & ~w3139;
assign w3321 = w3128 & ~w3320;
assign w3322 = ~w3128 & w3320;
assign w3323 = ~w3321 & ~w3322;
assign w3324 = w3319 & ~w3323;
assign w3325 = w1774 & ~w3222;
assign w3326 = ~w3315 & w6429;
assign w3327 = (~w3325 & w3315) | (~w3325 & w6430) | (w3315 & w6430);
assign w3328 = ~w3326 & ~w3327;
assign w3329 = ~w3324 & w3328;
assign w3330 = w3319 & w6431;
assign w3331 = ~w3329 & ~w3330;
assign w3332 = w3211 & ~w3331;
assign w3333 = ~w1556 & ~w3222;
assign w3334 = (~w3333 & w3324) | (~w3333 & w7034) | (w3324 & w7034);
assign w3335 = ~w3332 & w3334;
assign w3336 = ~w3324 & w7035;
assign w3337 = w3316 & w3333;
assign w3338 = w1774 & w7036;
assign w3339 = (~w3338 & w3324) | (~w3338 & w6432) | (w3324 & w6432);
assign w3340 = (~w3336 & ~w3211) | (~w3336 & w7037) | (~w3211 & w7037);
assign w3341 = ~w3151 & ~w3154;
assign w3342 = w3156 & ~w3341;
assign w3343 = ~w3156 & w3341;
assign w3344 = ~w3342 & ~w3343;
assign w3345 = ~w3335 & w6433;
assign w3346 = (~w3344 & w3335) | (~w3344 & w6434) | (w3335 & w6434);
assign w3347 = ~w3345 & ~w3346;
assign w3348 = ~w3211 & w3331;
assign w3349 = ~w3332 & ~w3348;
assign w3350 = ~w3319 & w3323;
assign w3351 = ~w3324 & ~w3350;
assign w3352 = w1561 & ~w3205;
assign w3353 = ~w3294 & ~w3303;
assign w3354 = ~w3304 & ~w3353;
assign w3355 = w1566 & ~w3205;
assign w3356 = ~w3275 & ~w3279;
assign w3357 = w1568 & ~w3205;
assign w3358 = w3277 & ~w3357;
assign w3359 = w3356 & ~w3358;
assign w3360 = ~w3277 & ~w3357;
assign w3361 = ~w3356 & ~w3360;
assign w3362 = ~w3359 & ~w3361;
assign w3363 = ~w3260 & ~w3268;
assign w3364 = ~w1572 & ~w3264;
assign w3365 = ~w1579 & ~w1584;
assign w3366 = (~w1012 & w1579) | (~w1012 & w7039) | (w1579 & w7039);
assign w3367 = ~w1584 & w3029;
assign w3368 = ~w4 & w6992;
assign w3369 = w3028 & ~w3368;
assign w3370 = w3221 & w3369;
assign w3371 = ~w3370 & w7488;
assign w3372 = ~w3366 & w3371;
assign w3373 = w1590 & w3372;
assign w3374 = ~w1590 & ~w3372;
assign w3375 = ~w3230 & w3232;
assign w3376 = w3228 & ~w3375;
assign w3377 = ~w3228 & w3375;
assign w3378 = ~w3376 & ~w3377;
assign w3379 = ~w3241 & w3245;
assign w3380 = ~w3246 & ~w3379;
assign w3381 = ~w1576 & w3380;
assign w3382 = (~w3373 & w3378) | (~w3373 & w7041) | (w3378 & w7041);
assign w3383 = ~w3381 & w3382;
assign w3384 = w1576 & ~w3380;
assign w3385 = (w1648 & w3383) | (w1648 & w7042) | (w3383 & w7042);
assign w3386 = ~w1572 & w3264;
assign w3387 = w3363 & w3386;
assign w3388 = ~w3383 & w7043;
assign w3389 = ~w3254 & ~w3258;
assign w3390 = w3255 & ~w3389;
assign w3391 = ~w3255 & w3389;
assign w3392 = ~w3390 & ~w3391;
assign w3393 = ~w3388 & w3392;
assign w3394 = ~w3205 & ~w3385;
assign w3395 = (w3394 & ~w3364) | (w3394 & w7044) | (~w3364 & w7044);
assign w3396 = ~w3387 & ~w3393;
assign w3397 = w3395 & w3396;
assign w3398 = w3264 & w3363;
assign w3399 = w1572 & ~w3205;
assign w3400 = (w3399 & w3363) | (w3399 & w6191) | (w3363 & w6191);
assign w3401 = ~w3398 & w3400;
assign w3402 = w1570 & ~w3205;
assign w3403 = ~w3397 & w7045;
assign w3404 = (w3402 & w3397) | (w3402 & w6192) | (w3397 & w6192);
assign w3405 = ~w3269 & ~w3271;
assign w3406 = w3273 & ~w3405;
assign w3407 = ~w3273 & w3405;
assign w3408 = ~w3406 & ~w3407;
assign w3409 = ~w3404 & ~w3408;
assign w3410 = ~w3403 & ~w3409;
assign w3411 = ~w3362 & w3410;
assign w3412 = w3277 & w3356;
assign w3413 = (w3357 & w3356) | (w3357 & w7046) | (w3356 & w7046);
assign w3414 = ~w3412 & w3413;
assign w3415 = ~w3411 & w7047;
assign w3416 = (w3355 & w3411) | (w3355 & w6193) | (w3411 & w6193);
assign w3417 = ~w3281 & ~w3287;
assign w3418 = w3283 & ~w3417;
assign w3419 = ~w3283 & w3417;
assign w3420 = ~w3418 & ~w3419;
assign w3421 = ~w3416 & w3420;
assign w3422 = (w3352 & w3354) | (w3352 & w6194) | (w3354 & w6194);
assign w3423 = (~w3352 & ~w3354) | (~w3352 & w6195) | (~w3354 & w6195);
assign w3424 = ~w3422 & ~w3423;
assign w3425 = ~w1563 & w3352;
assign w3426 = (w3425 & ~w3354) | (w3425 & w6196) | (~w3354 & w6196);
assign w3427 = ~w1559 & w1563;
assign w3428 = w1563 & w7048;
assign w3429 = (w3428 & w3354) | (w3428 & w6197) | (w3354 & w6197);
assign w3430 = ~w3426 & ~w3429;
assign w3431 = ~w3424 & w3430;
assign w3432 = ~w3306 & w3313;
assign w3433 = w3309 & ~w3432;
assign w3434 = ~w3309 & w3432;
assign w3435 = ~w3433 & ~w3434;
assign w3436 = ~w3431 & ~w3435;
assign w3437 = w1774 & ~w3205;
assign w3438 = w3436 & ~w3437;
assign w3439 = w3422 & ~w3426;
assign w3440 = ~w1774 & w3439;
assign w3441 = w3437 & ~w3439;
assign w3442 = ~w3440 & ~w3441;
assign w3443 = ~w3436 & ~w3442;
assign w3444 = ~w3438 & ~w3443;
assign w3445 = ~w3351 & ~w3444;
assign w3446 = w3437 & ~w3443;
assign w3447 = ~w3445 & ~w3446;
assign w3448 = w3349 & ~w3447;
assign w3449 = ~w3349 & w3447;
assign w3450 = ~w1556 & ~w3205;
assign w3451 = (w3450 & w3349) | (w3450 & w6435) | (w3349 & w6435);
assign w3452 = ~w3448 & ~w3451;
assign w3453 = w3347 & w3452;
assign w3454 = (~w3206 & w3453) | (~w3206 & w7049) | (w3453 & w7049);
assign w3455 = ~w1086 & ~w3222;
assign w3456 = ~w3188 & ~w3190;
assign w3457 = ~w3191 & ~w3456;
assign w3458 = ~w6433 & ~w3335;
assign w3459 = (~w3458 & ~w3457) | (~w3458 & w7050) | (~w3457 & w7050);
assign w3460 = w2513 & ~w3222;
assign w3461 = ~w3183 & w6198;
assign w3462 = ~w3186 & w3461;
assign w3463 = ~w3187 & ~w3462;
assign w3464 = w3459 & ~w3463;
assign w3465 = ~w3332 & w7051;
assign w3466 = (~w3465 & ~w6433) | (~w3465 & w7052) | (~w6433 & w7052);
assign w3467 = ~w3457 & w3466;
assign w3468 = w3457 & ~w3466;
assign w3469 = ~w3467 & ~w3468;
assign w3470 = ~w3464 & w3469;
assign w3471 = w3184 & ~w3186;
assign w3472 = ~w3187 & ~w3471;
assign w3473 = ~w3459 & w3472;
assign w3474 = (~w3473 & ~w3470) | (~w3473 & w6199) | (~w3470 & w6199);
assign w3475 = w3197 & ~w3474;
assign w3476 = (~w3195 & w3474) | (~w3195 & w7053) | (w3474 & w7053);
assign w3477 = w3015 & ~w3476;
assign w3478 = (~w3013 & w3476) | (~w3013 & w7054) | (w3476 & w7054);
assign w3479 = ~w2663 & w2837;
assign w3480 = ~w2838 & ~w3479;
assign w3481 = ~w3478 & w3480;
assign w3482 = (~w2838 & w3478) | (~w2838 & w7055) | (w3478 & w7055);
assign w3483 = w2661 & w3482;
assign w3484 = (~w2659 & ~w3482) | (~w2659 & w7056) | (~w3482 & w7056);
assign w3485 = ~w2504 & w2506;
assign w3486 = ~w2507 & ~w3485;
assign w3487 = w3484 & w3486;
assign w3488 = w2374 & w7489;
assign w3489 = (w2367 & ~w2366) | (w2367 & w7057) | (~w2366 & w7057);
assign w3490 = (~w2361 & ~w2363) | (~w2361 & w6201) | (~w2363 & w6201);
assign w3491 = ~w1974 & ~w1978;
assign w3492 = ~w1979 & ~w3491;
assign w3493 = w3490 & ~w3492;
assign w3494 = ~w3490 & w3492;
assign w3495 = ~w3493 & ~w3494;
assign w3496 = w177 & w3495;
assign w3497 = ~w177 & ~w3495;
assign w3498 = ~w3496 & ~w3497;
assign w3499 = ~w3489 & ~w3498;
assign w3500 = w3489 & w3498;
assign w3501 = ~w3499 & ~w3500;
assign w3502 = w3488 & w3501;
assign w3503 = w1886 & ~w1981;
assign w3504 = ~w1982 & ~w3503;
assign w3505 = (~w3493 & ~w3495) | (~w3493 & w7058) | (~w3495 & w7058);
assign w3506 = ~w3504 & w3505;
assign w3507 = w3504 & ~w3505;
assign w3508 = ~w3506 & ~w3507;
assign w3509 = (w2372 & ~w3498) | (w2372 & w6202) | (~w3498 & w6202);
assign w3510 = (w3508 & w3509) | (w3508 & w7059) | (w3509 & w7059);
assign w3511 = ~w3509 & w7060;
assign w3512 = ~w3510 & ~w3511;
assign w3513 = w3502 & w3512;
assign w3514 = ~w3506 & ~w3510;
assign w3515 = (w3514 & ~w3502) | (w3514 & w7061) | (~w3502 & w7061);
assign w3516 = (~w1086 & w3515) | (~w1086 & w7062) | (w3515 & w7062);
assign w3517 = ~w2507 & w7490;
assign w3518 = ~w3488 & ~w3517;
assign w3519 = ~w3454 & w3469;
assign w3520 = w3454 & ~w3469;
assign w3521 = ~w3519 & ~w3520;
assign w3522 = ~w3347 & ~w3452;
assign w3523 = ~w3453 & ~w3522;
assign w3524 = ~w3448 & ~w3449;
assign w3525 = w3431 & w3435;
assign w3526 = ~w3436 & ~w3525;
assign w3527 = w3351 & w3444;
assign w3528 = ~w3445 & ~w3527;
assign w3529 = ~w1556 & ~w3528;
assign w3530 = (w3207 & w3528) | (w3207 & w7064) | (w3528 & w7064);
assign w3531 = w3524 & ~w3530;
assign w3532 = ~w3351 & ~w3526;
assign w3533 = ~w3444 & w3532;
assign w3534 = w3351 & ~w3526;
assign w3535 = w3444 & w3534;
assign w3536 = ~w3533 & ~w3535;
assign w3537 = ~w3450 & ~w3536;
assign w3538 = ~w3536 & w6204;
assign w3539 = (w3207 & w3536) | (w3207 & w7065) | (w3536 & w7065);
assign w3540 = ~w3524 & w7066;
assign w3541 = ~w3531 & ~w3540;
assign w3542 = w3523 & ~w3541;
assign w3543 = ~w3523 & w3541;
assign w3544 = ~w3542 & ~w3543;
assign w3545 = w3450 & w3536;
assign w3546 = ~w3537 & ~w3545;
assign w3547 = w3524 & ~w3546;
assign w3548 = ~w3524 & w3546;
assign w3549 = ~w3547 & ~w3548;
assign w3550 = w3549 & w7067;
assign w3551 = ~w3544 & w3550;
assign w3552 = ~w3521 & w3551;
assign w3553 = ~w3464 & ~w3473;
assign w3554 = ~w3519 & w3553;
assign w3555 = w3519 & ~w3553;
assign w3556 = ~w3554 & ~w3555;
assign w3557 = w3552 & w3556;
assign w3558 = ~w3197 & w3474;
assign w3559 = ~w3475 & ~w3558;
assign w3560 = w3557 & ~w3559;
assign w3561 = ~w3015 & w3476;
assign w3562 = ~w3477 & ~w3561;
assign w3563 = w3560 & ~w3562;
assign w3564 = w3478 & ~w3480;
assign w3565 = ~w3481 & ~w3564;
assign w3566 = w3563 & ~w3565;
assign w3567 = ~w2661 & ~w3482;
assign w3568 = ~w3483 & ~w3567;
assign w3569 = w3566 & w3568;
assign w3570 = ~w3484 & ~w3486;
assign w3571 = ~w3487 & ~w3570;
assign w3572 = w3569 & ~w3571;
assign w3573 = ~w3518 & w3572;
assign w3574 = (w3501 & w3488) | (w3501 & w7068) | (w3488 & w7068);
assign w3575 = ~w3488 & w7069;
assign w3576 = ~w3574 & ~w3575;
assign w3577 = w3573 & ~w3576;
assign w3578 = ~w3502 & ~w3512;
assign w3579 = ~w3513 & ~w3578;
assign w3580 = w3577 & ~w3579;
assign w3581 = ~w3516 & ~w3580;
assign w3582 = ~w3580 & w7070;
assign w3583 = ~w3516 & w3580;
assign w3584 = w3516 & ~w3580;
assign w3585 = ~w3583 & ~w3584;
assign w3586 = ~w1584 & w3585;
assign w3587 = ~w3577 & w3579;
assign w3588 = ~w3580 & ~w3587;
assign w3589 = ~w1584 & w3588;
assign w3590 = ~w3566 & ~w3568;
assign w3591 = ~w3569 & ~w3590;
assign w3592 = ~w1584 & w3591;
assign w3593 = ~w3563 & w3565;
assign w3594 = ~w3566 & ~w3593;
assign w3595 = ~w1579 & w3594;
assign w3596 = ~w3557 & w3559;
assign w3597 = ~w3560 & ~w3596;
assign w3598 = w1590 & w3597;
assign w3599 = ~w3552 & ~w3556;
assign w3600 = ~w3557 & ~w3599;
assign w3601 = w1590 & w3600;
assign w3602 = w3521 & ~w3551;
assign w3603 = ~w3552 & ~w3602;
assign w3604 = w1590 & w3603;
assign w3605 = w1572 & w3526;
assign w3606 = w3351 & w3526;
assign w3607 = ~w3532 & ~w3606;
assign w3608 = w3444 & w3607;
assign w3609 = ~w3444 & ~w3607;
assign w3610 = ~w3608 & ~w3609;
assign w3611 = (~w3605 & ~w3610) | (~w3605 & w6205) | (~w3610 & w6205);
assign w3612 = ~w1648 & w3526;
assign w3613 = ~w1572 & ~w1576;
assign w3614 = w1572 & w1576;
assign w3615 = ~w3613 & ~w3614;
assign w3616 = ~w3528 & w6206;
assign w3617 = (~w1576 & w3528) | (~w1576 & w7071) | (w3528 & w7071);
assign w3618 = ~w3611 & w3617;
assign w3619 = ~w3549 & w3618;
assign w3620 = ~w3528 & w7072;
assign w3621 = (~w3620 & w3549) | (~w3620 & w6207) | (w3549 & w6207);
assign w3622 = ~w3544 & ~w3621;
assign w3623 = ~w1576 & w3621;
assign w3624 = w3544 & w3623;
assign w3625 = ~w3622 & ~w3624;
assign w3626 = w1570 & w3526;
assign w3627 = (~w3626 & ~w3610) | (~w3626 & w7073) | (~w3610 & w7073);
assign w3628 = w1569 & ~w1571;
assign w3629 = ~w3528 & w7074;
assign w3630 = ~w3627 & ~w3629;
assign w3631 = w3549 & ~w3630;
assign w3632 = w3526 & w7075;
assign w3633 = ~w3528 & w3632;
assign w3634 = (w1648 & w3627) | (w1648 & w7076) | (w3627 & w7076);
assign w3635 = ~w1648 & ~w3627;
assign w3636 = (~w3634 & w3549) | (~w3634 & w7077) | (w3549 & w7077);
assign w3637 = ~w3629 & ~w3636;
assign w3638 = ~w3631 & ~w3637;
assign w3639 = ~w3625 & ~w3638;
assign w3640 = w3625 & w3638;
assign w3641 = ~w3639 & ~w3640;
assign w3642 = ~w3604 & w3641;
assign w3643 = w3604 & ~w3641;
assign w3644 = (w3612 & ~w3610) | (w3612 & w7078) | (~w3610 & w7078);
assign w3645 = w3610 & w7079;
assign w3646 = ~w3644 & ~w3645;
assign w3647 = ~w3549 & w7080;
assign w3648 = (w3646 & w3549) | (w3646 & w7081) | (w3549 & w7081);
assign w3649 = ~w3647 & ~w3648;
assign w3650 = ~w1576 & w3526;
assign w3651 = w3610 & w7082;
assign w3652 = w3649 & w3651;
assign w3653 = (~w3647 & ~w3649) | (~w3647 & w6208) | (~w3649 & w6208);
assign w3654 = w1590 & w3544;
assign w3655 = w3653 & ~w3654;
assign w3656 = w3544 & ~w3653;
assign w3657 = ~w3611 & ~w3616;
assign w3658 = (~w3657 & w3549) | (~w3657 & w7083) | (w3549 & w7083);
assign w3659 = ~w3619 & ~w3658;
assign w3660 = ~w3656 & ~w3659;
assign w3661 = ~w3655 & ~w3660;
assign w3662 = ~w3643 & ~w3661;
assign w3663 = ~w3642 & ~w3662;
assign w3664 = (~w3601 & w3662) | (~w3601 & w7084) | (w3662 & w7084);
assign w3665 = ~w3662 & w6209;
assign w3666 = ~w1576 & w3603;
assign w3667 = (w3621 & ~w3544) | (w3621 & w7085) | (~w3544 & w7085);
assign w3668 = (~w3667 & w3625) | (~w3667 & w7086) | (w3625 & w7086);
assign w3669 = w3666 & w3668;
assign w3670 = ~w3666 & ~w3668;
assign w3671 = ~w3669 & ~w3670;
assign w3672 = (~w3629 & w3549) | (~w3629 & w7087) | (w3549 & w7087);
assign w3673 = (~w1648 & w3544) | (~w1648 & w6210) | (w3544 & w6210);
assign w3674 = w3544 & ~w3672;
assign w3675 = w3673 & ~w3674;
assign w3676 = w3526 & w7088;
assign w3677 = ~w3528 & w7089;
assign w3678 = w1568 & w3526;
assign w3679 = (~w3678 & ~w3610) | (~w3678 & w7090) | (~w3610 & w7090);
assign w3680 = ~w3528 & w3676;
assign w3681 = ~w3528 & w7091;
assign w3682 = ~w3677 & ~w3681;
assign w3683 = ~w3679 & w3682;
assign w3684 = (w3683 & w3549) | (w3683 & w7092) | (w3549 & w7092);
assign w3685 = ~w3549 & w7093;
assign w3686 = ~w3684 & ~w3685;
assign w3687 = w3675 & w3686;
assign w3688 = ~w3675 & ~w3686;
assign w3689 = ~w3687 & ~w3688;
assign w3690 = w3671 & ~w3689;
assign w3691 = ~w3671 & w3689;
assign w3692 = ~w3690 & ~w3691;
assign w3693 = ~w3665 & ~w3692;
assign w3694 = ~w3693 & w6211;
assign w3695 = (~w3598 & w3693) | (~w3598 & w6212) | (w3693 & w6212);
assign w3696 = ~w3694 & ~w3695;
assign w3697 = ~w1576 & w3600;
assign w3698 = ~w3669 & w3689;
assign w3699 = ~w3698 & w6213;
assign w3700 = (~w3697 & w3698) | (~w3697 & w6214) | (w3698 & w6214);
assign w3701 = ~w3699 & ~w3700;
assign w3702 = (w3686 & ~w3544) | (w3686 & w7094) | (~w3544 & w7094);
assign w3703 = w3673 & ~w3702;
assign w3704 = (~w3703 & ~w3603) | (~w3703 & w7095) | (~w3603 & w7095);
assign w3705 = w3603 & w3703;
assign w3706 = (w3610 & w7096) | (w3610 & w7097) | (w7096 & w7097);
assign w3707 = (~w3677 & w3549) | (~w3677 & w6216) | (w3549 & w6216);
assign w3708 = ~w3544 & ~w3707;
assign w3709 = (w3549 & w7098) | (w3549 & w7099) | (w7098 & w7099);
assign w3710 = w3544 & w3709;
assign w3711 = ~w3708 & ~w3710;
assign w3712 = w1566 & w3526;
assign w3713 = (w3712 & ~w3610) | (w3712 & w7100) | (~w3610 & w7100);
assign w3714 = w3610 & w7101;
assign w3715 = ~w3713 & ~w3714;
assign w3716 = ~w3549 & w3680;
assign w3717 = (~w3680 & w3549) | (~w3680 & w6217) | (w3549 & w6217);
assign w3718 = ~w3716 & ~w3717;
assign w3719 = w3715 & ~w3718;
assign w3720 = ~w3715 & w3718;
assign w3721 = ~w3719 & ~w3720;
assign w3722 = ~w3711 & ~w3721;
assign w3723 = w3711 & w3721;
assign w3724 = ~w3722 & ~w3723;
assign w3725 = ~w3704 & w3741;
assign w3726 = (~w3724 & w3704) | (~w3724 & w6218) | (w3704 & w6218);
assign w3727 = ~w3725 & ~w3726;
assign w3728 = w3701 & ~w3727;
assign w3729 = ~w3701 & w3727;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = w3696 & w3730;
assign w3732 = ~w3560 & w3562;
assign w3733 = ~w3563 & ~w3732;
assign w3734 = w1590 & w3733;
assign w3735 = (~w3734 & w3693) | (~w3734 & w6518) | (w3693 & w6518);
assign w3736 = (w3735 & ~w3696) | (w3735 & w7102) | (~w3696 & w7102);
assign w3737 = ~w3693 & w6519;
assign w3738 = (~w3737 & w3731) | (~w3737 & w6436) | (w3731 & w6436);
assign w3739 = w3696 & w6437;
assign w3740 = ~w1648 & w3600;
assign w3741 = ~w3705 & w3724;
assign w3742 = ~w3704 & ~w3741;
assign w3743 = w3740 & w3742;
assign w3744 = ~w3740 & ~w3742;
assign w3745 = ~w3743 & ~w3744;
assign w3746 = w1572 & w3603;
assign w3747 = (w3707 & ~w3544) | (w3707 & w7103) | (~w3544 & w7103);
assign w3748 = (~w3747 & w3711) | (~w3747 & w7104) | (w3711 & w7104);
assign w3749 = w3746 & w3748;
assign w3750 = ~w3746 & ~w3748;
assign w3751 = ~w3749 & ~w3750;
assign w3752 = w3610 & w7105;
assign w3753 = (~w3752 & w3549) | (~w3752 & w7106) | (w3549 & w7106);
assign w3754 = ~w3680 & w3715;
assign w3755 = ~w3753 & ~w3754;
assign w3756 = w3544 & w3755;
assign w3757 = w1570 & w3544;
assign w3758 = (~w3755 & ~w3544) | (~w3755 & w7107) | (~w3544 & w7107);
assign w3759 = w1568 & ~w3549;
assign w3760 = ~w3528 & w7108;
assign w3761 = ~w3528 & w7109;
assign w3762 = w1563 & w3526;
assign w3763 = (w3762 & w3528) | (w3762 & w7110) | (w3528 & w7110);
assign w3764 = w3610 & w7111;
assign w3765 = ~w3760 & ~w3763;
assign w3766 = ~w3764 & w3765;
assign w3767 = ~w3761 & ~w3766;
assign w3768 = w3759 & ~w3767;
assign w3769 = ~w3759 & w3767;
assign w3770 = ~w3768 & ~w3769;
assign w3771 = ~w3758 & w6219;
assign w3772 = (~w3770 & w3758) | (~w3770 & w6220) | (w3758 & w6220);
assign w3773 = ~w3771 & ~w3772;
assign w3774 = w3751 & ~w3773;
assign w3775 = ~w3751 & w3773;
assign w3776 = ~w3774 & ~w3775;
assign w3777 = w3745 & ~w3776;
assign w3778 = ~w3745 & w3776;
assign w3779 = ~w3777 & ~w3778;
assign w3780 = ~w3699 & w3727;
assign w3781 = ~w3700 & ~w3780;
assign w3782 = ~w1576 & w3597;
assign w3783 = (~w3782 & w3780) | (~w3782 & w6438) | (w3780 & w6438);
assign w3784 = ~w3700 & w3782;
assign w3785 = ~w3780 & w3784;
assign w3786 = ~w3783 & ~w3785;
assign w3787 = w3779 & w3786;
assign w3788 = ~w3779 & ~w3786;
assign w3789 = ~w3787 & ~w3788;
assign w3790 = ~w3739 & w3789;
assign w3791 = w3738 & w3790;
assign w3792 = (~w3789 & ~w3738) | (~w3789 & w6520) | (~w3738 & w6520);
assign w3793 = ~w3791 & ~w3792;
assign w3794 = ~w3696 & ~w3730;
assign w3795 = ~w3731 & ~w3794;
assign w3796 = ~w1579 & w3733;
assign w3797 = w3795 & w3796;
assign w3798 = ~w3795 & ~w3796;
assign w3799 = ~w3797 & ~w3798;
assign w3800 = ~w1579 & w3597;
assign w3801 = ~w1579 & w3600;
assign w3802 = ~w1579 & w3603;
assign w3803 = (~w3650 & ~w3610) | (~w3650 & w7112) | (~w3610 & w7112);
assign w3804 = ~w3651 & ~w3803;
assign w3805 = ~w1579 & ~w3549;
assign w3806 = (~w3804 & w3549) | (~w3804 & w7113) | (w3549 & w7113);
assign w3807 = w1590 & w3526;
assign w3808 = ~w3528 & w7114;
assign w3809 = ~w3549 & w7115;
assign w3810 = ~w3806 & ~w3809;
assign w3811 = ~w3808 & w3810;
assign w3812 = (~w3806 & ~w3810) | (~w3806 & w6221) | (~w3810 & w6221);
assign w3813 = ~w1579 & w3544;
assign w3814 = ~w3812 & ~w3813;
assign w3815 = w3544 & w3812;
assign w3816 = ~w3814 & ~w3815;
assign w3817 = ~w3649 & ~w3651;
assign w3818 = ~w3652 & ~w3817;
assign w3819 = ~w3814 & w7116;
assign w3820 = (~w3814 & ~w3816) | (~w3814 & w6439) | (~w3816 & w6439);
assign w3821 = w3802 & w3820;
assign w3822 = ~w3802 & ~w3820;
assign w3823 = ~w3821 & ~w3822;
assign w3824 = (w3659 & w3655) | (w3659 & w7117) | (w3655 & w7117);
assign w3825 = ~w3655 & w3660;
assign w3826 = ~w3824 & ~w3825;
assign w3827 = w3823 & ~w3826;
assign w3828 = (~w3821 & ~w3823) | (~w3821 & w6521) | (~w3823 & w6521);
assign w3829 = w3801 & ~w3828;
assign w3830 = ~w3801 & w3828;
assign w3831 = ~w3642 & ~w3643;
assign w3832 = ~w3661 & w3831;
assign w3833 = w3661 & ~w3831;
assign w3834 = ~w3832 & ~w3833;
assign w3835 = ~w3830 & ~w3834;
assign w3836 = ~w3835 & w7118;
assign w3837 = (w3800 & w3835) | (w3800 & w7119) | (w3835 & w7119);
assign w3838 = ~w3664 & ~w3665;
assign w3839 = ~w3692 & w3838;
assign w3840 = w3692 & ~w3838;
assign w3841 = ~w3839 & ~w3840;
assign w3842 = ~w3837 & w3841;
assign w3843 = ~w3836 & ~w3842;
assign w3844 = w3799 & w3843;
assign w3845 = (~w3797 & ~w3799) | (~w3797 & w6440) | (~w3799 & w6440);
assign w3846 = ~w3793 & ~w3845;
assign w3847 = w3793 & w3845;
assign w3848 = ~w3846 & ~w3847;
assign w3849 = w3595 & ~w3848;
assign w3850 = ~w3595 & w3848;
assign w3851 = ~w3849 & ~w3850;
assign w3852 = ~w3592 & w3851;
assign w3853 = ~w1584 & w3733;
assign w3854 = ~w1584 & w3600;
assign w3855 = (w3818 & w3814) | (w3818 & w7120) | (w3814 & w7120);
assign w3856 = ~w3819 & ~w3855;
assign w3857 = w3808 & ~w3810;
assign w3858 = ~w3811 & ~w3857;
assign w3859 = ~w3528 & w7121;
assign w3860 = ~w3549 & w3859;
assign w3861 = (~w3807 & ~w3610) | (~w3807 & w7122) | (~w3610 & w7122);
assign w3862 = ~w3808 & ~w3861;
assign w3863 = w3549 & ~w3859;
assign w3864 = (~w1584 & w3549) | (~w1584 & w6222) | (w3549 & w6222);
assign w3865 = ~w3863 & w3864;
assign w3866 = w3862 & w3865;
assign w3867 = (~w3860 & ~w3865) | (~w3860 & w7123) | (~w3865 & w7123);
assign w3868 = ~w3858 & ~w3867;
assign w3869 = ~w1584 & w3544;
assign w3870 = w3858 & w3867;
assign w3871 = ~w3868 & ~w3870;
assign w3872 = w3869 & w3871;
assign w3873 = (~w3868 & ~w3871) | (~w3868 & w6223) | (~w3871 & w6223);
assign w3874 = w3856 & w3873;
assign w3875 = ~w1584 & w3603;
assign w3876 = ~w3856 & ~w3873;
assign w3877 = ~w3874 & ~w3876;
assign w3878 = ~w3875 & w3877;
assign w3879 = (~w3874 & ~w3877) | (~w3874 & w6441) | (~w3877 & w6441);
assign w3880 = w3854 & w3879;
assign w3881 = ~w3823 & w3826;
assign w3882 = ~w3827 & ~w3881;
assign w3883 = ~w3854 & ~w3879;
assign w3884 = ~w3880 & ~w3883;
assign w3885 = w3882 & w3884;
assign w3886 = (~w3880 & ~w3884) | (~w3880 & w6522) | (~w3884 & w6522);
assign w3887 = w3597 & ~w3886;
assign w3888 = ~w1584 & w3597;
assign w3889 = w3886 & ~w3888;
assign w3890 = ~w3829 & ~w3830;
assign w3891 = ~w3834 & w3890;
assign w3892 = w3834 & ~w3890;
assign w3893 = ~w3891 & ~w3892;
assign w3894 = ~w3889 & w3893;
assign w3895 = (w3853 & w3894) | (w3853 & w7124) | (w3894 & w7124);
assign w3896 = ~w3894 & w7125;
assign w3897 = ~w3836 & ~w3837;
assign w3898 = w3841 & w3897;
assign w3899 = ~w3841 & ~w3897;
assign w3900 = ~w3898 & ~w3899;
assign w3901 = ~w3896 & ~w3900;
assign w3902 = (w3594 & w3901) | (w3594 & w7126) | (w3901 & w7126);
assign w3903 = ~w1584 & w3594;
assign w3904 = ~w3901 & w7127;
assign w3905 = ~w3799 & ~w3843;
assign w3906 = ~w3844 & ~w3905;
assign w3907 = (~w3902 & ~w3906) | (~w3902 & w7128) | (~w3906 & w7128);
assign w3908 = ~w3852 & ~w3907;
assign w3909 = w3592 & ~w3851;
assign w3910 = ~w3569 & w3571;
assign w3911 = ~w3572 & ~w3910;
assign w3912 = ~w1584 & w3911;
assign w3913 = (~w3912 & w3851) | (~w3912 & w6523) | (w3851 & w6523);
assign w3914 = ~w3908 & w3913;
assign w3915 = ~w1579 & w3591;
assign w3916 = (w3595 & ~w3845) | (w3595 & w6524) | (~w3845 & w6524);
assign w3917 = ~w3846 & ~w3916;
assign w3918 = ~w3915 & w3917;
assign w3919 = w3915 & ~w3917;
assign w3920 = ~w3918 & ~w3919;
assign w3921 = w1590 & w3594;
assign w3922 = ~w3736 & ~w3791;
assign w3923 = ~w1576 & w3733;
assign w3924 = w3779 & ~w3785;
assign w3925 = (~w3923 & w3924) | (~w3923 & w6224) | (w3924 & w6224);
assign w3926 = ~w3924 & w6225;
assign w3927 = ~w3925 & ~w3926;
assign w3928 = w1572 & w3600;
assign w3929 = ~w3750 & ~w3773;
assign w3930 = (w3928 & w3929) | (w3928 & w6226) | (w3929 & w6226);
assign w3931 = ~w3749 & ~w3928;
assign w3932 = ~w3929 & w3931;
assign w3933 = ~w3930 & ~w3932;
assign w3934 = w1570 & w3603;
assign w3935 = (~w3770 & w3757) | (~w3770 & w6227) | (w3757 & w6227);
assign w3936 = ~w3756 & ~w3935;
assign w3937 = ~w3934 & w3936;
assign w3938 = w3934 & ~w3936;
assign w3939 = ~w3937 & ~w3938;
assign w3940 = (~w3761 & ~w3759) | (~w3761 & w6228) | (~w3759 & w6228);
assign w3941 = w3544 & ~w3940;
assign w3942 = (w3940 & ~w3544) | (w3940 & w6229) | (~w3544 & w6229);
assign w3943 = ~w3941 & ~w3942;
assign w3944 = w1566 & ~w3549;
assign w3945 = w1561 & ~w3528;
assign w3946 = w3763 & w3945;
assign w3947 = ~w3528 & w7129;
assign w3948 = w1561 & w3526;
assign w3949 = (~w3948 & ~w3610) | (~w3948 & w6230) | (~w3610 & w6230);
assign w3950 = ~w3947 & ~w3949;
assign w3951 = ~w3946 & w3950;
assign w3952 = w3944 & w3951;
assign w3953 = ~w3944 & ~w3951;
assign w3954 = ~w3952 & ~w3953;
assign w3955 = ~w3943 & w3954;
assign w3956 = w3943 & ~w3954;
assign w3957 = ~w3955 & ~w3956;
assign w3958 = w3939 & w3957;
assign w3959 = ~w3939 & ~w3957;
assign w3960 = ~w3958 & ~w3959;
assign w3961 = w3933 & ~w3960;
assign w3962 = ~w3933 & w3960;
assign w3963 = ~w3961 & ~w3962;
assign w3964 = ~w1648 & w3597;
assign w3965 = (~w3964 & w3777) | (~w3964 & w6231) | (w3777 & w6231);
assign w3966 = ~w3777 & w6232;
assign w3967 = ~w3965 & ~w3966;
assign w3968 = w3963 & ~w3967;
assign w3969 = ~w3963 & w3967;
assign w3970 = ~w3968 & ~w3969;
assign w3971 = w3927 & w3970;
assign w3972 = ~w3927 & ~w3970;
assign w3973 = ~w3971 & ~w3972;
assign w3974 = w3922 & ~w3973;
assign w3975 = ~w3922 & w3973;
assign w3976 = ~w3974 & ~w3975;
assign w3977 = ~w3921 & ~w3976;
assign w3978 = w3921 & w3976;
assign w3979 = ~w3977 & ~w3978;
assign w3980 = w3920 & w3979;
assign w3981 = ~w3920 & ~w3979;
assign w3982 = ~w3980 & ~w3981;
assign w3983 = ~w3914 & w3982;
assign w3984 = w3518 & ~w3572;
assign w3985 = ~w3573 & ~w3984;
assign w3986 = ~w1584 & w3985;
assign w3987 = (w3907 & w3851) | (w3907 & w7130) | (w3851 & w7130);
assign w3988 = (w3911 & ~w3851) | (w3911 & w6525) | (~w3851 & w6525);
assign w3989 = ~w3987 & w3988;
assign w3990 = (~w3986 & w3987) | (~w3986 & w6526) | (w3987 & w6526);
assign w3991 = ~w3983 & w3990;
assign w3992 = ~w1579 & w3911;
assign w3993 = ~w3919 & ~w3979;
assign w3994 = (~w3992 & w3993) | (~w3992 & w7131) | (w3993 & w7131);
assign w3995 = ~w3993 & w7132;
assign w3996 = ~w3994 & ~w3995;
assign w3997 = ~w3921 & ~w3974;
assign w3998 = w1590 & w3591;
assign w3999 = ~w3975 & w3998;
assign w4000 = ~w3997 & w3999;
assign w4001 = w3921 & ~w3975;
assign w4002 = ~w3974 & ~w3998;
assign w4003 = ~w4001 & w4002;
assign w4004 = ~w4000 & ~w4003;
assign w4005 = ~w1576 & w3594;
assign w4006 = w4005 & ~w3925;
assign w4007 = ~w3971 & w4006;
assign w4008 = (~w4005 & w3971) | (~w4005 & w6442) | (w3971 & w6442);
assign w4009 = ~w4007 & ~w4008;
assign w4010 = ~w1648 & w3733;
assign w4011 = w3963 & ~w3965;
assign w4012 = (w4010 & w4011) | (w4010 & w6443) | (w4011 & w6443);
assign w4013 = ~w4011 & w6444;
assign w4014 = ~w4012 & ~w4013;
assign w4015 = w1572 & w3597;
assign w4016 = ~w3932 & w4015;
assign w4017 = ~w3960 & w4016;
assign w4018 = w3597 & w3930;
assign w4019 = ~w4017 & ~w4018;
assign w4020 = ~w3930 & ~w4015;
assign w4021 = ~w3961 & w4020;
assign w4022 = w4019 & ~w4021;
assign w4023 = w1570 & w3600;
assign w4024 = ~w3937 & ~w3957;
assign w4025 = (w4023 & w4024) | (w4023 & w6233) | (w4024 & w6233);
assign w4026 = ~w4024 & w6234;
assign w4027 = ~w4025 & ~w4026;
assign w4028 = (~w3947 & ~w3944) | (~w3947 & w6235) | (~w3944 & w6235);
assign w4029 = w3544 & ~w4028;
assign w4030 = ~w3528 & w7134;
assign w4031 = w1774 & w3526;
assign w4032 = w3610 & w7135;
assign w4033 = ~w4031 & ~w4032;
assign w4034 = w1563 & ~w3549;
assign w4035 = ~w3549 & w7136;
assign w4036 = (w4033 & w3549) | (w4033 & w7137) | (w3549 & w7137);
assign w4037 = (~w4030 & ~w4034) | (~w4030 & w6236) | (~w4034 & w6236);
assign w4038 = ~w4036 & w4037;
assign w4039 = ~w4029 & ~w4038;
assign w4040 = (w4028 & ~w3544) | (w4028 & w6237) | (~w3544 & w6237);
assign w4041 = w4039 & ~w4040;
assign w4042 = w3544 & w6238;
assign w4043 = ~w3544 & ~w4028;
assign w4044 = w4038 & ~w4043;
assign w4045 = ~w4042 & w4044;
assign w4046 = ~w4041 & ~w4045;
assign w4047 = ~w3941 & ~w3954;
assign w4048 = ~w3942 & ~w4047;
assign w4049 = w1568 & w3603;
assign w4050 = ~w4048 & ~w4049;
assign w4051 = w3603 & w4048;
assign w4052 = (w4046 & w4050) | (w4046 & w6239) | (w4050 & w6239);
assign w4053 = ~w4050 & w6240;
assign w4054 = ~w4052 & ~w4053;
assign w4055 = ~w4027 & w4054;
assign w4056 = w4027 & ~w4054;
assign w4057 = ~w4055 & ~w4056;
assign w4058 = ~w4022 & w4057;
assign w4059 = w4022 & ~w4057;
assign w4060 = ~w4058 & ~w4059;
assign w4061 = w4014 & ~w4060;
assign w4062 = ~w4014 & w4060;
assign w4063 = ~w4061 & ~w4062;
assign w4064 = w4009 & ~w4063;
assign w4065 = ~w4009 & w4063;
assign w4066 = ~w4064 & ~w4065;
assign w4067 = w4004 & ~w4066;
assign w4068 = ~w4004 & w4066;
assign w4069 = ~w4067 & ~w4068;
assign w4070 = w3996 & ~w4069;
assign w4071 = ~w3996 & w4069;
assign w4072 = ~w4070 & ~w4071;
assign w4073 = ~w3991 & w4072;
assign w4074 = ~w3573 & w3576;
assign w4075 = ~w3577 & ~w4074;
assign w4076 = ~w1584 & w4075;
assign w4077 = (w3986 & w3983) | (w3986 & w6527) | (w3983 & w6527);
assign w4078 = ~w4076 & ~w4077;
assign w4079 = ~w4073 & w4078;
assign w4080 = ~w1579 & w3985;
assign w4081 = ~w4000 & ~w4066;
assign w4082 = w1590 & w3911;
assign w4083 = ~w4003 & w4082;
assign w4084 = ~w4081 & w4083;
assign w4085 = ~w4003 & w4066;
assign w4086 = ~w4000 & ~w4082;
assign w4087 = ~w4085 & w4086;
assign w4088 = ~w4084 & ~w4087;
assign w4089 = w3594 & w7138;
assign w4090 = (~w4089 & w3971) | (~w4089 & w6445) | (w3971 & w6445);
assign w4091 = ~w4063 & ~w4090;
assign w4092 = ~w1576 & w3591;
assign w4093 = (~w4092 & w3971) | (~w4092 & w6528) | (w3971 & w6528);
assign w4094 = ~w4091 & w4093;
assign w4095 = ~w4007 & w4063;
assign w4096 = w4092 & ~w3925;
assign w4097 = w3594 & w7139;
assign w4098 = (~w4097 & w3971) | (~w4097 & w6446) | (w3971 & w6446);
assign w4099 = ~w4095 & ~w4098;
assign w4100 = ~w4094 & ~w4099;
assign w4101 = ~w4012 & ~w4060;
assign w4102 = ~w1648 & w3594;
assign w4103 = (w4102 & w4011) | (w4102 & w7140) | (w4011 & w7140);
assign w4104 = (w4103 & w4060) | (w4103 & w7141) | (w4060 & w7141);
assign w4105 = ~w4102 & ~w4012;
assign w4106 = (w4105 & ~w4060) | (w4105 & w7142) | (~w4060 & w7142);
assign w4107 = ~w4104 & ~w4106;
assign w4108 = w1572 & w3733;
assign w4109 = ~w3961 & w6447;
assign w4110 = ~w4017 & w6241;
assign w4111 = w4057 & w4110;
assign w4112 = ~w4109 & ~w4111;
assign w4113 = w4019 & w4057;
assign w4114 = (w4108 & w3961) | (w4108 & w6448) | (w3961 & w6448);
assign w4115 = ~w4113 & w4114;
assign w4116 = w4112 & ~w4115;
assign w4117 = ~w4025 & ~w4054;
assign w4118 = w1570 & w3597;
assign w4119 = ~w4026 & w4118;
assign w4120 = ~w4117 & w4119;
assign w4121 = ~w4026 & w4054;
assign w4122 = ~w4025 & ~w4118;
assign w4123 = ~w4121 & w4122;
assign w4124 = ~w4120 & ~w4123;
assign w4125 = w1566 & w3603;
assign w4126 = ~w4039 & ~w4040;
assign w4127 = ~w4125 & ~w4126;
assign w4128 = w4125 & w4126;
assign w4129 = ~w4127 & ~w4128;
assign w4130 = w3526 & w7143;
assign w4131 = ~w3528 & w7144;
assign w4132 = ~w4035 & ~w4131;
assign w4133 = (w4132 & ~w3544) | (w4132 & w7145) | (~w3544 & w7145);
assign w4134 = w3544 & ~w4132;
assign w4135 = ~w1556 & w3526;
assign w4136 = (~w4135 & ~w3610) | (~w4135 & w6242) | (~w3610 & w6242);
assign w4137 = w1555 & ~w1773;
assign w4138 = ~w3528 & w7146;
assign w4139 = ~w4136 & ~w4138;
assign w4140 = ~w3528 & w7147;
assign w4141 = ~w4139 & ~w4140;
assign w4142 = ~w4136 & w7148;
assign w4143 = ~w4141 & ~w4142;
assign w4144 = w1561 & ~w3549;
assign w4145 = ~w4143 & w4144;
assign w4146 = w4143 & ~w4144;
assign w4147 = ~w4145 & ~w4146;
assign w4148 = ~w4133 & w4240;
assign w4149 = (~w4147 & w4133) | (~w4147 & w6449) | (w4133 & w6449);
assign w4150 = ~w4148 & ~w4149;
assign w4151 = w4129 & w4150;
assign w4152 = ~w4129 & ~w4150;
assign w4153 = ~w4151 & ~w4152;
assign w4154 = w1568 & w3600;
assign w4155 = w4046 & ~w4051;
assign w4156 = ~w4050 & ~w4155;
assign w4157 = w4154 & w4156;
assign w4158 = ~w4154 & ~w4156;
assign w4159 = ~w4157 & ~w4158;
assign w4160 = w4153 & ~w4159;
assign w4161 = ~w4153 & w4159;
assign w4162 = ~w4160 & ~w4161;
assign w4163 = w4124 & w4162;
assign w4164 = ~w4124 & ~w4162;
assign w4165 = ~w4163 & ~w4164;
assign w4166 = ~w4116 & w4165;
assign w4167 = w4116 & ~w4165;
assign w4168 = ~w4166 & ~w4167;
assign w4169 = w4107 & ~w4168;
assign w4170 = ~w4107 & w4168;
assign w4171 = ~w4169 & ~w4170;
assign w4172 = w4100 & w4171;
assign w4173 = ~w4100 & ~w4171;
assign w4174 = ~w4172 & ~w4173;
assign w4175 = ~w4088 & w4174;
assign w4176 = w4088 & ~w4174;
assign w4177 = ~w4175 & ~w4176;
assign w4178 = w4080 & ~w4177;
assign w4179 = ~w4080 & w4177;
assign w4180 = ~w4178 & ~w4179;
assign w4181 = ~w3995 & w4069;
assign w4182 = ~w3994 & ~w4181;
assign w4183 = w4180 & w4182;
assign w4184 = ~w4180 & ~w4182;
assign w4185 = ~w4183 & ~w4184;
assign w4186 = ~w4079 & w4185;
assign w4187 = (w4076 & w3983) | (w4076 & w6529) | (w3983 & w6529);
assign w4188 = w4072 & w4187;
assign w4189 = (w3983 & w7149) | (w3983 & w7150) | (w7149 & w7150);
assign w4190 = ~w4188 & ~w4189;
assign w4191 = (w3589 & w4186) | (w3589 & w7151) | (w4186 & w7151);
assign w4192 = ~w3589 & w4190;
assign w4193 = ~w4186 & w4192;
assign w4194 = ~w1579 & w4075;
assign w4195 = w1590 & w3985;
assign w4196 = ~w4084 & ~w4174;
assign w4197 = ~w4087 & ~w4196;
assign w4198 = (~w4195 & w4196) | (~w4195 & w6530) | (w4196 & w6530);
assign w4199 = ~w4087 & w4195;
assign w4200 = ~w4196 & w4199;
assign w4201 = ~w4198 & ~w4200;
assign w4202 = ~w4094 & w4171;
assign w4203 = w4171 & w6450;
assign w4204 = ~w3571 & w3591;
assign w4205 = w4204 & ~w4008;
assign w4206 = ~w4095 & w4205;
assign w4207 = ~w1576 & w3911;
assign w4208 = (w3971 & w7152) | (w3971 & w7153) | (w7152 & w7153);
assign w4209 = (~w4207 & w3971) | (~w4207 & w7154) | (w3971 & w7154);
assign w4210 = w4063 & w4209;
assign w4211 = ~w4208 & ~w4210;
assign w4212 = ~w4206 & w4211;
assign w4213 = ~w4202 & ~w4212;
assign w4214 = ~w4203 & ~w4213;
assign w4215 = ~w1648 & w3591;
assign w4216 = ~w4106 & ~w4168;
assign w4217 = (w4215 & w4216) | (w4215 & w6451) | (w4216 & w6451);
assign w4218 = ~w4216 & w6452;
assign w4219 = ~w4217 & ~w4218;
assign w4220 = w1572 & w3594;
assign w4221 = w4112 & w4165;
assign w4222 = (w4220 & w4221) | (w4220 & w6453) | (w4221 & w6453);
assign w4223 = ~w4221 & w6454;
assign w4224 = ~w4222 & ~w4223;
assign w4225 = w1570 & w3733;
assign w4226 = (~w4120 & ~w4162) | (~w4120 & w6243) | (~w4162 & w6243);
assign w4227 = w4225 & ~w4226;
assign w4228 = ~w4225 & w4226;
assign w4229 = ~w4227 & ~w4228;
assign w4230 = w1568 & w3597;
assign w4231 = (w4230 & w4161) | (w4230 & w6244) | (w4161 & w6244);
assign w4232 = ~w4161 & w6245;
assign w4233 = ~w4231 & ~w4232;
assign w4234 = w1566 & w3600;
assign w4235 = (~w4127 & ~w4129) | (~w4127 & w6246) | (~w4129 & w6246);
assign w4236 = w4234 & w4235;
assign w4237 = ~w4234 & ~w4235;
assign w4238 = ~w4236 & ~w4237;
assign w4239 = w1563 & w3603;
assign w4240 = ~w4134 & w4147;
assign w4241 = ~w4133 & ~w4240;
assign w4242 = ~w4239 & ~w4241;
assign w4243 = w4239 & w4241;
assign w4244 = ~w4242 & ~w4243;
assign w4245 = w1774 & ~w3549;
assign w4246 = ~w1556 & ~w4137;
assign w4247 = w3526 & ~w4246;
assign w4248 = (~w4247 & ~w3528) | (~w4247 & w7155) | (~w3528 & w7155);
assign w4249 = w4245 & ~w4248;
assign w4250 = (w4248 & w3549) | (w4248 & w7156) | (w3549 & w7156);
assign w4251 = ~w4249 & ~w4250;
assign w4252 = (~w4141 & w4144) | (~w4141 & w6247) | (w4144 & w6247);
assign w4253 = w3544 & w4252;
assign w4254 = (w1561 & w3544) | (w1561 & w6248) | (w3544 & w6248);
assign w4255 = ~w4253 & w4254;
assign w4256 = w4251 & ~w4255;
assign w4257 = ~w4251 & w4255;
assign w4258 = ~w4256 & ~w4257;
assign w4259 = w4244 & ~w4258;
assign w4260 = ~w4244 & w4258;
assign w4261 = ~w4259 & ~w4260;
assign w4262 = w4238 & w4261;
assign w4263 = ~w4238 & ~w4261;
assign w4264 = ~w4262 & ~w4263;
assign w4265 = w4233 & w4264;
assign w4266 = ~w4233 & ~w4264;
assign w4267 = ~w4265 & ~w4266;
assign w4268 = ~w4229 & ~w4267;
assign w4269 = w4229 & w4267;
assign w4270 = ~w4268 & ~w4269;
assign w4271 = w4224 & w4270;
assign w4272 = ~w4224 & ~w4270;
assign w4273 = ~w4271 & ~w4272;
assign w4274 = w4219 & w4273;
assign w4275 = ~w4219 & ~w4273;
assign w4276 = ~w4274 & ~w4275;
assign w4277 = w4214 & w4276;
assign w4278 = ~w4214 & ~w4276;
assign w4279 = ~w4277 & ~w4278;
assign w4280 = w4201 & ~w4279;
assign w4281 = ~w4201 & w4279;
assign w4282 = ~w4280 & ~w4281;
assign w4283 = w4194 & ~w4282;
assign w4284 = ~w4194 & w4282;
assign w4285 = ~w4283 & ~w4284;
assign w4286 = (~w4178 & ~w4180) | (~w4178 & w6531) | (~w4180 & w6531);
assign w4287 = ~w4285 & w4286;
assign w4288 = w4285 & ~w4286;
assign w4289 = ~w4287 & ~w4288;
assign w4290 = ~w4193 & w4289;
assign w4291 = ~w4290 & w7157;
assign w4292 = (w3586 & w4290) | (w3586 & w7158) | (w4290 & w7158);
assign w4293 = ~w4291 & ~w4292;
assign w4294 = ~w4283 & w4286;
assign w4295 = ~w1579 & w3588;
assign w4296 = ~w1579 & w7512;
assign w4297 = ~w4294 & w4296;
assign w4298 = (~w4295 & w4294) | (~w4295 & w7159) | (w4294 & w7159);
assign w4299 = ~w4297 & ~w4298;
assign w4300 = ~w4200 & ~w4279;
assign w4301 = (~w4198 & w4279) | (~w4198 & w6532) | (w4279 & w6532);
assign w4302 = w1590 & w4075;
assign w4303 = ~w4198 & w7491;
assign w4304 = (~w4302 & w4300) | (~w4302 & w6455) | (w4300 & w6455);
assign w4305 = ~w4303 & ~w4304;
assign w4306 = ~w1576 & w3985;
assign w4307 = (~w4206 & ~w6450) | (~w4206 & w7161) | (~w6450 & w7161);
assign w4308 = (w4306 & w4203) | (w4306 & w6533) | (w4203 & w6533);
assign w4309 = ~w4202 & ~w4211;
assign w4310 = (w4306 & w4202) | (w4306 & w6456) | (w4202 & w6456);
assign w4311 = w4276 & w4310;
assign w4312 = ~w4308 & ~w4311;
assign w4313 = w4276 & ~w4309;
assign w4314 = ~w4203 & w6534;
assign w4315 = ~w4313 & w4314;
assign w4316 = w4312 & ~w4315;
assign w4317 = ~w1648 & w3911;
assign w4318 = ~w4217 & ~w4273;
assign w4319 = (~w4317 & w4318) | (~w4317 & w6535) | (w4318 & w6535);
assign w4320 = ~w4318 & w6536;
assign w4321 = ~w4319 & ~w4320;
assign w4322 = w1570 & w3594;
assign w4323 = (~w4322 & w4226) | (~w4322 & w7162) | (w4226 & w7162);
assign w4324 = ~w4269 & w4323;
assign w4325 = w1570 & w7513;
assign w4326 = (w4325 & w4267) | (w4325 & w7163) | (w4267 & w7163);
assign w4327 = ~w4324 & ~w4326;
assign w4328 = w1563 & w3600;
assign w4329 = ~w4243 & w4258;
assign w4330 = ~w4329 & w6249;
assign w4331 = (~w4328 & w4329) | (~w4328 & w6250) | (w4329 & w6250);
assign w4332 = ~w4330 & ~w4331;
assign w4333 = w1566 & w3597;
assign w4334 = ~w4251 & ~w4253;
assign w4335 = w4254 & ~w4334;
assign w4336 = w1561 & w3603;
assign w4337 = ~w4335 & ~w4336;
assign w4338 = w3603 & w4335;
assign w4339 = w3549 & w6251;
assign w4340 = (~w4135 & w3528) | (~w4135 & w7164) | (w3528 & w7164);
assign w4341 = w1556 & w3610;
assign w4342 = (~w4341 & w3549) | (~w4341 & w6252) | (w3549 & w6252);
assign w4343 = ~w4339 & w4342;
assign w4344 = w3544 & w4249;
assign w4345 = ~w3544 & ~w4249;
assign w4346 = (w1774 & ~w3544) | (w1774 & w6253) | (~w3544 & w6253);
assign w4347 = ~w4345 & w4346;
assign w4348 = w4343 & ~w4347;
assign w4349 = ~w4343 & w4347;
assign w4350 = ~w4348 & ~w4349;
assign w4351 = ~w4337 & w6254;
assign w4352 = (w4350 & w4337) | (w4350 & w6255) | (w4337 & w6255);
assign w4353 = ~w4351 & ~w4352;
assign w4354 = w4333 & w4353;
assign w4355 = w4332 & w4354;
assign w4356 = w4333 & ~w4353;
assign w4357 = ~w4332 & w4356;
assign w4358 = ~w4355 & ~w4357;
assign w4359 = ~w4333 & w4353;
assign w4360 = ~w4332 & w4359;
assign w4361 = ~w4333 & ~w4353;
assign w4362 = w4332 & w4361;
assign w4363 = ~w4360 & ~w4362;
assign w4364 = w4358 & w4363;
assign w4365 = w1568 & w3733;
assign w4366 = ~w4236 & ~w4261;
assign w4367 = ~w4237 & ~w4366;
assign w4368 = (~w4365 & w4366) | (~w4365 & w6457) | (w4366 & w6457);
assign w4369 = ~w4364 & w4368;
assign w4370 = w4363 & w4367;
assign w4371 = w4358 & ~w4365;
assign w4372 = w4370 & w4371;
assign w4373 = ~w4369 & ~w4372;
assign w4374 = ~w4366 & w6458;
assign w4375 = ~w4364 & w4374;
assign w4376 = w4358 & ~w4367;
assign w4377 = w4363 & w4365;
assign w4378 = w4376 & w4377;
assign w4379 = ~w4375 & ~w4378;
assign w4380 = w4373 & w4379;
assign w4381 = ~w4231 & ~w4265;
assign w4382 = w4380 & ~w4381;
assign w4383 = ~w4380 & w4381;
assign w4384 = ~w4382 & ~w4383;
assign w4385 = w4327 & w4384;
assign w4386 = ~w4327 & ~w4384;
assign w4387 = ~w4385 & ~w4386;
assign w4388 = w1572 & w3591;
assign w4389 = (~w4223 & w4270) | (~w4223 & w6459) | (w4270 & w6459);
assign w4390 = w4388 & w4389;
assign w4391 = ~w4388 & ~w4389;
assign w4392 = ~w4390 & ~w4391;
assign w4393 = w4387 & w4392;
assign w4394 = ~w4387 & ~w4392;
assign w4395 = ~w4393 & ~w4394;
assign w4396 = w4321 & ~w4395;
assign w4397 = ~w4321 & w4395;
assign w4398 = ~w4396 & ~w4397;
assign w4399 = ~w4316 & w4398;
assign w4400 = w4316 & ~w4398;
assign w4401 = ~w4399 & ~w4400;
assign w4402 = w4305 & ~w4401;
assign w4403 = ~w4305 & w4401;
assign w4404 = ~w4402 & ~w4403;
assign w4405 = w4299 & ~w4404;
assign w4406 = ~w4299 & w4404;
assign w4407 = ~w4405 & ~w4406;
assign w4408 = w4293 & ~w4407;
assign w4409 = ~w4293 & w4407;
assign w4410 = ~w4408 & ~w4409;
assign w4411 = w3582 & ~w4410;
assign w4412 = ~w3582 & w4410;
assign w4413 = ~w4411 & ~w4412;
assign w4414 = w1012 & w3585;
assign w4415 = w1012 & w3588;
assign w4416 = ~w4079 & w4190;
assign w4417 = w4185 & ~w4416;
assign w4418 = ~w4185 & w4416;
assign w4419 = ~w4417 & ~w4418;
assign w4420 = w4415 & ~w4419;
assign w4421 = ~w4415 & w4419;
assign w4422 = w1012 & w4075;
assign w4423 = ~w3991 & ~w4077;
assign w4424 = ~w4072 & w4423;
assign w4425 = w4072 & ~w4423;
assign w4426 = ~w4424 & ~w4425;
assign w4427 = w4422 & ~w4426;
assign w4428 = ~w4422 & w4426;
assign w4429 = w1012 & w3985;
assign w4430 = ~w3914 & w7165;
assign w4431 = (w3982 & w3914) | (w3982 & w7166) | (w3914 & w7166);
assign w4432 = ~w4430 & ~w4431;
assign w4433 = w4429 & ~w4432;
assign w4434 = ~w4429 & w4432;
assign w4435 = ~w3902 & ~w3904;
assign w4436 = w3906 & ~w4435;
assign w4437 = ~w3906 & w4435;
assign w4438 = ~w3895 & ~w3896;
assign w4439 = ~w3900 & w4438;
assign w4440 = w3900 & ~w4438;
assign w4441 = ~w4439 & ~w4440;
assign w4442 = w3875 & ~w3877;
assign w4443 = ~w3878 & ~w4442;
assign w4444 = w3600 & ~w4443;
assign w4445 = ~w3869 & ~w3871;
assign w4446 = ~w3872 & ~w4445;
assign w4447 = w3603 & w4446;
assign w4448 = ~w3549 & w7167;
assign w4449 = (w3610 & ~w3549) | (w3610 & w6256) | (~w3549 & w6256);
assign w4450 = (~w1584 & w3528) | (~w1584 & w7168) | (w3528 & w7168);
assign w4451 = w4449 & w4450;
assign w4452 = ~w4448 & ~w4451;
assign w4453 = w3544 & ~w4452;
assign w4454 = ~w3544 & w4452;
assign w4455 = ~w3862 & ~w3865;
assign w4456 = ~w3866 & ~w4455;
assign w4457 = ~w4454 & w4456;
assign w4458 = ~w4453 & ~w4457;
assign w4459 = (~w4458 & w4446) | (~w4458 & w7169) | (w4446 & w7169);
assign w4460 = ~w4447 & ~w4459;
assign w4461 = (~w4460 & ~w4443) | (~w4460 & w7170) | (~w4443 & w7170);
assign w4462 = ~w4444 & ~w4461;
assign w4463 = w3597 & ~w4462;
assign w4464 = ~w3597 & w4462;
assign w4465 = ~w3882 & ~w3884;
assign w4466 = ~w3885 & ~w4465;
assign w4467 = ~w4464 & w4466;
assign w4468 = ~w4467 & w7171;
assign w4469 = ~w3887 & ~w3889;
assign w4470 = ~w3893 & ~w4469;
assign w4471 = w3893 & w4469;
assign w4472 = ~w4468 & ~w4470;
assign w4473 = ~w4471 & w4472;
assign w4474 = w3594 & w4441;
assign w4475 = (w3733 & w4467) | (w3733 & w7172) | (w4467 & w7172);
assign w4476 = ~w4473 & ~w4475;
assign w4477 = ~w4474 & w4476;
assign w4478 = (w3591 & w4441) | (w3591 & w7173) | (w4441 & w7173);
assign w4479 = ~w4477 & w4478;
assign w4480 = ~w4436 & ~w4437;
assign w4481 = ~w4479 & w4480;
assign w4482 = ~w3852 & ~w3909;
assign w4483 = ~w3907 & w4482;
assign w4484 = w3907 & ~w4482;
assign w4485 = ~w4483 & ~w4484;
assign w4486 = ~w3591 & ~w3594;
assign w4487 = ~w4474 & w7174;
assign w4488 = (w1012 & w4441) | (w1012 & w7175) | (w4441 & w7175);
assign w4489 = ~w4487 & w4488;
assign w4490 = ~w4481 & w4489;
assign w4491 = (w4490 & w4485) | (w4490 & w7176) | (w4485 & w7176);
assign w4492 = w1012 & w3911;
assign w4493 = w4485 & w4492;
assign w4494 = ~w4491 & ~w4493;
assign w4495 = ~w4434 & ~w4494;
assign w4496 = ~w4433 & ~w4495;
assign w4497 = ~w4428 & ~w4496;
assign w4498 = ~w4427 & ~w4497;
assign w4499 = ~w4421 & ~w4498;
assign w4500 = (w4414 & w4499) | (w4414 & w7177) | (w4499 & w7177);
assign w4501 = ~w4499 & w7178;
assign w4502 = ~w4191 & ~w4193;
assign w4503 = ~w4289 & ~w4502;
assign w4504 = w4289 & w4502;
assign w4505 = ~w4503 & ~w4504;
assign w4506 = ~w4501 & w4505;
assign w4507 = ~w4500 & ~w4506;
assign w4508 = w4413 & w4507;
assign w4509 = ~w4413 & ~w4507;
assign w4510 = ~w4508 & ~w4509;
assign w4511 = ~w4297 & w4404;
assign w4512 = ~w4298 & ~w4511;
assign w4513 = ~w4304 & w4401;
assign w4514 = (~w4301 & ~w4401) | (~w4301 & w7179) | (~w4401 & w7179);
assign w4515 = (w3588 & w4401) | (w3588 & w6537) | (w4401 & w6537);
assign w4516 = ~w4514 & w4515;
assign w4517 = w1590 & w3588;
assign w4518 = ~w4303 & ~w4517;
assign w4519 = ~w4513 & w4518;
assign w4520 = ~w4516 & ~w4519;
assign w4521 = ~w1576 & w4075;
assign w4522 = w4312 & w4398;
assign w4523 = (~w4521 & w4522) | (~w4521 & w7180) | (w4522 & w7180);
assign w4524 = ~w3576 & w4306;
assign w4525 = ~w4522 & w4524;
assign w4526 = (w4307 & ~w4276) | (w4307 & w7181) | (~w4276 & w7181);
assign w4527 = w4521 & ~w4526;
assign w4528 = ~w4398 & w4527;
assign w4529 = ~w4525 & ~w4528;
assign w4530 = ~w4523 & w4529;
assign w4531 = ~w4319 & w4395;
assign w4532 = ~w1648 & w3985;
assign w4533 = ~w4320 & ~w4532;
assign w4534 = ~w4531 & w4533;
assign w4535 = w3911 & w7182;
assign w4536 = w4395 & w4535;
assign w4537 = w4387 & ~w4391;
assign w4538 = (~w3911 & ~w4389) | (~w3911 & w7183) | (~w4389 & w7183);
assign w4539 = w4387 & w7184;
assign w4540 = ~w3911 & ~w4387;
assign w4541 = ~w4392 & w4540;
assign w4542 = ~w4318 & w7185;
assign w4543 = ~w4541 & w7186;
assign w4544 = ~w4536 & ~w4543;
assign w4545 = ~w4534 & w4544;
assign w4546 = w1572 & w3911;
assign w4547 = (~w4390 & ~w4387) | (~w4390 & w6460) | (~w4387 & w6460);
assign w4548 = w4546 & ~w4547;
assign w4549 = (~w4546 & ~w4389) | (~w4546 & w7187) | (~w4389 & w7187);
assign w4550 = (w4549 & ~w4387) | (w4549 & w7188) | (~w4387 & w7188);
assign w4551 = ~w4548 & ~w4550;
assign w4552 = w1570 & w3591;
assign w4553 = (w4552 & w4269) | (w4552 & w7189) | (w4269 & w7189);
assign w4554 = (w4553 & w4384) | (w4553 & w7190) | (w4384 & w7190);
assign w4555 = ~w4326 & ~w4552;
assign w4556 = ~w4385 & w4555;
assign w4557 = ~w4554 & ~w4556;
assign w4558 = w1568 & w3594;
assign w4559 = w4379 & w4381;
assign w4560 = w4373 & ~w4559;
assign w4561 = w1566 & w3733;
assign w4562 = w4358 & ~w4561;
assign w4563 = ~w4370 & w4562;
assign w4564 = w4363 & w4561;
assign w4565 = ~w4376 & w4564;
assign w4566 = ~w4563 & ~w4565;
assign w4567 = w1561 & w3600;
assign w4568 = (~w4338 & w4337) | (~w4338 & w6254) | (w4337 & w6254);
assign w4569 = ~w4567 & w4568;
assign w4570 = w4567 & ~w4568;
assign w4571 = ~w4569 & ~w4570;
assign w4572 = w1563 & w3597;
assign w4573 = w1774 & ~w4343;
assign w4574 = ~w4344 & ~w4573;
assign w4575 = ~w4345 & ~w4574;
assign w4576 = w3603 & w4575;
assign w4577 = w1774 & w3603;
assign w4578 = ~w4575 & ~w4577;
assign w4579 = ~w1556 & w4449;
assign w4580 = ~w3544 & w4579;
assign w4581 = (w3549 & w7191) | (w3549 & w7192) | (w7191 & w7192);
assign w4582 = w3544 & w4581;
assign w4583 = ~w4580 & ~w4582;
assign w4584 = w3549 & w4583;
assign w4585 = ~w3549 & ~w4583;
assign w4586 = ~w4584 & ~w4585;
assign w4587 = ~w4578 & w4738;
assign w4588 = (w4586 & w4578) | (w4586 & w6257) | (w4578 & w6257);
assign w4589 = ~w4587 & ~w4588;
assign w4590 = ~w4572 & ~w4589;
assign w4591 = w4571 & w4590;
assign w4592 = ~w4572 & w4589;
assign w4593 = ~w4571 & w4592;
assign w4594 = ~w4591 & ~w4593;
assign w4595 = w4572 & ~w4589;
assign w4596 = ~w4571 & w4595;
assign w4597 = w4572 & w4589;
assign w4598 = w4571 & w4597;
assign w4599 = ~w4596 & ~w4598;
assign w4600 = w4594 & w4599;
assign w4601 = ~w4330 & w4353;
assign w4602 = ~w4331 & ~w4601;
assign w4603 = w4600 & ~w4602;
assign w4604 = ~w4600 & w4602;
assign w4605 = ~w4603 & ~w4604;
assign w4606 = w4566 & ~w4605;
assign w4607 = ~w4566 & w4605;
assign w4608 = ~w4606 & ~w4607;
assign w4609 = w4560 & w4608;
assign w4610 = ~w4560 & ~w4608;
assign w4611 = ~w4609 & ~w4610;
assign w4612 = w4558 & w4611;
assign w4613 = ~w4558 & ~w4611;
assign w4614 = ~w4612 & ~w4613;
assign w4615 = w4557 & w4614;
assign w4616 = ~w4557 & ~w4614;
assign w4617 = ~w4615 & ~w4616;
assign w4618 = w4551 & ~w4617;
assign w4619 = ~w4551 & w4617;
assign w4620 = ~w4618 & ~w4619;
assign w4621 = w4545 & ~w4620;
assign w4622 = ~w4545 & w4620;
assign w4623 = ~w4621 & ~w4622;
assign w4624 = ~w4530 & w4623;
assign w4625 = w4530 & ~w4623;
assign w4626 = ~w4624 & ~w4625;
assign w4627 = w4520 & ~w4626;
assign w4628 = ~w4520 & w4626;
assign w4629 = ~w4627 & ~w4628;
assign w4630 = ~w4512 & ~w4629;
assign w4631 = w4512 & w4629;
assign w4632 = ~w4630 & ~w4631;
assign w4633 = ~w1579 & w3585;
assign w4634 = ~w3580 & w7193;
assign w4635 = (~w4634 & ~w3585) | (~w4634 & w7194) | (~w3585 & w7194);
assign w4636 = ~w4632 & w4635;
assign w4637 = w3585 & w7195;
assign w4638 = w4632 & w4637;
assign w4639 = ~w4636 & ~w4638;
assign w4640 = w4632 & w4633;
assign w4641 = (w4634 & w4632) | (w4634 & w6538) | (w4632 & w6538);
assign w4642 = ~w4640 & w4641;
assign w4643 = w4639 & ~w4642;
assign w4644 = ~w4291 & w4407;
assign w4645 = ~w4292 & ~w4644;
assign w4646 = ~w4643 & w4645;
assign w4647 = w4643 & ~w4645;
assign w4648 = ~w4646 & ~w4647;
assign w4649 = ~w4412 & ~w4507;
assign w4650 = ~w4411 & ~w4649;
assign w4651 = ~w4648 & w4650;
assign w4652 = w4648 & ~w4650;
assign w4653 = ~w4651 & ~w4652;
assign w4654 = ~w3582 & ~w4653;
assign w4655 = w3582 & w4653;
assign w4656 = ~w4654 & ~w4655;
assign w4657 = w3582 & ~w4651;
assign w4658 = ~w3582 & ~w4652;
assign w4659 = ~w4657 & ~w4658;
assign w4660 = w4639 & ~w4645;
assign w4661 = ~w4642 & ~w4660;
assign w4662 = ~w3580 & w7196;
assign w4663 = ~w4629 & w6539;
assign w4664 = (~w4633 & ~w4629) | (~w4633 & w6540) | (~w4629 & w6540);
assign w4665 = ~w4663 & ~w4664;
assign w4666 = (w4662 & w4629) | (w4662 & w6541) | (w4629 & w6541);
assign w4667 = w4665 & ~w4666;
assign w4668 = w1590 & w3585;
assign w4669 = ~w4516 & ~w4668;
assign w4670 = ~w4627 & w4669;
assign w4671 = w4516 & w4668;
assign w4672 = (w4668 & w4513) | (w4668 & w7197) | (w4513 & w7197);
assign w4673 = ~w4626 & w4672;
assign w4674 = ~w4671 & ~w4673;
assign w4675 = ~w4670 & w4674;
assign w4676 = ~w1576 & w3588;
assign w4677 = w4523 & ~w4676;
assign w4678 = (~w4677 & ~w6542) | (~w4677 & w7198) | (~w6542 & w7198);
assign w4679 = w4529 & ~w4623;
assign w4680 = ~w4523 & w4676;
assign w4681 = ~w4679 & w4680;
assign w4682 = w4678 & ~w4681;
assign w4683 = w1572 & w3985;
assign w4684 = (w4683 & w4537) | (w4683 & w6461) | (w4537 & w6461);
assign w4685 = ~w4547 & w7199;
assign w4686 = (~w4685 & ~w4617) | (~w4685 & w7200) | (~w4617 & w7200);
assign w4687 = (~w4683 & w4547) | (~w4683 & w7201) | (w4547 & w7201);
assign w4688 = (w4687 & ~w4617) | (w4687 & w7202) | (~w4617 & w7202);
assign w4689 = w4686 & ~w4688;
assign w4690 = w1570 & w3911;
assign w4691 = w4554 & w4690;
assign w4692 = (w4690 & w4385) | (w4690 & w6462) | (w4385 & w6462);
assign w4693 = (~w4691 & ~w4614) | (~w4691 & w7203) | (~w4614 & w7203);
assign w4694 = ~w4554 & ~w4690;
assign w4695 = ~w4615 & w4694;
assign w4696 = w4693 & ~w4695;
assign w4697 = ~w4558 & ~w4609;
assign w4698 = w1568 & w3591;
assign w4699 = ~w4610 & w4698;
assign w4700 = ~w4697 & w4699;
assign w4701 = w4558 & ~w4610;
assign w4702 = ~w4609 & ~w4698;
assign w4703 = ~w4701 & w4702;
assign w4704 = ~w4700 & ~w4703;
assign w4705 = w3594 & w4565;
assign w4706 = w1566 & w3594;
assign w4707 = ~w4563 & w4706;
assign w4708 = ~w4605 & w4707;
assign w4709 = ~w4705 & ~w4708;
assign w4710 = ~w4565 & ~w4706;
assign w4711 = ~w4606 & w4710;
assign w4712 = w4709 & ~w4711;
assign w4713 = w4599 & ~w4602;
assign w4714 = w4594 & ~w4713;
assign w4715 = w1563 & w3733;
assign w4716 = ~w4569 & ~w4589;
assign w4717 = ~w4570 & ~w4716;
assign w4718 = (w3549 & ~w3544) | (w3549 & w6258) | (~w3544 & w6258);
assign w4719 = (~w4579 & ~w3544) | (~w4579 & w6543) | (~w3544 & w6543);
assign w4720 = ~w4718 & ~w4719;
assign w4721 = ~w1556 & ~w3469;
assign w4722 = w3454 & w4721;
assign w4723 = ~w1556 & w3469;
assign w4724 = ~w3454 & w4723;
assign w4725 = ~w4722 & ~w4724;
assign w4726 = w3549 & w7204;
assign w4727 = ~w3544 & ~w4726;
assign w4728 = w4725 & ~w4727;
assign w4729 = ~w4725 & w4727;
assign w4730 = ~w4728 & ~w4729;
assign w4731 = w4720 & ~w4730;
assign w4732 = ~w4720 & w4730;
assign w4733 = ~w4731 & ~w4732;
assign w4734 = w1774 & w3600;
assign w4735 = ~w4733 & ~w4734;
assign w4736 = w4733 & w4734;
assign w4737 = ~w4735 & ~w4736;
assign w4738 = ~w4576 & ~w4586;
assign w4739 = ~w4578 & ~w4738;
assign w4740 = w1561 & w3597;
assign w4741 = ~w4739 & w4740;
assign w4742 = w4739 & ~w4740;
assign w4743 = ~w4741 & ~w4742;
assign w4744 = w4737 & w4743;
assign w4745 = ~w4737 & ~w4743;
assign w4746 = ~w4744 & ~w4745;
assign w4747 = ~w4717 & w4746;
assign w4748 = w4717 & ~w4746;
assign w4749 = ~w4747 & ~w4748;
assign w4750 = w4715 & ~w4749;
assign w4751 = ~w4715 & w4749;
assign w4752 = ~w4750 & ~w4751;
assign w4753 = w4714 & w4752;
assign w4754 = ~w4714 & ~w4752;
assign w4755 = ~w4753 & ~w4754;
assign w4756 = ~w4712 & ~w4755;
assign w4757 = w4712 & w4755;
assign w4758 = ~w4756 & ~w4757;
assign w4759 = ~w4704 & w4758;
assign w4760 = w4704 & ~w4758;
assign w4761 = ~w4759 & ~w4760;
assign w4762 = ~w4696 & w4761;
assign w4763 = w4696 & ~w4761;
assign w4764 = ~w4762 & ~w4763;
assign w4765 = w4689 & w4764;
assign w4766 = ~w4689 & ~w4764;
assign w4767 = ~w4765 & ~w4766;
assign w4768 = ~w1648 & w4075;
assign w4769 = ~w4544 & w4768;
assign w4770 = (w4768 & w4531) | (w4768 & w7205) | (w4531 & w7205);
assign w4771 = ~w4620 & w4770;
assign w4772 = ~w4769 & ~w4771;
assign w4773 = w4544 & ~w4768;
assign w4774 = ~w4621 & w4773;
assign w4775 = w4772 & ~w4774;
assign w4776 = w4767 & w4775;
assign w4777 = ~w4767 & ~w4775;
assign w4778 = ~w4776 & ~w4777;
assign w4779 = ~w4682 & w4778;
assign w4780 = w4682 & ~w4778;
assign w4781 = ~w4779 & ~w4780;
assign w4782 = ~w4675 & w4781;
assign w4783 = w4675 & ~w4781;
assign w4784 = ~w4782 & ~w4783;
assign w4785 = ~w4667 & w4784;
assign w4786 = w4667 & ~w4784;
assign w4787 = ~w4785 & ~w4786;
assign w4788 = w4661 & w4787;
assign w4789 = ~w4661 & ~w4787;
assign w4790 = ~w4788 & ~w4789;
assign w4791 = ~w4634 & w4790;
assign w4792 = w4634 & ~w4790;
assign w4793 = ~w4791 & ~w4792;
assign w4794 = w4659 & ~w4793;
assign w4795 = ~w4659 & w4793;
assign w4796 = ~w4794 & ~w4795;
assign w4797 = ~w4657 & w4793;
assign w4798 = (w3581 & w4652) | (w3581 & w7206) | (w4652 & w7206);
assign w4799 = (w4798 & ~w4793) | (w4798 & w7207) | (~w4793 & w7207);
assign w4800 = (~w4658 & ~w4793) | (~w4658 & w6544) | (~w4793 & w6544);
assign w4801 = ~w4799 & w4800;
assign w4802 = w4634 & ~w4788;
assign w4803 = (~w4634 & w4661) | (~w4634 & w6545) | (w4661 & w6545);
assign w4804 = ~w4802 & ~w4803;
assign w4805 = ~w4662 & ~w4784;
assign w4806 = ~w4664 & w4666;
assign w4807 = ~w4784 & ~w4806;
assign w4808 = ~w3581 & w4665;
assign w4809 = ~w4807 & ~w4808;
assign w4810 = ~w4805 & ~w4809;
assign w4811 = ~w3580 & w7208;
assign w4812 = (w6463 & w6546) | (w6463 & w6547) | (w6546 & w6547);
assign w4813 = (~w6463 & w6548) | (~w6463 & w6549) | (w6548 & w6549);
assign w4814 = ~w4812 & ~w4813;
assign w4815 = w4678 & w4778;
assign w4816 = ~w1576 & w3585;
assign w4817 = (~w4816 & w4679) | (~w4816 & w7209) | (w4679 & w7209);
assign w4818 = (w4817 & ~w4778) | (w4817 & w7210) | (~w4778 & w7210);
assign w4819 = (~w4681 & ~w4778) | (~w4681 & w6550) | (~w4778 & w6550);
assign w4820 = (w3585 & w4815) | (w3585 & w6464) | (w4815 & w6464);
assign w4821 = ~w4818 & ~w4820;
assign w4822 = ~w1648 & w3588;
assign w4823 = w4767 & ~w4774;
assign w4824 = (w4822 & w4823) | (w4822 & w6465) | (w4823 & w6465);
assign w4825 = ~w4823 & w6466;
assign w4826 = ~w4824 & ~w4825;
assign w4827 = w4686 & ~w4764;
assign w4828 = w4075 & ~w4688;
assign w4829 = (w4828 & w4764) | (w4828 & w7211) | (w4764 & w7211);
assign w4830 = w1572 & w4075;
assign w4831 = w4686 & ~w4830;
assign w4832 = (w4831 & ~w4764) | (w4831 & w7212) | (~w4764 & w7212);
assign w4833 = ~w4829 & ~w4832;
assign w4834 = ~w4700 & ~w4758;
assign w4835 = w3911 & ~w4703;
assign w4836 = ~w4834 & w4835;
assign w4837 = ~w4703 & w4758;
assign w4838 = w1568 & w3911;
assign w4839 = ~w4700 & ~w4838;
assign w4840 = ~w4837 & w4839;
assign w4841 = ~w4836 & ~w4840;
assign w4842 = w1566 & w3591;
assign w4843 = ~w4708 & w7213;
assign w4844 = ~w4757 & w4843;
assign w4845 = w3594 & w7214;
assign w4846 = ~w4563 & w4845;
assign w4847 = ~w4605 & w4846;
assign w4848 = w4565 & w7215;
assign w4849 = ~w4847 & ~w4848;
assign w4850 = ~w4755 & w4849;
assign w4851 = (w4842 & w4606) | (w4842 & w6467) | (w4606 & w6467);
assign w4852 = (w4851 & w4755) | (w4851 & w6468) | (w4755 & w6468);
assign w4853 = ~w4844 & ~w4852;
assign w4854 = ~w4714 & ~w4750;
assign w4855 = ~w4854 & w6259;
assign w4856 = w1563 & w3594;
assign w4857 = (~w4856 & w4854) | (~w4856 & w6260) | (w4854 & w6260);
assign w4858 = ~w4855 & ~w4857;
assign w4859 = w1561 & w3733;
assign w4860 = ~w4740 & w4746;
assign w4861 = ~w4748 & ~w4860;
assign w4862 = w4859 & w4861;
assign w4863 = ~w4859 & ~w4861;
assign w4864 = ~w4862 & ~w4863;
assign w4865 = w3544 & ~w4725;
assign w4866 = (~w4865 & w4730) | (~w4865 & w6551) | (w4730 & w6551);
assign w4867 = ~w1086 & w3603;
assign w4868 = w3603 & w6552;
assign w4869 = w4866 & ~w4868;
assign w4870 = ~w1556 & w3600;
assign w4871 = ~w4867 & ~w4870;
assign w4872 = w4869 & ~w4871;
assign w4873 = w1774 & w3597;
assign w4874 = w4872 & w4873;
assign w4875 = (~w4868 & w4870) | (~w4868 & w6553) | (w4870 & w6553);
assign w4876 = w3597 & w6554;
assign w4877 = ~w4875 & w4876;
assign w4878 = ~w4874 & ~w4877;
assign w4879 = (~w4866 & w4871) | (~w4866 & w6261) | (w4871 & w6261);
assign w4880 = ~w4872 & ~w4873;
assign w4881 = ~w4879 & w4880;
assign w4882 = w4878 & ~w4881;
assign w4883 = ~w4736 & ~w4739;
assign w4884 = ~w4735 & ~w4883;
assign w4885 = ~w4882 & w4884;
assign w4886 = w4882 & ~w4884;
assign w4887 = ~w4885 & ~w4886;
assign w4888 = w4864 & w4887;
assign w4889 = ~w4864 & ~w4887;
assign w4890 = ~w4888 & ~w4889;
assign w4891 = w4858 & ~w4890;
assign w4892 = ~w4858 & w4890;
assign w4893 = ~w4891 & ~w4892;
assign w4894 = w4853 & ~w4893;
assign w4895 = ~w4853 & w4893;
assign w4896 = ~w4894 & ~w4895;
assign w4897 = ~w4841 & ~w4896;
assign w4898 = w4841 & w4896;
assign w4899 = ~w4897 & ~w4898;
assign w4900 = w1570 & w3985;
assign w4901 = w4693 & w4761;
assign w4902 = (~w4900 & w4901) | (~w4900 & w6469) | (w4901 & w6469);
assign w4903 = ~w4901 & w6470;
assign w4904 = ~w4902 & ~w4903;
assign w4905 = w4899 & ~w4904;
assign w4906 = ~w4899 & w4904;
assign w4907 = ~w4905 & ~w4906;
assign w4908 = w4833 & ~w4907;
assign w4909 = ~w4833 & w4907;
assign w4910 = ~w4908 & ~w4909;
assign w4911 = w4826 & ~w4910;
assign w4912 = ~w4826 & w4910;
assign w4913 = ~w4911 & ~w4912;
assign w4914 = w4821 & ~w4913;
assign w4915 = ~w4821 & w4913;
assign w4916 = ~w4914 & ~w4915;
assign w4917 = w4814 & ~w4916;
assign w4918 = ~w4814 & w4916;
assign w4919 = ~w4917 & ~w4918;
assign w4920 = w4810 & w4919;
assign w4921 = ~w4810 & ~w4919;
assign w4922 = ~w4920 & ~w4921;
assign w4923 = w4804 & ~w4922;
assign w4924 = ~w4804 & w4922;
assign w4925 = ~w4923 & ~w4924;
assign w4926 = ~w4801 & w4925;
assign w4927 = w4801 & ~w4925;
assign w4928 = ~w4926 & ~w4927;
assign w4929 = w4800 & ~w4925;
assign w4930 = w3580 & w7216;
assign w4931 = (~w2513 & w3515) | (~w2513 & w7217) | (w3515 & w7217);
assign w4932 = ~w3580 & ~w4931;
assign w4933 = ~w4930 & ~w4932;
assign w4934 = (w4933 & w4929) | (w4933 & w7218) | (w4929 & w7218);
assign w4935 = w1012 & w4933;
assign w4936 = (~w4935 & w4797) | (~w4935 & w6555) | (w4797 & w6555);
assign w4937 = ~w4929 & w4936;
assign w4938 = ~w4934 & ~w4937;
assign w4939 = w4665 & ~w4807;
assign w4940 = w4919 & w4939;
assign w4941 = ~w4662 & ~w4940;
assign w4942 = w4807 & ~w4919;
assign w4943 = (w3581 & w4919) | (w3581 & w7219) | (w4919 & w7219);
assign w4944 = ~w4941 & ~w4943;
assign w4945 = ~w3580 & w7220;
assign w4946 = ~w4945 & ~w4820;
assign w4947 = (w4946 & ~w4913) | (w4946 & w7221) | (~w4913 & w7221);
assign w4948 = (w3581 & w4815) | (w3581 & w6471) | (w4815 & w6471);
assign w4949 = w3581 & ~w4819;
assign w4950 = (~w4949 & ~w4913) | (~w4949 & w7222) | (~w4913 & w7222);
assign w4951 = ~w4947 & w4950;
assign w4952 = ~w1648 & w3585;
assign w4953 = ~w4824 & w7514;
assign w4954 = (~w6472 & w7224) | (~w6472 & w7225) | (w7224 & w7225);
assign w4955 = ~w4953 & ~w4954;
assign w4956 = ~w4832 & w4907;
assign w4957 = w1572 & w3588;
assign w4958 = (~w4957 & w4827) | (~w4957 & w6556) | (w4827 & w6556);
assign w4959 = ~w4956 & w4958;
assign w4960 = (w4764 & w7226) | (w4764 & w7227) | (w7226 & w7227);
assign w4961 = w4907 & w4960;
assign w4962 = ~w4827 & w6557;
assign w4963 = ~w4961 & ~w4962;
assign w4964 = ~w4959 & w4963;
assign w4965 = w4899 & ~w4903;
assign w4966 = w1570 & w4075;
assign w4967 = w4966 & ~w4902;
assign w4968 = ~w4965 & w4967;
assign w4969 = ~w4899 & ~w4902;
assign w4970 = (~w4966 & w4901) | (~w4966 & w6558) | (w4901 & w6558);
assign w4971 = ~w4969 & w4970;
assign w4972 = ~w4968 & ~w4971;
assign w4973 = w1568 & w3985;
assign w4974 = w4840 & ~w4973;
assign w4975 = ~w4836 & ~w4973;
assign w4976 = w4896 & w4975;
assign w4977 = ~w4974 & ~w4976;
assign w4978 = w3985 & ~w4840;
assign w4979 = ~w4898 & w4978;
assign w4980 = w4977 & ~w4979;
assign w4981 = ~w4852 & ~w4893;
assign w4982 = w1566 & w3911;
assign w4983 = (w4982 & w4757) | (w4982 & w6474) | (w4757 & w6474);
assign w4984 = ~w4981 & w4983;
assign w4985 = ~w4757 & w6475;
assign w4986 = (~w4982 & w4850) | (~w4982 & w6262) | (w4850 & w6262);
assign w4987 = ~w4893 & w4986;
assign w4988 = ~w4985 & ~w4987;
assign w4989 = ~w4984 & w4988;
assign w4990 = w1561 & w3594;
assign w4991 = ~w1774 & w3733;
assign w4992 = w4880 & w6559;
assign w4993 = ~w4884 & ~w4991;
assign w4994 = w4878 & w4993;
assign w4995 = ~w4992 & ~w4994;
assign w4996 = (~w3206 & ~w3600) | (~w3206 & w6263) | (~w3600 & w6263);
assign w4997 = ~w1556 & w3597;
assign w4998 = w4996 & ~w4997;
assign w4999 = ~w4996 & w4997;
assign w5000 = ~w4998 & ~w4999;
assign w5001 = ~w4869 & ~w4871;
assign w5002 = w3733 & w5001;
assign w5003 = ~w5000 & w5002;
assign w5004 = w3733 & ~w5001;
assign w5005 = w5000 & w5004;
assign w5006 = ~w5003 & ~w5005;
assign w5007 = ~w3733 & w5001;
assign w5008 = w5000 & w5007;
assign w5009 = ~w3733 & ~w5001;
assign w5010 = ~w5000 & w5009;
assign w5011 = ~w5008 & ~w5010;
assign w5012 = w5006 & w5011;
assign w5013 = w4995 & ~w5012;
assign w5014 = ~w4995 & w5012;
assign w5015 = ~w5013 & ~w5014;
assign w5016 = w4990 & ~w5015;
assign w5017 = ~w4990 & w5015;
assign w5018 = ~w5016 & ~w5017;
assign w5019 = ~w4863 & ~w4887;
assign w5020 = ~w4862 & ~w5019;
assign w5021 = w5018 & ~w5020;
assign w5022 = ~w5018 & w5020;
assign w5023 = ~w5021 & ~w5022;
assign w5024 = ~w4855 & w4890;
assign w5025 = (~w4854 & w7228) | (~w4854 & w7229) | (w7228 & w7229);
assign w5026 = (w5025 & ~w4890) | (w5025 & w7230) | (~w4890 & w7230);
assign w5027 = w1563 & w3591;
assign w5028 = (~w5027 & w4854) | (~w5027 & w7231) | (w4854 & w7231);
assign w5029 = (w5028 & w4890) | (w5028 & w7232) | (w4890 & w7232);
assign w5030 = ~w5026 & ~w5029;
assign w5031 = w5023 & w5030;
assign w5032 = ~w5023 & ~w5030;
assign w5033 = ~w5031 & ~w5032;
assign w5034 = ~w4989 & w5033;
assign w5035 = w4989 & ~w5033;
assign w5036 = ~w5034 & ~w5035;
assign w5037 = ~w4980 & w5036;
assign w5038 = w4980 & ~w5036;
assign w5039 = ~w5037 & ~w5038;
assign w5040 = w4972 & ~w5039;
assign w5041 = ~w4972 & w5039;
assign w5042 = ~w5040 & ~w5041;
assign w5043 = ~w4964 & w5042;
assign w5044 = w4964 & ~w5042;
assign w5045 = ~w5043 & ~w5044;
assign w5046 = ~w4955 & w5045;
assign w5047 = w4955 & ~w5045;
assign w5048 = ~w5046 & ~w5047;
assign w5049 = w4951 & w5048;
assign w5050 = ~w4951 & ~w5048;
assign w5051 = ~w5049 & ~w5050;
assign w5052 = ~w4916 & w6560;
assign w5053 = w4674 & w7492;
assign w5054 = w4916 & w5053;
assign w5055 = ~w5052 & ~w5054;
assign w5056 = w5051 & w5055;
assign w5057 = ~w5051 & ~w5055;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = w4944 & ~w5058;
assign w5060 = ~w4944 & w5058;
assign w5061 = ~w5059 & ~w5060;
assign w5062 = ~w4803 & w4922;
assign w5063 = ~w4802 & ~w5062;
assign w5064 = (w4634 & w5062) | (w4634 & w6561) | (w5062 & w6561);
assign w5065 = ~w4634 & ~w5062;
assign w5066 = ~w5064 & ~w5065;
assign w5067 = w5061 & ~w5066;
assign w5068 = ~w5061 & w5066;
assign w5069 = ~w5067 & ~w5068;
assign w5070 = w4938 & w5069;
assign w5071 = ~w4938 & ~w5069;
assign w5072 = ~w5070 & ~w5071;
assign w5073 = ~w4937 & w5069;
assign w5074 = ~w4934 & ~w5073;
assign w5075 = ~w5061 & ~w5063;
assign w5076 = ~w1584 & w4933;
assign w5077 = (~w4634 & ~w4933) | (~w4634 & w7234) | (~w4933 & w7234);
assign w5078 = ~w5075 & w5077;
assign w5079 = ~w5062 & w6562;
assign w5080 = w5061 & ~w5079;
assign w5081 = (w5076 & w5062) | (w5076 & w6563) | (w5062 & w6563);
assign w5082 = ~w5061 & ~w5081;
assign w5083 = ~w5080 & ~w5082;
assign w5084 = ~w5078 & ~w5083;
assign w5085 = (~w4813 & w4916) | (~w4813 & w6564) | (w4916 & w6564);
assign w5086 = w5051 & w5085;
assign w5087 = ~w5051 & ~w5085;
assign w5088 = ~w5086 & ~w5087;
assign w5089 = ~w3581 & ~w5088;
assign w5090 = ~w4941 & ~w5089;
assign w5091 = (w1579 & w4807) | (w1579 & w7235) | (w4807 & w7235);
assign w5092 = ~w4942 & ~w5091;
assign w5093 = ~w5058 & ~w5092;
assign w5094 = w3581 & ~w5093;
assign w5095 = w5090 & ~w5094;
assign w5096 = ~w5055 & ~w5088;
assign w5097 = w3581 & w5049;
assign w5098 = ~w3581 & ~w4947;
assign w5099 = ~w5049 & w5098;
assign w5100 = ~w5097 & ~w5099;
assign w5101 = ~w3580 & w7236;
assign w5102 = (~w5101 & w6565) | (~w5101 & w7493) | (w6565 & w7493);
assign w5103 = (w5102 & w5045) | (w5102 & w7439) | (w5045 & w7439);
assign w5104 = ~w5045 & w7237;
assign w5105 = ~w5103 & ~w5104;
assign w5106 = ~w4959 & ~w5042;
assign w5107 = (w3585 & w5106) | (w3585 & w6566) | (w5106 & w6566);
assign w5108 = w1572 & w3585;
assign w5109 = ~w4961 & w6567;
assign w5110 = ~w5106 & w5109;
assign w5111 = ~w5107 & ~w5110;
assign w5112 = w1570 & w3588;
assign w5113 = (~w4968 & ~w5039) | (~w4968 & w6476) | (~w5039 & w6476);
assign w5114 = ~w5112 & w5113;
assign w5115 = w5112 & ~w5113;
assign w5116 = ~w5114 & ~w5115;
assign w5117 = w4977 & ~w5036;
assign w5118 = w1568 & w4075;
assign w5119 = ~w5117 & w6477;
assign w5120 = (w4075 & w5117) | (w4075 & w6478) | (w5117 & w6478);
assign w5121 = ~w5119 & ~w5120;
assign w5122 = ~w4984 & ~w5033;
assign w5123 = w1566 & w3985;
assign w5124 = ~w4987 & w7238;
assign w5125 = ~w5122 & w5124;
assign w5126 = (~w6264 & w7239) | (~w6264 & w7240) | (w7239 & w7240);
assign w5127 = ~w5125 & ~w5126;
assign w5128 = ~w5016 & ~w5021;
assign w5129 = w1561 & w3591;
assign w5130 = ~w4881 & w5011;
assign w5131 = ~w4886 & w5130;
assign w5132 = ~w1774 & w3594;
assign w5133 = (~w5132 & w5006) | (~w5132 & w6568) | (w5006 & w6568);
assign w5134 = ~w5131 & w5133;
assign w5135 = ~w1086 & w3597;
assign w5136 = w2513 & w3600;
assign w5137 = ~w5135 & ~w5136;
assign w5138 = w3557 & w6569;
assign w5139 = w3562 & w5138;
assign w5140 = (~w1556 & ~w3557) | (~w1556 & w6570) | (~w3557 & w6570);
assign w5141 = ~w3562 & w5140;
assign w5142 = ~w5139 & ~w5141;
assign w5143 = w5137 & ~w5142;
assign w5144 = ~w5137 & w5142;
assign w5145 = ~w5143 & ~w5144;
assign w5146 = ~w4999 & ~w5001;
assign w5147 = ~w4998 & ~w5146;
assign w5148 = ~w5145 & ~w5147;
assign w5149 = w5145 & w5147;
assign w5150 = ~w5148 & ~w5149;
assign w5151 = w3594 & ~w5150;
assign w5152 = ~w3594 & w5150;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = w5134 & w5153;
assign w5155 = ~w5134 & ~w5153;
assign w5156 = ~w5154 & ~w5155;
assign w5157 = w5129 & ~w5156;
assign w5158 = ~w5129 & w5156;
assign w5159 = ~w5157 & ~w5158;
assign w5160 = w5128 & ~w5159;
assign w5161 = ~w5128 & w5159;
assign w5162 = ~w5160 & ~w5161;
assign w5163 = w5023 & ~w5029;
assign w5164 = w1563 & w3911;
assign w5165 = (~w5164 & w5024) | (~w5164 & w6265) | (w5024 & w6265);
assign w5166 = ~w5163 & w5165;
assign w5167 = ~w5024 & w6266;
assign w5168 = w3911 & w5023;
assign w5169 = ~w5029 & w5168;
assign w5170 = ~w5167 & ~w5169;
assign w5171 = w5170 & w5285;
assign w5172 = (~w5162 & ~w5170) | (~w5162 & w7241) | (~w5170 & w7241);
assign w5173 = ~w5171 & ~w5172;
assign w5174 = w5127 & ~w5173;
assign w5175 = ~w5127 & w5173;
assign w5176 = ~w5174 & ~w5175;
assign w5177 = w5121 & ~w5176;
assign w5178 = ~w5121 & w5176;
assign w5179 = ~w5177 & ~w5178;
assign w5180 = w5116 & ~w5179;
assign w5181 = ~w5116 & w5179;
assign w5182 = ~w5180 & ~w5181;
assign w5183 = w5111 & ~w5182;
assign w5184 = ~w5111 & w5182;
assign w5185 = ~w5183 & ~w5184;
assign w5186 = ~w5105 & w5185;
assign w5187 = w5105 & ~w5185;
assign w5188 = ~w5186 & ~w5187;
assign w5189 = w5100 & ~w5188;
assign w5190 = ~w5100 & w5188;
assign w5191 = ~w5189 & ~w5190;
assign w5192 = w5096 & w5191;
assign w5193 = ~w5096 & ~w5191;
assign w5194 = ~w5192 & ~w5193;
assign w5195 = ~w5095 & w5194;
assign w5196 = w5095 & ~w5194;
assign w5197 = ~w5195 & ~w5196;
assign w5198 = w5084 & w5197;
assign w5199 = ~w5084 & ~w5197;
assign w5200 = ~w5198 & ~w5199;
assign w5201 = ~w5074 & ~w5200;
assign w5202 = w5074 & w5200;
assign w5203 = ~w5201 & ~w5202;
assign w5204 = ~w5076 & ~w5084;
assign w5205 = ~w3581 & ~w5075;
assign w5206 = w5061 & w5063;
assign w5207 = w5076 & ~w5206;
assign w5208 = ~w5205 & w5207;
assign w5209 = w5197 & ~w5208;
assign w5210 = ~w5204 & ~w5209;
assign w5211 = (w5090 & w5194) | (w5090 & w6571) | (w5194 & w6571);
assign w5212 = w4933 & w5211;
assign w5213 = ~w1579 & w4933;
assign w5214 = ~w5211 & ~w5213;
assign w5215 = ~w5212 & ~w5214;
assign w5216 = (w4811 & ~w5189) | (w4811 & w7242) | (~w5189 & w7242);
assign w5217 = (~w5216 & w5192) | (~w5216 & w7243) | (w5192 & w7243);
assign w5218 = w5097 & ~w5188;
assign w5219 = w5099 & w5188;
assign w5220 = ~w5218 & ~w5219;
assign w5221 = (w5101 & w5045) | (w5101 & w7244) | (w5045 & w7244);
assign w5222 = (~w5221 & w5105) | (~w5221 & w6572) | (w5105 & w6572);
assign w5223 = ~w5110 & ~w5182;
assign w5224 = (w3581 & w5106) | (w3581 & w6573) | (w5106 & w6573);
assign w5225 = ~w5107 & ~w5224;
assign w5226 = ~w5223 & w5225;
assign w5227 = (w3581 & w5106) | (w3581 & w7245) | (w5106 & w7245);
assign w5228 = (~w5227 & w5182) | (~w5227 & w7440) | (w5182 & w7440);
assign w5229 = ~w5226 & w5228;
assign w5230 = w1570 & w3585;
assign w5231 = ~w5114 & w5179;
assign w5232 = (w5230 & w5231) | (w5230 & w6574) | (w5231 & w6574);
assign w5233 = ~w5231 & w6575;
assign w5234 = ~w5232 & ~w5233;
assign w5235 = w1568 & w3588;
assign w5236 = ~w5120 & w5176;
assign w5237 = (~w6479 & w7246) | (~w6479 & w7247) | (w7246 & w7247);
assign w5238 = (w3588 & w5117) | (w3588 & w7441) | (w5117 & w7441);
assign w5239 = ~w5236 & w5238;
assign w5240 = ~w5237 & ~w5239;
assign w5241 = ~w5125 & ~w5173;
assign w5242 = ~w5126 & ~w5241;
assign w5243 = w1566 & w4075;
assign w5244 = (~w5243 & w5241) | (~w5243 & w6267) | (w5241 & w6267);
assign w5245 = ~w5241 & w6268;
assign w5246 = ~w5244 & ~w5245;
assign w5247 = ~w5157 & ~w5161;
assign w5248 = w1774 & w3594;
assign w5249 = ~w5131 & w6269;
assign w5250 = (~w5150 & w5131) | (~w5150 & w7442) | (w5131 & w7442);
assign w5251 = w1774 & w3591;
assign w5252 = ~w5251 & w7494;
assign w5253 = ~w5250 & w5252;
assign w5254 = w3591 & ~w5150;
assign w5255 = ~w5249 & w5254;
assign w5256 = (w5131 & w7215) | (w5131 & w7443) | (w7215 & w7443);
assign w5257 = ~w5255 & ~w5256;
assign w5258 = ~w5253 & w5257;
assign w5259 = w1561 & w3911;
assign w5260 = ~w5142 & ~w5148;
assign w5261 = w4997 & ~w5146;
assign w5262 = (~w5261 & w5148) | (~w5261 & w7248) | (w5148 & w7248);
assign w5263 = w2513 & w3597;
assign w5264 = (~w5263 & ~w3733) | (~w5263 & w6271) | (~w3733 & w6271);
assign w5265 = ~w1556 & w3594;
assign w5266 = w5264 & ~w5265;
assign w5267 = ~w5264 & w5265;
assign w5268 = ~w5266 & ~w5267;
assign w5269 = w5262 & ~w5268;
assign w5270 = ~w5262 & w5268;
assign w5271 = ~w5269 & ~w5270;
assign w5272 = w5259 & ~w5271;
assign w5273 = ~w5259 & w5271;
assign w5274 = ~w5272 & ~w5273;
assign w5275 = w5258 & w5274;
assign w5276 = ~w5258 & ~w5274;
assign w5277 = ~w5275 & ~w5276;
assign w5278 = ~w5247 & ~w5277;
assign w5279 = w5247 & w5277;
assign w5280 = ~w5278 & ~w5279;
assign w5281 = (w3985 & w5169) | (w3985 & w6272) | (w5169 & w6272);
assign w5282 = w3985 & w5162;
assign w5283 = ~w5166 & w5282;
assign w5284 = ~w5281 & ~w5283;
assign w5285 = w5162 & ~w5166;
assign w5286 = w1563 & w3985;
assign w5287 = ~w5169 & w6273;
assign w5288 = ~w5285 & w5287;
assign w5289 = (w5280 & ~w5284) | (w5280 & w7249) | (~w5284 & w7249);
assign w5290 = w5284 & w7250;
assign w5291 = ~w5289 & ~w5290;
assign w5292 = w5246 & w5291;
assign w5293 = ~w5246 & ~w5291;
assign w5294 = ~w5292 & ~w5293;
assign w5295 = w5240 & ~w5294;
assign w5296 = ~w5240 & w5294;
assign w5297 = ~w5295 & ~w5296;
assign w5298 = w5234 & ~w5297;
assign w5299 = ~w5234 & w5297;
assign w5300 = ~w5298 & ~w5299;
assign w5301 = ~w5229 & ~w5300;
assign w5302 = w5229 & w5300;
assign w5303 = ~w5301 & ~w5302;
assign w5304 = ~w5222 & ~w5303;
assign w5305 = w5222 & w5303;
assign w5306 = ~w5304 & ~w5305;
assign w5307 = w5101 & ~w5306;
assign w5308 = ~w5101 & w5306;
assign w5309 = ~w5307 & ~w5308;
assign w5310 = ~w5220 & ~w5309;
assign w5311 = w5220 & w5309;
assign w5312 = ~w5310 & ~w5311;
assign w5313 = ~w5217 & w5312;
assign w5314 = w5217 & ~w5312;
assign w5315 = ~w5313 & ~w5314;
assign w5316 = w5215 & ~w5315;
assign w5317 = ~w5215 & w5315;
assign w5318 = ~w5316 & ~w5317;
assign w5319 = w5210 & w5318;
assign w5320 = ~w5210 & ~w5318;
assign w5321 = ~w5319 & ~w5320;
assign w5322 = w5201 & ~w5321;
assign w5323 = ~w5201 & w5321;
assign w5324 = ~w5322 & ~w5323;
assign w5325 = ~w4933 & ~w5216;
assign w5326 = w1590 & w4933;
assign w5327 = (w5326 & w5192) | (w5326 & w7251) | (w5192 & w7251);
assign w5328 = (w5327 & w5312) | (w5327 & w7444) | (w5312 & w7444);
assign w5329 = (w1590 & w5312) | (w1590 & w6480) | (w5312 & w6480);
assign w5330 = ~w5328 & w5329;
assign w5331 = (~w5101 & w5303) | (~w5101 & w7252) | (w5303 & w7252);
assign w5332 = (w5101 & ~w5303) | (w5101 & w7253) | (~w5303 & w7253);
assign w5333 = ~w5331 & ~w5332;
assign w5334 = w5229 & w6576;
assign w5335 = (~w3581 & w5223) | (~w3581 & w7254) | (w5223 & w7254);
assign w5336 = (w5335 & ~w5229) | (w5335 & w7255) | (~w5229 & w7255);
assign w5337 = ~w5334 & ~w5336;
assign w5338 = ~w5233 & w5297;
assign w5339 = ~w3580 & w7256;
assign w5340 = (~w5339 & w6481) | (~w5339 & w7495) | (w6481 & w7495);
assign w5341 = ~w5338 & w5340;
assign w5342 = (w5339 & w5297) | (w5339 & w6482) | (w5297 & w6482);
assign w5343 = ~w5341 & ~w5342;
assign w5344 = ~w5239 & w5294;
assign w5345 = ~w5237 & ~w5344;
assign w5346 = ~w5344 & w6483;
assign w5347 = w1568 & w3585;
assign w5348 = (~w5347 & w5344) | (~w5347 & w6484) | (w5344 & w6484);
assign w5349 = ~w5346 & ~w5348;
assign w5350 = ~w5245 & w5291;
assign w5351 = ~w5244 & ~w5350;
assign w5352 = w1566 & w3588;
assign w5353 = w5280 & ~w5288;
assign w5354 = w1563 & w4075;
assign w5355 = ~w5283 & w6274;
assign w5356 = ~w5353 & w5355;
assign w5357 = (w4075 & w5283) | (w4075 & w6275) | (w5283 & w6275);
assign w5358 = w4075 & w5280;
assign w5359 = ~w5288 & w5358;
assign w5360 = ~w5357 & ~w5359;
assign w5361 = w5259 & w5277;
assign w5362 = ~w5278 & ~w5361;
assign w5363 = w1561 & w3985;
assign w5364 = ~w5253 & w5271;
assign w5365 = w5257 & ~w5364;
assign w5366 = ~w1774 & w3911;
assign w5367 = ~w5364 & w6485;
assign w5368 = ~w1556 & w3591;
assign w5369 = ~w1086 & w3594;
assign w5370 = w2513 & w3733;
assign w5371 = ~w5369 & ~w5370;
assign w5372 = w5368 & ~w5371;
assign w5373 = ~w5368 & w5371;
assign w5374 = ~w5372 & ~w5373;
assign w5375 = (w5265 & w5261) | (w5265 & w5267) | (w5261 & w5267);
assign w5376 = ~w5260 & ~w5375;
assign w5377 = w5374 & ~w5376;
assign w5378 = ~w5374 & w5376;
assign w5379 = ~w5377 & ~w5378;
assign w5380 = ~w3911 & ~w5379;
assign w5381 = w3911 & w5379;
assign w5382 = ~w5380 & ~w5381;
assign w5383 = ~w5367 & w5382;
assign w5384 = w5367 & ~w5382;
assign w5385 = ~w5383 & ~w5384;
assign w5386 = w5363 & w5385;
assign w5387 = ~w5363 & ~w5385;
assign w5388 = ~w5386 & ~w5387;
assign w5389 = w5362 & ~w5388;
assign w5390 = ~w5362 & w5388;
assign w5391 = ~w5389 & ~w5390;
assign w5392 = w5360 & w5457;
assign w5393 = (~w5391 & ~w5360) | (~w5391 & w7257) | (~w5360 & w7257);
assign w5394 = ~w5392 & ~w5393;
assign w5395 = ~w5352 & w5394;
assign w5396 = w5352 & ~w5394;
assign w5397 = ~w5395 & ~w5396;
assign w5398 = w5351 & w5397;
assign w5399 = ~w5351 & ~w5397;
assign w5400 = ~w5398 & ~w5399;
assign w5401 = ~w5349 & w5400;
assign w5402 = w5349 & ~w5400;
assign w5403 = ~w5401 & ~w5402;
assign w5404 = ~w5343 & w5403;
assign w5405 = w5343 & ~w5403;
assign w5406 = ~w5404 & ~w5405;
assign w5407 = w5337 & w5406;
assign w5408 = ~w5337 & ~w5406;
assign w5409 = ~w5407 & ~w5408;
assign w5410 = w5333 & ~w5409;
assign w5411 = ~w5333 & w5409;
assign w5412 = ~w5410 & ~w5411;
assign w5413 = (~w4948 & w5309) | (~w4948 & w6486) | (w5309 & w6486);
assign w5414 = ~w5306 & w6487;
assign w5415 = (w4948 & w5188) | (w4948 & w7258) | (w5188 & w7258);
assign w5416 = (w4815 & w7259) | (w4815 & w7260) | (w7259 & w7260);
assign w5417 = (~w5415 & ~w5306) | (~w5415 & w7261) | (~w5306 & w7261);
assign w5418 = ~w5414 & w5417;
assign w5419 = ~w5413 & w5436;
assign w5420 = (~w5412 & w5413) | (~w5412 & w7262) | (w5413 & w7262);
assign w5421 = ~w5419 & ~w5420;
assign w5422 = ~w5328 & w7263;
assign w5423 = (w5421 & w5328) | (w5421 & w7264) | (w5328 & w7264);
assign w5424 = ~w5422 & ~w5423;
assign w5425 = (~w5212 & w5315) | (~w5212 & w7265) | (w5315 & w7265);
assign w5426 = ~w5424 & w5425;
assign w5427 = w5424 & ~w5425;
assign w5428 = ~w5426 & ~w5427;
assign w5429 = ~w5201 & ~w5319;
assign w5430 = ~w5320 & ~w5429;
assign w5431 = w5428 & w5430;
assign w5432 = ~w5428 & ~w5430;
assign w5433 = ~w5431 & ~w5432;
assign w5434 = (~w5427 & w5429) | (~w5427 & w6488) | (w5429 & w6488);
assign w5435 = (~w5328 & ~w5330) | (~w5328 & w6489) | (~w5330 & w6489);
assign w5436 = w5412 & w5418;
assign w5437 = ~w1576 & w4933;
assign w5438 = (~w5437 & w5436) | (~w5437 & w6490) | (w5436 & w6490);
assign w5439 = ~w5436 & w6491;
assign w5440 = ~w5438 & ~w5439;
assign w5441 = ~w5331 & ~w5410;
assign w5442 = (~w5339 & w5338) | (~w5339 & w6492) | (w5338 & w6492);
assign w5443 = w5403 & w5442;
assign w5444 = ~w6482 & w7266;
assign w5445 = ~w5403 & w5444;
assign w5446 = ~w5443 & ~w5445;
assign w5447 = w5397 & w6276;
assign w5448 = ~w5351 & w5395;
assign w5449 = w5242 & ~w5291;
assign w5450 = w4075 & w7267;
assign w5451 = ~w5350 & w5450;
assign w5452 = ~w5394 & ~w5449;
assign w5453 = ~w5451 & w5452;
assign w5454 = ~w5448 & ~w5453;
assign w5455 = ~w5447 & w5454;
assign w5456 = (~w3579 & w5359) | (~w3579 & w7268) | (w5359 & w7268);
assign w5457 = ~w5356 & w5391;
assign w5458 = ~w5356 & w6493;
assign w5459 = ~w5456 & ~w5458;
assign w5460 = w1563 & w3588;
assign w5461 = ~w5359 & w7269;
assign w5462 = ~w5457 & w5461;
assign w5463 = w5459 & ~w5462;
assign w5464 = w1566 & w3585;
assign w5465 = (w5379 & w7270) | (w5379 & w7271) | (w7270 & w7271);
assign w5466 = (~w5465 & w5365) | (~w5465 & w7272) | (w5365 & w7272);
assign w5467 = (~w5379 & w5365) | (~w5379 & w7273) | (w5365 & w7273);
assign w5468 = w1774 & w3911;
assign w5469 = ~w5364 & w7274;
assign w5470 = w3985 & ~w5469;
assign w5471 = ~w5467 & w5470;
assign w5472 = w1561 & w4075;
assign w5473 = ~w1556 & w3911;
assign w5474 = (~w4486 & w5260) | (~w4486 & w7275) | (w5260 & w7275);
assign w5475 = ~w1086 & w3591;
assign w5476 = w2513 & w3594;
assign w5477 = ~w5475 & ~w5476;
assign w5478 = ~w5474 & w6494;
assign w5479 = (~w5477 & w5474) | (~w5477 & w7276) | (w5474 & w7276);
assign w5480 = ~w5478 & ~w5479;
assign w5481 = w5473 & ~w5480;
assign w5482 = ~w5473 & w5480;
assign w5483 = ~w5481 & ~w5482;
assign w5484 = w5472 & w5483;
assign w5485 = ~w5472 & ~w5483;
assign w5486 = ~w5484 & ~w5485;
assign w5487 = ~w5471 & w7277;
assign w5488 = (~w5486 & w5471) | (~w5486 & w7278) | (w5471 & w7278);
assign w5489 = ~w5487 & ~w5488;
assign w5490 = (~w5387 & ~w5362) | (~w5387 & w7279) | (~w5362 & w7279);
assign w5491 = ~w5489 & w5490;
assign w5492 = w5489 & ~w5490;
assign w5493 = ~w5491 & ~w5492;
assign w5494 = w5464 & w5493;
assign w5495 = ~w5464 & ~w5493;
assign w5496 = ~w5494 & ~w5495;
assign w5497 = w5463 & w5496;
assign w5498 = ~w5463 & ~w5496;
assign w5499 = ~w5497 & ~w5498;
assign w5500 = w5455 & w5499;
assign w5501 = ~w5455 & ~w5499;
assign w5502 = ~w5500 & ~w5501;
assign w5503 = ~w5348 & ~w5400;
assign w5504 = ~w3580 & w7280;
assign w5505 = ~w5346 & ~w5504;
assign w5506 = ~w5503 & w5505;
assign w5507 = ~w5345 & w5400;
assign w5508 = w3581 & ~w5348;
assign w5509 = ~w5507 & w5508;
assign w5510 = ~w5506 & ~w5509;
assign w5511 = w5502 & ~w5510;
assign w5512 = ~w5502 & w5510;
assign w5513 = ~w5511 & ~w5512;
assign w5514 = w5446 & ~w5513;
assign w5515 = ~w5446 & w5513;
assign w5516 = ~w5514 & ~w5515;
assign w5517 = ~w5334 & w5406;
assign w5518 = ~w5336 & ~w5406;
assign w5519 = ~w5517 & ~w5518;
assign w5520 = w5516 & w5519;
assign w5521 = ~w5516 & ~w5519;
assign w5522 = ~w5520 & ~w5521;
assign w5523 = w5101 & ~w5522;
assign w5524 = ~w5101 & w5522;
assign w5525 = ~w5523 & ~w5524;
assign w5526 = w5441 & ~w5525;
assign w5527 = ~w5441 & w5525;
assign w5528 = ~w5526 & ~w5527;
assign w5529 = w5440 & ~w5528;
assign w5530 = ~w5440 & w5528;
assign w5531 = ~w5529 & ~w5530;
assign w5532 = ~w5435 & w5531;
assign w5533 = w5435 & ~w5531;
assign w5534 = ~w5532 & ~w5533;
assign w5535 = ~w5426 & w5534;
assign w5536 = ~w5434 & w5535;
assign w5537 = ~w5427 & ~w5534;
assign w5538 = ~w5431 & w5537;
assign w5539 = ~w5536 & ~w5538;
assign w5540 = ~w5516 & w5519;
assign w5541 = ~w5224 & ~w5540;
assign w5542 = w5224 & ~w5520;
assign w5543 = ~w5541 & ~w5542;
assign w5544 = ~w1648 & w4933;
assign w5545 = w5445 & w5513;
assign w5546 = w5443 & ~w5513;
assign w5547 = ~w5545 & ~w5546;
assign w5548 = w5502 & ~w5506;
assign w5549 = ~w5508 & ~w5548;
assign w5550 = w5502 & w5504;
assign w5551 = ~w5509 & ~w5550;
assign w5552 = ~w5549 & w5551;
assign w5553 = w5464 & ~w5499;
assign w5554 = w1563 & w3585;
assign w5555 = w5462 & ~w5554;
assign w5556 = ~w5493 & ~w5554;
assign w5557 = w5459 & w5556;
assign w5558 = ~w5555 & ~w5557;
assign w5559 = ~w5458 & w7281;
assign w5560 = w3585 & ~w5462;
assign w5561 = ~w5559 & w5560;
assign w5562 = w5472 & w5489;
assign w5563 = ~w5491 & ~w5562;
assign w5564 = (~w5365 & w7282) | (~w5365 & w7283) | (w7282 & w7283);
assign w5565 = ~w1774 & w4075;
assign w5566 = ~w5471 & w7284;
assign w5567 = w1561 & w3588;
assign w5568 = (w4075 & ~w3588) | (w4075 & w7285) | (~w3588 & w7285);
assign w5569 = w2513 & w3591;
assign w5570 = ~w1086 & w3911;
assign w5571 = ~w5569 & ~w5570;
assign w5572 = (w5473 & w5474) | (w5473 & w7286) | (w5474 & w7286);
assign w5573 = ~w5479 & ~w5572;
assign w5574 = ~w1556 & w3985;
assign w5575 = ~w5573 & w5574;
assign w5576 = w5573 & ~w5574;
assign w5577 = ~w5575 & ~w5576;
assign w5578 = w5571 & w5577;
assign w5579 = ~w5571 & ~w5577;
assign w5580 = ~w5578 & ~w5579;
assign w5581 = w5568 & ~w5580;
assign w5582 = ~w5568 & w5580;
assign w5583 = ~w5581 & ~w5582;
assign w5584 = w5566 & w5583;
assign w5585 = ~w5566 & ~w5583;
assign w5586 = ~w5584 & ~w5585;
assign w5587 = ~w5491 & w7287;
assign w5588 = (w5586 & w5491) | (w5586 & w7288) | (w5491 & w7288);
assign w5589 = ~w5587 & ~w5588;
assign w5590 = ~w3580 & w7289;
assign w5591 = w5589 & w5590;
assign w5592 = ~w5589 & ~w5590;
assign w5593 = ~w5591 & ~w5592;
assign w5594 = w5558 & w7290;
assign w5595 = (~w5593 & ~w5558) | (~w5593 & w7291) | (~w5558 & w7291);
assign w5596 = ~w5594 & ~w5595;
assign w5597 = (~w6495 & w7292) | (~w6495 & w7293) | (w7292 & w7293);
assign w5598 = (w6495 & w7294) | (w6495 & w7295) | (w7294 & w7295);
assign w5599 = ~w5597 & ~w5598;
assign w5600 = ~w5552 & w5599;
assign w5601 = w5552 & ~w5599;
assign w5602 = ~w5600 & ~w5601;
assign w5603 = w5547 & ~w5602;
assign w5604 = ~w5547 & w5602;
assign w5605 = ~w5603 & ~w5604;
assign w5606 = w5544 & ~w5605;
assign w5607 = w5543 & ~w5606;
assign w5608 = w5544 & w5605;
assign w5609 = ~w5543 & ~w5608;
assign w5610 = ~w5607 & ~w5609;
assign w5611 = ~w5544 & w5605;
assign w5612 = w5543 & w5611;
assign w5613 = ~w5544 & ~w5605;
assign w5614 = ~w5543 & w5613;
assign w5615 = ~w5612 & ~w5614;
assign w5616 = ~w5610 & w5615;
assign w5617 = w5441 & ~w5524;
assign w5618 = ~w5523 & ~w5617;
assign w5619 = ~w5616 & w5618;
assign w5620 = w5616 & ~w5618;
assign w5621 = ~w5619 & ~w5620;
assign w5622 = (~w5439 & w5528) | (~w5439 & w6496) | (w5528 & w6496);
assign w5623 = w5621 & ~w5622;
assign w5624 = ~w5621 & w5622;
assign w5625 = ~w5623 & ~w5624;
assign w5626 = ~w5536 & w7296;
assign w5627 = (w5625 & w5536) | (w5625 & w7297) | (w5536 & w7297);
assign w5628 = ~w5626 & ~w5627;
assign w5629 = ~w5610 & w5618;
assign w5630 = w5615 & ~w5629;
assign w5631 = ~w5542 & ~w5605;
assign w5632 = (w4933 & w5540) | (w4933 & w7298) | (w5540 & w7298);
assign w5633 = ~w5631 & w5632;
assign w5634 = w1572 & w4933;
assign w5635 = ~w5605 & ~w5634;
assign w5636 = ~w5540 & w7299;
assign w5637 = (~w5636 & ~w5635) | (~w5636 & w7300) | (~w5635 & w7300);
assign w5638 = w5545 & ~w5602;
assign w5639 = w5546 & w5602;
assign w5640 = ~w5638 & ~w5639;
assign w5641 = ~w5590 & w5596;
assign w5642 = ~w5598 & ~w5641;
assign w5643 = w3581 & ~w5586;
assign w5644 = w5563 & w5643;
assign w5645 = w3581 & w5586;
assign w5646 = ~w5563 & w5645;
assign w5647 = ~w5644 & ~w5646;
assign w5648 = ~w5555 & ~w5647;
assign w5649 = ~w5557 & w5648;
assign w5650 = w3581 & ~w5462;
assign w5651 = ~w5559 & w5650;
assign w5652 = ~w5649 & ~w5651;
assign w5653 = ~w5557 & w7301;
assign w5654 = ~w3580 & w7302;
assign w5655 = ~w5561 & ~w5654;
assign w5656 = ~w5653 & w5655;
assign w5657 = w5652 & ~w5656;
assign w5658 = w1561 & w3585;
assign w5659 = w1774 & w4075;
assign w5660 = ~w5471 & w7303;
assign w5661 = ~w5580 & ~w5660;
assign w5662 = (w4075 & w5471) | (w4075 & w7304) | (w5471 & w7304);
assign w5663 = (w3588 & w5661) | (w3588 & w7305) | (w5661 & w7305);
assign w5664 = w1774 & w3588;
assign w5665 = ~w5662 & ~w5664;
assign w5666 = ~w5661 & w5665;
assign w5667 = ~w1556 & w4075;
assign w5668 = ~w3985 & ~w5572;
assign w5669 = (w5577 & w7308) | (w5577 & w7309) | (w7308 & w7309);
assign w5670 = w5667 & w7496;
assign w5671 = ~w5669 & ~w5670;
assign w5672 = ~w5666 & w5671;
assign w5673 = (~w5658 & w5672) | (~w5658 & w7310) | (w5672 & w7310);
assign w5674 = w5658 & ~w5671;
assign w5675 = ~w5666 & w5674;
assign w5676 = ~w5663 & w5675;
assign w5677 = ~w5658 & w5671;
assign w5678 = w5666 & w7311;
assign w5679 = ~w5676 & ~w5678;
assign w5680 = ~w5673 & w5679;
assign w5681 = ~w5567 & w5586;
assign w5682 = ~w5587 & ~w5681;
assign w5683 = w5680 & ~w5682;
assign w5684 = ~w5680 & w5682;
assign w5685 = ~w5683 & ~w5684;
assign w5686 = ~w5657 & w5685;
assign w5687 = w5657 & ~w5685;
assign w5688 = ~w5686 & ~w5687;
assign w5689 = ~w5590 & ~w5688;
assign w5690 = w5590 & w5688;
assign w5691 = ~w5689 & ~w5690;
assign w5692 = w5642 & ~w5691;
assign w5693 = ~w5642 & w5691;
assign w5694 = ~w5692 & ~w5693;
assign w5695 = ~w3581 & ~w5599;
assign w5696 = w3581 & w5599;
assign w5697 = ~w5695 & ~w5696;
assign w5698 = w5552 & ~w5697;
assign w5699 = ~w5694 & w5698;
assign w5700 = w5694 & ~w5698;
assign w5701 = ~w5699 & ~w5700;
assign w5702 = ~w5640 & ~w5701;
assign w5703 = w5640 & w5701;
assign w5704 = ~w5702 & ~w5703;
assign w5705 = w5637 & w6497;
assign w5706 = (~w5704 & ~w5637) | (~w5704 & w6498) | (~w5637 & w6498);
assign w5707 = ~w5705 & ~w5706;
assign w5708 = w5630 & w5707;
assign w5709 = ~w5630 & ~w5707;
assign w5710 = ~w5708 & ~w5709;
assign w5711 = ~w5532 & ~w5623;
assign w5712 = (~w5624 & w5532) | (~w5624 & w7312) | (w5532 & w7312);
assign w5713 = w5427 & ~w5624;
assign w5714 = w5534 & w5713;
assign w5715 = ~w5320 & w5625;
assign w5716 = w5428 & w5715;
assign w5717 = ~w5429 & w5534;
assign w5718 = w5716 & w5717;
assign w5719 = ~w5712 & ~w5714;
assign w5720 = ~w5718 & w5719;
assign w5721 = w5710 & w5720;
assign w5722 = ~w5710 & ~w5720;
assign w5723 = ~w5721 & ~w5722;
assign w5724 = (~w5633 & ~w5637) | (~w5633 & w6499) | (~w5637 & w6499);
assign w5725 = (w5339 & w5602) | (w5339 & w7313) | (w5602 & w7313);
assign w5726 = (~w5725 & w5640) | (~w5725 & w7314) | (w5640 & w7314);
assign w5727 = w5508 & ~w5699;
assign w5728 = w5601 & w5694;
assign w5729 = ~w5508 & ~w5728;
assign w5730 = ~w5727 & ~w5729;
assign w5731 = w1570 & w4933;
assign w5732 = w5642 & w5689;
assign w5733 = w5598 & w5690;
assign w5734 = ~w5732 & ~w5733;
assign w5735 = ~w5676 & w7315;
assign w5736 = (~w5735 & w5680) | (~w5735 & w7316) | (w5680 & w7316);
assign w5737 = ~w3580 & w7317;
assign w5738 = w1774 & w3585;
assign w5739 = (~w5738 & w5666) | (~w5738 & w7318) | (w5666 & w7318);
assign w5740 = ~w5666 & w7319;
assign w5741 = ~w5739 & ~w5740;
assign w5742 = ~w1556 & w3588;
assign w5743 = (w5667 & w5572) | (w5667 & w7320) | (w5572 & w7320);
assign w5744 = (w5577 & w7321) | (w5577 & w7322) | (w7321 & w7322);
assign w5745 = (~w5742 & w5744) | (~w5742 & w7323) | (w5744 & w7323);
assign w5746 = ~w5741 & w5745;
assign w5747 = w5741 & ~w5745;
assign w5748 = ~w5746 & ~w5747;
assign w5749 = w5737 & w5748;
assign w5750 = ~w5737 & ~w5748;
assign w5751 = ~w5749 & ~w5750;
assign w5752 = ~w5736 & w5751;
assign w5753 = w5736 & ~w5751;
assign w5754 = ~w5752 & ~w5753;
assign w5755 = w5652 & ~w5685;
assign w5756 = ~w5656 & ~w5755;
assign w5757 = (~w5654 & w5755) | (~w5654 & w6279) | (w5755 & w6279);
assign w5758 = ~w5755 & w6280;
assign w5759 = ~w5757 & ~w5758;
assign w5760 = w5754 & w5759;
assign w5761 = ~w5754 & ~w5759;
assign w5762 = ~w5760 & ~w5761;
assign w5763 = w5734 & ~w5762;
assign w5764 = ~w5734 & w5762;
assign w5765 = ~w5763 & ~w5764;
assign w5766 = w5731 & ~w5765;
assign w5767 = ~w5731 & w5765;
assign w5768 = ~w5766 & ~w5767;
assign w5769 = w5730 & w5768;
assign w5770 = ~w5730 & ~w5768;
assign w5771 = ~w5769 & ~w5770;
assign w5772 = w5726 & ~w5771;
assign w5773 = ~w5726 & w5771;
assign w5774 = ~w5772 & ~w5773;
assign w5775 = w5724 & w5774;
assign w5776 = ~w5724 & ~w5774;
assign w5777 = ~w5775 & ~w5776;
assign w5778 = ~w5709 & w5777;
assign w5779 = w5709 & ~w5777;
assign w5780 = ~w5778 & ~w5779;
assign w5781 = (~w5780 & ~w5720) | (~w5780 & w6281) | (~w5720 & w6281);
assign w5782 = w5720 & w6282;
assign w5783 = ~w5781 & ~w5782;
assign w5784 = ~w5731 & w5771;
assign w5785 = ~w5772 & ~w5784;
assign w5786 = ~w1568 & w4933;
assign w5787 = ~w5729 & w5765;
assign w5788 = ~w5727 & ~w5787;
assign w5789 = ~w5787 & w6283;
assign w5790 = w5733 & ~w5762;
assign w5791 = w5732 & w5762;
assign w5792 = ~w5790 & ~w5791;
assign w5793 = w3581 & w5754;
assign w5794 = ~w5754 & w5756;
assign w5795 = ~w5757 & ~w5793;
assign w5796 = ~w5794 & w5795;
assign w5797 = (~w5749 & ~w5751) | (~w5749 & w7324) | (~w5751 & w7324);
assign w5798 = ~w3588 & ~w5743;
assign w5799 = ~w1556 & w3585;
assign w5800 = ~w5798 & w7497;
assign w5801 = w5798 & ~w5799;
assign w5802 = ~w5800 & ~w5801;
assign w5803 = w3585 & w7498;
assign w5804 = ~w5802 & ~w5803;
assign w5805 = (w5666 & w7329) | (w5666 & w7330) | (w7329 & w7330);
assign w5806 = ~w5739 & ~w5805;
assign w5807 = ~w3580 & w7331;
assign w5808 = ~w5806 & w5807;
assign w5809 = ~w3581 & w5806;
assign w5810 = ~w5808 & ~w5809;
assign w5811 = w5804 & ~w5810;
assign w5812 = ~w5804 & w5810;
assign w5813 = ~w5811 & ~w5812;
assign w5814 = w5737 & w5813;
assign w5815 = ~w5737 & ~w5813;
assign w5816 = ~w5814 & ~w5815;
assign w5817 = w5797 & w5816;
assign w5818 = ~w5797 & ~w5816;
assign w5819 = ~w5817 & ~w5818;
assign w5820 = w5796 & ~w5819;
assign w5821 = ~w5796 & w5819;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = ~w5792 & ~w5822;
assign w5824 = w5792 & w5822;
assign w5825 = ~w5823 & ~w5824;
assign w5826 = ~w4933 & ~w5825;
assign w5827 = w4933 & w5825;
assign w5828 = ~w5826 & ~w5827;
assign w5829 = w5789 & ~w5828;
assign w5830 = ~w5789 & w5828;
assign w5831 = ~w5829 & ~w5830;
assign w5832 = w5785 & w5831;
assign w5833 = ~w5785 & ~w5831;
assign w5834 = ~w5832 & ~w5833;
assign w5835 = w5777 & w5834;
assign w5836 = w5710 & w5835;
assign w5837 = ~w5624 & w5836;
assign w5838 = ~w5434 & w6285;
assign w5839 = ~w5776 & ~w5834;
assign w5840 = ~w5778 & w5839;
assign w5841 = ~w5711 & w5837;
assign w5842 = w5776 & w5834;
assign w5843 = w5708 & w5835;
assign w5844 = ~w5842 & ~w5843;
assign w5845 = ~w5708 & w5839;
assign w5846 = w5720 & w5845;
assign w5847 = ~w5841 & w7332;
assign w5848 = ~w5838 & w5847;
assign w5849 = ~w5846 & w5848;
assign w5850 = ~w5841 & w6286;
assign w5851 = w5536 & w5850;
assign w5852 = w1566 & w4933;
assign w5853 = w5590 & ~w5790;
assign w5854 = (w5852 & w5823) | (w5852 & w6287) | (w5823 & w6287);
assign w5855 = ~w5823 & w6288;
assign w5856 = ~w5854 & ~w5855;
assign w5857 = ~w5654 & ~w5758;
assign w5858 = (~w5857 & ~w5796) | (~w5857 & w6289) | (~w5796 & w6289);
assign w5859 = w5797 & w5813;
assign w5860 = ~w5797 & ~w5813;
assign w5861 = ~w5859 & ~w5860;
assign w5862 = w5759 & w7333;
assign w5863 = w5857 & ~w5862;
assign w5864 = ~w5858 & ~w5863;
assign w5865 = (~w5737 & w5797) | (~w5737 & w7334) | (w5797 & w7334);
assign w5866 = ~w5806 & w7335;
assign w5867 = w1086 & w2512;
assign w5868 = w3585 & ~w5867;
assign w5869 = w5800 & w5868;
assign w5870 = ~w5800 & ~w5868;
assign w5871 = ~w5869 & ~w5870;
assign w5872 = w5806 & w7337;
assign w5873 = ~w3580 & w7338;
assign w5874 = w5871 & w5873;
assign w5875 = ~w5871 & ~w5873;
assign w5876 = ~w5874 & ~w5875;
assign w5877 = (~w5876 & ~w5806) | (~w5876 & w7339) | (~w5806 & w7339);
assign w5878 = ~w5866 & ~w5872;
assign w5879 = ~w5877 & w5878;
assign w5880 = ~w5865 & ~w5879;
assign w5881 = (w5879 & w5861) | (w5879 & w7340) | (w5861 & w7340);
assign w5882 = ~w5880 & ~w5881;
assign w5883 = w5864 & w5882;
assign w5884 = ~w5864 & ~w5882;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = w5796 & w7341;
assign w5887 = ~w5885 & ~w5886;
assign w5888 = w5856 & w5887;
assign w5889 = ~w5856 & w5885;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = w5825 & w6290;
assign w5892 = (~w5826 & ~w5788) | (~w5826 & w6291) | (~w5788 & w6291);
assign w5893 = ~w5890 & ~w5892;
assign w5894 = w5890 & w5892;
assign w5895 = ~w5893 & ~w5894;
assign w5896 = w5832 & w5895;
assign w5897 = ~w5832 & ~w5895;
assign w5898 = ~w5896 & ~w5897;
assign w5899 = (~w5898 & w5841) | (~w5898 & w6292) | (w5841 & w6292);
assign w5900 = ~w5841 & w6293;
assign w5901 = ~w5899 & ~w5900;
assign w5902 = ~w5851 & ~w5901;
assign w5903 = w5851 & w5901;
assign w5904 = ~w5902 & ~w5903;
assign w5905 = (w5893 & ~w5785) | (w5893 & w7342) | (~w5785 & w7342);
assign w5906 = (~w5894 & ~w5832) | (~w5894 & w6294) | (~w5832 & w6294);
assign w5907 = ~w5842 & w5906;
assign w5908 = ~w5843 & w5907;
assign w5909 = ~w5905 & w5908;
assign w5910 = ~w5841 & w5909;
assign w5911 = ~w5806 & w7343;
assign w5912 = ~w5872 & ~w5911;
assign w5913 = ~w3580 & w7344;
assign w5914 = (~w5869 & ~w5871) | (~w5869 & w7345) | (~w5871 & w7345);
assign w5915 = ~w5913 & w5914;
assign w5916 = w5913 & ~w5914;
assign w5917 = ~w5915 & ~w5916;
assign w5918 = ~w5873 & w5917;
assign w5919 = (~w5911 & ~w5878) | (~w5911 & w7346) | (~w5878 & w7346);
assign w5920 = ~w5737 & w5919;
assign w5921 = w5737 & ~w5919;
assign w5922 = ~w5920 & ~w5921;
assign w5923 = ~w5861 & w7347;
assign w5924 = ~w5913 & ~w5918;
assign w5925 = w5912 & w5924;
assign w5926 = ~w5923 & w5925;
assign w5927 = (w1563 & w5923) | (w1563 & w7348) | (w5923 & w7348);
assign w5928 = (w4933 & w5862) | (w4933 & w7349) | (w5862 & w7349);
assign w5929 = (w5928 & ~w5864) | (w5928 & w7350) | (~w5864 & w7350);
assign w5930 = (w5926 & w5929) | (w5926 & w7351) | (w5929 & w7351);
assign w5931 = ~w5927 & ~w5930;
assign w5932 = (~w5854 & ~w5856) | (~w5854 & w7352) | (~w5856 & w7352);
assign w5933 = w5931 & ~w5932;
assign w5934 = w5863 & ~w5882;
assign w5935 = ~w5823 & w7353;
assign w5936 = w5852 & ~w5935;
assign w5937 = ~w5823 & w7354;
assign w5938 = ~w5859 & ~w5865;
assign w5939 = w5922 & w5938;
assign w5940 = ~w5881 & w7355;
assign w5941 = ~w5939 & ~w5940;
assign w5942 = (~w5864 & w5937) | (~w5864 & w7356) | (w5937 & w7356);
assign w5943 = w5864 & w5941;
assign w5944 = ~w5855 & ~w5943;
assign w5945 = ~w5942 & w5944;
assign w5946 = ~w5931 & ~w5936;
assign w5947 = ~w5945 & w5946;
assign w5948 = ~w5933 & ~w5947;
assign w5949 = w5910 & ~w5948;
assign w5950 = ~w5838 & w5949;
assign w5951 = w5905 & ~w5948;
assign w5952 = ~w5905 & w5948;
assign w5953 = ~w5951 & ~w5952;
assign w5954 = ~w5910 & ~w5953;
assign w5955 = w5836 & w7357;
assign w5956 = ~w5434 & w6295;
assign w5957 = ~w5954 & ~w5956;
assign w5958 = ~w5950 & w5957;
assign w5959 = (~w5933 & w5905) | (~w5933 & w7358) | (w5905 & w7358);
assign w5960 = (~w5959 & ~w5908) | (~w5959 & w6296) | (~w5908 & w6296);
assign w5961 = (~w5858 & ~w5864) | (~w5858 & w7359) | (~w5864 & w7359);
assign w5962 = w1563 & w4933;
assign w5963 = w5961 & ~w5962;
assign w5964 = (~w1561 & w3580) | (~w1561 & w7360) | (w3580 & w7360);
assign w5965 = ~w5737 & ~w5964;
assign w5966 = w5873 & ~w5917;
assign w5967 = ~w5918 & ~w5966;
assign w5968 = w5912 & ~w5967;
assign w5969 = ~w5912 & w5967;
assign w5970 = ~w5968 & ~w5969;
assign w5971 = ~w5923 & w5970;
assign w5972 = w5965 & w7499;
assign w5973 = ~w5963 & w5972;
assign w5974 = ~w5965 & ~w5927;
assign w5975 = ~w5929 & w5974;
assign w5976 = ~w5973 & ~w5975;
assign w5977 = w5720 & w6297;
assign w5978 = w5895 & w5948;
assign w5979 = w5836 & w7362;
assign w5980 = ~w5720 & w5979;
assign w5981 = (~w5976 & ~w5836) | (~w5976 & w7363) | (~w5836 & w7363);
assign w5982 = ~w5960 & w5981;
assign w5983 = w5976 & ~w5959;
assign w5984 = (w5983 & ~w5908) | (w5983 & w7364) | (~w5908 & w7364);
assign w5985 = ~w5982 & ~w5984;
assign w5986 = ~w5980 & w5985;
assign w5987 = ~w5977 & w5986;
assign w5988 = (w5737 & w4933) | (w5737 & w7365) | (w4933 & w7365);
assign w5989 = (~w1774 & w3580) | (~w1774 & w7366) | (w3580 & w7366);
assign w5990 = (~w5989 & w4933) | (~w5989 & w7367) | (w4933 & w7367);
assign w5991 = ~w5737 & ~w5990;
assign w5992 = ~w5988 & ~w5991;
assign w5993 = (~w1563 & w5961) | (~w1563 & w7368) | (w5961 & w7368);
assign w5994 = w5972 & ~w5993;
assign w5995 = ~w5992 & ~w5994;
assign w5996 = w5990 & w5994;
assign w5997 = ~w5995 & ~w5996;
assign w5998 = (w6298 & ~w5908) | (w6298 & w7369) | (~w5908 & w7369);
assign w5999 = (w5908 & w7370) | (w5908 & w7371) | (w7370 & w7371);
assign w6000 = ~w5998 & ~w5999;
assign w6001 = (w6000 & w5720) | (w6000 & w7372) | (w5720 & w7372);
assign w6002 = ~w5720 & w6300;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = (~w5737 & w4933) | (~w5737 & w7373) | (w4933 & w7373);
assign w6005 = w1556 & w3581;
assign w6006 = ~w1556 & w4933;
assign w6007 = ~w6005 & ~w6006;
assign w6008 = ~w6004 & ~w6007;
assign w6009 = w6004 & w6007;
assign w6010 = ~w6008 & ~w6009;
assign w6011 = (~w6010 & ~w5994) | (~w6010 & w7374) | (~w5994 & w7374);
assign w6012 = (w5908 & w7375) | (w5908 & w7376) | (w7375 & w7376);
assign w6013 = w5720 & ~w6012;
assign w6014 = (w6010 & w5994) | (w6010 & w7377) | (w5994 & w7377);
assign w6015 = w5836 & w7378;
assign w6016 = ~w5720 & ~w6015;
assign w6017 = ~w6013 & ~w6016;
assign w6018 = w5976 & ~w5995;
assign w6019 = w5836 & w7379;
assign w6020 = ~w5959 & w6018;
assign w6021 = (w6020 & ~w5908) | (w6020 & w7380) | (~w5908 & w7380);
assign w6022 = ~w6021 & w6301;
assign w6023 = w6014 & ~w5999;
assign w6024 = ~w6022 & ~w6023;
assign w6025 = ~w6017 & w6024;
assign w6026 = w2513 & ~w3580;
assign w6027 = (~w1086 & ~w3581) | (~w1086 & w7381) | (~w3581 & w7381);
assign w6028 = ~w6026 & ~w6027;
assign w6029 = ~w6028 & ~w6014;
assign w6030 = (w6028 & ~w6007) | (w6028 & w7382) | (~w6007 & w7382);
assign w6031 = (w5994 & w7384) | (w5994 & w7385) | (w7384 & w7385);
assign w6032 = ~w6029 & ~w6031;
assign w6033 = w5836 & w7386;
assign w6034 = (~w6028 & w6007) | (~w6028 & w7387) | (w6007 & w7387);
assign w6035 = ~w5996 & w6034;
assign w6036 = (w5908 & w7388) | (w5908 & w7389) | (w7388 & w7389);
assign w6037 = w6032 & ~w6036;
assign w6038 = (~w6037 & w5720) | (~w6037 & w7390) | (w5720 & w7390);
assign w6039 = (w6030 & w6021) | (w6030 & w6303) | (w6021 & w6303);
assign w6040 = (w6039 & ~w5720) | (w6039 & w7391) | (~w5720 & w7391);
assign w6041 = ~w6038 & ~w6040;
assign w6042 = (~w6028 & ~w6007) | (~w6028 & w7392) | (~w6007 & w7392);
assign w6043 = (w6042 & w6021) | (w6042 & w6304) | (w6021 & w6304);
assign w6044 = (w6043 & ~w5720) | (w6043 & w7393) | (~w5720 & w7393);
assign w6045 = w2513 & w3580;
assign w6046 = ~w6044 & ~w6045;
assign w6047 = w7 & w23;
assign w6048 = ~pi19 & pi09;
assign w6049 = w13 & w93;
assign w6050 = w11 & w7394;
assign w6051 = pi01 & w33;
assign w6052 = ~pi19 & pi10;
assign w6053 = pi15 & pi08;
assign w6054 = pi14 & w113;
assign w6055 = ~w119 & ~w10;
assign w6056 = pi07 & pi00;
assign w6057 = w23 & w72;
assign w6058 = w7 & pi14;
assign w6059 = ~pi19 & pi11;
assign w6060 = w23 & w113;
assign w6061 = pi15 & pi09;
assign w6062 = w23 & pi09;
assign w6063 = ~pi19 & pi13;
assign w6064 = ~w182 & w7395;
assign w6065 = pi07 & w31;
assign w6066 = ~pi06 & pi00;
assign w6067 = w20 & w231;
assign w6068 = pi15 & pi10;
assign w6069 = (~w10 & ~w249) | (~w10 & w7396) | (~w249 & w7396);
assign w6070 = w110 & pi12;
assign w6071 = ~pi19 & pi14;
assign w6072 = w299 & ~w268;
assign w6073 = ~pi19 & pi08;
assign w6074 = pi15 & pi06;
assign w6075 = pi14 & w70;
assign w6076 = ~w353 & ~w10;
assign w6077 = ~w301 & w365;
assign w6078 = w404 & w406;
assign w6079 = (~w364 & ~w406) | (~w364 & w6305) | (~w406 & w6305);
assign w6080 = ~w433 & w436;
assign w6081 = w366 & ~w457;
assign w6082 = ~w376 & w413;
assign w6083 = w525 & ~w513;
assign w6084 = ~w142 & ~w220;
assign w6085 = ~w556 & ~w566;
assign w6086 = w571 & w575;
assign w6087 = (w555 & w515) | (w555 & w6500) | (w515 & w6500);
assign w6088 = ~w515 & w6501;
assign w6089 = w406 & w6306;
assign w6090 = w301 & w342;
assign w6091 = w671 & ~w669;
assign w6092 = (~w342 & w6307) | (~w342 & w7500) | (w6307 & w7500);
assign w6093 = (w681 & w7397) | (w681 & w7398) | (w7397 & w7398);
assign w6094 = (~w699 & w6309) | (~w699 & w7500) | (w6309 & w7500);
assign w6095 = w703 & ~w696;
assign w6096 = w742 & ~w744;
assign w6097 = ~w608 & ~w746;
assign w6098 = w608 & ~w403;
assign w6099 = ~w754 & w649;
assign w6100 = ~w654 & ~w615;
assign w6101 = ~w598 & w553;
assign w6102 = ~w713 & ~w103;
assign w6103 = ~w707 & w754;
assign w6104 = ~w707 & ~w512;
assign w6105 = ~w856 & ~w858;
assign w6106 = w783 & ~w756;
assign w6107 = ~w876 & ~w904;
assign w6108 = w876 & w904;
assign w6109 = ~w798 & w797;
assign w6110 = w937 & ~w920;
assign w6111 = w907 & ~w180;
assign w6112 = ~w912 & w983;
assign w6113 = w912 & ~w983;
assign w6114 = w911 & w719;
assign w6115 = ~w988 & ~w994;
assign w6116 = ~w937 & w920;
assign w6117 = w981 & w1039;
assign w6118 = ~w981 & ~w1039;
assign w6119 = (w886 & w6310) | (w886 & w7501) | (w6310 & w7501);
assign w6120 = ~w886 & ~w1131;
assign w6121 = w719 & ~w633;
assign w6122 = ~w719 & ~w633;
assign w6123 = ~w1149 & ~w1143;
assign w6124 = w716 & ~w633;
assign w6125 = w1207 & ~w1203;
assign w6126 = w1231 & ~w1230;
assign w6127 = ~w707 & ~w1260;
assign w6128 = ~w1270 & ~w1268;
assign w6129 = w1291 & ~w1284;
assign w6130 = w821 & ~w817;
assign w6131 = w259 & w1331;
assign w6132 = ~w1337 & ~w1327;
assign w6133 = w1337 & w1327;
assign w6134 = w1345 & ~w1344;
assign w6135 = w1390 & ~w1425;
assign w6136 = w926 & w1455;
assign w6137 = ~w1462 & w6311;
assign w6138 = (~w1449 & w1462) | (~w1449 & w6312) | (w1462 & w6312);
assign w6139 = ~w1007 & ~w1503;
assign w6140 = ~w1003 & w6313;
assign w6141 = ~w1504 & w1511;
assign w6142 = w2018 & ~w2015;
assign w6143 = (~w141 & ~w2103) | (~w141 & w7399) | (~w2103 & w7399);
assign w6144 = (~w2185 & ~w1520) | (~w2185 & w7400) | (~w1520 & w7400);
assign w6145 = w1581 & ~w2199;
assign w6146 = w2201 & w7502;
assign w6147 = ~w2249 & w2251;
assign w6148 = w2253 & ~w1568;
assign w6149 = ~w2253 & w2260;
assign w6150 = ~w2271 & ~w2269;
assign w6151 = w2420 & ~w2409;
assign w6152 = w2426 & ~w364;
assign w6153 = ~w2449 & w2383;
assign w6154 = ~w2455 & w2382;
assign w6155 = w2455 & ~w2382;
assign w6156 = w2461 & ~w2460;
assign w6157 = w2465 & ~w2464;
assign w6158 = w2470 & ~w2469;
assign w6159 = ~w2478 & ~w2474;
assign w6160 = w2579 & w2538;
assign w6161 = ~w2579 & ~w2538;
assign w6162 = w2587 & ~w2586;
assign w6163 = ~w2700 & ~w2694;
assign w6164 = (~w2679 & w2552) | (~w2679 & w6314) | (w2552 & w6314);
assign w6165 = w2732 & ~w2745;
assign w6166 = ~w2679 & w7515;
assign w6167 = ~w2916 & ~w2859;
assign w6168 = ~w2925 & w6315;
assign w6169 = (~w2858 & w2925) | (~w2858 & w6316) | (w2925 & w6316);
assign w6170 = ~w2960 & ~w1988;
assign w6171 = (~w2996 & ~w2965) | (~w2996 & w7402) | (~w2965 & w7402);
assign w6172 = w2965 & w7403;
assign w6173 = w2994 & ~w2996;
assign w6174 = w1590 & ~w3029;
assign w6175 = ~w3088 & w3094;
assign w6176 = w3095 & ~w1570;
assign w6177 = ~w3033 & w3031;
assign w6178 = w3033 & w3113;
assign w6179 = w3033 & ~w3031;
assign w6180 = ~w3033 & w3119;
assign w6181 = (w3030 & w3148) | (w3030 & w7404) | (w3148 & w7404);
assign w6182 = (~w3030 & ~w3139) | (~w3030 & w7405) | (~w3139 & w7405);
assign w6183 = w3247 & ~w3255;
assign w6184 = ~w3247 & w3255;
assign w6185 = w3268 & ~w3226;
assign w6186 = ~w3269 & w3225;
assign w6187 = w3269 & ~w3225;
assign w6188 = w3275 & ~w3279;
assign w6189 = (~w3285 & w3279) | (~w3285 & w7406) | (w3279 & w7406);
assign w6190 = (w1563 & ~w3287) | (w1563 & w6317) | (~w3287 & w6317);
assign w6191 = w3264 & w3399;
assign w6192 = w3400 & w7407;
assign w6193 = w3413 & w6318;
assign w6194 = ~w3421 & w7408;
assign w6195 = (~w3352 & w3421) | (~w3352 & w7409) | (w3421 & w7409);
assign w6196 = (w3425 & w3421) | (w3425 & w7410) | (w3421 & w7410);
assign w6197 = ~w3421 & w7411;
assign w6198 = ~w3165 & ~w3460;
assign w6199 = w3454 & ~w3473;
assign w6200 = ~w3484 & ~w2507;
assign w6201 = ~w2357 & ~w2361;
assign w6202 = ~w3489 & w2372;
assign w6203 = ~w1556 & ~w3526;
assign w6204 = (~w3207 & w1556) | (~w3207 & w7412) | (w1556 & w7412);
assign w6205 = (w1648 & ~w3526) | (w1648 & w7413) | (~w3526 & w7413);
assign w6206 = w3526 & w7414;
assign w6207 = (~w3620 & w3611) | (~w3620 & w7415) | (w3611 & w7415);
assign w6208 = ~w3651 & ~w3647;
assign w6209 = ~w3642 & w3601;
assign w6210 = ~w3672 & ~w1648;
assign w6211 = (w3598 & w3663) | (w3598 & w6319) | (w3663 & w6319);
assign w6212 = ~w3663 & w6320;
assign w6213 = ~w3670 & w3697;
assign w6214 = w3670 & ~w3697;
assign w6215 = (~w1542 & ~w3526) | (~w1542 & w7416) | (~w3526 & w7416);
assign w6216 = ~w3706 & ~w3677;
assign w6217 = (~w1570 & w3528) | (~w1570 & w7417) | (w3528 & w7417);
assign w6218 = w3705 & ~w3724;
assign w6219 = ~w3756 & w3770;
assign w6220 = w3756 & ~w3770;
assign w6221 = (w3808 & w3805) | (w3808 & w6321) | (w3805 & w6321);
assign w6222 = (~w1584 & w3528) | (~w1584 & w7418) | (w3528 & w7418);
assign w6223 = (~w3869 & w3858) | (~w3869 & w6322) | (w3858 & w6322);
assign w6224 = ~w3781 & w6323;
assign w6225 = (w3923 & w3781) | (w3923 & w6324) | (w3781 & w6324);
assign w6226 = w3749 & w3928;
assign w6227 = w3755 & ~w3770;
assign w6228 = w3766 & ~w3761;
assign w6229 = ~w1568 & w3940;
assign w6230 = (~w1563 & ~w3526) | (~w1563 & w7419) | (~w3526 & w7419);
assign w6231 = w3744 & ~w3964;
assign w6232 = ~w3744 & w3964;
assign w6233 = w3938 & w4023;
assign w6234 = ~w3938 & ~w4023;
assign w6235 = (~w3947 & ~w3950) | (~w3947 & w7420) | (~w3950 & w7420);
assign w6236 = ~w4032 & w7421;
assign w6237 = ~w1566 & w4028;
assign w6238 = w1566 & w4028;
assign w6239 = w4051 & w4046;
assign w6240 = ~w4051 & ~w4046;
assign w6241 = ~w4018 & ~w4108;
assign w6242 = (~w1774 & ~w3526) | (~w1774 & w7422) | (~w3526 & w7422);
assign w6243 = w4123 & ~w4120;
assign w6244 = w4157 & w4230;
assign w6245 = ~w4157 & ~w4230;
assign w6246 = ~w4150 & ~w4127;
assign w6247 = w4142 & ~w4141;
assign w6248 = w4252 & w1561;
assign w6249 = ~w4242 & w4328;
assign w6250 = w4242 & ~w4328;
assign w6251 = ~w3526 & w3528;
assign w6252 = w4340 & ~w4341;
assign w6253 = (w6325 & w3549) | (w6325 & w7423) | (w3549 & w7423);
assign w6254 = ~w4338 & ~w4350;
assign w6255 = w4338 & w4350;
assign w6256 = w3526 & w3610;
assign w6257 = w4576 & w4586;
assign w6258 = ~w4449 & w3549;
assign w6259 = (w3594 & ~w4749) | (w3594 & w6326) | (~w4749 & w6326);
assign w6260 = w4749 & w6327;
assign w6261 = w4868 & ~w4866;
assign w6262 = ~w4851 & ~w4982;
assign w6263 = (w1086 & ~w2513) | (w1086 & w7424) | (~w2513 & w7424);
assign w6264 = w4984 & w4988;
assign w6265 = ~w5025 & ~w5164;
assign w6266 = w5025 & ~w3571;
assign w6267 = w5126 & ~w5243;
assign w6268 = ~w5126 & w5243;
assign w6269 = (~w5248 & w5006) | (~w5248 & w7425) | (w5006 & w7425);
assign w6270 = ~w5006 & w5248;
assign w6271 = w1086 & ~w5263;
assign w6272 = ~w5024 & w7426;
assign w6273 = (~w5286 & w5024) | (~w5286 & w7427) | (w5024 & w7427);
assign w6274 = ~w5354 & ~w5281;
assign w6275 = (w5169 & w7428) | (w5169 & w7429) | (w7428 & w7429);
assign w6276 = w5351 & ~w5394;
assign w6277 = ~w3911 & ~w3985;
assign w6278 = ~w5571 & w5574;
assign w6279 = w5656 & ~w5654;
assign w6280 = ~w5656 & w3581;
assign w6281 = ~w5710 & ~w5780;
assign w6282 = w5710 & w5780;
assign w6283 = (~w5786 & w5699) | (~w5786 & w7430) | (w5699 & w7430);
assign w6284 = ~w3585 & w5745;
assign w6285 = w5535 & w5837;
assign w6286 = w5844 & w5837;
assign w6287 = w5853 & w5852;
assign w6288 = ~w5853 & ~w5852;
assign w6289 = w5819 & ~w5857;
assign w6290 = w4933 & w1568;
assign w6291 = w5891 & ~w5826;
assign w6292 = ~w5844 & ~w5898;
assign w6293 = w5844 & w5898;
assign w6294 = ~w5895 & ~w5894;
assign w6295 = w5535 & w5955;
assign w6296 = w5933 & ~w5959;
assign w6297 = ~w5960 & ~w5976;
assign w6298 = w5983 & ~w5997;
assign w6299 = ~w5983 & w5997;
assign w6300 = w5979 & w5997;
assign w6301 = ~w6019 & w6011;
assign w6302 = ~w5983 & w6035;
assign w6303 = w6019 & w6030;
assign w6304 = w6019 & w6042;
assign w6305 = ~w403 & ~w364;
assign w6306 = w403 & ~w364;
assign w6307 = ~w688 & ~w342;
assign w6308 = w688 & w342;
assign w6309 = ~w688 & ~w699;
assign w6310 = w732 & w886;
assign w6311 = w1464 & w1449;
assign w6312 = ~w1464 & ~w1449;
assign w6313 = w1007 & w1503;
assign w6314 = w2546 & ~w2679;
assign w6315 = w2927 & w2858;
assign w6316 = ~w2927 & ~w2858;
assign w6317 = w3285 & w1563;
assign w6318 = ~w3412 & w3355;
assign w6319 = w1590 & w7503;
assign w6320 = ~w3601 & ~w3598;
assign w6321 = w3804 & w3808;
assign w6322 = w3867 & ~w3869;
assign w6323 = ~w3782 & ~w3923;
assign w6324 = ~w1576 & w7504;
assign w6325 = w4248 & w1774;
assign w6326 = w4715 & w3594;
assign w6327 = ~w4715 & ~w4856;
assign w6328 = ~pi05 & ~w31;
assign w6329 = pi10 & pi07;
assign w6330 = w263 & w39;
assign w6331 = w15 & ~w278;
assign w6332 = ~w296 & ~w299;
assign w6333 = pi19 & pi17;
assign w6334 = ~w146 & ~w95;
assign w6335 = pi09 & pi07;
assign w6336 = pi15 & pi13;
assign w6337 = w143 & pi12;
assign w6338 = w327 & w329;
assign w6339 = ~w335 & ~w341;
assign w6340 = w20 & w284;
assign w6341 = pi10 & ~w384;
assign w6342 = w134 & ~w386;
assign w6343 = w382 & w402;
assign w6344 = w142 & w404;
assign w6345 = w411 & w413;
assign w6346 = ~w411 & ~w413;
assign w6347 = ~w194 & ~w364;
assign w6348 = w142 & w421;
assign w6349 = w421 & ~w141;
assign w6350 = w253 & w7505;
assign w6351 = ~w141 & ~w364;
assign w6352 = ~w369 & ~w308;
assign w6353 = ~w463 & ~w452;
assign w6354 = w468 & w260;
assign w6355 = ~w468 & ~w260;
assign w6356 = ~w411 & w483;
assign w6357 = ~w424 & w512;
assign w6358 = ~w424 & ~w519;
assign w6359 = ~w525 & w253;
assign w6360 = w539 & ~w511;
assign w6361 = ~w539 & w511;
assign w6362 = ~w519 & w177;
assign w6363 = w564 & w558;
assign w6364 = w594 & w554;
assign w6365 = ~w594 & ~w554;
assign w6366 = w595 & w597;
assign w6367 = ~w599 & w602;
assign w6368 = ~w606 & ~w608;
assign w6369 = ~w549 & w610;
assign w6370 = ~w471 & w614;
assign w6371 = w469 & w616;
assign w6372 = ~w634 & ~w630;
assign w6373 = w693 & ~w342;
assign w6374 = w693 & ~w6093;
assign w6375 = ~w6094 & ~w693;
assign w6376 = ~w643 & ~w641;
assign w6377 = ~w711 & ~w803;
assign w6378 = w711 & w803;
assign w6379 = w809 & ~w745;
assign w6380 = w753 & ~w403;
assign w6381 = ~w410 & ~w253;
assign w6382 = w879 & ~w403;
assign w6383 = ~w879 & ~w972;
assign w6384 = w865 & ~w999;
assign w6385 = ~w1000 & ~w996;
assign w6386 = w633 & w1132;
assign w6387 = ~w1202 & ~w1233;
assign w6388 = w1280 & ~w1259;
assign w6389 = ~w1280 & w1259;
assign w6390 = ~w1301 & w1256;
assign w6391 = w1301 & ~w1256;
assign w6392 = w1326 & ~w1344;
assign w6393 = w1326 & ~w1347;
assign w6394 = ~w1326 & w1344;
assign w6395 = ~w1326 & w1347;
assign w6396 = ~w827 & ~w1391;
assign w6397 = w827 & w1391;
assign w6398 = ~w1386 & ~w1425;
assign w6399 = ~w1386 & w1423;
assign w6400 = w1386 & w1425;
assign w6401 = w1386 & ~w1423;
assign w6402 = ~w1511 & ~w1503;
assign w6403 = ~w1511 & ~w6140;
assign w6404 = w1088 & w7506;
assign w6405 = w1090 & w1503;
assign w6406 = w1090 & w6140;
assign w6407 = w1465 & w1472;
assign w6408 = ~w1465 & ~w1472;
assign w6409 = ~w1618 & ~w1623;
assign w6410 = w1500 & ~w1481;
assign w6411 = w1815 & ~w1811;
assign w6412 = w1807 & ~w253;
assign w6413 = ~w220 & ~w1616;
assign w6414 = w220 & w1616;
assign w6415 = w1912 & w1891;
assign w6416 = ~w1912 & ~w1891;
assign w6417 = w2047 & ~w2045;
assign w6418 = ~w1581 & ~w2100;
assign w6419 = w1581 & ~w2099;
assign w6420 = ~w2142 & ~w2085;
assign w6421 = w2142 & w2085;
assign w6422 = w1509 & ~w364;
assign w6423 = ~w2560 & w7445;
assign w6424 = w2571 & w2539;
assign w6425 = ~w2571 & ~w2539;
assign w6426 = ~w2746 & ~w2759;
assign w6427 = ~w2940 & w3129;
assign w6428 = ~w3310 & ~w3223;
assign w6429 = ~w3307 & w3325;
assign w6430 = w3307 & ~w3325;
assign w6431 = ~w3323 & w3325;
assign w6432 = ~w3337 & ~w3338;
assign w6433 = w3340 & w3344;
assign w6434 = ~w3340 & ~w3344;
assign w6435 = (w3450 & w3445) | (w3450 & w7446) | (w3445 & w7446);
assign w6436 = ~w3735 & ~w3737;
assign w6437 = w3730 & w3734;
assign w6438 = w3700 & ~w3782;
assign w6439 = w3818 & ~w3814;
assign w6440 = ~w3843 & ~w3797;
assign w6441 = w3875 & ~w3874;
assign w6442 = w3925 & ~w4005;
assign w6443 = ~w3777 & w6502;
assign w6444 = (~w4010 & w3777) | (~w4010 & w6503) | (w3777 & w6503);
assign w6445 = w3925 & ~w4089;
assign w6446 = ~w4096 & ~w4097;
assign w6447 = w4020 & ~w4108;
assign w6448 = ~w4020 & w4108;
assign w6449 = w4134 & ~w4147;
assign w6450 = ~w4094 & w3911;
assign w6451 = ~w4101 & w6504;
assign w6452 = (~w4215 & w4101) | (~w4215 & w6505) | (w4101 & w6505);
assign w6453 = ~w4113 & w6506;
assign w6454 = (~w4220 & w4113) | (~w4220 & w6507) | (w4113 & w6507);
assign w6455 = ~w4197 & w6508;
assign w6456 = ~w4210 & w6509;
assign w6457 = w4237 & ~w4365;
assign w6458 = ~w4237 & w4365;
assign w6459 = w4222 & ~w4223;
assign w6460 = w4391 & ~w4390;
assign w6461 = ~w4549 & w4683;
assign w6462 = ~w4555 & w4690;
assign w6463 = w4670 & w4674;
assign w6464 = ~w4679 & w7447;
assign w6465 = ~w4772 & w4822;
assign w6466 = w4772 & ~w4822;
assign w6467 = ~w4710 & w4842;
assign w6468 = ~w4849 & w4851;
assign w6469 = ~w4615 & w6510;
assign w6470 = (w4900 & w4615) | (w4900 & w6511) | (w4615 & w6511);
assign w6471 = (w3581 & w4681) | (w3581 & w6512) | (w4681 & w6512);
assign w6472 = w4825 & ~w4824;
assign w6473 = (w3588 & ~w4686) | (w3588 & w6513) | (~w4686 & w6513);
assign w6474 = ~w4843 & w4982;
assign w6475 = w4843 & ~w4982;
assign w6476 = w4971 & ~w4968;
assign w6477 = (~w5118 & w4898) | (~w5118 & w6514) | (w4898 & w6514);
assign w6478 = ~w4898 & w6515;
assign w6479 = w5120 & ~w5119;
assign w6480 = ~w5325 & w1590;
assign w6481 = ~w5230 & ~w5339;
assign w6482 = (w5339 & w5231) | (w5339 & w7448) | (w5231 & w7448);
assign w6483 = ~w5237 & w3585;
assign w6484 = w5237 & ~w5347;
assign w6485 = ~w5255 & w7449;
assign w6486 = w5220 & ~w4948;
assign w6487 = w5101 & ~w4947;
assign w6488 = w5320 & ~w5427;
assign w6489 = w5421 & ~w5328;
assign w6490 = (w5309 & w7450) | (w5309 & w7451) | (w7450 & w7451);
assign w6491 = w4933 & ~w5413;
assign w6492 = ~w5340 & ~w5339;
assign w6493 = w5391 & w3588;
assign w6494 = ~w5372 & w5477;
assign w6495 = ~w5499 & ~w5553;
assign w6496 = w5438 & ~w5439;
assign w6497 = ~w5633 & w5704;
assign w6498 = w5633 & ~w5704;
assign w6499 = ~w5704 & ~w5633;
assign w6500 = ~w6085 & w555;
assign w6501 = w6085 & ~w555;
assign w6502 = w6232 & w4010;
assign w6503 = ~w6232 & ~w4010;
assign w6504 = w4103 & w4215;
assign w6505 = ~w4103 & ~w4215;
assign w6506 = w4114 & w4220;
assign w6507 = ~w4114 & ~w4220;
assign w6508 = ~w4195 & ~w4302;
assign w6509 = ~w4208 & w4306;
assign w6510 = w4694 & ~w4900;
assign w6511 = ~w4694 & w4900;
assign w6512 = w4816 & w3581;
assign w6513 = w4830 & w3588;
assign w6514 = ~w4978 & ~w5118;
assign w6515 = w4978 & w4075;
assign w6516 = w6087 & ~w301;
assign w6517 = ~w6087 & ~w585;
assign w6518 = ~w6211 & ~w3734;
assign w6519 = w6211 & w3733;
assign w6520 = w3739 & ~w3789;
assign w6521 = w3826 & ~w3821;
assign w6522 = ~w3882 & ~w3880;
assign w6523 = ~w3592 & ~w3912;
assign w6524 = ~w3793 & w3595;
assign w6525 = w3592 & w3911;
assign w6526 = ~w3988 & ~w3986;
assign w6527 = w3989 & w3986;
assign w6528 = ~w4006 & ~w4092;
assign w6529 = ~w3990 & w4076;
assign w6530 = w4087 & ~w4195;
assign w6531 = ~w4182 & ~w4178;
assign w6532 = w4200 & ~w4198;
assign w6533 = w4206 & w4306;
assign w6534 = ~w4206 & ~w4306;
assign w6535 = ~w4216 & w7452;
assign w6536 = (w4317 & w4216) | (w4317 & w7453) | (w4216 & w7453);
assign w6537 = w4075 & w3588;
assign w6538 = w4633 & w4634;
assign w6539 = ~w4512 & ~w4662;
assign w6540 = ~w4512 & ~w4633;
assign w6541 = w4512 & w4662;
assign w6542 = ~w4525 & w7454;
assign w6543 = ~w4581 & ~w4579;
assign w6544 = w3582 & ~w4658;
assign w6545 = w4787 & ~w4634;
assign w6546 = ~w4811 & w4674;
assign w6547 = ~w4811 & w4781;
assign w6548 = w4811 & ~w4674;
assign w6549 = w4811 & ~w4781;
assign w6550 = ~w4678 & ~w4681;
assign w6551 = ~w4720 & ~w4865;
assign w6552 = w3556 & w7381;
assign w6553 = w4867 & ~w4868;
assign w6554 = w1774 & ~w4866;
assign w6555 = ~w4798 & ~w4935;
assign w6556 = ~w4828 & ~w4957;
assign w6557 = w4828 & ~w3579;
assign w6558 = ~w6470 & ~w4966;
assign w6559 = ~w4879 & ~w4991;
assign w6560 = ~w4812 & ~w4811;
assign w6561 = w4802 & w4634;
assign w6562 = ~w4802 & ~w5076;
assign w6563 = w4802 & w5076;
assign w6564 = w4812 & ~w4813;
assign w6565 = w4952 & ~w5101;
assign w6566 = (w3585 & w4961) | (w3585 & w7455) | (w4961 & w7455);
assign w6567 = (~w5108 & w4827) | (~w5108 & w7456) | (w4827 & w7456);
assign w6568 = ~w1774 & ~w5132;
assign w6569 = ~w3559 & ~w1556;
assign w6570 = w3559 & ~w1556;
assign w6571 = w5094 & w5090;
assign w6572 = ~w5185 & ~w5221;
assign w6573 = (w3581 & w4961) | (w3581 & w7457) | (w4961 & w7457);
assign w6574 = ~w5113 & w7458;
assign w6575 = (~w5230 & w5113) | (~w5230 & w7459) | (w5113 & w7459);
assign w6576 = w5300 & w3581;
assign w6577 = pi03 & ~pi04;
assign w6578 = ~pi06 & ~pi05;
assign w6579 = w13 & w15;
assign w6580 = w20 & ~w21;
assign w6581 = w27 & ~w30;
assign w6582 = w46 & w49;
assign w6583 = w46 & ~w48;
assign w6584 = w54 & ~w53;
assign w6585 = w13 & w2;
assign w6586 = w60 & ~pi19;
assign w6587 = w134 & w130;
assign w6588 = w13 & pi02;
assign w6589 = w143 & pi08;
assign w6590 = pi07 & pi01;
assign w6591 = ~pi19 & pi12;
assign w6592 = ~w142 & w253;
assign w6593 = pi13 & pi11;
assign w6594 = pi04 & pi02;
assign w6595 = pi01 & w95;
assign w6596 = w301 & w376;
assign w6597 = ~pi04 & ~pi02;
assign w6598 = ~pi19 & ~pi17;
assign w6599 = ~w396 & ~w395;
assign w6600 = ~w300 & w403;
assign w6601 = w447 & ~w255;
assign w6602 = ~w177 & w473;
assign w6603 = w177 & ~w473;
assign w6604 = ~w463 & ~w478;
assign w6605 = w495 & w499;
assign w6606 = ~w500 & ~w497;
assign w6607 = ~w512 & ~w528;
assign w6608 = w537 & ~w253;
assign w6609 = w537 & ~w6359;
assign w6610 = w569 & ~w177;
assign w6611 = ~w587 & w585;
assign w6612 = ~w6365 & ~w403;
assign w6613 = w6361 & w342;
assign w6614 = ~w6361 & ~w605;
assign w6615 = ~w403 & ~w621;
assign w6616 = w374 & w177;
assign w6617 = ~w374 & ~w177;
assign w6618 = w296 & ~w268;
assign w6619 = w142 & ~w220;
assign w6620 = ~w6602 & ~w648;
assign w6621 = w145 & ~w364;
assign w6622 = w252 & ~w364;
assign w6623 = ~w253 & w375;
assign w6624 = ~w665 & ~w220;
assign w6625 = w665 & w220;
assign w6626 = ~w6624 & w301;
assign w6627 = w676 & w682;
assign w6628 = w676 & ~w675;
assign w6629 = w689 & w694;
assign w6630 = w692 & w701;
assign w6631 = w253 & ~w180;
assign w6632 = ~w707 & w260;
assign w6633 = ~w734 & w259;
assign w6634 = w739 & ~w737;
assign w6635 = ~w180 & ~w742;
assign w6636 = w730 & ~w736;
assign w6637 = w374 & ~w177;
assign w6638 = ~w259 & w220;
assign w6639 = ~w815 & ~w813;
assign w6640 = w180 & ~w837;
assign w6641 = ~w737 & w731;
assign w6642 = ~w259 & w180;
assign w6643 = ~w707 & w857;
assign w6644 = w725 & w553;
assign w6645 = w845 & ~w865;
assign w6646 = ~w749 & ~w868;
assign w6647 = ~w753 & ~w871;
assign w6648 = ~w790 & w872;
assign w6649 = w772 & w882;
assign w6650 = ~w772 & ~w882;
assign w6651 = w778 & ~w305;
assign w6652 = ~w845 & w865;
assign w6653 = ~w707 & w568;
assign w6654 = w716 & w553;
assign w6655 = w935 & ~w931;
assign w6656 = w873 & ~w259;
assign w6657 = ~w891 & w253;
assign w6658 = w891 & ~w253;
assign w6659 = ~w6658 & ~w889;
assign w6660 = ~w894 & ~w883;
assign w6661 = w897 & w963;
assign w6662 = ~w897 & ~w963;
assign w6663 = w877 & w901;
assign w6664 = ~w969 & ~w971;
assign w6665 = w964 & w1014;
assign w6666 = ~w964 & ~w1014;
assign w6667 = ~w959 & ~w957;
assign w6668 = w949 & ~w253;
assign w6669 = w949 & ~w6657;
assign w6670 = ~w1021 & ~w1019;
assign w6671 = w1021 & w1019;
assign w6672 = w734 & ~w1031;
assign w6673 = ~w734 & w1031;
assign w6674 = w1024 & ~w1046;
assign w6675 = ~w1024 & ~w403;
assign w6676 = w301 & ~w6668;
assign w6677 = w301 & ~w6669;
assign w6678 = ~w220 & w1019;
assign w6679 = w1051 & w1050;
assign w6680 = ~w1051 & ~w1050;
assign w6681 = w1028 & ~w1016;
assign w6682 = ~w306 & w1058;
assign w6683 = w306 & ~w1058;
assign w6684 = w1013 & ~w1062;
assign w6685 = ~w1013 & w1062;
assign w6686 = w1050 & ~w6676;
assign w6687 = w1050 & ~w6677;
assign w6688 = ~w1072 & ~w1019;
assign w6689 = ~w1072 & ~w6678;
assign w6690 = ~w6675 & ~w1074;
assign w6691 = w1055 & w1075;
assign w6692 = w1071 & w633;
assign w6693 = ~w1078 & ~w1077;
assign w6694 = ~w1065 & ~w1081;
assign w6695 = ~w1069 & ~w1085;
assign w6696 = w1069 & w1085;
assign w6697 = w932 & w886;
assign w6698 = w932 & w1211;
assign w6699 = ~w707 & ~w732;
assign w6700 = ~w1098 & ~w1103;
assign w6701 = ~w1105 & ~w920;
assign w6702 = w886 & ~w1107;
assign w6703 = ~w886 & w1090;
assign w6704 = ~w716 & ~w886;
assign w6705 = ~w633 & w1131;
assign w6706 = ~w633 & ~w6120;
assign w6707 = w1146 & w1103;
assign w6708 = ~w1146 & ~w1103;
assign w6709 = ~w1115 & ~w1113;
assign w6710 = w1115 & w1113;
assign w6711 = ~w1124 & w1156;
assign w6712 = w1158 & ~w1121;
assign w6713 = w1170 & ~w1161;
assign w6714 = ~w1088 & ~w633;
assign w6715 = w1178 & ~w633;
assign w6716 = w1178 & w6714;
assign w6717 = w1183 & ~w6716;
assign w6718 = w1183 & ~w6715;
assign w6719 = ~w1111 & ~w6718;
assign w6720 = ~w1111 & ~w6717;
assign w6721 = w1188 & ~w342;
assign w6722 = ~w1181 & w1188;
assign w6723 = ~w6721 & ~w1191;
assign w6724 = ~w403 & ~w342;
assign w6725 = ~w707 & w1209;
assign w6726 = ~w707 & w1215;
assign w6727 = ~w1218 & ~w1210;
assign w6728 = w1223 & ~w1221;
assign w6729 = w1223 & ~w306;
assign w6730 = ~w1206 & w1228;
assign w6731 = ~w1207 & ~w1229;
assign w6732 = ~w1200 & w1188;
assign w6733 = w1242 & w1246;
assign w6734 = ~w810 & w738;
assign w6735 = ~w306 & w1221;
assign w6736 = w1294 & ~w1257;
assign w6737 = ~w1312 & w734;
assign w6738 = w1314 & w1317;
assign w6739 = ~w1183 & w6716;
assign w6740 = ~w1183 & w6715;
assign w6741 = ~w1317 & w1321;
assign w6742 = ~w734 & ~w1322;
assign w6743 = w1348 & w1356;
assign w6744 = ~w1251 & ~w259;
assign w6745 = ~w1249 & ~w1317;
assign w6746 = w1249 & w1317;
assign w6747 = w1428 & ~w1426;
assign w6748 = w1432 & w1088;
assign w6749 = ~w1438 & ~w1435;
assign w6750 = ~w1439 & ~w180;
assign w6751 = ~w1314 & ~w1251;
assign w6752 = ~w6138 & w1088;
assign w6753 = w1474 & w1478;
assign w6754 = w1385 & ~w1377;
assign w6755 = ~w103 & ~w1088;
assign w6756 = ~w103 & ~w1510;
assign w6757 = ~w1523 & w1515;
assign w6758 = w1523 & ~w1515;
assign w6759 = ~w1488 & ~w1385;
assign w6760 = ~w1540 & ~w1499;
assign w6761 = ~w1446 & ~w1444;
assign w6762 = w1383 & w1325;
assign w6763 = w1194 & w1325;
assign w6764 = w1194 & w6762;
assign w6765 = w1322 & w1194;
assign w6766 = ~w1551 & ~w6763;
assign w6767 = ~w1551 & ~w6764;
assign w6768 = ~w1192 & ~w6766;
assign w6769 = ~w1192 & ~w6767;
assign w6770 = ~w1190 & ~w886;
assign w6771 = ~w1322 & ~w1194;
assign w6772 = ~w1383 & ~w1325;
assign w6773 = ~w1547 & ~w1444;
assign w6774 = ~w1547 & w6761;
assign w6775 = w403 & ~w1012;
assign w6776 = ~w403 & ~w1595;
assign w6777 = w403 & w1595;
assign w6778 = ~w1591 & ~w1598;
assign w6779 = ~w403 & ~w1584;
assign w6780 = w342 & w1616;
assign w6781 = w301 & ~w1617;
assign w6782 = ~w342 & w1594;
assign w6783 = w342 & ~w1594;
assign w6784 = w1619 & ~w1618;
assign w6785 = ~w342 & ~w1631;
assign w6786 = ~w1630 & ~w1631;
assign w6787 = ~w1630 & w6785;
assign w6788 = w1633 & ~w1627;
assign w6789 = w1591 & w1598;
assign w6790 = w1638 & ~w1636;
assign w6791 = w1435 & ~w1487;
assign w6792 = w1649 & ~w1643;
assign w6793 = w1611 & ~w1601;
assign w6794 = ~w403 & ~w1606;
assign w6795 = w1669 & ~w1654;
assign w6796 = ~w1655 & ~w1664;
assign w6797 = ~w403 & ~w1659;
assign w6798 = w1689 & ~w1674;
assign w6799 = w1675 & ~w1684;
assign w6800 = ~w1710 & ~w1695;
assign w6801 = ~w403 & ~w1700;
assign w6802 = w403 & w1722;
assign w6803 = ~w403 & ~w1722;
assign w6804 = ~w1696 & ~w1705;
assign w6805 = ~w1716 & ~w1564;
assign w6806 = w1716 & w1563;
assign w6807 = ~w1719 & ~w1727;
assign w6808 = ~w1734 & w1561;
assign w6809 = ~w1736 & ~w1746;
assign w6810 = w1570 & w1737;
assign w6811 = ~w1720 & w1570;
assign w6812 = ~w1758 & ~w1737;
assign w6813 = ~w1758 & ~w6810;
assign w6814 = w1734 & ~w1769;
assign w6815 = ~w1753 & ~w1775;
assign w6816 = w1753 & w1774;
assign w6817 = ~w1754 & ~w1763;
assign w6818 = ~w1566 & ~w1737;
assign w6819 = ~w1566 & ~w6810;
assign w6820 = ~w1783 & ~w1781;
assign w6821 = w1783 & w1781;
assign w6822 = w220 & ~w301;
assign w6823 = ~w1805 & ~w1631;
assign w6824 = w1804 & w948;
assign w6825 = w1806 & ~w1808;
assign w6826 = w1820 & ~w1818;
assign w6827 = w1827 & ~w1825;
assign w6828 = ~w1833 & w1800;
assign w6829 = w1833 & ~w1800;
assign w6830 = w1840 & ~w1839;
assign w6831 = ~w1844 & w1798;
assign w6832 = w1844 & ~w1798;
assign w6833 = w1850 & w1797;
assign w6834 = ~w1850 & ~w1797;
assign w6835 = w1856 & w1796;
assign w6836 = ~w1856 & ~w1796;
assign w6837 = w1870 & ~w1864;
assign w6838 = ~w1876 & ~w1875;
assign w6839 = ~w1807 & w1896;
assign w6840 = w220 & w1806;
assign w6841 = w1806 & ~w1900;
assign w6842 = w1918 & w1890;
assign w6843 = ~w1918 & ~w1890;
assign w6844 = w1924 & w1889;
assign w6845 = ~w1924 & ~w1889;
assign w6846 = w1930 & w1568;
assign w6847 = ~w1930 & ~w1937;
assign w6848 = ~w1936 & ~w1945;
assign w6849 = w1936 & w1566;
assign w6850 = w1949 & ~w1946;
assign w6851 = w1951 & w1561;
assign w6852 = ~w1951 & ~w1961;
assign w6853 = w1958 & w1774;
assign w6854 = ~w1958 & ~w1966;
assign w6855 = ~w1192 & w1553;
assign w6856 = w1556 & ~w1971;
assign w6857 = ~w1981 & ~w253;
assign w6858 = w1782 & ~w1984;
assign w6859 = w1559 & ~w403;
assign w6860 = ~w1779 & ~w1787;
assign w6861 = ~w1995 & w1994;
assign w6862 = w1995 & ~w1994;
assign w6863 = w1776 & w1556;
assign w6864 = w1776 & ~w301;
assign w6865 = ~w1993 & ~w1983;
assign w6866 = w253 & ~w1804;
assign w6867 = ~w2017 & ~w1804;
assign w6868 = w1807 & w301;
assign w6869 = w1896 & w253;
assign w6870 = w1896 & ~w6412;
assign w6871 = w2026 & ~w2027;
assign w6872 = ~w2028 & ~w2025;
assign w6873 = w2035 & ~w2034;
assign w6874 = ~w2035 & w2034;
assign w6875 = ~w2058 & ~w2054;
assign w6876 = w2065 & ~w2061;
assign w6877 = ~w2070 & ~w2068;
assign w6878 = w1804 & w254;
assign w6879 = ~w2018 & ~w2088;
assign w6880 = ~w2129 & w2086;
assign w6881 = w2129 & ~w2086;
assign w6882 = w2134 & w2141;
assign w6883 = w2140 & w2145;
assign w6884 = ~w2148 & w2084;
assign w6885 = w2148 & ~w2084;
assign w6886 = ~w2154 & ~w2083;
assign w6887 = w2154 & w2083;
assign w6888 = w2160 & ~w2166;
assign w6889 = ~w2160 & w1563;
assign w6890 = ~w103 & w516;
assign w6891 = w2187 & w2201;
assign w6892 = ~w1525 & ~w103;
assign w6893 = ~w103 & w1532;
assign w6894 = w1576 & ~w2223;
assign w6895 = ~w2232 & ~w2228;
assign w6896 = ~w2237 & w2243;
assign w6897 = w2176 & ~w1560;
assign w6898 = w2175 & ~w2280;
assign w6899 = ~w2176 & ~w2173;
assign w6900 = w2175 & w2283;
assign w6901 = ~w2284 & ~w2172;
assign w6902 = w2173 & ~w1192;
assign w6903 = w2287 & w2010;
assign w6904 = w2167 & ~w2289;
assign w6905 = ~w2167 & w1561;
assign w6906 = ~w2079 & ~w2075;
assign w6907 = ~w2173 & ~w2010;
assign w6908 = w2307 & ~w2288;
assign w6909 = w2301 & ~w2295;
assign w6910 = ~w2290 & w1774;
assign w6911 = w2290 & ~w2325;
assign w6912 = w2330 & ~w2313;
assign w6913 = w2320 & ~w2316;
assign w6914 = w2324 & ~w1556;
assign w6915 = ~w2324 & ~w2346;
assign w6916 = ~w103 & ~w2352;
assign w6917 = w2335 & ~w2339;
assign w6918 = ~w2348 & ~w2345;
assign w6919 = ~w2200 & ~w2185;
assign w6920 = w1525 & ~w364;
assign w6921 = ~w1525 & ~w364;
assign w6922 = w2441 & ~w2384;
assign w6923 = ~w2441 & w2384;
assign w6924 = w2450 & ~w2449;
assign w6925 = ~w2381 & ~w2460;
assign w6926 = ~w2381 & w2463;
assign w6927 = w2381 & w2460;
assign w6928 = w2381 & ~w2463;
assign w6929 = w2481 & ~w2377;
assign w6930 = ~w364 & ~w1192;
assign w6931 = ~w1774 & ~w2490;
assign w6932 = w2487 & w2495;
assign w6933 = ~w2487 & ~w1556;
assign w6934 = ~w2499 & ~w2498;
assign w6935 = w301 & w2510;
assign w6936 = pi00 & w95;
assign w6937 = pi01 & w31;
assign w6938 = w23 & w89;
assign w6939 = ~pi19 & pi07;
assign w6940 = w10 & w2530;
assign w6941 = ~w1525 & ~w2531;
assign w6942 = w1525 & ~w2531;
assign w6943 = w2545 & w103;
assign w6944 = ~w2537 & w2591;
assign w6945 = ~w2606 & ~w2602;
assign w6946 = ~w2618 & w2535;
assign w6947 = ~w1561 & ~w1988;
assign w6948 = ~w2637 & ~w2628;
assign w6949 = w2640 & w2533;
assign w6950 = ~w2640 & ~w2533;
assign w6951 = w2499 & w2498;
assign w6952 = ~w2646 & w2654;
assign w6953 = ~w2646 & ~w2532;
assign w6954 = pi00 & w31;
assign w6955 = pi15 & pi04;
assign w6956 = ~pi19 & pi06;
assign w6957 = ~w2677 & ~w10;
assign w6958 = ~w2512 & ~w2679;
assign w6959 = ~w2531 & w364;
assign w6960 = ~w1509 & ~w2531;
assign w6961 = w2546 & ~w2554;
assign w6962 = ~w2679 & w1532;
assign w6963 = w103 & ~w2679;
assign w6964 = ~w103 & ~w2679;
assign w6965 = w2770 & w2773;
assign w6966 = ~w2762 & ~w2772;
assign w6967 = ~w2793 & w2790;
assign w6968 = w2793 & ~w2790;
assign w6969 = ~w2795 & ~w2807;
assign w6970 = ~w2808 & w2684;
assign w6971 = ~w2797 & w2807;
assign w6972 = w2796 & w2812;
assign w6973 = w2683 & w2818;
assign w6974 = ~w2820 & w2815;
assign w6975 = w2825 & w2833;
assign w6976 = w2825 & ~w2680;
assign w6977 = ~pi19 & pi05;
assign w6978 = pi15 & pi03;
assign w6979 = ~w2853 & ~w10;
assign w6980 = ~w103 & w2854;
assign w6981 = w103 & w2854;
assign w6982 = w2872 & w2531;
assign w6983 = w2875 & ~w2874;
assign w6984 = w2545 & w2679;
assign w6985 = ~w2882 & w2854;
assign w6986 = w2892 & w2871;
assign w6987 = ~w2892 & ~w2871;
assign w6988 = w2905 & ~w2904;
assign w6989 = ~w2940 & ~w2936;
assign w6990 = ~w2999 & w2996;
assign w6991 = ~w2857 & ~w3004;
assign w6992 = ~pi19 & pi04;
assign w6993 = pi15 & pi02;
assign w6994 = ~w3019 & ~w3024;
assign w6995 = w2872 & ~w2531;
assign w6996 = ~w3029 & w2872;
assign w6997 = ~w2854 & ~w3058;
assign w6998 = w3061 & ~w3057;
assign w6999 = ~w3029 & w1532;
assign w7000 = ~w3042 & w3078;
assign w7001 = w3042 & ~w3078;
assign w7002 = w103 & ~w3029;
assign w7003 = ~w103 & ~w3029;
assign w7004 = ~w3079 & ~w3094;
assign w7005 = w3079 & w3094;
assign w7006 = ~w3099 & w3041;
assign w7007 = w3088 & w3095;
assign w7008 = ~w3126 & ~w3115;
assign w7009 = ~w2512 & ~w3029;
assign w7010 = ~w3152 & ~w3161;
assign w7011 = ~w3190 & w3192;
assign w7012 = w3184 & w3193;
assign w7013 = pi15 & pi00;
assign w7014 = ~pi19 & pi02;
assign w7015 = ~w3202 & ~w3199;
assign w7016 = ~pi19 & pi03;
assign w7017 = pi15 & pi01;
assign w7018 = ~w3217 & ~w3212;
assign w7019 = w3029 & ~w2872;
assign w7020 = ~w3029 & w1012;
assign w7021 = ~w3229 & ~w3228;
assign w7022 = w3229 & ~w3222;
assign w7023 = w3245 & ~w3239;
assign w7024 = ~w3247 & w3257;
assign w7025 = w3247 & ~w3257;
assign w7026 = w3099 & ~w3041;
assign w7027 = ~w3288 & ~w3224;
assign w7028 = w3305 & ~w3223;
assign w7029 = w3288 & w1563;
assign w7030 = ~w3311 & ~w3310;
assign w7031 = ~w3314 & ~w3307;
assign w7032 = ~w3305 & w3223;
assign w7033 = ~w3313 & w3317;
assign w7034 = ~w3326 & ~w3333;
assign w7035 = w3326 & ~w1556;
assign w7036 = ~w3222 & w1553;
assign w7037 = w3339 & ~w3336;
assign w7038 = ~w1584 & ~w3222;
assign w7039 = ~w7038 & ~w1012;
assign w7040 = w3029 & ~w3367;
assign w7041 = w3374 & ~w3373;
assign w7042 = w3384 & w1648;
assign w7043 = ~w3384 & ~w1648;
assign w7044 = w3363 & w3394;
assign w7045 = ~w3401 & ~w3402;
assign w7046 = w3277 & w3357;
assign w7047 = ~w3414 & ~w3355;
assign w7048 = ~w1559 & ~w3205;
assign w7049 = ~w3207 & ~w3206;
assign w7050 = ~w3455 & ~w3458;
assign w7051 = w3334 & w3455;
assign w7052 = w3335 & ~w3465;
assign w7053 = ~w3197 & ~w3195;
assign w7054 = ~w3015 & ~w3013;
assign w7055 = ~w3480 & ~w2838;
assign w7056 = ~w2661 & ~w2659;
assign w7057 = w141 & w2367;
assign w7058 = ~w177 & ~w3493;
assign w7059 = w3499 & w3508;
assign w7060 = ~w3499 & ~w3508;
assign w7061 = ~w3512 & w3514;
assign w7062 = w2008 & ~w1086;
assign w7063 = ~w2374 & ~w3486;
assign w7064 = ~w6203 & w3207;
assign w7065 = ~w3205 & w7381;
assign w7066 = ~w3538 & ~w3539;
assign w7067 = ~w3526 & ~w3528;
assign w7068 = w2372 & w3501;
assign w7069 = ~w2372 & ~w3501;
assign w7070 = ~w3516 & w1012;
assign w7071 = ~w6206 & ~w1576;
assign w7072 = w3612 & w3613;
assign w7073 = ~w1572 & ~w3626;
assign w7074 = w3612 & w3628;
assign w7075 = w1572 & w1542;
assign w7076 = w3633 & w1648;
assign w7077 = ~w3635 & ~w3634;
assign w7078 = w1576 & w3612;
assign w7079 = ~w1576 & ~w3612;
assign w7080 = w1590 & ~w3646;
assign w7081 = ~w1590 & w3646;
assign w7082 = w1590 & w3650;
assign w7083 = w1576 & ~w3657;
assign w7084 = w3642 & ~w3601;
assign w7085 = ~w3623 & w3621;
assign w7086 = w3638 & ~w3667;
assign w7087 = ~w3635 & ~w3629;
assign w7088 = w1570 & w1568;
assign w7089 = w3632 & ~w3676;
assign w7090 = ~w1570 & ~w3678;
assign w7091 = w3676 & ~w3632;
assign w7092 = ~w1572 & w3683;
assign w7093 = w1572 & ~w3683;
assign w7094 = w3672 & w3686;
assign w7095 = w1648 & ~w3703;
assign w7096 = w1572 & w3678;
assign w7097 = w1572 & ~w6215;
assign w7098 = w1572 & ~w3677;
assign w7099 = w1572 & w6216;
assign w7100 = ~w1568 & w3712;
assign w7101 = w1568 & ~w3712;
assign w7102 = ~w3730 & w3735;
assign w7103 = ~w3709 & w3707;
assign w7104 = w3721 & ~w3747;
assign w7105 = w7101 & w3626;
assign w7106 = ~w1570 & ~w3752;
assign w7107 = ~w1570 & ~w3755;
assign w7108 = w3712 & w1568;
assign w7109 = w7108 & ~w1563;
assign w7110 = ~w3712 & w3762;
assign w7111 = ~w3762 & w1566;
assign w7112 = ~w1590 & ~w3650;
assign w7113 = w1579 & ~w3804;
assign w7114 = ~w1579 & w3807;
assign w7115 = ~w1579 & w3804;
assign w7116 = ~w3815 & ~w3818;
assign w7117 = w3656 & w3659;
assign w7118 = ~w3829 & ~w3800;
assign w7119 = w3829 & w3800;
assign w7120 = w3815 & w3818;
assign w7121 = w3526 & w3365;
assign w7122 = w1579 & ~w3807;
assign w7123 = ~w3862 & ~w3860;
assign w7124 = w3887 & w3853;
assign w7125 = ~w3887 & ~w3853;
assign w7126 = w3895 & w3594;
assign w7127 = ~w3895 & ~w3903;
assign w7128 = w3904 & ~w3902;
assign w7129 = w3712 & w3427;
assign w7130 = ~w3592 & w3907;
assign w7131 = w3918 & ~w3992;
assign w7132 = ~w3918 & w3992;
assign w7133 = w1561 & ~w1192;
assign w7134 = w7133 & ~w1563;
assign w7135 = ~w3762 & w1561;
assign w7136 = w1563 & ~w4033;
assign w7137 = ~w1563 & w4033;
assign w7138 = ~w1576 & ~w3568;
assign w7139 = ~w1576 & w3568;
assign w7140 = ~w6444 & w4102;
assign w7141 = w4012 & w4103;
assign w7142 = w4013 & w4105;
assign w7143 = w1563 & w1192;
assign w7144 = w1561 & w4130;
assign w7145 = ~w1563 & w4132;
assign w7146 = w3526 & w4137;
assign w7147 = w7133 & w3526;
assign w7148 = ~w4138 & w4140;
assign w7149 = w4075 & w3986;
assign w7150 = w4075 & w6527;
assign w7151 = ~w4190 & w3589;
assign w7152 = ~w4207 & ~w4097;
assign w7153 = ~w4207 & w6446;
assign w7154 = ~w4006 & ~w4207;
assign w7155 = w1556 & ~w4247;
assign w7156 = ~w1774 & w4248;
assign w7157 = ~w4191 & ~w3586;
assign w7158 = w4191 & w3586;
assign w7159 = w4284 & ~w4295;
assign w7160 = w4302 & w4279;
assign w7161 = ~w4171 & ~w4206;
assign w7162 = ~w4225 & ~w4322;
assign w7163 = w4227 & w4325;
assign w7164 = w1556 & ~w4135;
assign w7165 = ~w3989 & ~w3982;
assign w7166 = w3989 & w3982;
assign w7167 = ~w1579 & w3526;
assign w7168 = w1579 & ~w1584;
assign w7169 = w3603 & ~w4458;
assign w7170 = w3600 & ~w4460;
assign w7171 = ~w4463 & ~w3733;
assign w7172 = w4463 & w3733;
assign w7173 = w3594 & w3591;
assign w7174 = w4476 & ~w3591;
assign w7175 = ~w4486 & w1012;
assign w7176 = w3911 & w4490;
assign w7177 = w4420 & w4414;
assign w7178 = ~w4420 & ~w4414;
assign w7179 = w4304 & ~w4301;
assign w7180 = ~w4313 & w7460;
assign w7181 = w4309 & w4307;
assign w7182 = ~w1648 & ~w3518;
assign w7183 = ~w4388 & ~w3911;
assign w7184 = ~w4391 & w4538;
assign w7185 = (w4532 & w4216) | (w4532 & w7461) | (w4216 & w7461);
assign w7186 = ~w4539 & w4542;
assign w7187 = ~w4388 & ~w4546;
assign w7188 = w4391 & w4549;
assign w7189 = ~w4323 & w4552;
assign w7190 = w4326 & w4553;
assign w7191 = ~w1556 & ~w3610;
assign w7192 = ~w1556 & ~w6256;
assign w7193 = ~w3516 & ~w1584;
assign w7194 = w1579 & ~w4634;
assign w7195 = ~w1579 & ~w4634;
assign w7196 = ~w3516 & ~w1579;
assign w7197 = ~w4518 & w4668;
assign w7198 = w4623 & ~w4677;
assign w7199 = w4546 & w3985;
assign w7200 = ~w4684 & ~w4685;
assign w7201 = ~w4546 & ~w4683;
assign w7202 = w4550 & w4687;
assign w7203 = ~w4692 & ~w4691;
assign w7204 = ~w3526 & w3529;
assign w7205 = ~w4533 & w4768;
assign w7206 = ~w3580 & w7508;
assign w7207 = w4657 & w4798;
assign w7208 = ~w3516 & w1590;
assign w7209 = ~w4680 & ~w4816;
assign w7210 = ~w4678 & w4817;
assign w7211 = ~w4686 & w4828;
assign w7212 = ~w4689 & w4831;
assign w7213 = ~w4705 & ~w4842;
assign w7214 = w1566 & w3568;
assign w7215 = w3594 & w3568;
assign w7216 = ~w3516 & w50;
assign w7217 = w2008 & ~w2513;
assign w7218 = w4799 & w4933;
assign w7219 = ~w4807 & w3581;
assign w7220 = ~w3516 & ~w1576;
assign w7221 = w4818 & w4946;
assign w7222 = ~w4948 & ~w4949;
assign w7223 = ~w4952 & w4910;
assign w7224 = (w4823 & w7462) | (w4823 & w7463) | (w7462 & w7463);
assign w7225 = w4952 & ~w4910;
assign w7226 = w6473 & w3588;
assign w7227 = (w3588 & w6473) | (w3588 & w4689) | (w6473 & w4689);
assign w7228 = w3591 & w4856;
assign w7229 = (w3591 & ~w4749) | (w3591 & w7464) | (~w4749 & w7464);
assign w7230 = w4855 & w5025;
assign w7231 = (w4749 & w7465) | (w4749 & w7466) | (w7465 & w7466);
assign w7232 = w4857 & w5028;
assign w7233 = w4811 & w4781;
assign w7234 = w1584 & ~w4634;
assign w7235 = ~w4665 & w1579;
assign w7236 = ~w3516 & ~w1648;
assign w7237 = ~w4954 & w5101;
assign w7238 = ~w4985 & w5123;
assign w7239 = (~w5123 & w4987) | (~w5123 & w7467) | (w4987 & w7467);
assign w7240 = ~w5123 & ~w5033;
assign w7241 = w5166 & ~w5162;
assign w7242 = ~w5086 & w4811;
assign w7243 = w4811 & ~w5216;
assign w7244 = w4954 & w5101;
assign w7245 = ~w4963 & w3581;
assign w7246 = ~w5117 & w7468;
assign w7247 = ~w5235 & w5176;
assign w7248 = w5142 & ~w5261;
assign w7249 = w5288 & w5280;
assign w7250 = ~w5288 & ~w5280;
assign w7251 = w4811 & w5326;
assign w7252 = (w6572 & w7469) | (w6572 & w7470) | (w7469 & w7470);
assign w7253 = (~w6572 & w7471) | (~w6572 & w7472) | (w7471 & w7472);
assign w7254 = ~w5225 & ~w3581;
assign w7255 = ~w5300 & w5335;
assign w7256 = ~w3516 & w1570;
assign w7257 = w5356 & ~w5391;
assign w7258 = (w4948 & ~w5049) | (w4948 & w7473) | (~w5049 & w7473);
assign w7259 = w1648 & w3581;
assign w7260 = w1648 & w6471;
assign w7261 = ~w5416 & ~w5415;
assign w7262 = ~w5418 & ~w5412;
assign w7263 = w5329 & ~w5421;
assign w7264 = ~w5329 & w5421;
assign w7265 = ~w5212 & ~w5215;
assign w7266 = ~w5297 & w5339;
assign w7267 = w1566 & ~w3579;
assign w7268 = w5357 & ~w3579;
assign w7269 = ~w5357 & ~w5460;
assign w7270 = w1774 & w3985;
assign w7271 = w1774 & ~w6277;
assign w7272 = w5380 & ~w5465;
assign w7273 = w5380 & ~w5379;
assign w7274 = w5257 & ~w5468;
assign w7275 = w5375 & ~w4486;
assign w7276 = w5372 & ~w5477;
assign w7277 = ~w5466 & w5486;
assign w7278 = w5466 & ~w5486;
assign w7279 = w5386 & ~w5387;
assign w7280 = ~w3516 & w1568;
assign w7281 = ~w5456 & ~w5493;
assign w7282 = ~w5483 & w5465;
assign w7283 = ~w5483 & ~w7272;
assign w7284 = ~w5564 & ~w5565;
assign w7285 = ~w1561 & w4075;
assign w7286 = ~w6494 & w5473;
assign w7287 = ~w5562 & ~w5586;
assign w7288 = w5562 & w5586;
assign w7289 = ~w3516 & w1566;
assign w7290 = ~w5561 & w5593;
assign w7291 = w5561 & ~w5593;
assign w7292 = w5596 & w5553;
assign w7293 = w5596 & w5455;
assign w7294 = ~w5596 & ~w5553;
assign w7295 = ~w5596 & ~w5455;
assign w7296 = ~w5532 & ~w5625;
assign w7297 = w5532 & w5625;
assign w7298 = w5224 & w4933;
assign w7299 = ~w5224 & ~w5634;
assign w7300 = w5542 & ~w5636;
assign w7301 = ~w5555 & ~w5589;
assign w7302 = ~w3516 & w1563;
assign w7303 = ~w5564 & ~w5659;
assign w7304 = w5564 & w4075;
assign w7305 = w5662 & w3588;
assign w7306 = ~w5668 & ~w5574;
assign w7307 = ~w5668 & ~w6278;
assign w7308 = ~w5667 & w7307;
assign w7309 = ~w5667 & w7306;
assign w7310 = w5663 & ~w5658;
assign w7311 = ~w5674 & ~w5677;
assign w7312 = w5623 & ~w5624;
assign w7313 = ~w5545 & w5339;
assign w7314 = w5701 & ~w5725;
assign w7315 = ~w5678 & w5658;
assign w7316 = ~w5682 & ~w5735;
assign w7317 = ~w3516 & w1561;
assign w7318 = w5671 & ~w5738;
assign w7319 = ~w5671 & w3585;
assign w7320 = w3985 & w5667;
assign w7321 = ~w4075 & ~w5574;
assign w7322 = ~w4075 & ~w6278;
assign w7323 = w5743 & ~w5742;
assign w7324 = w5736 & ~w5749;
assign w7325 = w5742 & ~w7321;
assign w7326 = w5742 & ~w7322;
assign w7327 = ~w5799 & ~w7326;
assign w7328 = ~w5799 & ~w7325;
assign w7329 = w6284 | w5745;
assign w7330 = (w5745 & w6284) | (w5745 & w5671) | (w6284 & w5671);
assign w7331 = ~w3516 & w1774;
assign w7332 = w5844 & ~w5840;
assign w7333 = w5754 & w5861;
assign w7334 = w5813 & ~w5737;
assign w7335 = w5807 & w5804;
assign w7336 = ~w3581 & ~w5804;
assign w7337 = w7336 & w5871;
assign w7338 = ~w3516 & ~w1556;
assign w7339 = ~w7336 & ~w5876;
assign w7340 = w5816 & w5879;
assign w7341 = ~w5819 & w3581;
assign w7342 = ~w5831 & w5893;
assign w7343 = w7335 & ~w5876;
assign w7344 = ~w3516 & ~w50;
assign w7345 = ~w5873 & ~w5869;
assign w7346 = w5877 & ~w5911;
assign w7347 = ~w5816 & w5922;
assign w7348 = ~w5925 & w1563;
assign w7349 = ~w5857 & w4933;
assign w7350 = ~w5882 & w5928;
assign w7351 = ~w1563 & w5926;
assign w7352 = ~w5887 & ~w5854;
assign w7353 = ~w5853 & ~w5934;
assign w7354 = ~w5853 & ~w5858;
assign w7355 = ~w5880 & ~w5922;
assign w7356 = ~w5941 & ~w5864;
assign w7357 = ~w5624 & ~w5953;
assign w7358 = ~w5948 & ~w5933;
assign w7359 = ~w5941 & ~w5858;
assign w7360 = w3516 & ~w1561;
assign w7361 = ~w4933 & w5971;
assign w7362 = w5978 & w5976;
assign w7363 = ~w5978 & ~w5976;
assign w7364 = w5933 & w5983;
assign w7365 = ~w1774 & w5737;
assign w7366 = w3516 & ~w1774;
assign w7367 = ~w1774 & ~w5989;
assign w7368 = ~w4933 & ~w1563;
assign w7369 = w5933 & w6298;
assign w7370 = w6299 & w5997;
assign w7371 = (w5997 & w6299) | (w5997 & ~w5933) | (w6299 & ~w5933);
assign w7372 = ~w5979 & w6000;
assign w7373 = ~w1774 & ~w5737;
assign w7374 = ~w5990 & ~w6010;
assign w7375 = w6011 & w5959;
assign w7376 = w6011 & ~w6296;
assign w7377 = w5992 & w6010;
assign w7378 = w7362 & w6014;
assign w7379 = w5978 & w6018;
assign w7380 = w5933 & w6020;
assign w7381 = ~w1556 & ~w1086;
assign w7382 = ~w6004 & w6028;
assign w7383 = ~w5990 & ~w6008;
assign w7384 = w6030 & w6008;
assign w7385 = w6030 & ~w7383;
assign w7386 = w7362 & w6032;
assign w7387 = ~w5988 & ~w6028;
assign w7388 = w6302 & w6035;
assign w7389 = (w6035 & w6302) | (w6035 & ~w5933) | (w6302 & ~w5933);
assign w7390 = ~w6033 & ~w6037;
assign w7391 = w5960 & w6039;
assign w7392 = ~w6004 & ~w6028;
assign w7393 = w5960 & w6043;
assign w7394 = pi10 & pi02;
assign w7395 = ~w183 & ~w10;
assign w7396 = w247 & ~w10;
assign w7397 = w6308 & w675;
assign w7398 = w6308 & ~w6628;
assign w7399 = w2120 & ~w141;
assign w7400 = w1523 & ~w2185;
assign w7401 = ~w103 & ~w6144;
assign w7402 = ~w2966 & ~w2996;
assign w7403 = w2854 & w7510;
assign w7404 = w3149 & w3030;
assign w7405 = ~w1561 & ~w3030;
assign w7406 = ~w1568 & ~w3285;
assign w7407 = ~w3398 & w3402;
assign w7408 = ~w3415 & w3352;
assign w7409 = w3415 & ~w3352;
assign w7410 = w3415 & w3425;
assign w7411 = ~w3415 & w3428;
assign w7412 = w3205 & ~w3207;
assign w7413 = ~w1572 & w1648;
assign w7414 = ~w1648 & ~w3615;
assign w7415 = ~w3617 & ~w3620;
assign w7416 = ~w1568 & ~w1542;
assign w7417 = ~w3676 & ~w1570;
assign w7418 = ~w7121 & ~w1584;
assign w7419 = ~w1561 & ~w1563;
assign w7420 = w3946 & ~w3947;
assign w7421 = ~w4031 & ~w4030;
assign w7422 = w1556 & ~w1774;
assign w7423 = w1774 | w6325;
assign w7424 = w3205 & w1086;
assign w7425 = ~w1774 & ~w5248;
assign w7426 = w6266 & w3985;
assign w7427 = ~w6266 & ~w5286;
assign w7428 = w4075 & w3985;
assign w7429 = w4075 & w6272;
assign w7430 = ~w5508 & ~w5786;
assign w7431 = ~w6083 & w529;
assign w7432 = w530 & w538;
assign w7433 = w540 & w541;
assign w7434 = w6360 & ~w511;
assign w7435 = (~w511 & w6360) | (~w511 & w543) | (w6360 & w543);
assign w7436 = ~w543 & w6361;
assign w7437 = w1360 & w1369;
assign w7438 = w1590 & ~w3063;
assign w7439 = w4954 & w5102;
assign w7440 = ~w5224 & ~w5227;
assign w7441 = ~w6477 & w3588;
assign w7442 = ~w6269 & ~w5150;
assign w7443 = w3568 & w6270;
assign w7444 = w5216 & w5327;
assign w7445 = ~w2553 & ~w2531;
assign w7446 = w3446 & w3450;
assign w7447 = w4680 & w3585;
assign w7448 = w5115 & w5339;
assign w7449 = ~w5256 & ~w5366;
assign w7450 = ~w5437 & ~w4948;
assign w7451 = ~w5437 & w6486;
assign w7452 = w6452 & ~w4317;
assign w7453 = ~w6452 & w4317;
assign w7454 = ~w4528 & ~w4676;
assign w7455 = w4962 & w3585;
assign w7456 = ~w6557 & ~w5108;
assign w7457 = ~w6567 & w3581;
assign w7458 = w1570 & w7511;
assign w7459 = ~w5112 & ~w5230;
assign w7460 = w4314 & ~w4521;
assign w7461 = ~w6452 & w4532;
assign w7462 = ~w1648 & w7511;
assign w7463 = w4952 & w6465;
assign w7464 = ~w6327 & w3591;
assign w7465 = ~w5027 & ~w3594;
assign w7466 = ~w5027 & ~w6326;
assign w7467 = w4985 & ~w5123;
assign w7468 = w6477 & ~w5235;
assign w7469 = ~w5101 & ~w5221;
assign w7470 = ~w5101 & w5105;
assign w7471 = w5101 & w5221;
assign w7472 = w5101 & ~w5105;
assign w7473 = ~w3581 & w4948;
assign w7474 = (w511 & ~w6360) | (w511 & ~w546) | (~w6360 & ~w546);
assign w7475 = (w1230 & w1233) | (w1230 & ~w6126) | (w1233 & ~w6126);
assign w7476 = (w1231 & ~w1202) | (w1231 & w6387) | (~w1202 & w6387);
assign w7477 = (w633 & ~w6714) | (w633 & ~w1172) | (~w6714 & ~w1172);
assign w7478 = (~w1356 & ~w6743) | (~w1356 & ~w1355) | (~w6743 & ~w1355);
assign w7479 = (w1444 & ~w6761) | (w1444 & ~w1544) | (~w6761 & ~w1544);
assign w7480 = (w886 & ~w6770) | (w886 & ~w1189) | (~w6770 & ~w1189);
assign w7481 = ~w1551 & ~w1550;
assign w7482 = (w1500 & ~w103) | (w1500 & w6893) | (~w103 & w6893);
assign w7483 = (w2586 & ~w2591) | (w2586 & ~w6162) | (~w2591 & ~w6162);
assign w7484 = (w2587 & ~w2537) | (w2587 & w6944) | (~w2537 & w6944);
assign w7485 = (w1500 & ~w2679) | (w1500 & w6962) | (~w2679 & w6962);
assign w7486 = (w1500 & ~w3029) | (w1500 & w6999) | (~w3029 & w6999);
assign w7487 = (w3279 & ~w3277) | (w3279 & ~w6188) | (~w3277 & ~w6188);
assign w7488 = (w3367 & ~w7040) | (w3367 & ~w1579) | (~w7040 & ~w1579);
assign w7489 = (w2507 & w3486) | (w2507 & ~w6200) | (w3486 & ~w6200);
assign w7490 = (~w3484 & ~w2374) | (~w3484 & w7063) | (~w2374 & w7063);
assign w7491 = (w4200 & w4302) | (w4200 & w7160) | (w4302 & w7160);
assign w7492 = (w4670 & w4811) | (w4670 & w7233) | (w4811 & w7233);
assign w7493 = (w4824 & ~w4910) | (w4824 & ~w6472) | (~w4910 & ~w6472);
assign w7494 = (~w3594 & ~w6270) | (~w3594 & ~w5131) | (~w6270 & ~w5131);
assign w7495 = ~w5115 & ~w5231;
assign w7496 = (~w7307 & ~w7306) | (~w7307 & ~w5577) | (~w7306 & ~w5577);
assign w7497 = (~w7328 & ~w7327) | (~w7328 & ~w5577) | (~w7327 & ~w5577);
assign w7498 = w5742 & ~w5744;
assign w7499 = (~w5971 & ~w7361) | (~w5971 & ~w5961) | (~w7361 & ~w5961);
assign w7500 = (~w675 & w6628) | (~w675 & ~w681) | (w6628 & ~w681);
assign w7501 = w707 & ~w841;
assign w7502 = (w2187 & ~w103) | (w2187 & w7401) | (~w103 & w7401);
assign w7503 = w3597 & w3600;
assign w7504 = w3733 & w3597;
assign w7505 = ~w177 & ~w141;
assign w7506 = (w1502 & ~w6402) | (w1502 & ~w6403) | (~w6402 & ~w6403);
assign w7507 = w3594 & w3733;
assign w7508 = ~w3516 & w7070;
assign w7509 = w1566 & w1568;
assign w7510 = ~w1556 & w1774;
assign w7511 = w3585 & w3588;
assign w7512 = (w3588 & w6537) | (w3588 & ~w4282) | (w6537 & ~w4282);
assign w7513 = (w3594 & w7507) | (w3594 & ~w4226) | (w7507 & ~w4226);
assign w7514 = (w4825 & ~w4952) | (w4825 & w7223) | (~w4952 & w7223);
assign w7515 = (w1566 & w7509) | (w1566 & ~w2761) | (w7509 & ~w2761);
assign one = 1;
assign po00 = w51;// level 8
assign po01 = ~w59;// level 7
assign po02 = w64;// level 6
assign po03 = w65;// level 5
assign po04 = ~w25;// level 3
assign po05 = ~w4510;// level 127
assign po06 = w4656;// level 131
assign po07 = w4796;// level 132
assign po08 = w4928;// level 134
assign po09 = w5072;// level 136
assign po10 = w5203;// level 137
assign po11 = ~w5324;// level 139
assign po12 = w5433;// level 140
assign po13 = w5539;// level 141
assign po14 = w5628;// level 141
assign po15 = ~w5723;// level 142
assign po16 = w5783;// level 142
assign po17 = w5849;// level 142
assign po18 = ~w5904;// level 143
assign po19 = w5958;// level 143
assign po20 = w5987;// level 143
assign po21 = w6003;// level 143
assign po22 = w6025;// level 143
assign po23 = ~w6041;// level 143
assign po24 = ~w6046;// level 143
endmodule
