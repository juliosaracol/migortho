module top (
            a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27], a[28], a[29], a[30], a[31], a[32], a[33], a[34], a[35], a[36], a[37], a[38], a[39], a[40], a[41], a[42], a[43], a[44], a[45], a[46], a[47], a[48], a[49], a[50], a[51], a[52], a[53], a[54], a[55], a[56], a[57], a[58], a[59], a[60], a[61], a[62], a[63], b[0], b[1], b[2], b[3], b[4], b[5], b[6], b[7], b[8], b[9], b[10], b[11], b[12], b[13], b[14], b[15], b[16], b[17], b[18], b[19], b[20], b[21], b[22], b[23], b[24], b[25], b[26], b[27], b[28], b[29], b[30], b[31], b[32], b[33], b[34], b[35], b[36], b[37], b[38], b[39], b[40], b[41], b[42], b[43], b[44], b[45], b[46], b[47], b[48], b[49], b[50], b[51], b[52], b[53], b[54], b[55], b[56], b[57], b[58], b[59], b[60], b[61], b[62], b[63], 
            f[0], f[1], f[2], f[3], f[4], f[5], f[6], f[7], f[8], f[9], f[10], f[11], f[12], f[13], f[14], f[15], f[16], f[17], f[18], f[19], f[20], f[21], f[22], f[23], f[24], f[25], f[26], f[27], f[28], f[29], f[30], f[31], f[32], f[33], f[34], f[35], f[36], f[37], f[38], f[39], f[40], f[41], f[42], f[43], f[44], f[45], f[46], f[47], f[48], f[49], f[50], f[51], f[52], f[53], f[54], f[55], f[56], f[57], f[58], f[59], f[60], f[61], f[62], f[63], f[64], f[65], f[66], f[67], f[68], f[69], f[70], f[71], f[72], f[73], f[74], f[75], f[76], f[77], f[78], f[79], f[80], f[81], f[82], f[83], f[84], f[85], f[86], f[87], f[88], f[89], f[90], f[91], f[92], f[93], f[94], f[95], f[96], f[97], f[98], f[99], f[100], f[101], f[102], f[103], f[104], f[105], f[106], f[107], f[108], f[109], f[110], f[111], f[112], f[113], f[114], f[115], f[116], f[117], f[118], f[119], f[120], f[121], f[122], f[123], f[124], f[125], f[126], f[127]);
input a[0], a[1], a[2], a[3], a[4], a[5], a[6], a[7], a[8], a[9], a[10], a[11], a[12], a[13], a[14], a[15], a[16], a[17], a[18], a[19], a[20], a[21], a[22], a[23], a[24], a[25], a[26], a[27], a[28], a[29], a[30], a[31], a[32], a[33], a[34], a[35], a[36], a[37], a[38], a[39], a[40], a[41], a[42], a[43], a[44], a[45], a[46], a[47], a[48], a[49], a[50], a[51], a[52], a[53], a[54], a[55], a[56], a[57], a[58], a[59], a[60], a[61], a[62], a[63], b[0], b[1], b[2], b[3], b[4], b[5], b[6], b[7], b[8], b[9], b[10], b[11], b[12], b[13], b[14], b[15], b[16], b[17], b[18], b[19], b[20], b[21], b[22], b[23], b[24], b[25], b[26], b[27], b[28], b[29], b[30], b[31], b[32], b[33], b[34], b[35], b[36], b[37], b[38], b[39], b[40], b[41], b[42], b[43], b[44], b[45], b[46], b[47], b[48], b[49], b[50], b[51], b[52], b[53], b[54], b[55], b[56], b[57], b[58], b[59], b[60], b[61], b[62], b[63];
output f[0], f[1], f[2], f[3], f[4], f[5], f[6], f[7], f[8], f[9], f[10], f[11], f[12], f[13], f[14], f[15], f[16], f[17], f[18], f[19], f[20], f[21], f[22], f[23], f[24], f[25], f[26], f[27], f[28], f[29], f[30], f[31], f[32], f[33], f[34], f[35], f[36], f[37], f[38], f[39], f[40], f[41], f[42], f[43], f[44], f[45], f[46], f[47], f[48], f[49], f[50], f[51], f[52], f[53], f[54], f[55], f[56], f[57], f[58], f[59], f[60], f[61], f[62], f[63], f[64], f[65], f[66], f[67], f[68], f[69], f[70], f[71], f[72], f[73], f[74], f[75], f[76], f[77], f[78], f[79], f[80], f[81], f[82], f[83], f[84], f[85], f[86], f[87], f[88], f[89], f[90], f[91], f[92], f[93], f[94], f[95], f[96], f[97], f[98], f[99], f[100], f[101], f[102], f[103], f[104], f[105], f[106], f[107], f[108], f[109], f[110], f[111], f[112], f[113], f[114], f[115], f[116], f[117], f[118], f[119], f[120], f[121], f[122], f[123], f[124], f[125], f[126], f[127];
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771;
assign w0 = a[0] & b[0];
assign w1 = a[2] & w0;
assign w2 = a[1] & ~a[2];
assign w3 = ~a[1] & a[2];
assign w4 = ~w2 & ~w3;
assign w5 = a[0] & ~w4;
assign w6 = ~b[0] & b[1];
assign w7 = b[0] & ~b[1];
assign w8 = ~w6 & ~w7;
assign w9 = ~a[0] & a[1];
assign w10 = b[0] & w9;
assign w11 = a[0] & w4;
assign w12 = w4 & w24057;
assign w13 = (~w10 & ~w5) | (~w10 & w24058) | (~w5 & w24058);
assign w14 = w13 & w24059;
assign w15 = (w1 & ~w13) | (w1 & w24060) | (~w13 & w24060);
assign w16 = ~w14 & ~w15;
assign w17 = a[2] & ~w0;
assign w18 = w13 & w24061;
assign w19 = a[2] & ~w18;
assign w20 = ~b[2] & ~w6;
assign w21 = b[2] & w6;
assign w22 = ~w20 & ~w21;
assign w23 = w5 & w22;
assign w24 = ~a[0] & ~a[1];
assign w25 = a[2] & w24;
assign w26 = w24 & w24062;
assign w27 = b[1] & w9;
assign w28 = w4 & w24063;
assign w29 = ~w26 & ~w27;
assign w30 = ~w23 & w24064;
assign w31 = w19 & ~w30;
assign w32 = ~w19 & w30;
assign w33 = ~w31 & ~w32;
assign w34 = w18 & w30;
assign w35 = a[2] & ~a[3];
assign w36 = ~a[2] & a[3];
assign w37 = ~w35 & ~w36;
assign w38 = b[0] & ~w37;
assign w39 = w4 & w24065;
assign w40 = b[2] & w9;
assign w41 = ~b[1] & ~b[3];
assign w42 = b[1] & b[3];
assign w43 = ~w41 & ~w42;
assign w44 = ~w20 & w43;
assign w45 = w20 & ~w43;
assign w46 = ~w44 & ~w45;
assign w47 = w5 & w46;
assign w48 = ~w39 & ~w40;
assign w49 = (a[2] & ~w24) | (a[2] & w24066) | (~w24 & w24066);
assign w50 = ~w47 & w24353;
assign w51 = (~w38 & w50) | (~w38 & w24068) | (w50 & w24068);
assign w52 = ~w50 & w24069;
assign w53 = ~w51 & ~w52;
assign w54 = ~w34 & ~w53;
assign w55 = w34 & w53;
assign w56 = ~w54 & ~w55;
assign w57 = ~w37 & w24070;
assign w58 = a[3] & ~a[4];
assign w59 = ~a[3] & a[4];
assign w60 = ~w58 & ~w59;
assign w61 = w37 & ~w60;
assign w62 = b[0] & w61;
assign w63 = ~a[4] & ~a[5];
assign w64 = a[4] & a[5];
assign w65 = ~w63 & ~w64;
assign w66 = ~w37 & w65;
assign w67 = ~w8 & w66;
assign w68 = ~w37 & ~w65;
assign w69 = b[1] & w68;
assign w70 = ~w62 & ~w67;
assign w71 = w70 & w24071;
assign w72 = (w57 & ~w70) | (w57 & w24072) | (~w70 & w24072);
assign w73 = ~w71 & ~w72;
assign w74 = w4 & w24073;
assign w75 = b[3] & w9;
assign w76 = ~b[3] & ~b[4];
assign w77 = b[3] & b[4];
assign w78 = ~w76 & ~w77;
assign w79 = b[2] & ~w41;
assign w80 = b[0] & w42;
assign w81 = ~w79 & ~w80;
assign w82 = ~w78 & w81;
assign w83 = w78 & ~w81;
assign w84 = ~w82 & ~w83;
assign w85 = ~w74 & ~w75;
assign w86 = (w85 & ~w84) | (w85 & w24074) | (~w84 & w24074);
assign w87 = (a[2] & ~w24) | (a[2] & w24075) | (~w24 & w24075);
assign w88 = w86 & ~w87;
assign w89 = a[2] & ~w86;
assign w90 = ~w88 & ~w89;
assign w91 = w73 & w90;
assign w92 = ~w73 & ~w90;
assign w93 = ~w91 & ~w92;
assign w94 = (~w52 & ~w53) | (~w52 & w24076) | (~w53 & w24076);
assign w95 = w93 & ~w94;
assign w96 = ~w93 & w94;
assign w97 = ~w95 & ~w96;
assign w98 = a[5] & ~w71;
assign w99 = b[2] & w68;
assign w100 = w22 & w66;
assign w101 = b[1] & w61;
assign w102 = w37 & w60;
assign w103 = w65 & w102;
assign w104 = w102 & w24077;
assign w105 = ~w99 & ~w100;
assign w106 = w105 & w24078;
assign w107 = w98 & ~w106;
assign w108 = ~w98 & w106;
assign w109 = ~w107 & ~w108;
assign w110 = ~b[4] & ~b[5];
assign w111 = b[4] & b[5];
assign w112 = ~w110 & ~w111;
assign w113 = (~w77 & w81) | (~w77 & w24079) | (w81 & w24079);
assign w114 = w112 & ~w113;
assign w115 = ~w112 & w113;
assign w116 = ~w114 & ~w115;
assign w117 = a[0] & w3;
assign w118 = w4 & w24080;
assign w119 = b[4] & w9;
assign w120 = b[3] & w24;
assign w121 = ~w118 & w24081;
assign w122 = a[2] & ~w121;
assign w123 = ~w118 & w24082;
assign w124 = (w123 & ~w116) | (w123 & w24354) | (~w116 & w24354);
assign w125 = (~w122 & ~w116) | (~w122 & w24083) | (~w116 & w24083);
assign w126 = ~w124 & w125;
assign w127 = w109 & w126;
assign w128 = ~w109 & ~w126;
assign w129 = ~w127 & ~w128;
assign w130 = (~w91 & ~w93) | (~w91 & w24609) | (~w93 & w24609);
assign w131 = w129 & ~w130;
assign w132 = ~w129 & w130;
assign w133 = ~w131 & ~w132;
assign w134 = (~w127 & w130) | (~w127 & w24084) | (w130 & w24084);
assign w135 = ~a[5] & ~b[0];
assign w136 = ~a[6] & b[0];
assign w137 = ~w135 & ~w136;
assign w138 = w102 & w24085;
assign w139 = b[3] & w68;
assign w140 = b[2] & w61;
assign w141 = ~w139 & ~w140;
assign w142 = ~w138 & w141;
assign w143 = w142 & w24086;
assign w144 = (~w137 & ~w142) | (~w137 & w24087) | (~w142 & w24087);
assign w145 = ~w143 & ~w144;
assign w146 = ~w98 & w24088;
assign w147 = w145 & w146;
assign w148 = ~w145 & ~w146;
assign w149 = ~w147 & ~w148;
assign w150 = w4 & w24089;
assign w151 = b[5] & w9;
assign w152 = ~b[5] & ~b[6];
assign w153 = b[5] & b[6];
assign w154 = ~w152 & ~w153;
assign w155 = (w113 & w24091) | (w113 & w24092) | (w24091 & w24092);
assign w156 = w154 & w25717;
assign w157 = ~w155 & ~w156;
assign w158 = ~w150 & ~w151;
assign w159 = (w158 & ~w157) | (w158 & w24093) | (~w157 & w24093);
assign w160 = (a[2] & ~w24) | (a[2] & w24094) | (~w24 & w24094);
assign w161 = w159 & ~w160;
assign w162 = (w157 & w24095) | (w157 & w24096) | (w24095 & w24096);
assign w163 = ~w161 & ~w162;
assign w164 = ~w149 & w163;
assign w165 = w149 & ~w163;
assign w166 = ~w164 & ~w165;
assign w167 = ~w134 & w166;
assign w168 = w134 & ~w166;
assign w169 = ~w167 & ~w168;
assign w170 = (~w164 & w134) | (~w164 & w24097) | (w134 & w24097);
assign w171 = a[5] & a[6];
assign w172 = ~a[5] & ~a[6];
assign w173 = ~w171 & ~w172;
assign w174 = b[0] & w173;
assign w175 = w173 & w24098;
assign w176 = a[7] & ~a[8];
assign w177 = ~a[7] & a[8];
assign w178 = ~w176 & ~w177;
assign w179 = w173 & ~w178;
assign w180 = ~w8 & w179;
assign w181 = ~a[7] & ~w171;
assign w182 = a[7] & ~w172;
assign w183 = ~w181 & ~w182;
assign w184 = b[0] & w183;
assign w185 = w173 & w178;
assign w186 = b[1] & w185;
assign w187 = ~w180 & ~w184;
assign w188 = w187 & w24099;
assign w189 = (w175 & ~w187) | (w175 & w24100) | (~w187 & w24100);
assign w190 = ~w188 & ~w189;
assign w191 = w102 & w24101;
assign w192 = b[3] & w61;
assign w193 = b[4] & w68;
assign w194 = w66 & w84;
assign w195 = ~w192 & ~w193;
assign w196 = ~w191 & w195;
assign w197 = ~w194 & w196;
assign w198 = a[5] & ~w197;
assign w199 = ~a[5] & w197;
assign w200 = ~w198 & ~w199;
assign w201 = w190 & w200;
assign w202 = ~w190 & ~w200;
assign w203 = ~w201 & ~w202;
assign w204 = ~w143 & ~w174;
assign w205 = ~w148 & ~w204;
assign w206 = w203 & w205;
assign w207 = ~w203 & ~w205;
assign w208 = ~w206 & ~w207;
assign w209 = w4 & w24102;
assign w210 = b[6] & w9;
assign w211 = ~b[6] & ~b[7];
assign w212 = b[6] & b[7];
assign w213 = ~w211 & ~w212;
assign w214 = ~w156 & w24103;
assign w215 = (w213 & w156) | (w213 & w24104) | (w156 & w24104);
assign w216 = ~w214 & ~w215;
assign w217 = ~w209 & ~w210;
assign w218 = (w217 & ~w216) | (w217 & w24105) | (~w216 & w24105);
assign w219 = (a[2] & ~w24) | (a[2] & w24106) | (~w24 & w24106);
assign w220 = w218 & ~w219;
assign w221 = (w216 & w24107) | (w216 & w24108) | (w24107 & w24108);
assign w222 = ~w220 & ~w221;
assign w223 = w208 & w222;
assign w224 = ~w208 & ~w222;
assign w225 = ~w223 & ~w224;
assign w226 = w170 & ~w225;
assign w227 = ~w170 & w225;
assign w228 = ~w226 & ~w227;
assign w229 = (a[8] & ~w173) | (a[8] & w24109) | (~w173 & w24109);
assign w230 = w187 & w24110;
assign w231 = a[8] & ~w230;
assign w232 = b[1] & w183;
assign w233 = b[2] & w185;
assign w234 = w22 & w179;
assign w235 = w171 & w176;
assign w236 = w172 & w177;
assign w237 = ~w235 & ~w236;
assign w238 = b[0] & ~w237;
assign w239 = ~w232 & ~w233;
assign w240 = ~w234 & ~w238;
assign w241 = w239 & w240;
assign w242 = ~w231 & w241;
assign w243 = w231 & ~w241;
assign w244 = ~w242 & ~w243;
assign w245 = (~a[5] & ~w116) | (~a[5] & w24111) | (~w116 & w24111);
assign w246 = ~a[4] & ~w37;
assign w247 = w116 & w246;
assign w248 = ~w245 & ~w247;
assign w249 = b[4] & w61;
assign w250 = b[5] & w68;
assign w251 = w102 & w24112;
assign w252 = ~w249 & ~w250;
assign w253 = ~w251 & w252;
assign w254 = (a[5] & ~w252) | (a[5] & w24113) | (~w252 & w24113);
assign w255 = (~w254 & w248) | (~w254 & w24114) | (w248 & w24114);
assign w256 = w244 & w255;
assign w257 = ~w244 & ~w255;
assign w258 = ~w256 & ~w257;
assign w259 = (~w201 & ~w203) | (~w201 & w24115) | (~w203 & w24115);
assign w260 = ~w258 & w259;
assign w261 = w258 & ~w259;
assign w262 = ~w260 & ~w261;
assign w263 = w4 & w24116;
assign w264 = b[7] & w9;
assign w265 = ~b[7] & ~b[8];
assign w266 = b[7] & b[8];
assign w267 = ~w265 & ~w266;
assign w268 = (w156 & w24119) | (w156 & w24120) | (w24119 & w24120);
assign w269 = ~w267 & w25718;
assign w270 = ~w268 & ~w269;
assign w271 = ~w263 & ~w264;
assign w272 = (w271 & ~w270) | (w271 & w24121) | (~w270 & w24121);
assign w273 = (a[2] & ~w24) | (a[2] & w24122) | (~w24 & w24122);
assign w274 = w272 & ~w273;
assign w275 = (w270 & w24123) | (w270 & w24124) | (w24123 & w24124);
assign w276 = ~w274 & ~w275;
assign w277 = w262 & w276;
assign w278 = ~w262 & ~w276;
assign w279 = ~w277 & ~w278;
assign w280 = (~w223 & ~w225) | (~w223 & w24125) | (~w225 & w24125);
assign w281 = w279 & ~w280;
assign w282 = ~w279 & w280;
assign w283 = ~w281 & ~w282;
assign w284 = w230 & w241;
assign w285 = ~a[8] & ~b[0];
assign w286 = ~a[9] & b[0];
assign w287 = ~w285 & ~w286;
assign w288 = b[2] & w183;
assign w289 = b[3] & w185;
assign w290 = b[1] & ~w237;
assign w291 = ~w288 & ~w289;
assign w292 = ~w290 & w291;
assign w293 = w292 & w24126;
assign w294 = (~w287 & ~w292) | (~w287 & w24127) | (~w292 & w24127);
assign w295 = ~w293 & ~w294;
assign w296 = w284 & w295;
assign w297 = ~w284 & ~w295;
assign w298 = ~w296 & ~w297;
assign w299 = w102 & w24128;
assign w300 = b[6] & w68;
assign w301 = b[5] & w61;
assign w302 = w66 & w157;
assign w303 = ~w300 & ~w301;
assign w304 = ~w299 & w303;
assign w305 = (a[5] & w302) | (a[5] & w24129) | (w302 & w24129);
assign w306 = ~w302 & w24130;
assign w307 = ~w305 & ~w306;
assign w308 = ~w298 & w307;
assign w309 = w298 & ~w307;
assign w310 = ~w308 & ~w309;
assign w311 = (~w256 & w259) | (~w256 & w24131) | (w259 & w24131);
assign w312 = ~w310 & w311;
assign w313 = w310 & ~w311;
assign w314 = ~w312 & ~w313;
assign w315 = w4 & w24132;
assign w316 = b[8] & w9;
assign w317 = ~b[8] & ~b[9];
assign w318 = b[8] & b[9];
assign w319 = ~w317 & ~w318;
assign w320 = ~w268 & w24133;
assign w321 = (w319 & w268) | (w319 & w24134) | (w268 & w24134);
assign w322 = ~w320 & ~w321;
assign w323 = ~w315 & ~w316;
assign w324 = (w323 & ~w322) | (w323 & w24135) | (~w322 & w24135);
assign w325 = (a[2] & ~w24) | (a[2] & w24136) | (~w24 & w24136);
assign w326 = w324 & ~w325;
assign w327 = (w322 & w24137) | (w322 & w24138) | (w24137 & w24138);
assign w328 = ~w326 & ~w327;
assign w329 = w314 & w328;
assign w330 = ~w314 & ~w328;
assign w331 = ~w329 & ~w330;
assign w332 = ~w277 & ~w281;
assign w333 = w331 & w332;
assign w334 = ~w331 & ~w332;
assign w335 = ~w333 & ~w334;
assign w336 = b[4] & w185;
assign w337 = b[2] & ~w237;
assign w338 = b[3] & w183;
assign w339 = w84 & w179;
assign w340 = ~w336 & ~w337;
assign w341 = ~w338 & w340;
assign w342 = ~w339 & w341;
assign w343 = a[8] & ~w342;
assign w344 = ~a[8] & w342;
assign w345 = ~w343 & ~w344;
assign w346 = a[8] & a[9];
assign w347 = ~a[8] & ~a[9];
assign w348 = ~w346 & ~w347;
assign w349 = b[0] & w348;
assign w350 = w348 & w24139;
assign w351 = a[10] & ~a[11];
assign w352 = ~a[10] & a[11];
assign w353 = ~w351 & ~w352;
assign w354 = w348 & ~w353;
assign w355 = ~w8 & w354;
assign w356 = ~a[10] & ~w346;
assign w357 = a[10] & ~w347;
assign w358 = ~w356 & ~w357;
assign w359 = b[0] & w358;
assign w360 = w348 & w353;
assign w361 = b[1] & w360;
assign w362 = ~w355 & ~w359;
assign w363 = w362 & w24140;
assign w364 = (w350 & ~w362) | (w350 & w24141) | (~w362 & w24141);
assign w365 = ~w363 & ~w364;
assign w366 = ~w345 & ~w365;
assign w367 = w345 & w365;
assign w368 = ~w366 & ~w367;
assign w369 = ~w293 & ~w349;
assign w370 = ~w297 & ~w369;
assign w371 = w368 & w370;
assign w372 = ~w368 & ~w370;
assign w373 = ~w371 & ~w372;
assign w374 = w102 & w24142;
assign w375 = b[7] & w68;
assign w376 = b[6] & w61;
assign w377 = ~w375 & ~w376;
assign w378 = ~w374 & w377;
assign w379 = (w378 & ~w216) | (w378 & w24143) | (~w216 & w24143);
assign w380 = a[5] & ~w379;
assign w381 = ~a[5] & w379;
assign w382 = ~w380 & ~w381;
assign w383 = w373 & w382;
assign w384 = ~w373 & ~w382;
assign w385 = ~w383 & ~w384;
assign w386 = (~w308 & w311) | (~w308 & w24144) | (w311 & w24144);
assign w387 = w385 & w386;
assign w388 = ~w385 & ~w386;
assign w389 = ~w387 & ~w388;
assign w390 = w4 & w24145;
assign w391 = b[9] & w9;
assign w392 = ~b[9] & ~b[10];
assign w393 = b[9] & b[10];
assign w394 = ~w392 & ~w393;
assign w395 = ~w394 & w25719;
assign w396 = (w268 & w24148) | (w268 & w24149) | (w24148 & w24149);
assign w397 = ~w395 & ~w396;
assign w398 = ~w390 & ~w391;
assign w399 = (w398 & ~w397) | (w398 & w24150) | (~w397 & w24150);
assign w400 = (a[2] & ~w24) | (a[2] & w24151) | (~w24 & w24151);
assign w401 = w399 & ~w400;
assign w402 = (w397 & w24152) | (w397 & w24153) | (w24152 & w24153);
assign w403 = ~w401 & ~w402;
assign w404 = w389 & ~w403;
assign w405 = ~w389 & w403;
assign w406 = ~w404 & ~w405;
assign w407 = (~w330 & ~w332) | (~w330 & w24154) | (~w332 & w24154);
assign w408 = w406 & w407;
assign w409 = ~w406 & ~w407;
assign w410 = ~w408 & ~w409;
assign w411 = ~w405 & ~w408;
assign w412 = (~w367 & ~w368) | (~w367 & w24155) | (~w368 & w24155);
assign w413 = (a[11] & ~w348) | (a[11] & w24156) | (~w348 & w24156);
assign w414 = w362 & w24157;
assign w415 = a[11] & ~w414;
assign w416 = w22 & w354;
assign w417 = w346 & w351;
assign w418 = w347 & w352;
assign w419 = ~w417 & ~w418;
assign w420 = b[0] & ~w419;
assign w421 = b[2] & w360;
assign w422 = b[1] & w358;
assign w423 = ~w416 & ~w420;
assign w424 = ~w421 & ~w422;
assign w425 = w423 & w424;
assign w426 = ~w415 & w425;
assign w427 = w415 & ~w425;
assign w428 = ~w426 & ~w427;
assign w429 = b[3] & ~w237;
assign w430 = b[4] & w183;
assign w431 = b[5] & w185;
assign w432 = ~w429 & ~w430;
assign w433 = ~w431 & w432;
assign w434 = (~a[8] & ~w116) | (~a[8] & w24158) | (~w116 & w24158);
assign w435 = w116 & w24159;
assign w436 = ~w434 & ~w435;
assign w437 = (a[8] & ~w432) | (a[8] & w24160) | (~w432 & w24160);
assign w438 = (~w437 & w436) | (~w437 & w24161) | (w436 & w24161);
assign w439 = w428 & w438;
assign w440 = ~w428 & ~w438;
assign w441 = ~w439 & ~w440;
assign w442 = w412 & w441;
assign w443 = ~w412 & ~w441;
assign w444 = ~w442 & ~w443;
assign w445 = w102 & w24162;
assign w446 = b[8] & w68;
assign w447 = b[7] & w61;
assign w448 = ~w446 & ~w447;
assign w449 = ~w445 & w448;
assign w450 = (w449 & ~w270) | (w449 & w24163) | (~w270 & w24163);
assign w451 = a[5] & ~w450;
assign w452 = ~a[5] & w450;
assign w453 = ~w451 & ~w452;
assign w454 = w444 & ~w453;
assign w455 = ~w444 & w453;
assign w456 = ~w454 & ~w455;
assign w457 = (~w384 & ~w385) | (~w384 & w24164) | (~w385 & w24164);
assign w458 = w456 & w457;
assign w459 = ~w456 & ~w457;
assign w460 = ~w458 & ~w459;
assign w461 = w4 & w24165;
assign w462 = b[10] & w9;
assign w463 = ~b[10] & ~b[11];
assign w464 = b[10] & b[11];
assign w465 = ~w463 & ~w464;
assign w466 = (~w268 & w24166) | (~w268 & w24167) | (w24166 & w24167);
assign w467 = w465 & ~w466;
assign w468 = ~w465 & w466;
assign w469 = ~w467 & ~w468;
assign w470 = ~w461 & ~w462;
assign w471 = (w470 & ~w469) | (w470 & w24168) | (~w469 & w24168);
assign w472 = (a[2] & ~w24) | (a[2] & w24169) | (~w24 & w24169);
assign w473 = w471 & ~w472;
assign w474 = (w469 & w24170) | (w469 & w24171) | (w24170 & w24171);
assign w475 = ~w473 & ~w474;
assign w476 = w460 & w475;
assign w477 = ~w460 & ~w475;
assign w478 = ~w476 & ~w477;
assign w479 = w411 & ~w478;
assign w480 = ~w411 & w478;
assign w481 = ~w479 & ~w480;
assign w482 = w414 & w425;
assign w483 = ~a[11] & ~b[0];
assign w484 = ~a[12] & b[0];
assign w485 = ~w483 & ~w484;
assign w486 = b[1] & ~w419;
assign w487 = b[3] & w360;
assign w488 = b[2] & w358;
assign w489 = ~w486 & ~w487;
assign w490 = ~w488 & w489;
assign w491 = w490 & w24172;
assign w492 = (~w485 & ~w490) | (~w485 & w24173) | (~w490 & w24173);
assign w493 = ~w491 & ~w492;
assign w494 = w482 & w493;
assign w495 = ~w482 & ~w493;
assign w496 = ~w494 & ~w495;
assign w497 = b[6] & w185;
assign w498 = b[5] & w183;
assign w499 = b[4] & ~w237;
assign w500 = w157 & w179;
assign w501 = ~w497 & ~w498;
assign w502 = ~w499 & w501;
assign w503 = (a[8] & w500) | (a[8] & w24174) | (w500 & w24174);
assign w504 = ~w500 & w24175;
assign w505 = ~w503 & ~w504;
assign w506 = ~w496 & w505;
assign w507 = w496 & ~w505;
assign w508 = ~w506 & ~w507;
assign w509 = (~w440 & ~w412) | (~w440 & w24176) | (~w412 & w24176);
assign w510 = ~w508 & ~w509;
assign w511 = w508 & w509;
assign w512 = ~w510 & ~w511;
assign w513 = w102 & w24177;
assign w514 = b[8] & w61;
assign w515 = b[9] & w68;
assign w516 = ~w514 & ~w515;
assign w517 = ~w513 & w516;
assign w518 = (w517 & ~w322) | (w517 & w24178) | (~w322 & w24178);
assign w519 = a[5] & ~w518;
assign w520 = ~a[5] & w518;
assign w521 = ~w519 & ~w520;
assign w522 = ~w512 & ~w521;
assign w523 = w512 & w521;
assign w524 = ~w522 & ~w523;
assign w525 = ~w455 & ~w458;
assign w526 = w524 & ~w525;
assign w527 = ~w524 & w525;
assign w528 = ~w526 & ~w527;
assign w529 = w4 & w24179;
assign w530 = b[11] & w9;
assign w531 = ~b[11] & ~b[12];
assign w532 = b[11] & b[12];
assign w533 = ~w531 & ~w532;
assign w534 = (w466 & w24181) | (w466 & w24182) | (w24181 & w24182);
assign w535 = w533 & w25720;
assign w536 = ~w534 & ~w535;
assign w537 = ~w529 & ~w530;
assign w538 = (w537 & ~w536) | (w537 & w24184) | (~w536 & w24184);
assign w539 = (a[2] & ~w24) | (a[2] & w24185) | (~w24 & w24185);
assign w540 = w538 & ~w539;
assign w541 = (w536 & w24186) | (w536 & w24187) | (w24186 & w24187);
assign w542 = ~w540 & ~w541;
assign w543 = w528 & w542;
assign w544 = ~w528 & ~w542;
assign w545 = ~w543 & ~w544;
assign w546 = (~w476 & w411) | (~w476 & w24188) | (w411 & w24188);
assign w547 = w545 & ~w546;
assign w548 = ~w545 & w546;
assign w549 = ~w547 & ~w548;
assign w550 = ~w543 & ~w547;
assign w551 = b[2] & ~w419;
assign w552 = b[3] & w358;
assign w553 = b[4] & w360;
assign w554 = w84 & w354;
assign w555 = ~w551 & ~w552;
assign w556 = ~w553 & w555;
assign w557 = ~w554 & w556;
assign w558 = a[11] & ~w557;
assign w559 = ~a[11] & w557;
assign w560 = ~w558 & ~w559;
assign w561 = a[11] & a[12];
assign w562 = ~a[11] & ~a[12];
assign w563 = ~w561 & ~w562;
assign w564 = b[0] & w563;
assign w565 = w563 & w24189;
assign w566 = a[13] & ~a[14];
assign w567 = ~a[13] & a[14];
assign w568 = ~w566 & ~w567;
assign w569 = w563 & ~w568;
assign w570 = ~w8 & w569;
assign w571 = ~a[13] & ~w561;
assign w572 = a[13] & ~w562;
assign w573 = ~w571 & ~w572;
assign w574 = b[0] & w573;
assign w575 = w563 & w568;
assign w576 = b[1] & w575;
assign w577 = ~w570 & ~w574;
assign w578 = w577 & w24190;
assign w579 = (w565 & ~w577) | (w565 & w24191) | (~w577 & w24191);
assign w580 = ~w578 & ~w579;
assign w581 = ~w560 & ~w580;
assign w582 = w560 & w580;
assign w583 = ~w581 & ~w582;
assign w584 = ~w491 & ~w564;
assign w585 = ~w495 & ~w584;
assign w586 = w583 & w585;
assign w587 = ~w583 & ~w585;
assign w588 = ~w586 & ~w587;
assign w589 = b[7] & w185;
assign w590 = b[5] & ~w237;
assign w591 = b[6] & w183;
assign w592 = ~w589 & ~w590;
assign w593 = ~w591 & w592;
assign w594 = (w593 & ~w216) | (w593 & w24192) | (~w216 & w24192);
assign w595 = a[8] & ~w594;
assign w596 = ~a[8] & w594;
assign w597 = ~w595 & ~w596;
assign w598 = w588 & w597;
assign w599 = ~w588 & ~w597;
assign w600 = ~w598 & ~w599;
assign w601 = (~w506 & ~w509) | (~w506 & w24193) | (~w509 & w24193);
assign w602 = ~w600 & w601;
assign w603 = w600 & ~w601;
assign w604 = ~w602 & ~w603;
assign w605 = w102 & w24194;
assign w606 = b[10] & w68;
assign w607 = b[9] & w61;
assign w608 = ~w606 & ~w607;
assign w609 = ~w605 & w608;
assign w610 = (w609 & ~w397) | (w609 & w24195) | (~w397 & w24195);
assign w611 = a[5] & ~w610;
assign w612 = ~a[5] & w610;
assign w613 = ~w611 & ~w612;
assign w614 = w604 & w613;
assign w615 = ~w604 & ~w613;
assign w616 = ~w614 & ~w615;
assign w617 = (~w523 & w525) | (~w523 & w24196) | (w525 & w24196);
assign w618 = w616 & ~w617;
assign w619 = ~w616 & w617;
assign w620 = ~w618 & ~w619;
assign w621 = w4 & w24197;
assign w622 = b[12] & w9;
assign w623 = ~b[12] & ~b[13];
assign w624 = b[12] & b[13];
assign w625 = ~w623 & ~w624;
assign w626 = w625 & w25721;
assign w627 = (w466 & w24202) | (w466 & w24203) | (w24202 & w24203);
assign w628 = ~w626 & ~w627;
assign w629 = ~w621 & ~w622;
assign w630 = (w629 & ~w628) | (w629 & w24204) | (~w628 & w24204);
assign w631 = (a[2] & ~w24) | (a[2] & w24205) | (~w24 & w24205);
assign w632 = w630 & ~w631;
assign w633 = (w628 & w24206) | (w628 & w24207) | (w24206 & w24207);
assign w634 = ~w632 & ~w633;
assign w635 = w620 & w634;
assign w636 = ~w620 & ~w634;
assign w637 = ~w635 & ~w636;
assign w638 = w550 & w637;
assign w639 = ~w550 & ~w637;
assign w640 = ~w638 & ~w639;
assign w641 = ~w614 & ~w618;
assign w642 = (a[14] & ~w563) | (a[14] & w24208) | (~w563 & w24208);
assign w643 = w577 & w24209;
assign w644 = a[14] & ~w643;
assign w645 = b[1] & w573;
assign w646 = w22 & w569;
assign w647 = w561 & w566;
assign w648 = w562 & w567;
assign w649 = ~w647 & ~w648;
assign w650 = b[0] & ~w649;
assign w651 = b[2] & w575;
assign w652 = ~w645 & ~w646;
assign w653 = ~w650 & ~w651;
assign w654 = w652 & w653;
assign w655 = ~w644 & w654;
assign w656 = w644 & ~w654;
assign w657 = ~w655 & ~w656;
assign w658 = b[4] & w358;
assign w659 = b[5] & w360;
assign w660 = b[3] & ~w419;
assign w661 = ~w658 & ~w659;
assign w662 = ~w660 & w661;
assign w663 = (~a[11] & ~w116) | (~a[11] & w24210) | (~w116 & w24210);
assign w664 = w116 & w24211;
assign w665 = ~w663 & ~w664;
assign w666 = (a[11] & ~w661) | (a[11] & w24212) | (~w661 & w24212);
assign w667 = (~w666 & w665) | (~w666 & w24213) | (w665 & w24213);
assign w668 = w657 & w667;
assign w669 = ~w657 & ~w667;
assign w670 = ~w668 & ~w669;
assign w671 = (~w582 & ~w583) | (~w582 & w24214) | (~w583 & w24214);
assign w672 = ~w670 & w671;
assign w673 = w670 & ~w671;
assign w674 = ~w672 & ~w673;
assign w675 = b[6] & ~w237;
assign w676 = b[7] & w183;
assign w677 = b[8] & w185;
assign w678 = ~w675 & ~w676;
assign w679 = ~w677 & w678;
assign w680 = (w679 & ~w270) | (w679 & w24215) | (~w270 & w24215);
assign w681 = a[8] & ~w680;
assign w682 = ~a[8] & w680;
assign w683 = ~w681 & ~w682;
assign w684 = ~w674 & ~w683;
assign w685 = w674 & w683;
assign w686 = ~w684 & ~w685;
assign w687 = (~w598 & ~w600) | (~w598 & w24216) | (~w600 & w24216);
assign w688 = w686 & ~w687;
assign w689 = ~w686 & w687;
assign w690 = ~w688 & ~w689;
assign w691 = w102 & w24217;
assign w692 = b[11] & w68;
assign w693 = b[10] & w61;
assign w694 = ~w692 & ~w693;
assign w695 = ~w691 & w694;
assign w696 = (w695 & ~w469) | (w695 & w24218) | (~w469 & w24218);
assign w697 = a[5] & ~w696;
assign w698 = ~a[5] & w696;
assign w699 = ~w697 & ~w698;
assign w700 = ~w690 & ~w699;
assign w701 = w690 & w699;
assign w702 = ~w700 & ~w701;
assign w703 = w641 & ~w702;
assign w704 = ~w641 & w702;
assign w705 = ~w703 & ~w704;
assign w706 = w4 & w24219;
assign w707 = b[13] & w9;
assign w708 = ~b[13] & ~b[14];
assign w709 = b[13] & b[14];
assign w710 = ~w708 & ~w709;
assign w711 = (w466 & w24220) | (w466 & w24221) | (w24220 & w24221);
assign w712 = ~w710 & w711;
assign w713 = w710 & ~w711;
assign w714 = ~w712 & ~w713;
assign w715 = ~w706 & ~w707;
assign w716 = (w715 & ~w714) | (w715 & w24222) | (~w714 & w24222);
assign w717 = (a[2] & ~w24) | (a[2] & w24223) | (~w24 & w24223);
assign w718 = w716 & ~w717;
assign w719 = (w714 & w24224) | (w714 & w24225) | (w24224 & w24225);
assign w720 = ~w718 & ~w719;
assign w721 = ~w705 & ~w720;
assign w722 = w705 & w720;
assign w723 = ~w721 & ~w722;
assign w724 = (~w636 & ~w550) | (~w636 & w24226) | (~w550 & w24226);
assign w725 = w723 & w724;
assign w726 = ~w723 & ~w724;
assign w727 = ~w725 & ~w726;
assign w728 = ~w722 & ~w725;
assign w729 = w102 & w24227;
assign w730 = b[12] & w68;
assign w731 = b[11] & w61;
assign w732 = ~w730 & ~w731;
assign w733 = ~w729 & w732;
assign w734 = (w733 & ~w536) | (w733 & w24228) | (~w536 & w24228);
assign w735 = a[5] & ~w734;
assign w736 = ~a[5] & w734;
assign w737 = ~w735 & ~w736;
assign w738 = ~w685 & ~w688;
assign w739 = w643 & w654;
assign w740 = ~a[14] & ~b[0];
assign w741 = ~a[15] & b[0];
assign w742 = ~w740 & ~w741;
assign w743 = b[2] & w573;
assign w744 = b[1] & ~w649;
assign w745 = b[3] & w575;
assign w746 = ~w743 & ~w744;
assign w747 = ~w745 & w746;
assign w748 = w747 & w24229;
assign w749 = (~w742 & ~w747) | (~w742 & w24230) | (~w747 & w24230);
assign w750 = ~w748 & ~w749;
assign w751 = w739 & w750;
assign w752 = ~w739 & ~w750;
assign w753 = ~w751 & ~w752;
assign w754 = b[5] & w358;
assign w755 = b[4] & ~w419;
assign w756 = b[6] & w360;
assign w757 = w157 & w354;
assign w758 = ~w754 & ~w755;
assign w759 = ~w756 & w758;
assign w760 = (a[11] & w757) | (a[11] & w24231) | (w757 & w24231);
assign w761 = ~w757 & w24232;
assign w762 = ~w760 & ~w761;
assign w763 = ~w753 & w762;
assign w764 = w753 & ~w762;
assign w765 = ~w763 & ~w764;
assign w766 = (~w668 & w671) | (~w668 & w24233) | (w671 & w24233);
assign w767 = w765 & ~w766;
assign w768 = ~w765 & w766;
assign w769 = ~w767 & ~w768;
assign w770 = b[9] & w185;
assign w771 = b[8] & w183;
assign w772 = b[7] & ~w237;
assign w773 = ~w770 & ~w771;
assign w774 = ~w772 & w773;
assign w775 = (w774 & ~w322) | (w774 & w24234) | (~w322 & w24234);
assign w776 = a[8] & ~w775;
assign w777 = ~a[8] & w775;
assign w778 = ~w776 & ~w777;
assign w779 = ~w769 & ~w778;
assign w780 = w769 & w778;
assign w781 = ~w779 & ~w780;
assign w782 = w738 & ~w781;
assign w783 = ~w738 & w781;
assign w784 = ~w782 & ~w783;
assign w785 = ~w737 & ~w784;
assign w786 = w737 & w784;
assign w787 = ~w785 & ~w786;
assign w788 = (~w701 & w641) | (~w701 & w24235) | (w641 & w24235);
assign w789 = w787 & ~w788;
assign w790 = ~w787 & w788;
assign w791 = ~w789 & ~w790;
assign w792 = w4 & w24236;
assign w793 = b[14] & w9;
assign w794 = ~b[14] & ~b[15];
assign w795 = b[14] & b[15];
assign w796 = ~w794 & ~w795;
assign w797 = ~w796 & w25722;
assign w798 = (w711 & w24238) | (w711 & w24239) | (w24238 & w24239);
assign w799 = ~w797 & ~w798;
assign w800 = ~w792 & ~w793;
assign w801 = (w800 & w799) | (w800 & w24240) | (w799 & w24240);
assign w802 = (a[2] & ~w24) | (a[2] & w24241) | (~w24 & w24241);
assign w803 = w801 & ~w802;
assign w804 = a[2] & ~w801;
assign w805 = ~w803 & ~w804;
assign w806 = ~w791 & ~w805;
assign w807 = w791 & w805;
assign w808 = ~w806 & ~w807;
assign w809 = w728 & w808;
assign w810 = ~w728 & ~w808;
assign w811 = ~w809 & ~w810;
assign w812 = ~w786 & ~w789;
assign w813 = (~w763 & w766) | (~w763 & w24242) | (w766 & w24242);
assign w814 = b[4] & w575;
assign w815 = b[3] & w573;
assign w816 = b[2] & ~w649;
assign w817 = w84 & w569;
assign w818 = ~w814 & ~w815;
assign w819 = ~w816 & w818;
assign w820 = ~w817 & w819;
assign w821 = a[14] & ~w820;
assign w822 = ~a[14] & w820;
assign w823 = ~w821 & ~w822;
assign w824 = a[14] & a[15];
assign w825 = ~a[14] & ~a[15];
assign w826 = ~w824 & ~w825;
assign w827 = b[0] & w826;
assign w828 = w826 & w24243;
assign w829 = ~a[16] & a[17];
assign w830 = a[16] & ~a[17];
assign w831 = ~w829 & ~w830;
assign w832 = w826 & ~w831;
assign w833 = ~w8 & w832;
assign w834 = w826 & w831;
assign w835 = b[1] & w834;
assign w836 = ~a[16] & ~w824;
assign w837 = a[16] & ~w825;
assign w838 = ~w836 & ~w837;
assign w839 = b[0] & w838;
assign w840 = ~w833 & ~w835;
assign w841 = w840 & w24244;
assign w842 = (w828 & ~w840) | (w828 & w24245) | (~w840 & w24245);
assign w843 = ~w841 & ~w842;
assign w844 = ~w823 & ~w843;
assign w845 = w823 & w843;
assign w846 = ~w844 & ~w845;
assign w847 = ~w748 & ~w827;
assign w848 = ~w752 & ~w847;
assign w849 = w846 & w848;
assign w850 = ~w846 & ~w848;
assign w851 = ~w849 & ~w850;
assign w852 = b[5] & ~w419;
assign w853 = b[7] & w360;
assign w854 = b[6] & w358;
assign w855 = ~w852 & ~w853;
assign w856 = ~w854 & w855;
assign w857 = (w856 & ~w216) | (w856 & w24246) | (~w216 & w24246);
assign w858 = a[11] & ~w857;
assign w859 = ~a[11] & w857;
assign w860 = ~w858 & ~w859;
assign w861 = ~w851 & ~w860;
assign w862 = w851 & w860;
assign w863 = ~w861 & ~w862;
assign w864 = w813 & w863;
assign w865 = ~w813 & ~w863;
assign w866 = ~w864 & ~w865;
assign w867 = b[8] & ~w237;
assign w868 = b[10] & w185;
assign w869 = b[9] & w183;
assign w870 = ~w867 & ~w868;
assign w871 = ~w869 & w870;
assign w872 = (w871 & ~w397) | (w871 & w24247) | (~w397 & w24247);
assign w873 = a[8] & ~w872;
assign w874 = ~a[8] & w872;
assign w875 = ~w873 & ~w874;
assign w876 = w866 & ~w875;
assign w877 = ~w866 & w875;
assign w878 = ~w876 & ~w877;
assign w879 = (~w780 & w738) | (~w780 & w24248) | (w738 & w24248);
assign w880 = w878 & ~w879;
assign w881 = ~w878 & w879;
assign w882 = ~w880 & ~w881;
assign w883 = w102 & w24249;
assign w884 = b[12] & w61;
assign w885 = b[13] & w68;
assign w886 = ~w884 & ~w885;
assign w887 = ~w883 & w886;
assign w888 = (w887 & ~w628) | (w887 & w24250) | (~w628 & w24250);
assign w889 = a[5] & ~w888;
assign w890 = ~a[5] & w888;
assign w891 = ~w889 & ~w890;
assign w892 = ~w882 & ~w891;
assign w893 = w882 & w891;
assign w894 = ~w892 & ~w893;
assign w895 = w812 & w894;
assign w896 = ~w812 & ~w894;
assign w897 = ~w895 & ~w896;
assign w898 = w4 & w24251;
assign w899 = b[15] & w9;
assign w900 = ~b[15] & ~b[16];
assign w901 = b[15] & b[16];
assign w902 = ~w900 & ~w901;
assign w903 = (w711 & w24254) | (w711 & w24255) | (w24254 & w24255);
assign w904 = w902 & w25723;
assign w905 = ~w903 & ~w904;
assign w906 = ~w898 & ~w899;
assign w907 = (w906 & ~w905) | (w906 & w24256) | (~w905 & w24256);
assign w908 = (a[2] & ~w24) | (a[2] & w24257) | (~w24 & w24257);
assign w909 = w907 & ~w908;
assign w910 = (w905 & w24258) | (w905 & w24259) | (w24258 & w24259);
assign w911 = ~w909 & ~w910;
assign w912 = w897 & ~w911;
assign w913 = ~w897 & w911;
assign w914 = ~w912 & ~w913;
assign w915 = (~w806 & ~w728) | (~w806 & w24260) | (~w728 & w24260);
assign w916 = w914 & w915;
assign w917 = ~w914 & ~w915;
assign w918 = ~w916 & ~w917;
assign w919 = w102 & w24261;
assign w920 = b[13] & w61;
assign w921 = b[14] & w68;
assign w922 = ~w920 & ~w921;
assign w923 = ~w919 & w922;
assign w924 = (w923 & ~w714) | (w923 & w24262) | (~w714 & w24262);
assign w925 = a[5] & ~w924;
assign w926 = ~a[5] & w924;
assign w927 = ~w925 & ~w926;
assign w928 = ~w877 & ~w880;
assign w929 = (a[17] & ~w826) | (a[17] & w24263) | (~w826 & w24263);
assign w930 = w840 & w24264;
assign w931 = a[17] & ~w930;
assign w932 = w824 & w830;
assign w933 = w825 & w829;
assign w934 = ~w932 & ~w933;
assign w935 = b[0] & ~w934;
assign w936 = b[1] & w838;
assign w937 = b[2] & w834;
assign w938 = w22 & w832;
assign w939 = ~w935 & ~w936;
assign w940 = ~w937 & ~w938;
assign w941 = w939 & w940;
assign w942 = ~w931 & w941;
assign w943 = w931 & ~w941;
assign w944 = ~w942 & ~w943;
assign w945 = b[3] & ~w649;
assign w946 = b[5] & w575;
assign w947 = b[4] & w573;
assign w948 = ~w945 & ~w946;
assign w949 = ~w947 & w948;
assign w950 = (~a[14] & ~w116) | (~a[14] & w24265) | (~w116 & w24265);
assign w951 = w116 & w24266;
assign w952 = ~w950 & ~w951;
assign w953 = (a[14] & ~w948) | (a[14] & w24267) | (~w948 & w24267);
assign w954 = (~w953 & w952) | (~w953 & w24268) | (w952 & w24268);
assign w955 = w944 & w954;
assign w956 = ~w944 & ~w954;
assign w957 = ~w955 & ~w956;
assign w958 = (~w845 & ~w846) | (~w845 & w24269) | (~w846 & w24269);
assign w959 = ~w957 & w958;
assign w960 = w957 & ~w958;
assign w961 = ~w959 & ~w960;
assign w962 = b[6] & ~w419;
assign w963 = b[8] & w360;
assign w964 = b[7] & w358;
assign w965 = ~w962 & ~w963;
assign w966 = ~w964 & w965;
assign w967 = (w966 & ~w270) | (w966 & w24270) | (~w270 & w24270);
assign w968 = a[11] & ~w967;
assign w969 = ~a[11] & w967;
assign w970 = ~w968 & ~w969;
assign w971 = ~w961 & ~w970;
assign w972 = w961 & w970;
assign w973 = ~w971 & ~w972;
assign w974 = (~w861 & ~w863) | (~w861 & w24271) | (~w863 & w24271);
assign w975 = w973 & w974;
assign w976 = ~w973 & ~w974;
assign w977 = ~w975 & ~w976;
assign w978 = b[11] & w185;
assign w979 = b[10] & w183;
assign w980 = b[9] & ~w237;
assign w981 = ~w978 & ~w979;
assign w982 = ~w980 & w981;
assign w983 = (w982 & ~w469) | (w982 & w24272) | (~w469 & w24272);
assign w984 = a[8] & ~w983;
assign w985 = ~a[8] & w983;
assign w986 = ~w984 & ~w985;
assign w987 = ~w977 & ~w986;
assign w988 = w977 & w986;
assign w989 = ~w987 & ~w988;
assign w990 = w928 & w989;
assign w991 = ~w928 & ~w989;
assign w992 = ~w990 & ~w991;
assign w993 = ~w927 & w992;
assign w994 = w927 & ~w992;
assign w995 = ~w993 & ~w994;
assign w996 = (~w892 & ~w812) | (~w892 & w24273) | (~w812 & w24273);
assign w997 = w995 & w996;
assign w998 = ~w995 & ~w996;
assign w999 = ~w997 & ~w998;
assign w1000 = w4 & w24274;
assign w1001 = b[16] & w9;
assign w1002 = ~b[16] & ~b[17];
assign w1003 = b[16] & b[17];
assign w1004 = ~w1002 & ~w1003;
assign w1005 = (w711 & w24275) | (w711 & w24276) | (w24275 & w24276);
assign w1006 = (~w1004 & w1005) | (~w1004 & w24277) | (w1005 & w24277);
assign w1007 = ~w1005 & w24278;
assign w1008 = ~w1006 & ~w1007;
assign w1009 = ~w1000 & ~w1001;
assign w1010 = (w1009 & ~w1008) | (w1009 & w24279) | (~w1008 & w24279);
assign w1011 = (a[2] & ~w24) | (a[2] & w24280) | (~w24 & w24280);
assign w1012 = w1010 & ~w1011;
assign w1013 = (w1008 & w24281) | (w1008 & w24282) | (w24281 & w24282);
assign w1014 = ~w1012 & ~w1013;
assign w1015 = w999 & w1014;
assign w1016 = ~w999 & ~w1014;
assign w1017 = ~w1015 & ~w1016;
assign w1018 = ~w913 & ~w916;
assign w1019 = ~w1017 & ~w1018;
assign w1020 = w1017 & w1018;
assign w1021 = ~w1019 & ~w1020;
assign w1022 = ~w994 & ~w997;
assign w1023 = b[11] & w183;
assign w1024 = b[12] & w185;
assign w1025 = b[10] & ~w237;
assign w1026 = ~w1023 & ~w1024;
assign w1027 = ~w1025 & w1026;
assign w1028 = (w1027 & ~w536) | (w1027 & w24283) | (~w536 & w24283);
assign w1029 = a[8] & ~w1028;
assign w1030 = ~a[8] & w1028;
assign w1031 = ~w1029 & ~w1030;
assign w1032 = ~w972 & ~w975;
assign w1033 = w930 & w941;
assign w1034 = ~a[17] & ~b[0];
assign w1035 = ~a[18] & b[0];
assign w1036 = ~w1034 & ~w1035;
assign w1037 = b[3] & w834;
assign w1038 = b[2] & w838;
assign w1039 = b[1] & ~w934;
assign w1040 = ~w1037 & ~w1038;
assign w1041 = ~w1039 & w1040;
assign w1042 = w1041 & w24284;
assign w1043 = (~w1036 & ~w1041) | (~w1036 & w24285) | (~w1041 & w24285);
assign w1044 = ~w1042 & ~w1043;
assign w1045 = w1033 & w1044;
assign w1046 = ~w1033 & ~w1044;
assign w1047 = ~w1045 & ~w1046;
assign w1048 = b[6] & w575;
assign w1049 = b[5] & w573;
assign w1050 = b[4] & ~w649;
assign w1051 = w157 & w569;
assign w1052 = ~w1048 & ~w1049;
assign w1053 = ~w1050 & w1052;
assign w1054 = (a[14] & w1051) | (a[14] & w24286) | (w1051 & w24286);
assign w1055 = ~w1051 & w24287;
assign w1056 = ~w1054 & ~w1055;
assign w1057 = ~w1047 & w1056;
assign w1058 = w1047 & ~w1056;
assign w1059 = ~w1057 & ~w1058;
assign w1060 = (~w955 & w958) | (~w955 & w24288) | (w958 & w24288);
assign w1061 = w1059 & ~w1060;
assign w1062 = ~w1059 & w1060;
assign w1063 = ~w1061 & ~w1062;
assign w1064 = b[8] & w358;
assign w1065 = b[9] & w360;
assign w1066 = b[7] & ~w419;
assign w1067 = ~w1064 & ~w1065;
assign w1068 = ~w1066 & w1067;
assign w1069 = (w1068 & ~w322) | (w1068 & w24289) | (~w322 & w24289);
assign w1070 = a[11] & ~w1069;
assign w1071 = ~a[11] & w1069;
assign w1072 = ~w1070 & ~w1071;
assign w1073 = w1063 & w1072;
assign w1074 = ~w1063 & ~w1072;
assign w1075 = ~w1073 & ~w1074;
assign w1076 = w1032 & ~w1075;
assign w1077 = ~w1032 & w1075;
assign w1078 = ~w1076 & ~w1077;
assign w1079 = ~w1031 & ~w1078;
assign w1080 = w1031 & w1078;
assign w1081 = ~w1079 & ~w1080;
assign w1082 = (~w987 & ~w928) | (~w987 & w24290) | (~w928 & w24290);
assign w1083 = w1081 & w1082;
assign w1084 = ~w1081 & ~w1082;
assign w1085 = ~w1083 & ~w1084;
assign w1086 = w102 & w24291;
assign w1087 = b[15] & w68;
assign w1088 = b[14] & w61;
assign w1089 = ~w1087 & ~w1088;
assign w1090 = ~w1086 & w1089;
assign w1091 = (w1090 & w799) | (w1090 & w24292) | (w799 & w24292);
assign w1092 = a[5] & ~w1091;
assign w1093 = (w799 & w24293) | (w799 & w24294) | (w24293 & w24294);
assign w1094 = ~w1092 & ~w1093;
assign w1095 = w1085 & w1094;
assign w1096 = ~w1085 & ~w1094;
assign w1097 = ~w1095 & ~w1096;
assign w1098 = w1022 & w1097;
assign w1099 = ~w1022 & ~w1097;
assign w1100 = ~w1098 & ~w1099;
assign w1101 = w4 & w24295;
assign w1102 = b[17] & w9;
assign w1103 = ~b[17] & ~b[18];
assign w1104 = b[17] & b[18];
assign w1105 = ~w1103 & ~w1104;
assign w1106 = ~w1105 & w25724;
assign w1107 = (w1005 & w24297) | (w1005 & w24298) | (w24297 & w24298);
assign w1108 = ~w1106 & ~w1107;
assign w1109 = ~w1101 & ~w1102;
assign w1110 = (w1109 & w1108) | (w1109 & w24299) | (w1108 & w24299);
assign w1111 = (a[2] & ~w24) | (a[2] & w24300) | (~w24 & w24300);
assign w1112 = w1110 & ~w1111;
assign w1113 = a[2] & ~w1110;
assign w1114 = ~w1112 & ~w1113;
assign w1115 = ~w1100 & w1114;
assign w1116 = w1100 & ~w1114;
assign w1117 = ~w1115 & ~w1116;
assign w1118 = (~w1016 & ~w1018) | (~w1016 & w24301) | (~w1018 & w24301);
assign w1119 = w1117 & w1118;
assign w1120 = ~w1117 & ~w1118;
assign w1121 = ~w1119 & ~w1120;
assign w1122 = w102 & w24302;
assign w1123 = b[16] & w68;
assign w1124 = b[15] & w61;
assign w1125 = ~w1123 & ~w1124;
assign w1126 = ~w1122 & w1125;
assign w1127 = (w1126 & ~w905) | (w1126 & w24303) | (~w905 & w24303);
assign w1128 = a[5] & ~w1127;
assign w1129 = ~a[5] & w1127;
assign w1130 = ~w1128 & ~w1129;
assign w1131 = (~w1057 & w1060) | (~w1057 & w24304) | (w1060 & w24304);
assign w1132 = b[4] & w834;
assign w1133 = b[3] & w838;
assign w1134 = b[2] & ~w934;
assign w1135 = w84 & w832;
assign w1136 = ~w1132 & ~w1133;
assign w1137 = ~w1134 & w1136;
assign w1138 = ~w1135 & w1137;
assign w1139 = a[17] & ~w1138;
assign w1140 = ~a[17] & w1138;
assign w1141 = ~w1139 & ~w1140;
assign w1142 = a[17] & a[18];
assign w1143 = ~a[17] & ~a[18];
assign w1144 = ~w1142 & ~w1143;
assign w1145 = b[0] & w1144;
assign w1146 = w1144 & w24305;
assign w1147 = ~a[19] & a[20];
assign w1148 = a[19] & ~a[20];
assign w1149 = ~w1147 & ~w1148;
assign w1150 = w1144 & ~w1149;
assign w1151 = ~w8 & w1150;
assign w1152 = ~a[19] & ~w1142;
assign w1153 = a[19] & ~w1143;
assign w1154 = ~w1152 & ~w1153;
assign w1155 = b[0] & w1154;
assign w1156 = w1144 & w1149;
assign w1157 = b[1] & w1156;
assign w1158 = ~w1151 & ~w1155;
assign w1159 = w1158 & w24306;
assign w1160 = (w1146 & ~w1158) | (w1146 & w24307) | (~w1158 & w24307);
assign w1161 = ~w1159 & ~w1160;
assign w1162 = ~w1141 & ~w1161;
assign w1163 = w1141 & w1161;
assign w1164 = ~w1162 & ~w1163;
assign w1165 = ~w1042 & ~w1145;
assign w1166 = ~w1046 & ~w1165;
assign w1167 = w1164 & w1166;
assign w1168 = ~w1164 & ~w1166;
assign w1169 = ~w1167 & ~w1168;
assign w1170 = b[7] & w575;
assign w1171 = b[6] & w573;
assign w1172 = b[5] & ~w649;
assign w1173 = ~w1170 & ~w1171;
assign w1174 = ~w1172 & w1173;
assign w1175 = (w1174 & ~w216) | (w1174 & w24308) | (~w216 & w24308);
assign w1176 = a[14] & ~w1175;
assign w1177 = ~a[14] & w1175;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = w1169 & w1178;
assign w1180 = ~w1169 & ~w1178;
assign w1181 = ~w1179 & ~w1180;
assign w1182 = w1131 & w1181;
assign w1183 = ~w1131 & ~w1181;
assign w1184 = ~w1182 & ~w1183;
assign w1185 = b[9] & w358;
assign w1186 = b[10] & w360;
assign w1187 = b[8] & ~w419;
assign w1188 = ~w1185 & ~w1186;
assign w1189 = ~w1187 & w1188;
assign w1190 = (w1189 & ~w397) | (w1189 & w24309) | (~w397 & w24309);
assign w1191 = a[11] & ~w1190;
assign w1192 = ~a[11] & w1190;
assign w1193 = ~w1191 & ~w1192;
assign w1194 = ~w1184 & w1193;
assign w1195 = w1184 & ~w1193;
assign w1196 = ~w1194 & ~w1195;
assign w1197 = (~w1073 & w1032) | (~w1073 & w24310) | (w1032 & w24310);
assign w1198 = ~w1196 & w1197;
assign w1199 = w1196 & ~w1197;
assign w1200 = ~w1198 & ~w1199;
assign w1201 = b[12] & w183;
assign w1202 = b[13] & w185;
assign w1203 = b[11] & ~w237;
assign w1204 = ~w1201 & ~w1202;
assign w1205 = ~w1203 & w1204;
assign w1206 = (w1205 & ~w628) | (w1205 & w24311) | (~w628 & w24311);
assign w1207 = a[8] & ~w1206;
assign w1208 = ~a[8] & w1206;
assign w1209 = ~w1207 & ~w1208;
assign w1210 = ~w1200 & ~w1209;
assign w1211 = w1200 & w1209;
assign w1212 = ~w1210 & ~w1211;
assign w1213 = ~w1080 & ~w1083;
assign w1214 = w1212 & w1213;
assign w1215 = ~w1212 & ~w1213;
assign w1216 = ~w1214 & ~w1215;
assign w1217 = w1130 & ~w1216;
assign w1218 = ~w1130 & w1216;
assign w1219 = ~w1217 & ~w1218;
assign w1220 = (~w1096 & ~w1022) | (~w1096 & w24312) | (~w1022 & w24312);
assign w1221 = ~w1219 & ~w1220;
assign w1222 = w1219 & w1220;
assign w1223 = ~w1221 & ~w1222;
assign w1224 = w4 & w24313;
assign w1225 = b[18] & w9;
assign w1226 = ~b[18] & ~b[19];
assign w1227 = b[18] & b[19];
assign w1228 = ~w1226 & ~w1227;
assign w1229 = ~w1228 & w25725;
assign w1230 = (w1005 & w24316) | (w1005 & w24317) | (w24316 & w24317);
assign w1231 = ~w1229 & ~w1230;
assign w1232 = ~w1224 & ~w1225;
assign w1233 = (w1232 & w1231) | (w1232 & w24318) | (w1231 & w24318);
assign w1234 = (a[2] & ~w24) | (a[2] & w24319) | (~w24 & w24319);
assign w1235 = w1233 & ~w1234;
assign w1236 = a[2] & ~w1233;
assign w1237 = ~w1235 & ~w1236;
assign w1238 = w1223 & w1237;
assign w1239 = ~w1223 & ~w1237;
assign w1240 = ~w1238 & ~w1239;
assign w1241 = ~w1115 & ~w1119;
assign w1242 = w1240 & w1241;
assign w1243 = ~w1240 & ~w1241;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = ~w1217 & ~w1222;
assign w1246 = b[14] & w185;
assign w1247 = b[12] & ~w237;
assign w1248 = b[13] & w183;
assign w1249 = ~w1246 & ~w1247;
assign w1250 = ~w1248 & w1249;
assign w1251 = (w1250 & ~w714) | (w1250 & w24320) | (~w714 & w24320);
assign w1252 = a[8] & ~w1251;
assign w1253 = ~a[8] & w1251;
assign w1254 = ~w1252 & ~w1253;
assign w1255 = ~w1194 & ~w1199;
assign w1256 = b[3] & ~w934;
assign w1257 = b[5] & w834;
assign w1258 = b[4] & w838;
assign w1259 = w116 & w832;
assign w1260 = ~w1256 & ~w1257;
assign w1261 = (a[17] & w1259) | (a[17] & w24321) | (w1259 & w24321);
assign w1262 = ~w1259 & w24322;
assign w1263 = ~w1261 & ~w1262;
assign w1264 = (a[20] & ~w1144) | (a[20] & w24323) | (~w1144 & w24323);
assign w1265 = w1158 & w24324;
assign w1266 = a[20] & ~w1265;
assign w1267 = b[2] & w1156;
assign w1268 = w22 & w1150;
assign w1269 = b[1] & w1154;
assign w1270 = w1142 & w1148;
assign w1271 = w1143 & w1147;
assign w1272 = ~w1270 & ~w1271;
assign w1273 = b[0] & ~w1272;
assign w1274 = ~w1267 & ~w1268;
assign w1275 = ~w1269 & ~w1273;
assign w1276 = w1274 & w1275;
assign w1277 = ~w1266 & w1276;
assign w1278 = w1266 & ~w1276;
assign w1279 = ~w1277 & ~w1278;
assign w1280 = w1263 & w1279;
assign w1281 = ~w1263 & ~w1279;
assign w1282 = ~w1280 & ~w1281;
assign w1283 = (~w1163 & ~w1164) | (~w1163 & w24325) | (~w1164 & w24325);
assign w1284 = ~w1282 & w1283;
assign w1285 = w1282 & ~w1283;
assign w1286 = ~w1284 & ~w1285;
assign w1287 = b[6] & ~w649;
assign w1288 = b[8] & w575;
assign w1289 = b[7] & w573;
assign w1290 = ~w1287 & ~w1288;
assign w1291 = ~w1289 & w1290;
assign w1292 = (w1291 & ~w270) | (w1291 & w24326) | (~w270 & w24326);
assign w1293 = a[14] & ~w1292;
assign w1294 = ~a[14] & w1292;
assign w1295 = ~w1293 & ~w1294;
assign w1296 = ~w1286 & ~w1295;
assign w1297 = w1286 & w1295;
assign w1298 = ~w1296 & ~w1297;
assign w1299 = (~w1180 & ~w1181) | (~w1180 & w24327) | (~w1181 & w24327);
assign w1300 = w1298 & w1299;
assign w1301 = ~w1298 & ~w1299;
assign w1302 = ~w1300 & ~w1301;
assign w1303 = b[10] & w358;
assign w1304 = b[11] & w360;
assign w1305 = b[9] & ~w419;
assign w1306 = ~w1303 & ~w1304;
assign w1307 = ~w1305 & w1306;
assign w1308 = (w1307 & ~w469) | (w1307 & w24328) | (~w469 & w24328);
assign w1309 = a[11] & ~w1308;
assign w1310 = ~a[11] & w1308;
assign w1311 = ~w1309 & ~w1310;
assign w1312 = ~w1302 & ~w1311;
assign w1313 = w1302 & w1311;
assign w1314 = ~w1312 & ~w1313;
assign w1315 = w1255 & w1314;
assign w1316 = ~w1255 & ~w1314;
assign w1317 = ~w1315 & ~w1316;
assign w1318 = w1254 & ~w1317;
assign w1319 = ~w1254 & w1317;
assign w1320 = ~w1318 & ~w1319;
assign w1321 = (~w1210 & ~w1213) | (~w1210 & w24329) | (~w1213 & w24329);
assign w1322 = w1320 & w1321;
assign w1323 = ~w1320 & ~w1321;
assign w1324 = ~w1322 & ~w1323;
assign w1325 = w102 & w24330;
assign w1326 = b[17] & w68;
assign w1327 = b[16] & w61;
assign w1328 = ~w1326 & ~w1327;
assign w1329 = ~w1325 & w1328;
assign w1330 = (w1329 & ~w1008) | (w1329 & w24331) | (~w1008 & w24331);
assign w1331 = a[5] & ~w1330;
assign w1332 = ~a[5] & w1330;
assign w1333 = ~w1331 & ~w1332;
assign w1334 = ~w1324 & ~w1333;
assign w1335 = w1324 & w1333;
assign w1336 = ~w1334 & ~w1335;
assign w1337 = w1245 & w1336;
assign w1338 = ~w1245 & ~w1336;
assign w1339 = ~w1337 & ~w1338;
assign w1340 = w4 & w24332;
assign w1341 = b[19] & w9;
assign w1342 = ~b[19] & ~b[20];
assign w1343 = b[19] & b[20];
assign w1344 = ~w1342 & ~w1343;
assign w1345 = (w1005 & w24335) | (w1005 & w24336) | (w24335 & w24336);
assign w1346 = (~w1005 & w24337) | (~w1005 & w24338) | (w24337 & w24338);
assign w1347 = ~w1345 & ~w1346;
assign w1348 = ~w1340 & ~w1341;
assign w1349 = (w1348 & ~w1347) | (w1348 & w24339) | (~w1347 & w24339);
assign w1350 = (a[2] & ~w24) | (a[2] & w24340) | (~w24 & w24340);
assign w1351 = w1349 & ~w1350;
assign w1352 = (w1347 & w24341) | (w1347 & w24342) | (w24341 & w24342);
assign w1353 = ~w1351 & ~w1352;
assign w1354 = ~w1339 & w1353;
assign w1355 = w1339 & ~w1353;
assign w1356 = ~w1354 & ~w1355;
assign w1357 = (~w1239 & ~w1241) | (~w1239 & w24343) | (~w1241 & w24343);
assign w1358 = w1356 & w1357;
assign w1359 = ~w1356 & ~w1357;
assign w1360 = ~w1358 & ~w1359;
assign w1361 = w102 & w24344;
assign w1362 = b[18] & w68;
assign w1363 = b[17] & w61;
assign w1364 = ~w1362 & ~w1363;
assign w1365 = ~w1361 & w1364;
assign w1366 = (w1365 & w1108) | (w1365 & w24345) | (w1108 & w24345);
assign w1367 = a[5] & ~w1366;
assign w1368 = (w1108 & w24346) | (w1108 & w24347) | (w24346 & w24347);
assign w1369 = ~w1367 & ~w1368;
assign w1370 = ~w1318 & ~w1322;
assign w1371 = ~w1297 & ~w1300;
assign w1372 = w1265 & w1276;
assign w1373 = ~a[20] & ~b[0];
assign w1374 = ~a[21] & b[0];
assign w1375 = ~w1373 & ~w1374;
assign w1376 = b[3] & w1156;
assign w1377 = b[1] & ~w1272;
assign w1378 = b[2] & w1154;
assign w1379 = ~w1376 & ~w1377;
assign w1380 = ~w1378 & w1379;
assign w1381 = w1380 & w24348;
assign w1382 = (~w1375 & ~w1380) | (~w1375 & w24349) | (~w1380 & w24349);
assign w1383 = ~w1381 & ~w1382;
assign w1384 = w1372 & w1383;
assign w1385 = ~w1372 & ~w1383;
assign w1386 = ~w1384 & ~w1385;
assign w1387 = b[5] & w838;
assign w1388 = b[6] & w834;
assign w1389 = b[4] & ~w934;
assign w1390 = w157 & w832;
assign w1391 = ~w1387 & ~w1388;
assign w1392 = ~w1389 & w1391;
assign w1393 = (a[17] & w1390) | (a[17] & w24350) | (w1390 & w24350);
assign w1394 = ~w1390 & w24351;
assign w1395 = ~w1393 & ~w1394;
assign w1396 = ~w1386 & w1395;
assign w1397 = w1386 & ~w1395;
assign w1398 = ~w1396 & ~w1397;
assign w1399 = (~w1280 & w1283) | (~w1280 & w24352) | (w1283 & w24352);
assign w1400 = w1398 & ~w1399;
assign w1401 = ~w1398 & w1399;
assign w1402 = ~w1400 & ~w1401;
assign w1403 = b[8] & w573;
assign w1404 = b[7] & ~w649;
assign w1405 = b[9] & w575;
assign w1406 = w322 & w569;
assign w1407 = ~w1403 & ~w1404;
assign w1408 = ~w1405 & w1407;
assign w1409 = ~w1406 & w1408;
assign w1410 = a[14] & ~w1409;
assign w1411 = ~a[14] & w1409;
assign w1412 = ~w1410 & ~w1411;
assign w1413 = w1402 & w1412;
assign w1414 = ~w1402 & ~w1412;
assign w1415 = ~w1413 & ~w1414;
assign w1416 = ~w1371 & w1415;
assign w1417 = w1371 & ~w1415;
assign w1418 = ~w1416 & ~w1417;
assign w1419 = b[11] & w358;
assign w1420 = b[12] & w360;
assign w1421 = b[10] & ~w419;
assign w1422 = w354 & w536;
assign w1423 = ~w1419 & ~w1420;
assign w1424 = ~w1421 & w1423;
assign w1425 = ~w1422 & w1424;
assign w1426 = a[11] & ~w1425;
assign w1427 = ~a[11] & w1425;
assign w1428 = ~w1426 & ~w1427;
assign w1429 = ~w1418 & ~w1428;
assign w1430 = w1418 & w1428;
assign w1431 = ~w1429 & ~w1430;
assign w1432 = (~w1312 & ~w1255) | (~w1312 & w24610) | (~w1255 & w24610);
assign w1433 = w1431 & w1432;
assign w1434 = ~w1431 & ~w1432;
assign w1435 = ~w1433 & ~w1434;
assign w1436 = b[13] & ~w237;
assign w1437 = b[14] & w183;
assign w1438 = b[15] & w185;
assign w1439 = w179 & ~w799;
assign w1440 = ~w1436 & ~w1437;
assign w1441 = ~w1438 & w1440;
assign w1442 = ~w1439 & w1441;
assign w1443 = a[8] & ~w1442;
assign w1444 = ~a[8] & w1442;
assign w1445 = ~w1443 & ~w1444;
assign w1446 = w1435 & w1445;
assign w1447 = ~w1435 & ~w1445;
assign w1448 = ~w1446 & ~w1447;
assign w1449 = w1370 & w1448;
assign w1450 = ~w1370 & ~w1448;
assign w1451 = ~w1449 & ~w1450;
assign w1452 = w1369 & ~w1451;
assign w1453 = ~w1369 & w1451;
assign w1454 = ~w1452 & ~w1453;
assign w1455 = (~w1334 & ~w1245) | (~w1334 & w24355) | (~w1245 & w24355);
assign w1456 = ~w1454 & ~w1455;
assign w1457 = w1454 & w1455;
assign w1458 = ~w1456 & ~w1457;
assign w1459 = b[21] & w11;
assign w1460 = b[20] & w9;
assign w1461 = ~w1343 & ~w1346;
assign w1462 = ~b[20] & ~b[21];
assign w1463 = b[20] & b[21];
assign w1464 = ~w1462 & ~w1463;
assign w1465 = w1461 & ~w1464;
assign w1466 = ~w1461 & w1464;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = w5 & w1467;
assign w1469 = ~w1459 & ~w1460;
assign w1470 = ~w1468 & w1469;
assign w1471 = b[19] & w24;
assign w1472 = a[2] & ~w1471;
assign w1473 = w1470 & ~w1472;
assign w1474 = a[2] & ~w1470;
assign w1475 = ~w1473 & ~w1474;
assign w1476 = w1458 & w1475;
assign w1477 = ~w1458 & ~w1475;
assign w1478 = ~w1476 & ~w1477;
assign w1479 = ~w1354 & ~w1358;
assign w1480 = w1478 & w1479;
assign w1481 = ~w1478 & ~w1479;
assign w1482 = ~w1480 & ~w1481;
assign w1483 = b[16] & w185;
assign w1484 = b[14] & ~w237;
assign w1485 = b[15] & w183;
assign w1486 = w179 & w905;
assign w1487 = ~w1483 & ~w1484;
assign w1488 = ~w1485 & w1487;
assign w1489 = ~w1486 & w1488;
assign w1490 = a[8] & ~w1489;
assign w1491 = ~a[8] & w1489;
assign w1492 = ~w1490 & ~w1491;
assign w1493 = ~w1430 & ~w1433;
assign w1494 = (~w1396 & w1399) | (~w1396 & w24611) | (w1399 & w24611);
assign w1495 = b[3] & w1154;
assign w1496 = b[2] & ~w1272;
assign w1497 = b[4] & w1156;
assign w1498 = w84 & w1150;
assign w1499 = ~w1495 & ~w1496;
assign w1500 = ~w1497 & w1499;
assign w1501 = ~w1498 & w1500;
assign w1502 = a[20] & ~w1501;
assign w1503 = ~a[20] & w1501;
assign w1504 = ~w1502 & ~w1503;
assign w1505 = a[20] & a[21];
assign w1506 = ~a[20] & ~a[21];
assign w1507 = ~w1505 & ~w1506;
assign w1508 = b[0] & w1507;
assign w1509 = a[23] & w1508;
assign w1510 = a[22] & ~a[23];
assign w1511 = ~a[22] & a[23];
assign w1512 = ~w1510 & ~w1511;
assign w1513 = w1507 & ~w1512;
assign w1514 = ~w8 & w1513;
assign w1515 = ~a[22] & ~w1505;
assign w1516 = a[22] & ~w1506;
assign w1517 = ~w1515 & ~w1516;
assign w1518 = b[0] & w1517;
assign w1519 = w1507 & w1512;
assign w1520 = b[1] & w1519;
assign w1521 = ~w1514 & ~w1518;
assign w1522 = ~w1520 & w1521;
assign w1523 = ~w1509 & w1522;
assign w1524 = w1509 & ~w1522;
assign w1525 = ~w1523 & ~w1524;
assign w1526 = ~w1504 & ~w1525;
assign w1527 = w1504 & w1525;
assign w1528 = ~w1526 & ~w1527;
assign w1529 = ~w1381 & ~w1508;
assign w1530 = ~w1385 & ~w1529;
assign w1531 = w1528 & w1530;
assign w1532 = ~w1528 & ~w1530;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = b[6] & w838;
assign w1535 = b[5] & ~w934;
assign w1536 = b[7] & w834;
assign w1537 = w216 & w832;
assign w1538 = ~w1534 & ~w1535;
assign w1539 = ~w1536 & w1538;
assign w1540 = ~w1537 & w1539;
assign w1541 = a[17] & ~w1540;
assign w1542 = ~a[17] & w1540;
assign w1543 = ~w1541 & ~w1542;
assign w1544 = w1533 & w1543;
assign w1545 = ~w1533 & ~w1543;
assign w1546 = ~w1544 & ~w1545;
assign w1547 = w1494 & w1546;
assign w1548 = ~w1494 & ~w1546;
assign w1549 = ~w1547 & ~w1548;
assign w1550 = b[10] & w575;
assign w1551 = b[8] & ~w649;
assign w1552 = b[9] & w573;
assign w1553 = w397 & w569;
assign w1554 = ~w1550 & ~w1551;
assign w1555 = ~w1552 & w1554;
assign w1556 = ~w1553 & w1555;
assign w1557 = a[14] & ~w1556;
assign w1558 = ~a[14] & w1556;
assign w1559 = ~w1557 & ~w1558;
assign w1560 = ~w1549 & w1559;
assign w1561 = w1549 & ~w1559;
assign w1562 = ~w1560 & ~w1561;
assign w1563 = (~w1413 & w1371) | (~w1413 & w24612) | (w1371 & w24612);
assign w1564 = ~w1562 & w1563;
assign w1565 = w1562 & ~w1563;
assign w1566 = ~w1564 & ~w1565;
assign w1567 = b[12] & w358;
assign w1568 = b[13] & w360;
assign w1569 = b[11] & ~w419;
assign w1570 = w354 & w628;
assign w1571 = ~w1567 & ~w1568;
assign w1572 = ~w1569 & w1571;
assign w1573 = ~w1570 & w1572;
assign w1574 = a[11] & ~w1573;
assign w1575 = ~a[11] & w1573;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = ~w1566 & ~w1576;
assign w1578 = w1566 & w1576;
assign w1579 = ~w1577 & ~w1578;
assign w1580 = w1493 & w1579;
assign w1581 = ~w1493 & ~w1579;
assign w1582 = ~w1580 & ~w1581;
assign w1583 = w1492 & ~w1582;
assign w1584 = ~w1492 & w1582;
assign w1585 = ~w1583 & ~w1584;
assign w1586 = (~w1447 & ~w1370) | (~w1447 & w24613) | (~w1370 & w24613);
assign w1587 = w1585 & w1586;
assign w1588 = ~w1585 & ~w1586;
assign w1589 = ~w1587 & ~w1588;
assign w1590 = b[17] & w103;
assign w1591 = b[18] & w61;
assign w1592 = b[19] & w68;
assign w1593 = w66 & ~w1231;
assign w1594 = ~w1591 & ~w1592;
assign w1595 = ~w1590 & w1594;
assign w1596 = ~w1593 & w1595;
assign w1597 = a[5] & ~w1596;
assign w1598 = ~a[5] & w1596;
assign w1599 = ~w1597 & ~w1598;
assign w1600 = w1589 & w1599;
assign w1601 = ~w1589 & ~w1599;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = ~w1452 & ~w1457;
assign w1604 = w1602 & w1603;
assign w1605 = ~w1602 & ~w1603;
assign w1606 = ~w1604 & ~w1605;
assign w1607 = b[22] & w11;
assign w1608 = b[21] & w9;
assign w1609 = ~w1463 & ~w1466;
assign w1610 = ~b[21] & ~b[22];
assign w1611 = b[21] & b[22];
assign w1612 = ~w1610 & ~w1611;
assign w1613 = ~w1609 & w1612;
assign w1614 = w1609 & ~w1612;
assign w1615 = ~w1613 & ~w1614;
assign w1616 = w5 & w1615;
assign w1617 = ~w1607 & ~w1608;
assign w1618 = ~w1616 & w1617;
assign w1619 = b[20] & w24;
assign w1620 = a[2] & ~w1619;
assign w1621 = w1618 & ~w1620;
assign w1622 = a[2] & ~w1618;
assign w1623 = ~w1621 & ~w1622;
assign w1624 = w1606 & ~w1623;
assign w1625 = ~w1606 & w1623;
assign w1626 = ~w1624 & ~w1625;
assign w1627 = (~w1477 & ~w1479) | (~w1477 & w24356) | (~w1479 & w24356);
assign w1628 = w1626 & w1627;
assign w1629 = ~w1626 & ~w1627;
assign w1630 = ~w1628 & ~w1629;
assign w1631 = b[18] & w103;
assign w1632 = b[20] & w68;
assign w1633 = b[19] & w61;
assign w1634 = w66 & w1347;
assign w1635 = ~w1632 & ~w1633;
assign w1636 = ~w1631 & w1635;
assign w1637 = ~w1634 & w1636;
assign w1638 = a[5] & ~w1637;
assign w1639 = ~a[5] & w1637;
assign w1640 = ~w1638 & ~w1639;
assign w1641 = ~w1583 & ~w1587;
assign w1642 = b[17] & w185;
assign w1643 = b[15] & ~w237;
assign w1644 = b[16] & w183;
assign w1645 = w179 & w1008;
assign w1646 = ~w1642 & ~w1643;
assign w1647 = ~w1644 & w1646;
assign w1648 = ~w1645 & w1647;
assign w1649 = a[8] & ~w1648;
assign w1650 = ~a[8] & w1648;
assign w1651 = ~w1649 & ~w1650;
assign w1652 = b[14] & w360;
assign w1653 = b[13] & w358;
assign w1654 = b[12] & ~w419;
assign w1655 = w354 & w714;
assign w1656 = ~w1652 & ~w1653;
assign w1657 = ~w1654 & w1656;
assign w1658 = ~w1655 & w1657;
assign w1659 = a[11] & ~w1658;
assign w1660 = ~a[11] & w1658;
assign w1661 = ~w1659 & ~w1660;
assign w1662 = ~w1560 & ~w1565;
assign w1663 = b[4] & w1154;
assign w1664 = b[3] & ~w1272;
assign w1665 = b[5] & w1156;
assign w1666 = w116 & w1150;
assign w1667 = ~w1663 & ~w1664;
assign w1668 = (a[20] & w1666) | (a[20] & w24756) | (w1666 & w24756);
assign w1669 = ~w1666 & w24757;
assign w1670 = ~w1668 & ~w1669;
assign w1671 = (a[23] & ~w1507) | (a[23] & w24915) | (~w1507 & w24915);
assign w1672 = w1521 & w24758;
assign w1673 = a[23] & ~w1672;
assign w1674 = w1505 & w1510;
assign w1675 = w1506 & w1511;
assign w1676 = ~w1674 & ~w1675;
assign w1677 = b[0] & ~w1676;
assign w1678 = b[1] & w1517;
assign w1679 = w22 & w1513;
assign w1680 = b[2] & w1519;
assign w1681 = ~w1677 & ~w1678;
assign w1682 = ~w1679 & ~w1680;
assign w1683 = w1681 & w1682;
assign w1684 = ~w1673 & w1683;
assign w1685 = w1673 & ~w1683;
assign w1686 = ~w1684 & ~w1685;
assign w1687 = w1670 & w1686;
assign w1688 = ~w1670 & ~w1686;
assign w1689 = ~w1687 & ~w1688;
assign w1690 = (~w1527 & ~w1528) | (~w1527 & w24614) | (~w1528 & w24614);
assign w1691 = ~w1689 & w1690;
assign w1692 = w1689 & ~w1690;
assign w1693 = ~w1691 & ~w1692;
assign w1694 = b[7] & w838;
assign w1695 = b[6] & ~w934;
assign w1696 = b[8] & w834;
assign w1697 = w270 & w832;
assign w1698 = ~w1694 & ~w1695;
assign w1699 = ~w1696 & w1698;
assign w1700 = ~w1697 & w1699;
assign w1701 = a[17] & ~w1700;
assign w1702 = ~a[17] & w1700;
assign w1703 = ~w1701 & ~w1702;
assign w1704 = ~w1693 & ~w1703;
assign w1705 = w1693 & w1703;
assign w1706 = ~w1704 & ~w1705;
assign w1707 = (~w1545 & ~w1546) | (~w1545 & w24615) | (~w1546 & w24615);
assign w1708 = w1706 & w1707;
assign w1709 = ~w1706 & ~w1707;
assign w1710 = ~w1708 & ~w1709;
assign w1711 = b[11] & w575;
assign w1712 = b[10] & w573;
assign w1713 = b[9] & ~w649;
assign w1714 = w469 & w569;
assign w1715 = ~w1711 & ~w1712;
assign w1716 = ~w1713 & w1715;
assign w1717 = ~w1714 & w1716;
assign w1718 = a[14] & ~w1717;
assign w1719 = ~a[14] & w1717;
assign w1720 = ~w1718 & ~w1719;
assign w1721 = ~w1710 & ~w1720;
assign w1722 = w1710 & w1720;
assign w1723 = ~w1721 & ~w1722;
assign w1724 = w1662 & w1723;
assign w1725 = ~w1662 & ~w1723;
assign w1726 = ~w1724 & ~w1725;
assign w1727 = w1661 & ~w1726;
assign w1728 = ~w1661 & w1726;
assign w1729 = ~w1727 & ~w1728;
assign w1730 = (~w1577 & ~w1493) | (~w1577 & w24357) | (~w1493 & w24357);
assign w1731 = w1729 & w1730;
assign w1732 = ~w1729 & ~w1730;
assign w1733 = ~w1731 & ~w1732;
assign w1734 = ~w1651 & ~w1733;
assign w1735 = w1651 & w1733;
assign w1736 = ~w1734 & ~w1735;
assign w1737 = ~w1641 & ~w1736;
assign w1738 = w1641 & w1736;
assign w1739 = ~w1737 & ~w1738;
assign w1740 = w1640 & ~w1739;
assign w1741 = ~w1640 & w1739;
assign w1742 = ~w1740 & ~w1741;
assign w1743 = (~w1601 & ~w1603) | (~w1601 & w24616) | (~w1603 & w24616);
assign w1744 = ~w1742 & ~w1743;
assign w1745 = w1742 & w1743;
assign w1746 = ~w1744 & ~w1745;
assign w1747 = b[23] & w11;
assign w1748 = b[22] & w9;
assign w1749 = ~b[22] & ~b[23];
assign w1750 = b[22] & b[23];
assign w1751 = ~w1749 & ~w1750;
assign w1752 = ~w1611 & ~w1613;
assign w1753 = w1751 & ~w1752;
assign w1754 = ~w1751 & w1752;
assign w1755 = ~w1753 & ~w1754;
assign w1756 = w5 & w1755;
assign w1757 = ~w1747 & ~w1748;
assign w1758 = ~w1756 & w1757;
assign w1759 = b[21] & w24;
assign w1760 = a[2] & ~w1759;
assign w1761 = w1758 & ~w1760;
assign w1762 = a[2] & ~w1758;
assign w1763 = ~w1761 & ~w1762;
assign w1764 = w1746 & w1763;
assign w1765 = ~w1746 & ~w1763;
assign w1766 = ~w1764 & ~w1765;
assign w1767 = ~w1625 & ~w1628;
assign w1768 = ~w1766 & ~w1767;
assign w1769 = w1766 & w1767;
assign w1770 = ~w1768 & ~w1769;
assign w1771 = ~w1740 & ~w1745;
assign w1772 = b[19] & w103;
assign w1773 = b[20] & w61;
assign w1774 = b[21] & w68;
assign w1775 = w66 & w1467;
assign w1776 = ~w1773 & ~w1774;
assign w1777 = ~w1772 & w1776;
assign w1778 = ~w1775 & w1777;
assign w1779 = a[5] & ~w1778;
assign w1780 = ~a[5] & w1778;
assign w1781 = ~w1779 & ~w1780;
assign w1782 = b[16] & ~w237;
assign w1783 = b[18] & w185;
assign w1784 = b[17] & w183;
assign w1785 = w179 & ~w1108;
assign w1786 = ~w1782 & ~w1783;
assign w1787 = ~w1784 & w1786;
assign w1788 = ~w1785 & w1787;
assign w1789 = a[8] & ~w1788;
assign w1790 = ~a[8] & w1788;
assign w1791 = ~w1789 & ~w1790;
assign w1792 = b[11] & w573;
assign w1793 = b[12] & w575;
assign w1794 = b[10] & ~w649;
assign w1795 = w536 & w569;
assign w1796 = ~w1792 & ~w1793;
assign w1797 = ~w1794 & w1796;
assign w1798 = ~w1795 & w1797;
assign w1799 = a[14] & ~w1798;
assign w1800 = ~a[14] & w1798;
assign w1801 = ~w1799 & ~w1800;
assign w1802 = ~w1705 & ~w1708;
assign w1803 = w1672 & w1683;
assign w1804 = ~a[23] & ~b[0];
assign w1805 = ~a[24] & b[0];
assign w1806 = ~w1804 & ~w1805;
assign w1807 = b[1] & ~w1676;
assign w1808 = b[3] & w1519;
assign w1809 = b[2] & w1517;
assign w1810 = ~w1807 & ~w1808;
assign w1811 = ~w1809 & w1810;
assign w1812 = w1811 & w24617;
assign w1813 = (~w1806 & ~w1811) | (~w1806 & w24618) | (~w1811 & w24618);
assign w1814 = ~w1812 & ~w1813;
assign w1815 = w1803 & w1814;
assign w1816 = ~w1803 & ~w1814;
assign w1817 = ~w1815 & ~w1816;
assign w1818 = b[4] & ~w1272;
assign w1819 = b[5] & w1154;
assign w1820 = b[6] & w1156;
assign w1821 = w157 & w1150;
assign w1822 = ~w1818 & ~w1819;
assign w1823 = ~w1820 & w1822;
assign w1824 = (a[20] & w1821) | (a[20] & w25101) | (w1821 & w25101);
assign w1825 = ~w1821 & w25102;
assign w1826 = ~w1824 & ~w1825;
assign w1827 = ~w1817 & w1826;
assign w1828 = w1817 & ~w1826;
assign w1829 = ~w1827 & ~w1828;
assign w1830 = (~w1687 & w1690) | (~w1687 & w24759) | (w1690 & w24759);
assign w1831 = w1829 & ~w1830;
assign w1832 = ~w1829 & w1830;
assign w1833 = ~w1831 & ~w1832;
assign w1834 = b[7] & ~w934;
assign w1835 = b[8] & w838;
assign w1836 = b[9] & w834;
assign w1837 = w322 & w832;
assign w1838 = ~w1834 & ~w1835;
assign w1839 = ~w1836 & w1838;
assign w1840 = ~w1837 & w1839;
assign w1841 = a[17] & ~w1840;
assign w1842 = ~a[17] & w1840;
assign w1843 = ~w1841 & ~w1842;
assign w1844 = w1833 & w1843;
assign w1845 = ~w1833 & ~w1843;
assign w1846 = ~w1844 & ~w1845;
assign w1847 = w1802 & ~w1846;
assign w1848 = ~w1802 & w1846;
assign w1849 = ~w1847 & ~w1848;
assign w1850 = ~w1801 & ~w1849;
assign w1851 = w1801 & w1849;
assign w1852 = ~w1850 & ~w1851;
assign w1853 = (~w1721 & ~w1662) | (~w1721 & w24760) | (~w1662 & w24760);
assign w1854 = w1852 & w1853;
assign w1855 = ~w1852 & ~w1853;
assign w1856 = ~w1854 & ~w1855;
assign w1857 = b[13] & ~w419;
assign w1858 = b[14] & w358;
assign w1859 = b[15] & w360;
assign w1860 = w354 & ~w799;
assign w1861 = ~w1857 & ~w1858;
assign w1862 = ~w1859 & w1861;
assign w1863 = ~w1860 & w1862;
assign w1864 = a[11] & ~w1863;
assign w1865 = ~a[11] & w1863;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = w1856 & w1866;
assign w1868 = ~w1856 & ~w1866;
assign w1869 = ~w1867 & ~w1868;
assign w1870 = ~w1727 & ~w1731;
assign w1871 = w1869 & w1870;
assign w1872 = ~w1869 & ~w1870;
assign w1873 = ~w1871 & ~w1872;
assign w1874 = ~w1791 & w1873;
assign w1875 = w1791 & ~w1873;
assign w1876 = ~w1874 & ~w1875;
assign w1877 = (~w1734 & ~w1641) | (~w1734 & w24358) | (~w1641 & w24358);
assign w1878 = w1876 & w1877;
assign w1879 = ~w1876 & ~w1877;
assign w1880 = ~w1878 & ~w1879;
assign w1881 = ~w1781 & ~w1880;
assign w1882 = w1781 & w1880;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = w1771 & w1883;
assign w1885 = ~w1771 & ~w1883;
assign w1886 = ~w1884 & ~w1885;
assign w1887 = b[24] & w11;
assign w1888 = b[23] & w9;
assign w1889 = ~w1750 & ~w1753;
assign w1890 = ~b[23] & ~b[24];
assign w1891 = b[23] & b[24];
assign w1892 = ~w1890 & ~w1891;
assign w1893 = w1889 & ~w1892;
assign w1894 = ~w1889 & w1892;
assign w1895 = ~w1893 & ~w1894;
assign w1896 = w5 & w1895;
assign w1897 = ~w1887 & ~w1888;
assign w1898 = ~w1896 & w1897;
assign w1899 = b[22] & w24;
assign w1900 = a[2] & ~w1899;
assign w1901 = w1898 & ~w1900;
assign w1902 = a[2] & ~w1898;
assign w1903 = ~w1901 & ~w1902;
assign w1904 = ~w1886 & w1903;
assign w1905 = w1886 & ~w1903;
assign w1906 = ~w1904 & ~w1905;
assign w1907 = (~w1765 & ~w1767) | (~w1765 & w24619) | (~w1767 & w24619);
assign w1908 = w1906 & w1907;
assign w1909 = ~w1906 & ~w1907;
assign w1910 = ~w1908 & ~w1909;
assign w1911 = ~w1904 & ~w1908;
assign w1912 = b[20] & w103;
assign w1913 = b[21] & w61;
assign w1914 = b[22] & w68;
assign w1915 = w66 & w1615;
assign w1916 = ~w1913 & ~w1914;
assign w1917 = ~w1912 & w1916;
assign w1918 = ~w1915 & w1917;
assign w1919 = a[5] & ~w1918;
assign w1920 = ~a[5] & w1918;
assign w1921 = ~w1919 & ~w1920;
assign w1922 = b[14] & ~w419;
assign w1923 = b[16] & w360;
assign w1924 = b[15] & w358;
assign w1925 = w354 & w905;
assign w1926 = ~w1922 & ~w1923;
assign w1927 = ~w1924 & w1926;
assign w1928 = ~w1925 & w1927;
assign w1929 = a[11] & ~w1928;
assign w1930 = ~a[11] & w1928;
assign w1931 = ~w1929 & ~w1930;
assign w1932 = (~w1827 & w1830) | (~w1827 & w24916) | (w1830 & w24916);
assign w1933 = b[2] & ~w1676;
assign w1934 = b[3] & w1517;
assign w1935 = b[4] & w1519;
assign w1936 = w84 & w1513;
assign w1937 = ~w1933 & ~w1934;
assign w1938 = ~w1935 & w1937;
assign w1939 = ~w1936 & w1938;
assign w1940 = a[23] & ~w1939;
assign w1941 = ~a[23] & w1939;
assign w1942 = ~w1940 & ~w1941;
assign w1943 = a[23] & a[24];
assign w1944 = ~a[23] & ~a[24];
assign w1945 = ~w1943 & ~w1944;
assign w1946 = b[0] & w1945;
assign w1947 = a[26] & w1946;
assign w1948 = a[25] & ~a[26];
assign w1949 = ~a[25] & a[26];
assign w1950 = ~w1948 & ~w1949;
assign w1951 = w1945 & ~w1950;
assign w1952 = ~w8 & w1951;
assign w1953 = ~a[25] & ~w1943;
assign w1954 = a[25] & ~w1944;
assign w1955 = ~w1953 & ~w1954;
assign w1956 = b[0] & w1955;
assign w1957 = w1945 & w1950;
assign w1958 = b[1] & w1957;
assign w1959 = ~w1952 & ~w1956;
assign w1960 = ~w1958 & w1959;
assign w1961 = ~w1947 & w1960;
assign w1962 = w1947 & ~w1960;
assign w1963 = ~w1961 & ~w1962;
assign w1964 = ~w1942 & ~w1963;
assign w1965 = w1942 & w1963;
assign w1966 = ~w1964 & ~w1965;
assign w1967 = ~w1812 & ~w1946;
assign w1968 = ~w1816 & ~w1967;
assign w1969 = w1966 & w1968;
assign w1970 = ~w1966 & ~w1968;
assign w1971 = ~w1969 & ~w1970;
assign w1972 = b[5] & ~w1272;
assign w1973 = b[7] & w1156;
assign w1974 = b[6] & w1154;
assign w1975 = w216 & w1150;
assign w1976 = ~w1972 & ~w1973;
assign w1977 = ~w1974 & w1976;
assign w1978 = ~w1975 & w1977;
assign w1979 = a[20] & ~w1978;
assign w1980 = ~a[20] & w1978;
assign w1981 = ~w1979 & ~w1980;
assign w1982 = w1971 & w1981;
assign w1983 = ~w1971 & ~w1981;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = w1932 & ~w1984;
assign w1986 = ~w1932 & w1984;
assign w1987 = ~w1985 & ~w1986;
assign w1988 = b[10] & w834;
assign w1989 = b[9] & w838;
assign w1990 = b[8] & ~w934;
assign w1991 = w397 & w832;
assign w1992 = ~w1988 & ~w1989;
assign w1993 = ~w1990 & w1992;
assign w1994 = ~w1991 & w1993;
assign w1995 = a[17] & ~w1994;
assign w1996 = ~a[17] & w1994;
assign w1997 = ~w1995 & ~w1996;
assign w1998 = w1987 & w1997;
assign w1999 = ~w1987 & ~w1997;
assign w2000 = ~w1998 & ~w1999;
assign w2001 = (~w1844 & w1802) | (~w1844 & w24761) | (w1802 & w24761);
assign w2002 = ~w2000 & w2001;
assign w2003 = w2000 & ~w2001;
assign w2004 = ~w2002 & ~w2003;
assign w2005 = b[12] & w573;
assign w2006 = b[13] & w575;
assign w2007 = b[11] & ~w649;
assign w2008 = w569 & w628;
assign w2009 = ~w2005 & ~w2006;
assign w2010 = ~w2007 & w2009;
assign w2011 = ~w2008 & w2010;
assign w2012 = a[14] & ~w2011;
assign w2013 = ~a[14] & w2011;
assign w2014 = ~w2012 & ~w2013;
assign w2015 = ~w2004 & ~w2014;
assign w2016 = w2004 & w2014;
assign w2017 = ~w2015 & ~w2016;
assign w2018 = ~w1851 & ~w1854;
assign w2019 = w2017 & w2018;
assign w2020 = ~w2017 & ~w2018;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = w1931 & ~w2021;
assign w2023 = ~w1931 & w2021;
assign w2024 = ~w2022 & ~w2023;
assign w2025 = (~w1868 & ~w1870) | (~w1868 & w24762) | (~w1870 & w24762);
assign w2026 = ~w2024 & ~w2025;
assign w2027 = w2024 & w2025;
assign w2028 = ~w2026 & ~w2027;
assign w2029 = b[19] & w185;
assign w2030 = b[17] & ~w237;
assign w2031 = b[18] & w183;
assign w2032 = w179 & ~w1231;
assign w2033 = ~w2029 & ~w2030;
assign w2034 = ~w2031 & w2033;
assign w2035 = ~w2032 & w2034;
assign w2036 = a[8] & ~w2035;
assign w2037 = ~a[8] & w2035;
assign w2038 = ~w2036 & ~w2037;
assign w2039 = w2028 & w2038;
assign w2040 = ~w2028 & ~w2038;
assign w2041 = ~w2039 & ~w2040;
assign w2042 = ~w1875 & ~w1878;
assign w2043 = w2041 & w2042;
assign w2044 = ~w2041 & ~w2042;
assign w2045 = ~w2043 & ~w2044;
assign w2046 = w1921 & ~w2045;
assign w2047 = ~w1921 & w2045;
assign w2048 = ~w2046 & ~w2047;
assign w2049 = (~w1881 & ~w1771) | (~w1881 & w24359) | (~w1771 & w24359);
assign w2050 = w2048 & w2049;
assign w2051 = ~w2048 & ~w2049;
assign w2052 = ~w2050 & ~w2051;
assign w2053 = b[25] & w11;
assign w2054 = b[24] & w9;
assign w2055 = ~b[24] & ~b[25];
assign w2056 = b[24] & b[25];
assign w2057 = ~w2055 & ~w2056;
assign w2058 = ~w1891 & ~w1894;
assign w2059 = w2057 & ~w2058;
assign w2060 = ~w2057 & w2058;
assign w2061 = ~w2059 & ~w2060;
assign w2062 = w5 & w2061;
assign w2063 = ~w2053 & ~w2054;
assign w2064 = ~w2062 & w2063;
assign w2065 = b[23] & w24;
assign w2066 = a[2] & ~w2065;
assign w2067 = w2064 & ~w2066;
assign w2068 = a[2] & ~w2064;
assign w2069 = ~w2067 & ~w2068;
assign w2070 = w2052 & w2069;
assign w2071 = ~w2052 & ~w2069;
assign w2072 = ~w2070 & ~w2071;
assign w2073 = w1911 & ~w2072;
assign w2074 = ~w1911 & w2072;
assign w2075 = ~w2073 & ~w2074;
assign w2076 = ~w2046 & ~w2050;
assign w2077 = b[18] & ~w237;
assign w2078 = b[20] & w185;
assign w2079 = b[19] & w183;
assign w2080 = w179 & w1347;
assign w2081 = ~w2077 & ~w2078;
assign w2082 = ~w2079 & w2081;
assign w2083 = ~w2080 & w2082;
assign w2084 = a[8] & ~w2083;
assign w2085 = ~a[8] & w2083;
assign w2086 = ~w2084 & ~w2085;
assign w2087 = ~w2022 & ~w2027;
assign w2088 = b[15] & ~w419;
assign w2089 = b[17] & w360;
assign w2090 = b[16] & w358;
assign w2091 = w354 & w1008;
assign w2092 = ~w2088 & ~w2089;
assign w2093 = ~w2090 & w2092;
assign w2094 = ~w2091 & w2093;
assign w2095 = a[11] & ~w2094;
assign w2096 = ~a[11] & w2094;
assign w2097 = ~w2095 & ~w2096;
assign w2098 = b[12] & ~w649;
assign w2099 = b[13] & w573;
assign w2100 = b[14] & w575;
assign w2101 = w569 & w714;
assign w2102 = ~w2098 & ~w2099;
assign w2103 = ~w2100 & w2102;
assign w2104 = ~w2101 & w2103;
assign w2105 = a[14] & ~w2104;
assign w2106 = ~a[14] & w2104;
assign w2107 = ~w2105 & ~w2106;
assign w2108 = ~w1998 & ~w2003;
assign w2109 = a[26] & ~w1946;
assign w2110 = w1959 & w24763;
assign w2111 = a[26] & ~w2110;
assign w2112 = w1943 & w1948;
assign w2113 = w1944 & w1949;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = b[0] & ~w2114;
assign w2116 = w22 & w1951;
assign w2117 = b[2] & w1957;
assign w2118 = b[1] & w1955;
assign w2119 = ~w2115 & ~w2116;
assign w2120 = ~w2117 & ~w2118;
assign w2121 = w2119 & w2120;
assign w2122 = ~w2111 & w2121;
assign w2123 = w2111 & ~w2121;
assign w2124 = ~w2122 & ~w2123;
assign w2125 = b[3] & ~w1676;
assign w2126 = b[5] & w1519;
assign w2127 = b[4] & w1517;
assign w2128 = ~w2125 & ~w2126;
assign w2129 = ~w2127 & w2128;
assign w2130 = (~a[23] & ~w116) | (~a[23] & w24620) | (~w116 & w24620);
assign w2131 = w116 & w24621;
assign w2132 = ~w2130 & ~w2131;
assign w2133 = a[23] & ~w2129;
assign w2134 = (~w2133 & w2132) | (~w2133 & w24764) | (w2132 & w24764);
assign w2135 = w2124 & w2134;
assign w2136 = ~w2124 & ~w2134;
assign w2137 = ~w2135 & ~w2136;
assign w2138 = (~w1965 & ~w1966) | (~w1965 & w24622) | (~w1966 & w24622);
assign w2139 = ~w2137 & w2138;
assign w2140 = w2137 & ~w2138;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = b[6] & ~w1272;
assign w2143 = b[7] & w1154;
assign w2144 = b[8] & w1156;
assign w2145 = w270 & w1150;
assign w2146 = ~w2142 & ~w2143;
assign w2147 = ~w2144 & w2146;
assign w2148 = ~w2145 & w2147;
assign w2149 = a[20] & ~w2148;
assign w2150 = ~a[20] & w2148;
assign w2151 = ~w2149 & ~w2150;
assign w2152 = ~w2141 & ~w2151;
assign w2153 = w2141 & w2151;
assign w2154 = ~w2152 & ~w2153;
assign w2155 = (~w1982 & ~w1984) | (~w1982 & w24917) | (~w1984 & w24917);
assign w2156 = w2154 & ~w2155;
assign w2157 = ~w2154 & w2155;
assign w2158 = ~w2156 & ~w2157;
assign w2159 = b[10] & w838;
assign w2160 = b[11] & w834;
assign w2161 = b[9] & ~w934;
assign w2162 = w469 & w832;
assign w2163 = ~w2159 & ~w2160;
assign w2164 = ~w2161 & w2163;
assign w2165 = ~w2162 & w2164;
assign w2166 = a[17] & ~w2165;
assign w2167 = ~a[17] & w2165;
assign w2168 = ~w2166 & ~w2167;
assign w2169 = ~w2158 & ~w2168;
assign w2170 = w2158 & w2168;
assign w2171 = ~w2169 & ~w2170;
assign w2172 = w2108 & ~w2171;
assign w2173 = ~w2108 & w2171;
assign w2174 = ~w2172 & ~w2173;
assign w2175 = w2107 & w2174;
assign w2176 = ~w2107 & ~w2174;
assign w2177 = ~w2175 & ~w2176;
assign w2178 = (~w2015 & ~w2018) | (~w2015 & w24918) | (~w2018 & w24918);
assign w2179 = w2177 & w2178;
assign w2180 = ~w2177 & ~w2178;
assign w2181 = ~w2179 & ~w2180;
assign w2182 = w2097 & w2181;
assign w2183 = ~w2097 & ~w2181;
assign w2184 = ~w2182 & ~w2183;
assign w2185 = w2087 & w2184;
assign w2186 = ~w2087 & ~w2184;
assign w2187 = ~w2185 & ~w2186;
assign w2188 = w2086 & ~w2187;
assign w2189 = ~w2086 & w2187;
assign w2190 = ~w2188 & ~w2189;
assign w2191 = (~w2040 & ~w2042) | (~w2040 & w24765) | (~w2042 & w24765);
assign w2192 = ~w2190 & ~w2191;
assign w2193 = w2190 & w2191;
assign w2194 = ~w2192 & ~w2193;
assign w2195 = b[21] & w103;
assign w2196 = b[22] & w61;
assign w2197 = b[23] & w68;
assign w2198 = w66 & w1755;
assign w2199 = ~w2196 & ~w2197;
assign w2200 = ~w2195 & w2199;
assign w2201 = ~w2198 & w2200;
assign w2202 = a[5] & ~w2201;
assign w2203 = ~a[5] & w2201;
assign w2204 = ~w2202 & ~w2203;
assign w2205 = w2194 & w2204;
assign w2206 = ~w2194 & ~w2204;
assign w2207 = ~w2205 & ~w2206;
assign w2208 = w2076 & w2207;
assign w2209 = ~w2076 & ~w2207;
assign w2210 = ~w2208 & ~w2209;
assign w2211 = b[26] & w11;
assign w2212 = b[25] & w9;
assign w2213 = ~b[25] & ~b[26];
assign w2214 = b[25] & b[26];
assign w2215 = ~w2213 & ~w2214;
assign w2216 = ~w2056 & ~w2059;
assign w2217 = ~w2215 & w2216;
assign w2218 = w2215 & ~w2216;
assign w2219 = ~w2217 & ~w2218;
assign w2220 = w5 & w2219;
assign w2221 = ~w2211 & ~w2212;
assign w2222 = ~w2220 & w2221;
assign w2223 = b[24] & w24;
assign w2224 = a[2] & ~w2223;
assign w2225 = w2222 & ~w2224;
assign w2226 = a[2] & ~w2222;
assign w2227 = ~w2225 & ~w2226;
assign w2228 = ~w2210 & w2227;
assign w2229 = w2210 & ~w2227;
assign w2230 = ~w2228 & ~w2229;
assign w2231 = (~w2070 & w1911) | (~w2070 & w24360) | (w1911 & w24360);
assign w2232 = w2230 & ~w2231;
assign w2233 = ~w2230 & w2231;
assign w2234 = ~w2232 & ~w2233;
assign w2235 = ~w2228 & ~w2232;
assign w2236 = b[22] & w103;
assign w2237 = b[24] & w68;
assign w2238 = b[23] & w61;
assign w2239 = w66 & w1895;
assign w2240 = ~w2237 & ~w2238;
assign w2241 = ~w2236 & w2240;
assign w2242 = ~w2239 & w2241;
assign w2243 = a[5] & ~w2242;
assign w2244 = ~a[5] & w2242;
assign w2245 = ~w2243 & ~w2244;
assign w2246 = b[18] & w360;
assign w2247 = b[17] & w358;
assign w2248 = b[16] & ~w419;
assign w2249 = w354 & ~w1108;
assign w2250 = ~w2246 & ~w2247;
assign w2251 = ~w2248 & w2250;
assign w2252 = ~w2249 & w2251;
assign w2253 = a[11] & ~w2252;
assign w2254 = ~a[11] & w2252;
assign w2255 = ~w2253 & ~w2254;
assign w2256 = ~w2153 & ~w2156;
assign w2257 = w2110 & w2121;
assign w2258 = ~a[26] & ~b[0];
assign w2259 = ~a[27] & b[0];
assign w2260 = ~w2258 & ~w2259;
assign w2261 = b[1] & ~w2114;
assign w2262 = b[2] & w1955;
assign w2263 = b[3] & w1957;
assign w2264 = ~w2261 & ~w2262;
assign w2265 = ~w2263 & w2264;
assign w2266 = w2265 & w24623;
assign w2267 = (~w2260 & ~w2265) | (~w2260 & w24624) | (~w2265 & w24624);
assign w2268 = ~w2266 & ~w2267;
assign w2269 = w2257 & w2268;
assign w2270 = ~w2257 & ~w2268;
assign w2271 = ~w2269 & ~w2270;
assign w2272 = b[6] & w1519;
assign w2273 = b[5] & w1517;
assign w2274 = b[4] & ~w1676;
assign w2275 = w157 & w1513;
assign w2276 = ~w2272 & ~w2273;
assign w2277 = ~w2274 & w2276;
assign w2278 = ~w2275 & w2277;
assign w2279 = a[23] & ~w2278;
assign w2280 = ~a[23] & w2278;
assign w2281 = ~w2279 & ~w2280;
assign w2282 = ~w2271 & w2281;
assign w2283 = w2271 & ~w2281;
assign w2284 = ~w2282 & ~w2283;
assign w2285 = (~w2135 & w2138) | (~w2135 & w24766) | (w2138 & w24766);
assign w2286 = w2284 & ~w2285;
assign w2287 = ~w2284 & w2285;
assign w2288 = ~w2286 & ~w2287;
assign w2289 = b[7] & ~w1272;
assign w2290 = b[8] & w1154;
assign w2291 = b[9] & w1156;
assign w2292 = w322 & w1150;
assign w2293 = ~w2289 & ~w2290;
assign w2294 = ~w2291 & w2293;
assign w2295 = ~w2292 & w2294;
assign w2296 = a[20] & ~w2295;
assign w2297 = ~a[20] & w2295;
assign w2298 = ~w2296 & ~w2297;
assign w2299 = w2288 & w2298;
assign w2300 = ~w2288 & ~w2298;
assign w2301 = ~w2299 & ~w2300;
assign w2302 = w2256 & w2301;
assign w2303 = ~w2256 & ~w2301;
assign w2304 = ~w2302 & ~w2303;
assign w2305 = b[12] & w834;
assign w2306 = b[10] & ~w934;
assign w2307 = b[11] & w838;
assign w2308 = w536 & w832;
assign w2309 = ~w2305 & ~w2306;
assign w2310 = ~w2307 & w2309;
assign w2311 = ~w2308 & w2310;
assign w2312 = a[17] & ~w2311;
assign w2313 = ~a[17] & w2311;
assign w2314 = ~w2312 & ~w2313;
assign w2315 = w2304 & ~w2314;
assign w2316 = ~w2304 & w2314;
assign w2317 = ~w2315 & ~w2316;
assign w2318 = (~w2170 & w2108) | (~w2170 & w24919) | (w2108 & w24919);
assign w2319 = w2317 & ~w2318;
assign w2320 = ~w2317 & w2318;
assign w2321 = ~w2319 & ~w2320;
assign w2322 = b[14] & w573;
assign w2323 = b[15] & w575;
assign w2324 = b[13] & ~w649;
assign w2325 = w569 & ~w799;
assign w2326 = ~w2322 & ~w2323;
assign w2327 = ~w2324 & w2326;
assign w2328 = ~w2325 & w2327;
assign w2329 = a[14] & ~w2328;
assign w2330 = ~a[14] & w2328;
assign w2331 = ~w2329 & ~w2330;
assign w2332 = w2321 & w2331;
assign w2333 = ~w2321 & ~w2331;
assign w2334 = ~w2332 & ~w2333;
assign w2335 = (~w2175 & ~w2178) | (~w2175 & w24361) | (~w2178 & w24361);
assign w2336 = w2334 & w2335;
assign w2337 = ~w2334 & ~w2335;
assign w2338 = ~w2336 & ~w2337;
assign w2339 = w2255 & ~w2338;
assign w2340 = ~w2255 & w2338;
assign w2341 = ~w2339 & ~w2340;
assign w2342 = (~w2183 & ~w2087) | (~w2183 & w24920) | (~w2087 & w24920);
assign w2343 = ~w2341 & ~w2342;
assign w2344 = w2341 & w2342;
assign w2345 = ~w2343 & ~w2344;
assign w2346 = b[19] & ~w237;
assign w2347 = b[21] & w185;
assign w2348 = b[20] & w183;
assign w2349 = w179 & w1467;
assign w2350 = ~w2346 & ~w2347;
assign w2351 = ~w2348 & w2350;
assign w2352 = ~w2349 & w2351;
assign w2353 = a[8] & ~w2352;
assign w2354 = ~a[8] & w2352;
assign w2355 = ~w2353 & ~w2354;
assign w2356 = ~w2345 & ~w2355;
assign w2357 = w2345 & w2355;
assign w2358 = ~w2356 & ~w2357;
assign w2359 = ~w2188 & ~w2193;
assign w2360 = w2358 & w2359;
assign w2361 = ~w2358 & ~w2359;
assign w2362 = ~w2360 & ~w2361;
assign w2363 = w2245 & ~w2362;
assign w2364 = ~w2245 & w2362;
assign w2365 = ~w2363 & ~w2364;
assign w2366 = (~w2206 & ~w2076) | (~w2206 & w24767) | (~w2076 & w24767);
assign w2367 = ~w2365 & ~w2366;
assign w2368 = w2365 & w2366;
assign w2369 = ~w2367 & ~w2368;
assign w2370 = b[27] & w11;
assign w2371 = b[26] & w9;
assign w2372 = ~w2214 & ~w2218;
assign w2373 = ~b[26] & ~b[27];
assign w2374 = b[26] & b[27];
assign w2375 = ~w2373 & ~w2374;
assign w2376 = w2372 & ~w2375;
assign w2377 = ~w2372 & w2375;
assign w2378 = ~w2376 & ~w2377;
assign w2379 = w5 & w2378;
assign w2380 = ~w2370 & ~w2371;
assign w2381 = ~w2379 & w2380;
assign w2382 = b[25] & w24;
assign w2383 = a[2] & ~w2382;
assign w2384 = w2381 & ~w2383;
assign w2385 = a[2] & ~w2381;
assign w2386 = ~w2384 & ~w2385;
assign w2387 = ~w2369 & ~w2386;
assign w2388 = w2369 & w2386;
assign w2389 = ~w2387 & ~w2388;
assign w2390 = w2235 & ~w2389;
assign w2391 = ~w2235 & w2389;
assign w2392 = ~w2390 & ~w2391;
assign w2393 = b[20] & ~w237;
assign w2394 = b[22] & w185;
assign w2395 = b[21] & w183;
assign w2396 = w179 & w1615;
assign w2397 = ~w2393 & ~w2394;
assign w2398 = ~w2395 & w2397;
assign w2399 = ~w2396 & w2398;
assign w2400 = a[8] & ~w2399;
assign w2401 = ~a[8] & w2399;
assign w2402 = ~w2400 & ~w2401;
assign w2403 = b[14] & ~w649;
assign w2404 = b[16] & w575;
assign w2405 = b[15] & w573;
assign w2406 = w569 & w905;
assign w2407 = ~w2403 & ~w2404;
assign w2408 = ~w2405 & w2407;
assign w2409 = ~w2406 & w2408;
assign w2410 = a[14] & ~w2409;
assign w2411 = ~a[14] & w2409;
assign w2412 = ~w2410 & ~w2411;
assign w2413 = ~w2282 & ~w2286;
assign w2414 = b[3] & w1955;
assign w2415 = b[4] & w1957;
assign w2416 = b[2] & ~w2114;
assign w2417 = w84 & w1951;
assign w2418 = ~w2414 & ~w2415;
assign w2419 = ~w2416 & w2418;
assign w2420 = ~w2417 & w2419;
assign w2421 = a[26] & ~w2420;
assign w2422 = ~a[26] & w2420;
assign w2423 = ~w2421 & ~w2422;
assign w2424 = a[26] & a[27];
assign w2425 = ~a[26] & ~a[27];
assign w2426 = ~w2424 & ~w2425;
assign w2427 = b[0] & w2426;
assign w2428 = a[29] & w2427;
assign w2429 = a[28] & ~a[29];
assign w2430 = ~a[28] & a[29];
assign w2431 = ~w2429 & ~w2430;
assign w2432 = w2426 & ~w2431;
assign w2433 = ~w8 & w2432;
assign w2434 = ~a[28] & ~w2424;
assign w2435 = a[28] & ~w2425;
assign w2436 = ~w2434 & ~w2435;
assign w2437 = b[0] & w2436;
assign w2438 = w2426 & w2431;
assign w2439 = b[1] & w2438;
assign w2440 = ~w2433 & ~w2437;
assign w2441 = ~w2439 & w2440;
assign w2442 = ~w2428 & w2441;
assign w2443 = w2428 & ~w2441;
assign w2444 = ~w2442 & ~w2443;
assign w2445 = ~w2423 & ~w2444;
assign w2446 = w2423 & w2444;
assign w2447 = ~w2445 & ~w2446;
assign w2448 = ~w2266 & ~w2427;
assign w2449 = ~w2270 & ~w2448;
assign w2450 = w2447 & w2449;
assign w2451 = ~w2447 & ~w2449;
assign w2452 = ~w2450 & ~w2451;
assign w2453 = b[7] & w1519;
assign w2454 = b[6] & w1517;
assign w2455 = b[5] & ~w1676;
assign w2456 = w216 & w1513;
assign w2457 = ~w2453 & ~w2454;
assign w2458 = ~w2455 & w2457;
assign w2459 = ~w2456 & w2458;
assign w2460 = a[23] & ~w2459;
assign w2461 = ~a[23] & w2459;
assign w2462 = ~w2460 & ~w2461;
assign w2463 = w2452 & w2462;
assign w2464 = ~w2452 & ~w2462;
assign w2465 = ~w2463 & ~w2464;
assign w2466 = w2413 & w2465;
assign w2467 = ~w2413 & ~w2465;
assign w2468 = ~w2466 & ~w2467;
assign w2469 = b[10] & w1156;
assign w2470 = b[8] & ~w1272;
assign w2471 = b[9] & w1154;
assign w2472 = w397 & w1150;
assign w2473 = ~w2469 & ~w2470;
assign w2474 = ~w2471 & w2473;
assign w2475 = ~w2472 & w2474;
assign w2476 = a[20] & ~w2475;
assign w2477 = ~a[20] & w2475;
assign w2478 = ~w2476 & ~w2477;
assign w2479 = ~w2468 & w2478;
assign w2480 = w2468 & ~w2478;
assign w2481 = ~w2479 & ~w2480;
assign w2482 = (~w2300 & ~w2256) | (~w2300 & w25103) | (~w2256 & w25103);
assign w2483 = ~w2481 & ~w2482;
assign w2484 = w2481 & w2482;
assign w2485 = ~w2483 & ~w2484;
assign w2486 = b[11] & ~w934;
assign w2487 = b[12] & w838;
assign w2488 = b[13] & w834;
assign w2489 = w628 & w832;
assign w2490 = ~w2486 & ~w2487;
assign w2491 = ~w2488 & w2490;
assign w2492 = ~w2489 & w2491;
assign w2493 = a[17] & ~w2492;
assign w2494 = ~a[17] & w2492;
assign w2495 = ~w2493 & ~w2494;
assign w2496 = w2485 & w2495;
assign w2497 = ~w2485 & ~w2495;
assign w2498 = ~w2496 & ~w2497;
assign w2499 = ~w2316 & ~w2319;
assign w2500 = w2498 & w2499;
assign w2501 = ~w2498 & ~w2499;
assign w2502 = ~w2500 & ~w2501;
assign w2503 = w2412 & ~w2502;
assign w2504 = ~w2412 & w2502;
assign w2505 = ~w2503 & ~w2504;
assign w2506 = (~w2333 & ~w2335) | (~w2333 & w24921) | (~w2335 & w24921);
assign w2507 = ~w2505 & ~w2506;
assign w2508 = w2505 & w2506;
assign w2509 = ~w2507 & ~w2508;
assign w2510 = b[18] & w358;
assign w2511 = b[17] & ~w419;
assign w2512 = b[19] & w360;
assign w2513 = w354 & ~w1231;
assign w2514 = ~w2510 & ~w2511;
assign w2515 = ~w2512 & w2514;
assign w2516 = ~w2513 & w2515;
assign w2517 = a[11] & ~w2516;
assign w2518 = ~a[11] & w2516;
assign w2519 = ~w2517 & ~w2518;
assign w2520 = w2509 & w2519;
assign w2521 = ~w2509 & ~w2519;
assign w2522 = ~w2520 & ~w2521;
assign w2523 = (~w2339 & ~w2342) | (~w2339 & w24362) | (~w2342 & w24362);
assign w2524 = w2522 & w2523;
assign w2525 = ~w2522 & ~w2523;
assign w2526 = ~w2524 & ~w2525;
assign w2527 = ~w2402 & w2526;
assign w2528 = w2402 & ~w2526;
assign w2529 = ~w2527 & ~w2528;
assign w2530 = (~w2356 & ~w2359) | (~w2356 & w24922) | (~w2359 & w24922);
assign w2531 = w2529 & w2530;
assign w2532 = ~w2529 & ~w2530;
assign w2533 = ~w2531 & ~w2532;
assign w2534 = b[23] & w103;
assign w2535 = b[25] & w68;
assign w2536 = b[24] & w61;
assign w2537 = w66 & w2061;
assign w2538 = ~w2535 & ~w2536;
assign w2539 = ~w2534 & w2538;
assign w2540 = ~w2537 & w2539;
assign w2541 = a[5] & ~w2540;
assign w2542 = ~a[5] & w2540;
assign w2543 = ~w2541 & ~w2542;
assign w2544 = w2533 & w2543;
assign w2545 = ~w2533 & ~w2543;
assign w2546 = ~w2544 & ~w2545;
assign w2547 = ~w2363 & ~w2368;
assign w2548 = w2546 & w2547;
assign w2549 = ~w2546 & ~w2547;
assign w2550 = ~w2548 & ~w2549;
assign w2551 = b[28] & w11;
assign w2552 = b[27] & w9;
assign w2553 = ~b[27] & ~b[28];
assign w2554 = b[27] & b[28];
assign w2555 = ~w2553 & ~w2554;
assign w2556 = ~w2374 & ~w2377;
assign w2557 = w2555 & ~w2556;
assign w2558 = ~w2555 & w2556;
assign w2559 = ~w2557 & ~w2558;
assign w2560 = w5 & w2559;
assign w2561 = ~w2551 & ~w2552;
assign w2562 = ~w2560 & w2561;
assign w2563 = b[26] & w24;
assign w2564 = a[2] & ~w2563;
assign w2565 = w2562 & ~w2564;
assign w2566 = a[2] & ~w2562;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = w2550 & ~w2567;
assign w2569 = ~w2550 & w2567;
assign w2570 = ~w2568 & ~w2569;
assign w2571 = (~w2388 & w2235) | (~w2388 & w24768) | (w2235 & w24768);
assign w2572 = w2570 & ~w2571;
assign w2573 = ~w2570 & w2571;
assign w2574 = ~w2572 & ~w2573;
assign w2575 = ~w2569 & ~w2572;
assign w2576 = b[24] & w103;
assign w2577 = b[26] & w68;
assign w2578 = b[25] & w61;
assign w2579 = w66 & w2219;
assign w2580 = ~w2577 & ~w2578;
assign w2581 = ~w2576 & w2580;
assign w2582 = ~w2579 & w2581;
assign w2583 = a[5] & ~w2582;
assign w2584 = ~a[5] & w2582;
assign w2585 = ~w2583 & ~w2584;
assign w2586 = (~w2528 & ~w2530) | (~w2528 & w24363) | (~w2530 & w24363);
assign w2587 = b[23] & w185;
assign w2588 = b[21] & ~w237;
assign w2589 = b[22] & w183;
assign w2590 = w179 & w1755;
assign w2591 = ~w2587 & ~w2588;
assign w2592 = ~w2589 & w2591;
assign w2593 = ~w2590 & w2592;
assign w2594 = a[8] & ~w2593;
assign w2595 = ~a[8] & w2593;
assign w2596 = ~w2594 & ~w2595;
assign w2597 = b[19] & w358;
assign w2598 = b[18] & ~w419;
assign w2599 = b[20] & w360;
assign w2600 = w354 & w1347;
assign w2601 = ~w2597 & ~w2598;
assign w2602 = ~w2599 & w2601;
assign w2603 = ~w2600 & w2602;
assign w2604 = a[11] & ~w2603;
assign w2605 = ~a[11] & w2603;
assign w2606 = ~w2604 & ~w2605;
assign w2607 = b[14] & w834;
assign w2608 = b[13] & w838;
assign w2609 = b[12] & ~w934;
assign w2610 = w714 & w832;
assign w2611 = ~w2607 & ~w2608;
assign w2612 = ~w2609 & w2611;
assign w2613 = ~w2610 & w2612;
assign w2614 = a[17] & ~w2613;
assign w2615 = ~a[17] & w2613;
assign w2616 = ~w2614 & ~w2615;
assign w2617 = (a[29] & ~w2426) | (a[29] & w24923) | (~w2426 & w24923);
assign w2618 = w2440 & w24769;
assign w2619 = a[29] & ~w2618;
assign w2620 = w2424 & w2429;
assign w2621 = w2425 & w2430;
assign w2622 = ~w2620 & ~w2621;
assign w2623 = b[0] & ~w2622;
assign w2624 = w22 & w2432;
assign w2625 = b[1] & w2436;
assign w2626 = b[2] & w2438;
assign w2627 = ~w2623 & ~w2624;
assign w2628 = ~w2625 & ~w2626;
assign w2629 = w2627 & w2628;
assign w2630 = ~w2619 & w2629;
assign w2631 = w2619 & ~w2629;
assign w2632 = ~w2630 & ~w2631;
assign w2633 = b[4] & w1955;
assign w2634 = b[3] & ~w2114;
assign w2635 = b[5] & w1957;
assign w2636 = ~w2633 & ~w2634;
assign w2637 = ~w2635 & w2636;
assign w2638 = (~a[26] & ~w116) | (~a[26] & w24625) | (~w116 & w24625);
assign w2639 = w116 & w24626;
assign w2640 = ~w2638 & ~w2639;
assign w2641 = (a[26] & ~w2636) | (a[26] & w24924) | (~w2636 & w24924);
assign w2642 = (~w2641 & w2640) | (~w2641 & w24770) | (w2640 & w24770);
assign w2643 = w2632 & w2642;
assign w2644 = ~w2632 & ~w2642;
assign w2645 = ~w2643 & ~w2644;
assign w2646 = (~w2446 & ~w2447) | (~w2446 & w24627) | (~w2447 & w24627);
assign w2647 = ~w2645 & w2646;
assign w2648 = w2645 & ~w2646;
assign w2649 = ~w2647 & ~w2648;
assign w2650 = b[8] & w1519;
assign w2651 = b[6] & ~w1676;
assign w2652 = b[7] & w1517;
assign w2653 = w270 & w1513;
assign w2654 = ~w2650 & ~w2651;
assign w2655 = ~w2652 & w2654;
assign w2656 = ~w2653 & w2655;
assign w2657 = a[23] & ~w2656;
assign w2658 = ~a[23] & w2656;
assign w2659 = ~w2657 & ~w2658;
assign w2660 = ~w2649 & ~w2659;
assign w2661 = w2649 & w2659;
assign w2662 = ~w2660 & ~w2661;
assign w2663 = (~w2464 & ~w2413) | (~w2464 & w24628) | (~w2413 & w24628);
assign w2664 = w2662 & w2663;
assign w2665 = ~w2662 & ~w2663;
assign w2666 = ~w2664 & ~w2665;
assign w2667 = b[9] & ~w1272;
assign w2668 = b[10] & w1154;
assign w2669 = b[11] & w1156;
assign w2670 = w469 & w1150;
assign w2671 = ~w2667 & ~w2668;
assign w2672 = ~w2669 & w2671;
assign w2673 = ~w2670 & w2672;
assign w2674 = a[20] & ~w2673;
assign w2675 = ~a[20] & w2673;
assign w2676 = ~w2674 & ~w2675;
assign w2677 = ~w2666 & ~w2676;
assign w2678 = w2666 & w2676;
assign w2679 = ~w2677 & ~w2678;
assign w2680 = ~w2679 & w25104;
assign w2681 = (w2679 & w2484) | (w2679 & w24629) | (w2484 & w24629);
assign w2682 = ~w2681 & w25105;
assign w2683 = (~w2616 & w2681) | (~w2616 & w25106) | (w2681 & w25106);
assign w2684 = ~w2682 & ~w2683;
assign w2685 = ~w2497 & ~w2500;
assign w2686 = ~w2684 & ~w2685;
assign w2687 = w2684 & w2685;
assign w2688 = ~w2686 & ~w2687;
assign w2689 = b[15] & ~w649;
assign w2690 = b[16] & w573;
assign w2691 = b[17] & w575;
assign w2692 = w569 & w1008;
assign w2693 = ~w2689 & ~w2690;
assign w2694 = ~w2691 & w2693;
assign w2695 = ~w2692 & w2694;
assign w2696 = a[14] & ~w2695;
assign w2697 = ~a[14] & w2695;
assign w2698 = ~w2696 & ~w2697;
assign w2699 = w2688 & w2698;
assign w2700 = ~w2688 & ~w2698;
assign w2701 = ~w2699 & ~w2700;
assign w2702 = ~w2503 & ~w2508;
assign w2703 = w2701 & w2702;
assign w2704 = ~w2701 & ~w2702;
assign w2705 = ~w2703 & ~w2704;
assign w2706 = w2606 & ~w2705;
assign w2707 = ~w2606 & w2705;
assign w2708 = ~w2706 & ~w2707;
assign w2709 = (~w2521 & ~w2523) | (~w2521 & w24925) | (~w2523 & w24925);
assign w2710 = w2708 & w2709;
assign w2711 = ~w2708 & ~w2709;
assign w2712 = ~w2710 & ~w2711;
assign w2713 = w2596 & w2712;
assign w2714 = ~w2596 & ~w2712;
assign w2715 = ~w2713 & ~w2714;
assign w2716 = w2586 & w2715;
assign w2717 = ~w2586 & ~w2715;
assign w2718 = ~w2716 & ~w2717;
assign w2719 = ~w2585 & w2718;
assign w2720 = w2585 & ~w2718;
assign w2721 = ~w2719 & ~w2720;
assign w2722 = (~w2545 & ~w2547) | (~w2545 & w24926) | (~w2547 & w24926);
assign w2723 = w2721 & w2722;
assign w2724 = ~w2721 & ~w2722;
assign w2725 = ~w2723 & ~w2724;
assign w2726 = b[29] & w11;
assign w2727 = b[28] & w9;
assign w2728 = ~b[28] & ~b[29];
assign w2729 = b[28] & b[29];
assign w2730 = ~w2728 & ~w2729;
assign w2731 = (~w2554 & w2556) | (~w2554 & w24630) | (w2556 & w24630);
assign w2732 = ~w2730 & w2731;
assign w2733 = w2730 & ~w2731;
assign w2734 = ~w2732 & ~w2733;
assign w2735 = w5 & w2734;
assign w2736 = ~w2726 & ~w2727;
assign w2737 = ~w2735 & w2736;
assign w2738 = b[27] & w24;
assign w2739 = a[2] & ~w2738;
assign w2740 = w2737 & ~w2739;
assign w2741 = a[2] & ~w2737;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = w2725 & w2742;
assign w2744 = ~w2725 & ~w2742;
assign w2745 = ~w2743 & ~w2744;
assign w2746 = w2575 & ~w2745;
assign w2747 = ~w2575 & w2745;
assign w2748 = ~w2746 & ~w2747;
assign w2749 = b[22] & ~w237;
assign w2750 = b[23] & w183;
assign w2751 = b[24] & w185;
assign w2752 = w179 & w1895;
assign w2753 = ~w2749 & ~w2750;
assign w2754 = ~w2751 & w2753;
assign w2755 = ~w2752 & w2754;
assign w2756 = a[8] & ~w2755;
assign w2757 = ~a[8] & w2755;
assign w2758 = ~w2756 & ~w2757;
assign w2759 = ~w2706 & ~w2710;
assign w2760 = b[16] & ~w649;
assign w2761 = b[17] & w573;
assign w2762 = b[18] & w575;
assign w2763 = w569 & ~w1108;
assign w2764 = ~w2760 & ~w2761;
assign w2765 = ~w2762 & w2764;
assign w2766 = ~w2763 & w2765;
assign w2767 = a[14] & ~w2766;
assign w2768 = ~a[14] & w2766;
assign w2769 = ~w2767 & ~w2768;
assign w2770 = (~w2661 & ~w2663) | (~w2661 & w24771) | (~w2663 & w24771);
assign w2771 = b[5] & w1955;
assign w2772 = b[4] & ~w2114;
assign w2773 = b[6] & w1957;
assign w2774 = w157 & w1951;
assign w2775 = ~w2771 & ~w2772;
assign w2776 = ~w2773 & w2775;
assign w2777 = (a[26] & w2774) | (a[26] & w24927) | (w2774 & w24927);
assign w2778 = ~w2774 & w24928;
assign w2779 = ~w2777 & ~w2778;
assign w2780 = w2618 & w2629;
assign w2781 = ~a[29] & ~b[0];
assign w2782 = ~a[30] & b[0];
assign w2783 = ~w2781 & ~w2782;
assign w2784 = b[3] & w2438;
assign w2785 = b[2] & w2436;
assign w2786 = b[1] & ~w2622;
assign w2787 = w46 & w2432;
assign w2788 = ~w2784 & ~w2785;
assign w2789 = ~w2786 & w2788;
assign w2790 = w2789 & w24631;
assign w2791 = (~w2783 & ~w2789) | (~w2783 & w24772) | (~w2789 & w24772);
assign w2792 = ~w2790 & ~w2791;
assign w2793 = w2780 & ~w2792;
assign w2794 = ~w2780 & w2792;
assign w2795 = ~w2793 & ~w2794;
assign w2796 = w2779 & w2795;
assign w2797 = ~w2779 & ~w2795;
assign w2798 = ~w2796 & ~w2797;
assign w2799 = (~w2643 & w2646) | (~w2643 & w24773) | (w2646 & w24773);
assign w2800 = w2798 & ~w2799;
assign w2801 = ~w2798 & w2799;
assign w2802 = ~w2800 & ~w2801;
assign w2803 = b[9] & w1519;
assign w2804 = b[8] & w1517;
assign w2805 = b[7] & ~w1676;
assign w2806 = w322 & w1513;
assign w2807 = ~w2803 & ~w2804;
assign w2808 = ~w2805 & w2807;
assign w2809 = ~w2806 & w2808;
assign w2810 = a[23] & ~w2809;
assign w2811 = ~a[23] & w2809;
assign w2812 = ~w2810 & ~w2811;
assign w2813 = w2802 & w2812;
assign w2814 = ~w2802 & ~w2812;
assign w2815 = ~w2813 & ~w2814;
assign w2816 = w2770 & ~w2815;
assign w2817 = ~w2770 & w2815;
assign w2818 = ~w2816 & ~w2817;
assign w2819 = b[10] & ~w1272;
assign w2820 = b[12] & w1156;
assign w2821 = b[11] & w1154;
assign w2822 = w536 & w1150;
assign w2823 = ~w2819 & ~w2820;
assign w2824 = ~w2821 & w2823;
assign w2825 = ~w2822 & w2824;
assign w2826 = a[20] & ~w2825;
assign w2827 = ~a[20] & w2825;
assign w2828 = ~w2826 & ~w2827;
assign w2829 = ~w2818 & ~w2828;
assign w2830 = w2818 & w2828;
assign w2831 = ~w2829 & ~w2830;
assign w2832 = ~w2678 & ~w2681;
assign w2833 = w2831 & ~w2832;
assign w2834 = ~w2831 & w2832;
assign w2835 = ~w2833 & ~w2834;
assign w2836 = b[14] & w838;
assign w2837 = b[15] & w834;
assign w2838 = b[13] & ~w934;
assign w2839 = ~w799 & w832;
assign w2840 = ~w2836 & ~w2837;
assign w2841 = ~w2838 & w2840;
assign w2842 = ~w2839 & w2841;
assign w2843 = a[17] & ~w2842;
assign w2844 = ~a[17] & w2842;
assign w2845 = ~w2843 & ~w2844;
assign w2846 = w2835 & w2845;
assign w2847 = ~w2835 & ~w2845;
assign w2848 = ~w2846 & ~w2847;
assign w2849 = (~w2682 & ~w2685) | (~w2682 & w24632) | (~w2685 & w24632);
assign w2850 = w2848 & w2849;
assign w2851 = ~w2848 & ~w2849;
assign w2852 = ~w2850 & ~w2851;
assign w2853 = w2769 & ~w2852;
assign w2854 = ~w2769 & w2852;
assign w2855 = ~w2853 & ~w2854;
assign w2856 = ~w2700 & ~w2703;
assign w2857 = ~w2855 & ~w2856;
assign w2858 = w2855 & w2856;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = b[19] & ~w419;
assign w2861 = b[20] & w358;
assign w2862 = b[21] & w360;
assign w2863 = w354 & w1467;
assign w2864 = ~w2860 & ~w2861;
assign w2865 = ~w2862 & w2864;
assign w2866 = ~w2863 & w2865;
assign w2867 = a[11] & ~w2866;
assign w2868 = ~a[11] & w2866;
assign w2869 = ~w2867 & ~w2868;
assign w2870 = w2859 & w2869;
assign w2871 = ~w2859 & ~w2869;
assign w2872 = ~w2870 & ~w2871;
assign w2873 = w2759 & w2872;
assign w2874 = ~w2759 & ~w2872;
assign w2875 = ~w2873 & ~w2874;
assign w2876 = w2758 & ~w2875;
assign w2877 = ~w2758 & w2875;
assign w2878 = ~w2876 & ~w2877;
assign w2879 = (~w2714 & ~w2586) | (~w2714 & w24929) | (~w2586 & w24929);
assign w2880 = ~w2878 & ~w2879;
assign w2881 = w2878 & w2879;
assign w2882 = ~w2880 & ~w2881;
assign w2883 = b[25] & w103;
assign w2884 = b[26] & w61;
assign w2885 = b[27] & w68;
assign w2886 = w66 & w2378;
assign w2887 = ~w2884 & ~w2885;
assign w2888 = ~w2883 & w2887;
assign w2889 = ~w2886 & w2888;
assign w2890 = a[5] & ~w2889;
assign w2891 = ~a[5] & w2889;
assign w2892 = ~w2890 & ~w2891;
assign w2893 = w2882 & w2892;
assign w2894 = ~w2882 & ~w2892;
assign w2895 = ~w2893 & ~w2894;
assign w2896 = (~w2720 & ~w2722) | (~w2720 & w24364) | (~w2722 & w24364);
assign w2897 = w2895 & w2896;
assign w2898 = ~w2895 & ~w2896;
assign w2899 = ~w2897 & ~w2898;
assign w2900 = b[30] & w11;
assign w2901 = b[29] & w9;
assign w2902 = ~w2729 & ~w2733;
assign w2903 = ~b[29] & ~b[30];
assign w2904 = b[29] & b[30];
assign w2905 = ~w2903 & ~w2904;
assign w2906 = ~w2902 & ~w2905;
assign w2907 = w2902 & w2905;
assign w2908 = ~w2906 & ~w2907;
assign w2909 = w5 & ~w2908;
assign w2910 = ~w2900 & ~w2901;
assign w2911 = ~w2909 & w2910;
assign w2912 = b[28] & w24;
assign w2913 = a[2] & ~w2912;
assign w2914 = w2911 & ~w2913;
assign w2915 = a[2] & ~w2911;
assign w2916 = ~w2914 & ~w2915;
assign w2917 = ~w2899 & w2916;
assign w2918 = w2899 & ~w2916;
assign w2919 = ~w2917 & ~w2918;
assign w2920 = (~w2743 & w2575) | (~w2743 & w24930) | (w2575 & w24930);
assign w2921 = w2919 & ~w2920;
assign w2922 = ~w2919 & w2920;
assign w2923 = ~w2921 & ~w2922;
assign w2924 = b[26] & w103;
assign w2925 = b[28] & w68;
assign w2926 = b[27] & w61;
assign w2927 = w66 & w2559;
assign w2928 = ~w2925 & ~w2926;
assign w2929 = ~w2924 & w2928;
assign w2930 = ~w2927 & w2929;
assign w2931 = a[5] & ~w2930;
assign w2932 = ~a[5] & w2930;
assign w2933 = ~w2931 & ~w2932;
assign w2934 = b[22] & w360;
assign w2935 = b[21] & w358;
assign w2936 = b[20] & ~w419;
assign w2937 = w354 & w1615;
assign w2938 = ~w2934 & ~w2935;
assign w2939 = ~w2936 & w2938;
assign w2940 = ~w2937 & w2939;
assign w2941 = a[11] & ~w2940;
assign w2942 = ~a[11] & w2940;
assign w2943 = ~w2941 & ~w2942;
assign w2944 = b[14] & ~w934;
assign w2945 = b[15] & w838;
assign w2946 = b[16] & w834;
assign w2947 = w832 & w905;
assign w2948 = ~w2944 & ~w2945;
assign w2949 = ~w2946 & w2948;
assign w2950 = ~w2947 & w2949;
assign w2951 = a[17] & ~w2950;
assign w2952 = ~a[17] & w2950;
assign w2953 = ~w2951 & ~w2952;
assign w2954 = (~w2796 & w2799) | (~w2796 & w24633) | (w2799 & w24633);
assign w2955 = b[4] & w2438;
assign w2956 = b[3] & w2436;
assign w2957 = b[2] & ~w2622;
assign w2958 = w84 & w2432;
assign w2959 = ~w2955 & ~w2956;
assign w2960 = ~w2957 & w2959;
assign w2961 = ~w2958 & w2960;
assign w2962 = a[29] & ~w2961;
assign w2963 = ~a[29] & w2961;
assign w2964 = ~w2962 & ~w2963;
assign w2965 = a[29] & ~a[30];
assign w2966 = ~a[29] & a[30];
assign w2967 = ~w2965 & ~w2966;
assign w2968 = b[0] & ~w2967;
assign w2969 = a[32] & w2968;
assign w2970 = a[30] & ~a[31];
assign w2971 = ~a[30] & a[31];
assign w2972 = ~w2970 & ~w2971;
assign w2973 = w2967 & ~w2972;
assign w2974 = b[0] & w2973;
assign w2975 = a[31] & ~a[32];
assign w2976 = ~a[31] & a[32];
assign w2977 = ~w2975 & ~w2976;
assign w2978 = ~w2967 & w2977;
assign w2979 = b[1] & w2978;
assign w2980 = ~w2967 & ~w2977;
assign w2981 = ~w8 & w2980;
assign w2982 = ~w2974 & ~w2979;
assign w2983 = ~w2981 & w2982;
assign w2984 = w2969 & ~w2983;
assign w2985 = ~w2969 & w2983;
assign w2986 = ~w2984 & ~w2985;
assign w2987 = ~w2964 & ~w2986;
assign w2988 = w2964 & w2986;
assign w2989 = ~w2987 & ~w2988;
assign w2990 = (~w2968 & ~w2789) | (~w2968 & w24774) | (~w2789 & w24774);
assign w2991 = w2780 & ~w2990;
assign w2992 = w2789 & w24775;
assign w2993 = (w2789 & w24931) | (w2789 & w24932) | (w24931 & w24932);
assign w2994 = ~w2992 & w2993;
assign w2995 = ~w2991 & ~w2994;
assign w2996 = w2989 & ~w2995;
assign w2997 = ~w2989 & w2995;
assign w2998 = ~w2996 & ~w2997;
assign w2999 = b[7] & w1957;
assign w3000 = b[5] & ~w2114;
assign w3001 = b[6] & w1955;
assign w3002 = w216 & w1951;
assign w3003 = ~w2999 & ~w3000;
assign w3004 = ~w3001 & w3003;
assign w3005 = ~w3002 & w3004;
assign w3006 = a[26] & ~w3005;
assign w3007 = ~a[26] & w3005;
assign w3008 = ~w3006 & ~w3007;
assign w3009 = w2998 & w3008;
assign w3010 = ~w2998 & ~w3008;
assign w3011 = ~w3009 & ~w3010;
assign w3012 = w2954 & ~w3011;
assign w3013 = ~w2954 & w3011;
assign w3014 = ~w3012 & ~w3013;
assign w3015 = b[8] & ~w1676;
assign w3016 = b[9] & w1517;
assign w3017 = b[10] & w1519;
assign w3018 = w397 & w1513;
assign w3019 = ~w3015 & ~w3016;
assign w3020 = ~w3017 & w3019;
assign w3021 = ~w3018 & w3020;
assign w3022 = a[23] & ~w3021;
assign w3023 = ~a[23] & w3021;
assign w3024 = ~w3022 & ~w3023;
assign w3025 = w3014 & w3024;
assign w3026 = ~w3014 & ~w3024;
assign w3027 = ~w3025 & ~w3026;
assign w3028 = (~w2813 & w2770) | (~w2813 & w24933) | (w2770 & w24933);
assign w3029 = ~w3027 & w3028;
assign w3030 = w3027 & ~w3028;
assign w3031 = ~w3029 & ~w3030;
assign w3032 = b[11] & ~w1272;
assign w3033 = b[12] & w1154;
assign w3034 = b[13] & w1156;
assign w3035 = w628 & w1150;
assign w3036 = ~w3032 & ~w3033;
assign w3037 = ~w3034 & w3036;
assign w3038 = ~w3035 & w3037;
assign w3039 = a[20] & ~w3038;
assign w3040 = ~a[20] & w3038;
assign w3041 = ~w3039 & ~w3040;
assign w3042 = ~w3031 & ~w3041;
assign w3043 = w3031 & w3041;
assign w3044 = ~w3042 & ~w3043;
assign w3045 = (~w2830 & w2832) | (~w2830 & w25107) | (w2832 & w25107);
assign w3046 = ~w3044 & w3045;
assign w3047 = w3044 & ~w3045;
assign w3048 = ~w3046 & ~w3047;
assign w3049 = w2953 & w3048;
assign w3050 = ~w2953 & ~w3048;
assign w3051 = ~w3049 & ~w3050;
assign w3052 = (~w2847 & ~w2849) | (~w2847 & w24934) | (~w2849 & w24934);
assign w3053 = ~w3051 & ~w3052;
assign w3054 = w3051 & w3052;
assign w3055 = ~w3053 & ~w3054;
assign w3056 = b[17] & ~w649;
assign w3057 = b[18] & w573;
assign w3058 = b[19] & w575;
assign w3059 = w569 & ~w1231;
assign w3060 = ~w3056 & ~w3057;
assign w3061 = ~w3058 & w3060;
assign w3062 = ~w3059 & w3061;
assign w3063 = a[14] & ~w3062;
assign w3064 = ~a[14] & w3062;
assign w3065 = ~w3063 & ~w3064;
assign w3066 = w3055 & w3065;
assign w3067 = ~w3055 & ~w3065;
assign w3068 = ~w3066 & ~w3067;
assign w3069 = (~w2853 & ~w2856) | (~w2853 & w24635) | (~w2856 & w24635);
assign w3070 = w3068 & w3069;
assign w3071 = ~w3068 & ~w3069;
assign w3072 = ~w3070 & ~w3071;
assign w3073 = w2943 & ~w3072;
assign w3074 = ~w2943 & w3072;
assign w3075 = ~w3073 & ~w3074;
assign w3076 = ~w2871 & ~w2873;
assign w3077 = ~w3075 & ~w3076;
assign w3078 = w3075 & w3076;
assign w3079 = ~w3077 & ~w3078;
assign w3080 = b[23] & ~w237;
assign w3081 = b[25] & w185;
assign w3082 = b[24] & w183;
assign w3083 = w179 & w2061;
assign w3084 = ~w3080 & ~w3081;
assign w3085 = ~w3082 & w3084;
assign w3086 = ~w3083 & w3085;
assign w3087 = a[8] & ~w3086;
assign w3088 = ~a[8] & w3086;
assign w3089 = ~w3087 & ~w3088;
assign w3090 = w3079 & w3089;
assign w3091 = ~w3079 & ~w3089;
assign w3092 = ~w3090 & ~w3091;
assign w3093 = ~w2876 & ~w2881;
assign w3094 = w3092 & w3093;
assign w3095 = ~w3092 & ~w3093;
assign w3096 = ~w3094 & ~w3095;
assign w3097 = w2933 & ~w3096;
assign w3098 = ~w2933 & w3096;
assign w3099 = ~w3097 & ~w3098;
assign w3100 = (~w2894 & ~w2896) | (~w2894 & w24935) | (~w2896 & w24935);
assign w3101 = ~w3099 & ~w3100;
assign w3102 = w3099 & w3100;
assign w3103 = ~w3101 & ~w3102;
assign w3104 = b[31] & w11;
assign w3105 = b[30] & w9;
assign w3106 = ~b[30] & ~b[31];
assign w3107 = b[30] & b[31];
assign w3108 = ~w3106 & ~w3107;
assign w3109 = ~w2903 & ~w2907;
assign w3110 = ~w3108 & w3109;
assign w3111 = w3108 & ~w3109;
assign w3112 = ~w3110 & ~w3111;
assign w3113 = w5 & ~w3112;
assign w3114 = ~w3104 & ~w3105;
assign w3115 = ~w3113 & w3114;
assign w3116 = b[29] & w24;
assign w3117 = a[2] & ~w3116;
assign w3118 = w3115 & ~w3117;
assign w3119 = a[2] & ~w3115;
assign w3120 = ~w3118 & ~w3119;
assign w3121 = w3103 & w3120;
assign w3122 = ~w3103 & ~w3120;
assign w3123 = ~w3121 & ~w3122;
assign w3124 = (~w2917 & w2920) | (~w2917 & w24365) | (w2920 & w24365);
assign w3125 = w3123 & w3124;
assign w3126 = ~w3123 & ~w3124;
assign w3127 = ~w3125 & ~w3126;
assign w3128 = ~w3097 & ~w3102;
assign w3129 = b[25] & w183;
assign w3130 = b[24] & ~w237;
assign w3131 = b[26] & w185;
assign w3132 = w179 & w2219;
assign w3133 = ~w3129 & ~w3130;
assign w3134 = ~w3131 & w3133;
assign w3135 = ~w3132 & w3134;
assign w3136 = a[8] & ~w3135;
assign w3137 = ~a[8] & w3135;
assign w3138 = ~w3136 & ~w3137;
assign w3139 = (~w3073 & ~w3076) | (~w3073 & w24636) | (~w3076 & w24636);
assign w3140 = b[23] & w360;
assign w3141 = b[22] & w358;
assign w3142 = b[21] & ~w419;
assign w3143 = w354 & w1755;
assign w3144 = ~w3140 & ~w3141;
assign w3145 = ~w3142 & w3144;
assign w3146 = ~w3143 & w3145;
assign w3147 = a[11] & ~w3146;
assign w3148 = ~a[11] & w3146;
assign w3149 = ~w3147 & ~w3148;
assign w3150 = b[20] & w575;
assign w3151 = b[18] & ~w649;
assign w3152 = b[19] & w573;
assign w3153 = w569 & w1347;
assign w3154 = ~w3150 & ~w3151;
assign w3155 = ~w3152 & w3154;
assign w3156 = ~w3153 & w3155;
assign w3157 = a[14] & ~w3156;
assign w3158 = ~a[14] & w3156;
assign w3159 = ~w3157 & ~w3158;
assign w3160 = b[12] & ~w1272;
assign w3161 = b[13] & w1154;
assign w3162 = b[14] & w1156;
assign w3163 = w714 & w1150;
assign w3164 = ~w3160 & ~w3161;
assign w3165 = ~w3162 & w3164;
assign w3166 = ~w3163 & w3165;
assign w3167 = a[20] & ~w3166;
assign w3168 = ~a[20] & w3166;
assign w3169 = ~w3167 & ~w3168;
assign w3170 = (a[32] & w2967) | (a[32] & w24936) | (w2967 & w24936);
assign w3171 = w2982 & w24776;
assign w3172 = a[32] & ~w3171;
assign w3173 = w22 & w2980;
assign w3174 = b[1] & w2973;
assign w3175 = b[2] & w2978;
assign w3176 = w2967 & w2972;
assign w3177 = ~w2977 & w3176;
assign w3178 = b[0] & w3177;
assign w3179 = ~w3173 & ~w3174;
assign w3180 = ~w3175 & w3179;
assign w3181 = ~w3178 & w3180;
assign w3182 = ~w3172 & w3181;
assign w3183 = w3172 & ~w3181;
assign w3184 = ~w3182 & ~w3183;
assign w3185 = b[5] & w2438;
assign w3186 = b[3] & ~w2622;
assign w3187 = b[4] & w2436;
assign w3188 = ~w3185 & ~w3186;
assign w3189 = ~w3187 & w3188;
assign w3190 = (~a[29] & ~w116) | (~a[29] & w24637) | (~w116 & w24637);
assign w3191 = w116 & w24638;
assign w3192 = ~w3190 & ~w3191;
assign w3193 = (a[29] & ~w3188) | (a[29] & w24937) | (~w3188 & w24937);
assign w3194 = (~w3193 & w3192) | (~w3193 & w24777) | (w3192 & w24777);
assign w3195 = w3184 & w3194;
assign w3196 = ~w3184 & ~w3194;
assign w3197 = ~w3195 & ~w3196;
assign w3198 = (~w2988 & ~w2989) | (~w2988 & w24639) | (~w2989 & w24639);
assign w3199 = ~w3197 & w3198;
assign w3200 = w3197 & ~w3198;
assign w3201 = ~w3199 & ~w3200;
assign w3202 = b[8] & w1957;
assign w3203 = b[6] & ~w2114;
assign w3204 = b[7] & w1955;
assign w3205 = w270 & w1951;
assign w3206 = ~w3202 & ~w3203;
assign w3207 = ~w3204 & w3206;
assign w3208 = ~w3205 & w3207;
assign w3209 = a[26] & ~w3208;
assign w3210 = ~a[26] & w3208;
assign w3211 = ~w3209 & ~w3210;
assign w3212 = w3201 & w3211;
assign w3213 = ~w3201 & ~w3211;
assign w3214 = ~w3212 & ~w3213;
assign w3215 = (~w3009 & ~w3011) | (~w3009 & w24778) | (~w3011 & w24778);
assign w3216 = ~w3214 & w3215;
assign w3217 = w3214 & ~w3215;
assign w3218 = ~w3216 & ~w3217;
assign w3219 = b[10] & w1517;
assign w3220 = b[11] & w1519;
assign w3221 = b[9] & ~w1676;
assign w3222 = w469 & w1513;
assign w3223 = ~w3219 & ~w3220;
assign w3224 = ~w3221 & w3223;
assign w3225 = ~w3222 & w3224;
assign w3226 = a[23] & ~w3225;
assign w3227 = ~a[23] & w3225;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = w3218 & w3228;
assign w3230 = ~w3218 & ~w3228;
assign w3231 = ~w3229 & ~w3230;
assign w3232 = ~w3025 & ~w3030;
assign w3233 = w3231 & w3232;
assign w3234 = ~w3231 & ~w3232;
assign w3235 = ~w3233 & ~w3234;
assign w3236 = ~w3169 & w3235;
assign w3237 = w3169 & ~w3235;
assign w3238 = ~w3236 & ~w3237;
assign w3239 = (~w3043 & w3045) | (~w3043 & w24366) | (w3045 & w24366);
assign w3240 = w3238 & ~w3239;
assign w3241 = ~w3238 & w3239;
assign w3242 = ~w3240 & ~w3241;
assign w3243 = b[15] & ~w934;
assign w3244 = b[16] & w838;
assign w3245 = b[17] & w834;
assign w3246 = w832 & w1008;
assign w3247 = ~w3243 & ~w3244;
assign w3248 = ~w3245 & w3247;
assign w3249 = ~w3246 & w3248;
assign w3250 = a[17] & ~w3249;
assign w3251 = ~a[17] & w3249;
assign w3252 = ~w3250 & ~w3251;
assign w3253 = w3242 & w3252;
assign w3254 = ~w3242 & ~w3252;
assign w3255 = ~w3253 & ~w3254;
assign w3256 = (~w3049 & ~w3052) | (~w3049 & w25108) | (~w3052 & w25108);
assign w3257 = w3255 & w3256;
assign w3258 = ~w3255 & ~w3256;
assign w3259 = ~w3257 & ~w3258;
assign w3260 = w3159 & ~w3259;
assign w3261 = ~w3159 & w3259;
assign w3262 = ~w3260 & ~w3261;
assign w3263 = (~w3067 & ~w3069) | (~w3067 & w24938) | (~w3069 & w24938);
assign w3264 = w3262 & w3263;
assign w3265 = ~w3262 & ~w3263;
assign w3266 = ~w3264 & ~w3265;
assign w3267 = ~w3149 & ~w3266;
assign w3268 = w3149 & w3266;
assign w3269 = ~w3267 & ~w3268;
assign w3270 = w3139 & w3269;
assign w3271 = ~w3139 & ~w3269;
assign w3272 = ~w3270 & ~w3271;
assign w3273 = w3138 & ~w3272;
assign w3274 = ~w3138 & w3272;
assign w3275 = ~w3273 & ~w3274;
assign w3276 = ~w3091 & ~w3094;
assign w3277 = ~w3275 & ~w3276;
assign w3278 = w3275 & w3276;
assign w3279 = ~w3277 & ~w3278;
assign w3280 = b[27] & w103;
assign w3281 = b[29] & w68;
assign w3282 = b[28] & w61;
assign w3283 = w66 & w2734;
assign w3284 = ~w3281 & ~w3282;
assign w3285 = ~w3280 & w3284;
assign w3286 = ~w3283 & w3285;
assign w3287 = a[5] & ~w3286;
assign w3288 = ~a[5] & w3286;
assign w3289 = ~w3287 & ~w3288;
assign w3290 = w3279 & w3289;
assign w3291 = ~w3279 & ~w3289;
assign w3292 = ~w3290 & ~w3291;
assign w3293 = w3128 & w3292;
assign w3294 = ~w3128 & ~w3292;
assign w3295 = ~w3293 & ~w3294;
assign w3296 = b[32] & w11;
assign w3297 = b[31] & w9;
assign w3298 = ~b[31] & ~b[32];
assign w3299 = b[31] & b[32];
assign w3300 = ~w3298 & ~w3299;
assign w3301 = ~w3106 & ~w3111;
assign w3302 = w3300 & w3301;
assign w3303 = ~w3300 & ~w3301;
assign w3304 = ~w3302 & ~w3303;
assign w3305 = w5 & w3304;
assign w3306 = ~w3296 & ~w3297;
assign w3307 = ~w3305 & w3306;
assign w3308 = b[30] & w24;
assign w3309 = a[2] & ~w3308;
assign w3310 = w3307 & ~w3309;
assign w3311 = a[2] & ~w3307;
assign w3312 = ~w3310 & ~w3311;
assign w3313 = ~w3295 & w3312;
assign w3314 = w3295 & ~w3312;
assign w3315 = ~w3313 & ~w3314;
assign w3316 = (~w3122 & ~w3124) | (~w3122 & w24939) | (~w3124 & w24939);
assign w3317 = w3315 & w3316;
assign w3318 = ~w3315 & ~w3316;
assign w3319 = ~w3317 & ~w3318;
assign w3320 = ~w3313 & ~w3317;
assign w3321 = b[28] & w103;
assign w3322 = b[30] & w68;
assign w3323 = b[29] & w61;
assign w3324 = w66 & ~w2908;
assign w3325 = ~w3322 & ~w3323;
assign w3326 = ~w3321 & w3325;
assign w3327 = ~w3324 & w3326;
assign w3328 = a[5] & ~w3327;
assign w3329 = ~a[5] & w3327;
assign w3330 = ~w3328 & ~w3329;
assign w3331 = b[24] & w360;
assign w3332 = b[23] & w358;
assign w3333 = b[22] & ~w419;
assign w3334 = w354 & w1895;
assign w3335 = ~w3331 & ~w3332;
assign w3336 = ~w3333 & w3335;
assign w3337 = ~w3334 & w3336;
assign w3338 = a[11] & ~w3337;
assign w3339 = ~a[11] & w3337;
assign w3340 = ~w3338 & ~w3339;
assign w3341 = (~w3260 & ~w3263) | (~w3260 & w25109) | (~w3263 & w25109);
assign w3342 = b[16] & ~w934;
assign w3343 = b[17] & w838;
assign w3344 = b[18] & w834;
assign w3345 = w832 & ~w1108;
assign w3346 = ~w3342 & ~w3343;
assign w3347 = ~w3344 & w3346;
assign w3348 = ~w3345 & w3347;
assign w3349 = a[17] & ~w3348;
assign w3350 = ~a[17] & w3348;
assign w3351 = ~w3349 & ~w3350;
assign w3352 = ~w3212 & ~w3217;
assign w3353 = w3176 & w24940;
assign w3354 = b[3] & w2978;
assign w3355 = b[2] & w2973;
assign w3356 = ~w3354 & ~w3355;
assign w3357 = ~w3353 & w3356;
assign w3358 = (a[32] & ~w3357) | (a[32] & w24941) | (~w3357 & w24941);
assign w3359 = w3357 & w24942;
assign w3360 = ~w3358 & ~w3359;
assign w3361 = a[32] & ~a[33];
assign w3362 = ~a[32] & a[33];
assign w3363 = ~w3361 & ~w3362;
assign w3364 = b[0] & ~w3363;
assign w3365 = w3181 & w24779;
assign w3366 = (~w3364 & ~w3181) | (~w3364 & w24780) | (~w3181 & w24780);
assign w3367 = ~w3365 & ~w3366;
assign w3368 = w3360 & w3367;
assign w3369 = ~w3360 & ~w3367;
assign w3370 = ~w3368 & ~w3369;
assign w3371 = b[5] & w2436;
assign w3372 = b[6] & w2438;
assign w3373 = b[4] & ~w2622;
assign w3374 = w157 & w2432;
assign w3375 = ~w3371 & ~w3372;
assign w3376 = ~w3373 & w3375;
assign w3377 = ~w3374 & w3376;
assign w3378 = a[29] & ~w3377;
assign w3379 = ~a[29] & w3377;
assign w3380 = ~w3378 & ~w3379;
assign w3381 = w3370 & w3380;
assign w3382 = ~w3370 & ~w3380;
assign w3383 = ~w3381 & ~w3382;
assign w3384 = (~w3195 & w3198) | (~w3195 & w24781) | (w3198 & w24781);
assign w3385 = w3383 & ~w3384;
assign w3386 = ~w3383 & w3384;
assign w3387 = ~w3385 & ~w3386;
assign w3388 = b[7] & ~w2114;
assign w3389 = b[9] & w1957;
assign w3390 = b[8] & w1955;
assign w3391 = w322 & w1951;
assign w3392 = ~w3388 & ~w3389;
assign w3393 = ~w3390 & w3392;
assign w3394 = ~w3391 & w3393;
assign w3395 = a[26] & ~w3394;
assign w3396 = ~a[26] & w3394;
assign w3397 = ~w3395 & ~w3396;
assign w3398 = w3387 & w3397;
assign w3399 = ~w3387 & ~w3397;
assign w3400 = ~w3398 & ~w3399;
assign w3401 = ~w3352 & ~w3400;
assign w3402 = w3352 & w3400;
assign w3403 = ~w3401 & ~w3402;
assign w3404 = b[11] & w1517;
assign w3405 = b[10] & ~w1676;
assign w3406 = b[12] & w1519;
assign w3407 = w536 & w1513;
assign w3408 = ~w3404 & ~w3405;
assign w3409 = ~w3406 & w3408;
assign w3410 = ~w3407 & w3409;
assign w3411 = a[23] & ~w3410;
assign w3412 = ~a[23] & w3410;
assign w3413 = ~w3411 & ~w3412;
assign w3414 = w3403 & ~w3413;
assign w3415 = ~w3403 & w3413;
assign w3416 = ~w3414 & ~w3415;
assign w3417 = (~w3230 & ~w3232) | (~w3230 & w24782) | (~w3232 & w24782);
assign w3418 = w3416 & w3417;
assign w3419 = ~w3416 & ~w3417;
assign w3420 = ~w3418 & ~w3419;
assign w3421 = b[15] & w1156;
assign w3422 = b[13] & ~w1272;
assign w3423 = b[14] & w1154;
assign w3424 = ~w799 & w1150;
assign w3425 = ~w3421 & ~w3422;
assign w3426 = ~w3423 & w3425;
assign w3427 = ~w3424 & w3426;
assign w3428 = a[20] & ~w3427;
assign w3429 = ~a[20] & w3427;
assign w3430 = ~w3428 & ~w3429;
assign w3431 = w3420 & w3430;
assign w3432 = ~w3420 & ~w3430;
assign w3433 = ~w3431 & ~w3432;
assign w3434 = (w3433 & w3240) | (w3433 & w24783) | (w3240 & w24783);
assign w3435 = ~w3240 & w24784;
assign w3436 = ~w3434 & ~w3435;
assign w3437 = w3351 & w3436;
assign w3438 = ~w3351 & ~w3436;
assign w3439 = ~w3437 & ~w3438;
assign w3440 = (~w3254 & ~w3256) | (~w3254 & w24367) | (~w3256 & w24367);
assign w3441 = ~w3439 & ~w3440;
assign w3442 = w3439 & w3440;
assign w3443 = ~w3441 & ~w3442;
assign w3444 = b[20] & w573;
assign w3445 = b[19] & ~w649;
assign w3446 = b[21] & w575;
assign w3447 = w569 & w1467;
assign w3448 = ~w3444 & ~w3445;
assign w3449 = ~w3446 & w3448;
assign w3450 = ~w3447 & w3449;
assign w3451 = a[14] & ~w3450;
assign w3452 = ~a[14] & w3450;
assign w3453 = ~w3451 & ~w3452;
assign w3454 = w3443 & w3453;
assign w3455 = ~w3443 & ~w3453;
assign w3456 = ~w3454 & ~w3455;
assign w3457 = ~w3341 & ~w3456;
assign w3458 = w3341 & w3456;
assign w3459 = ~w3457 & ~w3458;
assign w3460 = ~w3340 & w3459;
assign w3461 = w3340 & ~w3459;
assign w3462 = ~w3460 & ~w3461;
assign w3463 = (~w3267 & ~w3139) | (~w3267 & w24943) | (~w3139 & w24943);
assign w3464 = w3462 & w3463;
assign w3465 = ~w3462 & ~w3463;
assign w3466 = ~w3464 & ~w3465;
assign w3467 = b[25] & ~w237;
assign w3468 = b[26] & w183;
assign w3469 = b[27] & w185;
assign w3470 = w179 & w2378;
assign w3471 = ~w3467 & ~w3468;
assign w3472 = ~w3469 & w3471;
assign w3473 = ~w3470 & w3472;
assign w3474 = a[8] & ~w3473;
assign w3475 = ~a[8] & w3473;
assign w3476 = ~w3474 & ~w3475;
assign w3477 = w3466 & w3476;
assign w3478 = ~w3466 & ~w3476;
assign w3479 = ~w3477 & ~w3478;
assign w3480 = (~w3273 & ~w3276) | (~w3273 & w24640) | (~w3276 & w24640);
assign w3481 = ~w3479 & ~w3480;
assign w3482 = w3479 & w3480;
assign w3483 = ~w3481 & ~w3482;
assign w3484 = w3330 & ~w3483;
assign w3485 = ~w3330 & w3483;
assign w3486 = ~w3484 & ~w3485;
assign w3487 = ~w3291 & ~w3293;
assign w3488 = w3486 & w3487;
assign w3489 = ~w3486 & ~w3487;
assign w3490 = ~w3488 & ~w3489;
assign w3491 = b[33] & w11;
assign w3492 = b[32] & w9;
assign w3493 = (~w3299 & ~w3301) | (~w3299 & w24785) | (~w3301 & w24785);
assign w3494 = ~b[32] & ~b[33];
assign w3495 = b[32] & b[33];
assign w3496 = ~w3494 & ~w3495;
assign w3497 = w3493 & ~w3496;
assign w3498 = ~w3493 & w3496;
assign w3499 = ~w3497 & ~w3498;
assign w3500 = w5 & w3499;
assign w3501 = ~w3491 & ~w3492;
assign w3502 = ~w3500 & w3501;
assign w3503 = b[31] & w24;
assign w3504 = a[2] & ~w3503;
assign w3505 = w3502 & ~w3504;
assign w3506 = a[2] & ~w3502;
assign w3507 = ~w3505 & ~w3506;
assign w3508 = w3490 & w3507;
assign w3509 = ~w3490 & ~w3507;
assign w3510 = ~w3508 & ~w3509;
assign w3511 = w3320 & ~w3510;
assign w3512 = ~w3320 & w3510;
assign w3513 = ~w3511 & ~w3512;
assign w3514 = (~w3484 & ~w3487) | (~w3484 & w24641) | (~w3487 & w24641);
assign w3515 = b[28] & w185;
assign w3516 = b[26] & ~w237;
assign w3517 = b[27] & w183;
assign w3518 = w179 & w2559;
assign w3519 = ~w3515 & ~w3516;
assign w3520 = ~w3517 & w3519;
assign w3521 = ~w3518 & w3520;
assign w3522 = a[8] & ~w3521;
assign w3523 = ~a[8] & w3521;
assign w3524 = ~w3522 & ~w3523;
assign w3525 = (~w3461 & ~w3463) | (~w3461 & w25110) | (~w3463 & w25110);
assign w3526 = b[20] & ~w649;
assign w3527 = b[22] & w575;
assign w3528 = b[21] & w573;
assign w3529 = w569 & w1615;
assign w3530 = ~w3526 & ~w3527;
assign w3531 = ~w3528 & w3530;
assign w3532 = ~w3529 & w3531;
assign w3533 = a[14] & ~w3532;
assign w3534 = ~a[14] & w3532;
assign w3535 = ~w3533 & ~w3534;
assign w3536 = b[19] & w834;
assign w3537 = b[17] & ~w934;
assign w3538 = b[18] & w838;
assign w3539 = w832 & ~w1231;
assign w3540 = ~w3536 & ~w3537;
assign w3541 = ~w3538 & w3540;
assign w3542 = ~w3539 & w3541;
assign w3543 = a[17] & ~w3542;
assign w3544 = ~a[17] & w3542;
assign w3545 = ~w3543 & ~w3544;
assign w3546 = b[15] & w1154;
assign w3547 = b[14] & ~w1272;
assign w3548 = b[16] & w1156;
assign w3549 = w905 & w1150;
assign w3550 = ~w3546 & ~w3547;
assign w3551 = ~w3548 & w3550;
assign w3552 = ~w3549 & w3551;
assign w3553 = a[20] & ~w3552;
assign w3554 = ~a[20] & w3552;
assign w3555 = ~w3553 & ~w3554;
assign w3556 = ~w3415 & ~w3418;
assign w3557 = ~w3381 & ~w3385;
assign w3558 = (~w3365 & ~w3367) | (~w3365 & w24944) | (~w3367 & w24944);
assign w3559 = w3176 & w24786;
assign w3560 = b[3] & w2973;
assign w3561 = b[4] & w2978;
assign w3562 = w84 & w2980;
assign w3563 = ~w3560 & ~w3561;
assign w3564 = ~w3559 & w3563;
assign w3565 = ~w3562 & w3564;
assign w3566 = a[32] & ~w3565;
assign w3567 = ~a[32] & w3565;
assign w3568 = ~w3566 & ~w3567;
assign w3569 = a[35] & w3364;
assign w3570 = a[34] & ~a[35];
assign w3571 = ~a[34] & a[35];
assign w3572 = ~w3570 & ~w3571;
assign w3573 = ~w3363 & ~w3572;
assign w3574 = ~w8 & w3573;
assign w3575 = a[33] & ~a[34];
assign w3576 = ~a[33] & a[34];
assign w3577 = ~w3575 & ~w3576;
assign w3578 = w3363 & ~w3577;
assign w3579 = b[0] & w3578;
assign w3580 = ~w3363 & w3572;
assign w3581 = b[1] & w3580;
assign w3582 = ~w3574 & ~w3579;
assign w3583 = ~w3581 & w3582;
assign w3584 = ~w3569 & w3583;
assign w3585 = w3569 & ~w3583;
assign w3586 = ~w3584 & ~w3585;
assign w3587 = ~w3568 & ~w3586;
assign w3588 = w3568 & w3586;
assign w3589 = ~w3587 & ~w3588;
assign w3590 = ~w3558 & w3589;
assign w3591 = w3558 & ~w3589;
assign w3592 = ~w3590 & ~w3591;
assign w3593 = b[5] & ~w2622;
assign w3594 = b[6] & w2436;
assign w3595 = b[7] & w2438;
assign w3596 = w216 & w2432;
assign w3597 = ~w3593 & ~w3594;
assign w3598 = ~w3595 & w3597;
assign w3599 = ~w3596 & w3598;
assign w3600 = a[29] & ~w3599;
assign w3601 = ~a[29] & w3599;
assign w3602 = ~w3600 & ~w3601;
assign w3603 = ~w3592 & ~w3602;
assign w3604 = w3592 & w3602;
assign w3605 = ~w3603 & ~w3604;
assign w3606 = w3557 & ~w3605;
assign w3607 = ~w3557 & w3605;
assign w3608 = ~w3606 & ~w3607;
assign w3609 = b[9] & w1955;
assign w3610 = b[8] & ~w2114;
assign w3611 = b[10] & w1957;
assign w3612 = w397 & w1951;
assign w3613 = ~w3609 & ~w3610;
assign w3614 = ~w3611 & w3613;
assign w3615 = ~w3612 & w3614;
assign w3616 = a[26] & ~w3615;
assign w3617 = ~a[26] & w3615;
assign w3618 = ~w3616 & ~w3617;
assign w3619 = w3608 & w3618;
assign w3620 = ~w3608 & ~w3618;
assign w3621 = ~w3619 & ~w3620;
assign w3622 = (~w3399 & ~w3352) | (~w3399 & w24787) | (~w3352 & w24787);
assign w3623 = ~w3621 & ~w3622;
assign w3624 = w3621 & w3622;
assign w3625 = ~w3623 & ~w3624;
assign w3626 = b[11] & ~w1676;
assign w3627 = b[13] & w1519;
assign w3628 = b[12] & w1517;
assign w3629 = w628 & w1513;
assign w3630 = ~w3626 & ~w3627;
assign w3631 = ~w3628 & w3630;
assign w3632 = ~w3629 & w3631;
assign w3633 = a[23] & ~w3632;
assign w3634 = ~a[23] & w3632;
assign w3635 = ~w3633 & ~w3634;
assign w3636 = w3625 & w3635;
assign w3637 = ~w3625 & ~w3635;
assign w3638 = ~w3636 & ~w3637;
assign w3639 = w3556 & w3638;
assign w3640 = ~w3556 & ~w3638;
assign w3641 = ~w3639 & ~w3640;
assign w3642 = w3555 & ~w3641;
assign w3643 = ~w3555 & w3641;
assign w3644 = ~w3642 & ~w3643;
assign w3645 = ~w3431 & ~w3434;
assign w3646 = w3644 & ~w3645;
assign w3647 = ~w3644 & w3645;
assign w3648 = ~w3646 & ~w3647;
assign w3649 = w3545 & w3648;
assign w3650 = ~w3545 & ~w3648;
assign w3651 = ~w3649 & ~w3650;
assign w3652 = (~w3437 & ~w3440) | (~w3437 & w24788) | (~w3440 & w24788);
assign w3653 = ~w3651 & ~w3652;
assign w3654 = w3651 & w3652;
assign w3655 = ~w3653 & ~w3654;
assign w3656 = w3535 & ~w3655;
assign w3657 = ~w3535 & w3655;
assign w3658 = ~w3656 & ~w3657;
assign w3659 = (~w3455 & ~w3341) | (~w3455 & w24368) | (~w3341 & w24368);
assign w3660 = ~w3658 & ~w3659;
assign w3661 = w3658 & w3659;
assign w3662 = ~w3660 & ~w3661;
assign w3663 = b[25] & w360;
assign w3664 = b[23] & ~w419;
assign w3665 = b[24] & w358;
assign w3666 = w354 & w2061;
assign w3667 = ~w3663 & ~w3664;
assign w3668 = ~w3665 & w3667;
assign w3669 = ~w3666 & w3668;
assign w3670 = a[11] & ~w3669;
assign w3671 = ~a[11] & w3669;
assign w3672 = ~w3670 & ~w3671;
assign w3673 = w3662 & w3672;
assign w3674 = ~w3662 & ~w3672;
assign w3675 = ~w3673 & ~w3674;
assign w3676 = ~w3525 & ~w3675;
assign w3677 = w3525 & w3675;
assign w3678 = ~w3676 & ~w3677;
assign w3679 = w3524 & ~w3678;
assign w3680 = ~w3524 & w3678;
assign w3681 = ~w3679 & ~w3680;
assign w3682 = (~w3478 & ~w3480) | (~w3478 & w24945) | (~w3480 & w24945);
assign w3683 = ~w3681 & ~w3682;
assign w3684 = w3681 & w3682;
assign w3685 = ~w3683 & ~w3684;
assign w3686 = b[29] & w103;
assign w3687 = b[30] & w61;
assign w3688 = b[31] & w68;
assign w3689 = w66 & ~w3112;
assign w3690 = ~w3687 & ~w3688;
assign w3691 = ~w3686 & w3690;
assign w3692 = ~w3689 & w3691;
assign w3693 = a[5] & ~w3692;
assign w3694 = ~a[5] & w3692;
assign w3695 = ~w3693 & ~w3694;
assign w3696 = ~w3685 & ~w3695;
assign w3697 = w3685 & w3695;
assign w3698 = ~w3696 & ~w3697;
assign w3699 = w3514 & w3698;
assign w3700 = ~w3514 & ~w3698;
assign w3701 = ~w3699 & ~w3700;
assign w3702 = b[34] & w11;
assign w3703 = b[33] & w9;
assign w3704 = ~b[33] & ~b[34];
assign w3705 = b[33] & b[34];
assign w3706 = ~w3704 & ~w3705;
assign w3707 = ~w3495 & ~w3498;
assign w3708 = ~w3706 & ~w3707;
assign w3709 = w3706 & w3707;
assign w3710 = ~w3708 & ~w3709;
assign w3711 = w5 & ~w3710;
assign w3712 = ~w3702 & ~w3703;
assign w3713 = ~w3711 & w3712;
assign w3714 = b[32] & w24;
assign w3715 = a[2] & ~w3714;
assign w3716 = w3713 & ~w3715;
assign w3717 = a[2] & ~w3713;
assign w3718 = ~w3716 & ~w3717;
assign w3719 = ~w3701 & w3718;
assign w3720 = w3701 & ~w3718;
assign w3721 = ~w3719 & ~w3720;
assign w3722 = ~w3508 & ~w3512;
assign w3723 = w3721 & ~w3722;
assign w3724 = ~w3721 & w3722;
assign w3725 = ~w3723 & ~w3724;
assign w3726 = (~w3719 & w3722) | (~w3719 & w24642) | (w3722 & w24642);
assign w3727 = b[30] & w103;
assign w3728 = b[32] & w68;
assign w3729 = b[31] & w61;
assign w3730 = w66 & w3304;
assign w3731 = ~w3728 & ~w3729;
assign w3732 = ~w3727 & w3731;
assign w3733 = ~w3730 & w3732;
assign w3734 = a[5] & ~w3733;
assign w3735 = ~a[5] & w3733;
assign w3736 = ~w3734 & ~w3735;
assign w3737 = b[24] & ~w419;
assign w3738 = b[26] & w360;
assign w3739 = b[25] & w358;
assign w3740 = w354 & w2219;
assign w3741 = ~w3737 & ~w3738;
assign w3742 = ~w3739 & w3741;
assign w3743 = ~w3740 & w3742;
assign w3744 = a[11] & ~w3743;
assign w3745 = ~a[11] & w3743;
assign w3746 = ~w3744 & ~w3745;
assign w3747 = (~w3656 & ~w3659) | (~w3656 & w24789) | (~w3659 & w24789);
assign w3748 = b[18] & ~w934;
assign w3749 = b[19] & w838;
assign w3750 = b[20] & w834;
assign w3751 = w832 & w1347;
assign w3752 = ~w3748 & ~w3749;
assign w3753 = ~w3750 & w3752;
assign w3754 = ~w3751 & w3753;
assign w3755 = a[17] & ~w3754;
assign w3756 = ~a[17] & w3754;
assign w3757 = ~w3755 & ~w3756;
assign w3758 = b[14] & w1519;
assign w3759 = b[12] & ~w1676;
assign w3760 = b[13] & w1517;
assign w3761 = w714 & w1513;
assign w3762 = ~w3758 & ~w3759;
assign w3763 = ~w3760 & w3762;
assign w3764 = ~w3761 & w3763;
assign w3765 = a[23] & ~w3764;
assign w3766 = ~a[23] & w3764;
assign w3767 = ~w3765 & ~w3766;
assign w3768 = ~w3619 & ~w3624;
assign w3769 = ~w3604 & ~w3607;
assign w3770 = w3176 & w25111;
assign w3771 = b[5] & w2978;
assign w3772 = b[4] & w2973;
assign w3773 = w116 & w2980;
assign w3774 = ~w3771 & ~w3772;
assign w3775 = (a[32] & w3773) | (a[32] & w24946) | (w3773 & w24946);
assign w3776 = ~w3773 & w24947;
assign w3777 = ~w3775 & ~w3776;
assign w3778 = (a[35] & w3363) | (a[35] & w24790) | (w3363 & w24790);
assign w3779 = w3582 & w24643;
assign w3780 = a[35] & ~w3779;
assign w3781 = b[1] & w3578;
assign w3782 = w22 & w3573;
assign w3783 = b[2] & w3580;
assign w3784 = w3363 & ~w3572;
assign w3785 = w3577 & w3784;
assign w3786 = b[0] & w3785;
assign w3787 = ~w3781 & ~w3782;
assign w3788 = ~w3783 & w3787;
assign w3789 = ~w3786 & w3788;
assign w3790 = ~w3780 & w3789;
assign w3791 = w3780 & ~w3789;
assign w3792 = ~w3790 & ~w3791;
assign w3793 = w3777 & w3792;
assign w3794 = ~w3777 & ~w3792;
assign w3795 = ~w3793 & ~w3794;
assign w3796 = (~w3588 & ~w3589) | (~w3588 & w24948) | (~w3589 & w24948);
assign w3797 = ~w3795 & w3796;
assign w3798 = w3795 & ~w3796;
assign w3799 = ~w3797 & ~w3798;
assign w3800 = b[6] & ~w2622;
assign w3801 = b[8] & w2438;
assign w3802 = b[7] & w2436;
assign w3803 = w270 & w2432;
assign w3804 = ~w3800 & ~w3801;
assign w3805 = ~w3802 & w3804;
assign w3806 = ~w3803 & w3805;
assign w3807 = a[29] & ~w3806;
assign w3808 = ~a[29] & w3806;
assign w3809 = ~w3807 & ~w3808;
assign w3810 = w3799 & w3809;
assign w3811 = ~w3799 & ~w3809;
assign w3812 = ~w3810 & ~w3811;
assign w3813 = ~w3769 & w3812;
assign w3814 = w3769 & ~w3812;
assign w3815 = ~w3813 & ~w3814;
assign w3816 = b[9] & ~w2114;
assign w3817 = b[10] & w1955;
assign w3818 = b[11] & w1957;
assign w3819 = w469 & w1951;
assign w3820 = ~w3816 & ~w3817;
assign w3821 = ~w3818 & w3820;
assign w3822 = ~w3819 & w3821;
assign w3823 = a[26] & ~w3822;
assign w3824 = ~a[26] & w3822;
assign w3825 = ~w3823 & ~w3824;
assign w3826 = ~w3815 & ~w3825;
assign w3827 = w3815 & w3825;
assign w3828 = ~w3826 & ~w3827;
assign w3829 = ~w3768 & w3828;
assign w3830 = w3768 & ~w3828;
assign w3831 = ~w3829 & ~w3830;
assign w3832 = ~w3767 & ~w3831;
assign w3833 = w3767 & w3831;
assign w3834 = ~w3832 & ~w3833;
assign w3835 = (~w3637 & ~w3556) | (~w3637 & w25112) | (~w3556 & w25112);
assign w3836 = w3834 & w3835;
assign w3837 = ~w3834 & ~w3835;
assign w3838 = ~w3836 & ~w3837;
assign w3839 = b[15] & ~w1272;
assign w3840 = b[17] & w1156;
assign w3841 = b[16] & w1154;
assign w3842 = w1008 & w1150;
assign w3843 = ~w3839 & ~w3840;
assign w3844 = ~w3841 & w3843;
assign w3845 = ~w3842 & w3844;
assign w3846 = a[20] & ~w3845;
assign w3847 = ~a[20] & w3845;
assign w3848 = ~w3846 & ~w3847;
assign w3849 = w3838 & w3848;
assign w3850 = ~w3838 & ~w3848;
assign w3851 = ~w3849 & ~w3850;
assign w3852 = ~w3642 & ~w3646;
assign w3853 = w3851 & ~w3852;
assign w3854 = ~w3851 & w3852;
assign w3855 = ~w3853 & ~w3854;
assign w3856 = w3757 & w3855;
assign w3857 = ~w3757 & ~w3855;
assign w3858 = ~w3856 & ~w3857;
assign w3859 = (~w3650 & ~w3652) | (~w3650 & w25113) | (~w3652 & w25113);
assign w3860 = w3858 & w3859;
assign w3861 = ~w3858 & ~w3859;
assign w3862 = ~w3860 & ~w3861;
assign w3863 = b[23] & w575;
assign w3864 = b[21] & ~w649;
assign w3865 = b[22] & w573;
assign w3866 = w569 & w1755;
assign w3867 = ~w3863 & ~w3864;
assign w3868 = ~w3865 & w3867;
assign w3869 = ~w3866 & w3868;
assign w3870 = a[14] & ~w3869;
assign w3871 = ~a[14] & w3869;
assign w3872 = ~w3870 & ~w3871;
assign w3873 = ~w3862 & ~w3872;
assign w3874 = w3862 & w3872;
assign w3875 = ~w3873 & ~w3874;
assign w3876 = w3747 & ~w3875;
assign w3877 = ~w3747 & w3875;
assign w3878 = ~w3876 & ~w3877;
assign w3879 = ~w3746 & ~w3878;
assign w3880 = w3746 & w3878;
assign w3881 = ~w3879 & ~w3880;
assign w3882 = (~w3674 & ~w3525) | (~w3674 & w24369) | (~w3525 & w24369);
assign w3883 = w3881 & w3882;
assign w3884 = ~w3881 & ~w3882;
assign w3885 = ~w3883 & ~w3884;
assign w3886 = b[27] & ~w237;
assign w3887 = b[29] & w185;
assign w3888 = b[28] & w183;
assign w3889 = w179 & w2734;
assign w3890 = ~w3886 & ~w3887;
assign w3891 = ~w3888 & w3890;
assign w3892 = ~w3889 & w3891;
assign w3893 = a[8] & ~w3892;
assign w3894 = ~a[8] & w3892;
assign w3895 = ~w3893 & ~w3894;
assign w3896 = w3885 & w3895;
assign w3897 = ~w3885 & ~w3895;
assign w3898 = ~w3896 & ~w3897;
assign w3899 = (~w3679 & ~w3682) | (~w3679 & w25114) | (~w3682 & w25114);
assign w3900 = ~w3898 & ~w3899;
assign w3901 = w3898 & w3899;
assign w3902 = ~w3900 & ~w3901;
assign w3903 = w3736 & ~w3902;
assign w3904 = ~w3736 & w3902;
assign w3905 = ~w3903 & ~w3904;
assign w3906 = (~w3696 & ~w3514) | (~w3696 & w24949) | (~w3514 & w24949);
assign w3907 = w3905 & w3906;
assign w3908 = ~w3905 & ~w3906;
assign w3909 = ~w3907 & ~w3908;
assign w3910 = b[35] & w11;
assign w3911 = b[34] & w9;
assign w3912 = ~b[34] & ~b[35];
assign w3913 = b[34] & b[35];
assign w3914 = ~w3912 & ~w3913;
assign w3915 = ~w3704 & ~w3709;
assign w3916 = ~w3914 & ~w3915;
assign w3917 = w3914 & w3915;
assign w3918 = ~w3916 & ~w3917;
assign w3919 = w5 & w3918;
assign w3920 = ~w3910 & ~w3911;
assign w3921 = ~w3919 & w3920;
assign w3922 = b[33] & w24;
assign w3923 = a[2] & ~w3922;
assign w3924 = w3921 & ~w3923;
assign w3925 = a[2] & ~w3921;
assign w3926 = ~w3924 & ~w3925;
assign w3927 = w3909 & w3926;
assign w3928 = ~w3909 & ~w3926;
assign w3929 = ~w3927 & ~w3928;
assign w3930 = w3726 & ~w3929;
assign w3931 = ~w3726 & w3929;
assign w3932 = ~w3930 & ~w3931;
assign w3933 = (~w3903 & ~w3906) | (~w3903 & w25115) | (~w3906 & w25115);
assign w3934 = b[31] & w103;
assign w3935 = b[33] & w68;
assign w3936 = b[32] & w61;
assign w3937 = w66 & w3499;
assign w3938 = ~w3935 & ~w3936;
assign w3939 = ~w3934 & w3938;
assign w3940 = ~w3937 & w3939;
assign w3941 = a[5] & ~w3940;
assign w3942 = ~a[5] & w3940;
assign w3943 = ~w3941 & ~w3942;
assign w3944 = b[28] & ~w237;
assign w3945 = b[30] & w185;
assign w3946 = b[29] & w183;
assign w3947 = w179 & ~w2908;
assign w3948 = ~w3944 & ~w3945;
assign w3949 = ~w3946 & w3948;
assign w3950 = ~w3947 & w3949;
assign w3951 = a[8] & ~w3950;
assign w3952 = ~a[8] & w3950;
assign w3953 = ~w3951 & ~w3952;
assign w3954 = (~w3880 & ~w3882) | (~w3880 & w24791) | (~w3882 & w24791);
assign w3955 = b[24] & w575;
assign w3956 = b[22] & ~w649;
assign w3957 = b[23] & w573;
assign w3958 = w569 & w1895;
assign w3959 = ~w3955 & ~w3956;
assign w3960 = ~w3957 & w3959;
assign w3961 = ~w3958 & w3960;
assign w3962 = a[14] & ~w3961;
assign w3963 = ~a[14] & w3961;
assign w3964 = ~w3962 & ~w3963;
assign w3965 = ~w3856 & ~w3860;
assign w3966 = (~w3849 & w3852) | (~w3849 & w25255) | (w3852 & w25255);
assign w3967 = b[16] & ~w1272;
assign w3968 = b[18] & w1156;
assign w3969 = b[17] & w1154;
assign w3970 = ~w1108 & w1150;
assign w3971 = ~w3967 & ~w3968;
assign w3972 = ~w3969 & w3971;
assign w3973 = ~w3970 & w3972;
assign w3974 = a[20] & ~w3973;
assign w3975 = ~a[20] & w3973;
assign w3976 = ~w3974 & ~w3975;
assign w3977 = ~w3833 & ~w3836;
assign w3978 = (~w3810 & w3769) | (~w3810 & w24950) | (w3769 & w24950);
assign w3979 = w3784 & w24792;
assign w3980 = b[2] & w3578;
assign w3981 = b[3] & w3580;
assign w3982 = ~w3980 & ~w3981;
assign w3983 = ~w3979 & w3982;
assign w3984 = (a[35] & ~w3983) | (a[35] & w24793) | (~w3983 & w24793);
assign w3985 = w3983 & w24794;
assign w3986 = ~w3984 & ~w3985;
assign w3987 = a[35] & ~a[36];
assign w3988 = ~a[35] & a[36];
assign w3989 = ~w3987 & ~w3988;
assign w3990 = b[0] & ~w3989;
assign w3991 = w3789 & w24644;
assign w3992 = (~w3990 & ~w3789) | (~w3990 & w24645) | (~w3789 & w24645);
assign w3993 = ~w3991 & ~w3992;
assign w3994 = w3986 & w3993;
assign w3995 = ~w3986 & ~w3993;
assign w3996 = ~w3994 & ~w3995;
assign w3997 = b[4] & w3177;
assign w3998 = b[6] & w2978;
assign w3999 = b[5] & w2973;
assign w4000 = w157 & w2980;
assign w4001 = ~w3998 & ~w3999;
assign w4002 = ~w3997 & w4001;
assign w4003 = ~w4000 & w4002;
assign w4004 = a[32] & ~w4003;
assign w4005 = ~a[32] & w4003;
assign w4006 = ~w4004 & ~w4005;
assign w4007 = w3996 & w4006;
assign w4008 = ~w3996 & ~w4006;
assign w4009 = ~w4007 & ~w4008;
assign w4010 = (~w3793 & w3796) | (~w3793 & w24795) | (w3796 & w24795);
assign w4011 = w4009 & ~w4010;
assign w4012 = ~w4009 & w4010;
assign w4013 = ~w4011 & ~w4012;
assign w4014 = b[7] & ~w2622;
assign w4015 = b[8] & w2436;
assign w4016 = b[9] & w2438;
assign w4017 = w322 & w2432;
assign w4018 = ~w4014 & ~w4015;
assign w4019 = ~w4016 & w4018;
assign w4020 = ~w4017 & w4019;
assign w4021 = a[29] & ~w4020;
assign w4022 = ~a[29] & w4020;
assign w4023 = ~w4021 & ~w4022;
assign w4024 = w4013 & w4023;
assign w4025 = ~w4013 & ~w4023;
assign w4026 = ~w4024 & ~w4025;
assign w4027 = w3978 & ~w4026;
assign w4028 = ~w3978 & w4026;
assign w4029 = ~w4027 & ~w4028;
assign w4030 = b[12] & w1957;
assign w4031 = b[11] & w1955;
assign w4032 = b[10] & ~w2114;
assign w4033 = w536 & w1951;
assign w4034 = ~w4030 & ~w4031;
assign w4035 = ~w4032 & w4034;
assign w4036 = ~w4033 & w4035;
assign w4037 = a[26] & ~w4036;
assign w4038 = ~a[26] & w4036;
assign w4039 = ~w4037 & ~w4038;
assign w4040 = ~w4029 & ~w4039;
assign w4041 = w4029 & w4039;
assign w4042 = ~w4040 & ~w4041;
assign w4043 = ~w3827 & ~w3829;
assign w4044 = w4042 & ~w4043;
assign w4045 = ~w4042 & w4043;
assign w4046 = ~w4044 & ~w4045;
assign w4047 = b[15] & w1519;
assign w4048 = b[13] & ~w1676;
assign w4049 = b[14] & w1517;
assign w4050 = ~w799 & w1513;
assign w4051 = ~w4047 & ~w4048;
assign w4052 = ~w4049 & w4051;
assign w4053 = ~w4050 & w4052;
assign w4054 = a[23] & ~w4053;
assign w4055 = ~a[23] & w4053;
assign w4056 = ~w4054 & ~w4055;
assign w4057 = w4046 & w4056;
assign w4058 = ~w4046 & ~w4056;
assign w4059 = ~w4057 & ~w4058;
assign w4060 = w3977 & w4059;
assign w4061 = ~w3977 & ~w4059;
assign w4062 = ~w4060 & ~w4061;
assign w4063 = w3976 & ~w4062;
assign w4064 = ~w3976 & w4062;
assign w4065 = ~w4063 & ~w4064;
assign w4066 = w3966 & ~w4065;
assign w4067 = ~w3966 & w4065;
assign w4068 = ~w4066 & ~w4067;
assign w4069 = b[19] & ~w934;
assign w4070 = b[20] & w838;
assign w4071 = b[21] & w834;
assign w4072 = w832 & w1467;
assign w4073 = ~w4069 & ~w4070;
assign w4074 = ~w4071 & w4073;
assign w4075 = ~w4072 & w4074;
assign w4076 = a[17] & ~w4075;
assign w4077 = ~a[17] & w4075;
assign w4078 = ~w4076 & ~w4077;
assign w4079 = w4068 & w4078;
assign w4080 = ~w4068 & ~w4078;
assign w4081 = ~w4079 & ~w4080;
assign w4082 = ~w3965 & w4081;
assign w4083 = w3965 & ~w4081;
assign w4084 = ~w4082 & ~w4083;
assign w4085 = ~w3964 & ~w4084;
assign w4086 = w3964 & w4084;
assign w4087 = ~w4085 & ~w4086;
assign w4088 = (~w3874 & w3747) | (~w3874 & w25116) | (w3747 & w25116);
assign w4089 = w4087 & ~w4088;
assign w4090 = ~w4087 & w4088;
assign w4091 = ~w4089 & ~w4090;
assign w4092 = b[26] & w358;
assign w4093 = b[27] & w360;
assign w4094 = b[25] & ~w419;
assign w4095 = w354 & w2378;
assign w4096 = ~w4092 & ~w4093;
assign w4097 = ~w4094 & w4096;
assign w4098 = ~w4095 & w4097;
assign w4099 = a[11] & ~w4098;
assign w4100 = ~a[11] & w4098;
assign w4101 = ~w4099 & ~w4100;
assign w4102 = w4091 & w4101;
assign w4103 = ~w4091 & ~w4101;
assign w4104 = ~w4102 & ~w4103;
assign w4105 = w3954 & w4104;
assign w4106 = ~w3954 & ~w4104;
assign w4107 = ~w4105 & ~w4106;
assign w4108 = ~w3953 & w4107;
assign w4109 = w3953 & ~w4107;
assign w4110 = ~w4108 & ~w4109;
assign w4111 = (~w3897 & ~w3899) | (~w3897 & w24370) | (~w3899 & w24370);
assign w4112 = w4110 & w4111;
assign w4113 = ~w4110 & ~w4111;
assign w4114 = ~w4112 & ~w4113;
assign w4115 = w3943 & w4114;
assign w4116 = ~w3943 & ~w4114;
assign w4117 = ~w4115 & ~w4116;
assign w4118 = w3933 & w4117;
assign w4119 = ~w3933 & ~w4117;
assign w4120 = ~w4118 & ~w4119;
assign w4121 = b[36] & w11;
assign w4122 = b[35] & w9;
assign w4123 = ~w3913 & ~w3917;
assign w4124 = ~b[35] & ~b[36];
assign w4125 = b[35] & b[36];
assign w4126 = ~w4124 & ~w4125;
assign w4127 = w4123 & ~w4126;
assign w4128 = ~w4123 & w4126;
assign w4129 = ~w4127 & ~w4128;
assign w4130 = w5 & w4129;
assign w4131 = ~w4121 & ~w4122;
assign w4132 = ~w4130 & w4131;
assign w4133 = b[34] & w24;
assign w4134 = a[2] & ~w4133;
assign w4135 = w4132 & ~w4134;
assign w4136 = a[2] & ~w4132;
assign w4137 = ~w4135 & ~w4136;
assign w4138 = ~w4120 & w4137;
assign w4139 = w4120 & ~w4137;
assign w4140 = ~w4138 & ~w4139;
assign w4141 = (~w3927 & w3726) | (~w3927 & w24951) | (w3726 & w24951);
assign w4142 = w4140 & ~w4141;
assign w4143 = ~w4140 & w4141;
assign w4144 = ~w4142 & ~w4143;
assign w4145 = (~w4138 & w4141) | (~w4138 & w25117) | (w4141 & w25117);
assign w4146 = b[32] & w103;
assign w4147 = b[34] & w68;
assign w4148 = b[33] & w61;
assign w4149 = w66 & ~w3710;
assign w4150 = ~w4147 & ~w4148;
assign w4151 = ~w4146 & w4150;
assign w4152 = ~w4149 & w4151;
assign w4153 = a[5] & ~w4152;
assign w4154 = ~a[5] & w4152;
assign w4155 = ~w4153 & ~w4154;
assign w4156 = (~w4109 & ~w4111) | (~w4109 & w24796) | (~w4111 & w24796);
assign w4157 = b[29] & ~w237;
assign w4158 = b[30] & w183;
assign w4159 = b[31] & w185;
assign w4160 = w179 & ~w3112;
assign w4161 = ~w4157 & ~w4158;
assign w4162 = ~w4159 & w4161;
assign w4163 = ~w4160 & w4162;
assign w4164 = a[8] & ~w4163;
assign w4165 = ~a[8] & w4163;
assign w4166 = ~w4164 & ~w4165;
assign w4167 = b[28] & w360;
assign w4168 = b[26] & ~w419;
assign w4169 = b[27] & w358;
assign w4170 = w354 & w2559;
assign w4171 = ~w4167 & ~w4168;
assign w4172 = ~w4169 & w4171;
assign w4173 = ~w4170 & w4172;
assign w4174 = a[11] & ~w4173;
assign w4175 = ~a[11] & w4173;
assign w4176 = ~w4174 & ~w4175;
assign w4177 = ~w4086 & ~w4089;
assign w4178 = ~w4079 & ~w4082;
assign w4179 = b[20] & ~w934;
assign w4180 = b[21] & w838;
assign w4181 = b[22] & w834;
assign w4182 = w832 & w1615;
assign w4183 = ~w4179 & ~w4180;
assign w4184 = ~w4181 & w4183;
assign w4185 = ~w4182 & w4184;
assign w4186 = a[17] & ~w4185;
assign w4187 = ~a[17] & w4185;
assign w4188 = ~w4186 & ~w4187;
assign w4189 = b[14] & ~w1676;
assign w4190 = b[15] & w1517;
assign w4191 = b[16] & w1519;
assign w4192 = w905 & w1513;
assign w4193 = ~w4189 & ~w4190;
assign w4194 = ~w4191 & w4193;
assign w4195 = ~w4192 & w4194;
assign w4196 = a[23] & ~w4195;
assign w4197 = ~a[23] & w4195;
assign w4198 = ~w4196 & ~w4197;
assign w4199 = (~w4041 & w4043) | (~w4041 & w24952) | (w4043 & w24952);
assign w4200 = b[13] & w1957;
assign w4201 = b[12] & w1955;
assign w4202 = b[11] & ~w2114;
assign w4203 = w628 & w1951;
assign w4204 = ~w4200 & ~w4201;
assign w4205 = ~w4202 & w4204;
assign w4206 = ~w4203 & w4205;
assign w4207 = a[26] & ~w4206;
assign w4208 = ~a[26] & w4206;
assign w4209 = ~w4207 & ~w4208;
assign w4210 = b[9] & w2436;
assign w4211 = b[10] & w2438;
assign w4212 = b[8] & ~w2622;
assign w4213 = w397 & w2432;
assign w4214 = ~w4210 & ~w4211;
assign w4215 = ~w4212 & w4214;
assign w4216 = ~w4213 & w4215;
assign w4217 = a[29] & ~w4216;
assign w4218 = ~a[29] & w4216;
assign w4219 = ~w4217 & ~w4218;
assign w4220 = ~w4007 & ~w4011;
assign w4221 = (~w3991 & ~w3993) | (~w3991 & w24797) | (~w3993 & w24797);
assign w4222 = w3784 & w24798;
assign w4223 = b[3] & w3578;
assign w4224 = b[4] & w3580;
assign w4225 = w84 & w3573;
assign w4226 = ~w4223 & ~w4224;
assign w4227 = ~w4222 & w4226;
assign w4228 = ~w4225 & w4227;
assign w4229 = a[35] & ~w4228;
assign w4230 = ~a[35] & w4228;
assign w4231 = ~w4229 & ~w4230;
assign w4232 = a[38] & w3990;
assign w4233 = a[37] & ~a[38];
assign w4234 = ~a[37] & a[38];
assign w4235 = ~w4233 & ~w4234;
assign w4236 = ~w3989 & ~w4235;
assign w4237 = ~w8 & w4236;
assign w4238 = a[36] & ~a[37];
assign w4239 = ~a[36] & a[37];
assign w4240 = ~w4238 & ~w4239;
assign w4241 = w3989 & ~w4240;
assign w4242 = b[0] & w4241;
assign w4243 = ~w3989 & w4235;
assign w4244 = b[1] & w4243;
assign w4245 = ~w4237 & ~w4242;
assign w4246 = ~w4244 & w4245;
assign w4247 = ~w4232 & w4246;
assign w4248 = w4232 & ~w4246;
assign w4249 = ~w4247 & ~w4248;
assign w4250 = ~w4231 & ~w4249;
assign w4251 = w4231 & w4249;
assign w4252 = ~w4250 & ~w4251;
assign w4253 = w4221 & ~w4252;
assign w4254 = ~w4221 & w4252;
assign w4255 = ~w4253 & ~w4254;
assign w4256 = b[5] & w3177;
assign w4257 = b[6] & w2973;
assign w4258 = b[7] & w2978;
assign w4259 = w216 & w2980;
assign w4260 = ~w4257 & ~w4258;
assign w4261 = ~w4256 & w4260;
assign w4262 = ~w4259 & w4261;
assign w4263 = a[32] & ~w4262;
assign w4264 = ~a[32] & w4262;
assign w4265 = ~w4263 & ~w4264;
assign w4266 = ~w4255 & ~w4265;
assign w4267 = w4255 & w4265;
assign w4268 = ~w4266 & ~w4267;
assign w4269 = w4220 & ~w4268;
assign w4270 = ~w4220 & w4268;
assign w4271 = ~w4269 & ~w4270;
assign w4272 = ~w4219 & ~w4271;
assign w4273 = w4219 & w4271;
assign w4274 = ~w4272 & ~w4273;
assign w4275 = (~w4024 & w3978) | (~w4024 & w24799) | (w3978 & w24799);
assign w4276 = w4274 & ~w4275;
assign w4277 = ~w4274 & w4275;
assign w4278 = ~w4276 & ~w4277;
assign w4279 = ~w4209 & ~w4278;
assign w4280 = w4209 & w4278;
assign w4281 = ~w4279 & ~w4280;
assign w4282 = w4199 & w4281;
assign w4283 = ~w4199 & ~w4281;
assign w4284 = ~w4282 & ~w4283;
assign w4285 = w4198 & ~w4284;
assign w4286 = ~w4198 & w4284;
assign w4287 = ~w4285 & ~w4286;
assign w4288 = (~w4058 & ~w3977) | (~w4058 & w24953) | (~w3977 & w24953);
assign w4289 = ~w4287 & ~w4288;
assign w4290 = w4287 & w4288;
assign w4291 = ~w4289 & ~w4290;
assign w4292 = b[17] & ~w1272;
assign w4293 = b[18] & w1154;
assign w4294 = b[19] & w1156;
assign w4295 = w1150 & ~w1231;
assign w4296 = ~w4292 & ~w4293;
assign w4297 = ~w4294 & w4296;
assign w4298 = ~w4295 & w4297;
assign w4299 = a[20] & ~w4298;
assign w4300 = ~a[20] & w4298;
assign w4301 = ~w4299 & ~w4300;
assign w4302 = w4291 & w4301;
assign w4303 = ~w4291 & ~w4301;
assign w4304 = ~w4302 & ~w4303;
assign w4305 = ~w4304 & w25256;
assign w4306 = (w4304 & w4067) | (w4304 & w24954) | (w4067 & w24954);
assign w4307 = (~w4188 & w4306) | (~w4188 & w25257) | (w4306 & w25257);
assign w4308 = ~w4306 & w25258;
assign w4309 = ~w4307 & ~w4308;
assign w4310 = w4178 & ~w4309;
assign w4311 = ~w4178 & w4309;
assign w4312 = ~w4310 & ~w4311;
assign w4313 = b[24] & w573;
assign w4314 = b[23] & ~w649;
assign w4315 = b[25] & w575;
assign w4316 = w569 & w2061;
assign w4317 = ~w4313 & ~w4314;
assign w4318 = ~w4315 & w4317;
assign w4319 = ~w4316 & w4318;
assign w4320 = a[14] & ~w4319;
assign w4321 = ~a[14] & w4319;
assign w4322 = ~w4320 & ~w4321;
assign w4323 = ~w4312 & ~w4322;
assign w4324 = w4312 & w4322;
assign w4325 = ~w4323 & ~w4324;
assign w4326 = ~w4177 & w4325;
assign w4327 = w4177 & ~w4325;
assign w4328 = ~w4326 & ~w4327;
assign w4329 = ~w4176 & ~w4328;
assign w4330 = w4176 & w4328;
assign w4331 = ~w4329 & ~w4330;
assign w4332 = (~w4103 & ~w3954) | (~w4103 & w25118) | (~w3954 & w25118);
assign w4333 = w4331 & w4332;
assign w4334 = ~w4331 & ~w4332;
assign w4335 = ~w4333 & ~w4334;
assign w4336 = ~w4166 & ~w4335;
assign w4337 = w4166 & w4335;
assign w4338 = ~w4336 & ~w4337;
assign w4339 = ~w4156 & ~w4338;
assign w4340 = w4156 & w4338;
assign w4341 = ~w4339 & ~w4340;
assign w4342 = w4155 & ~w4341;
assign w4343 = ~w4155 & w4341;
assign w4344 = ~w4342 & ~w4343;
assign w4345 = (~w4116 & ~w3933) | (~w4116 & w24371) | (~w3933 & w24371);
assign w4346 = ~w4344 & ~w4345;
assign w4347 = w4344 & w4345;
assign w4348 = ~w4346 & ~w4347;
assign w4349 = b[37] & w11;
assign w4350 = b[36] & w9;
assign w4351 = ~b[36] & ~b[37];
assign w4352 = b[36] & b[37];
assign w4353 = ~w4351 & ~w4352;
assign w4354 = (~w4125 & w4123) | (~w4125 & w24955) | (w4123 & w24955);
assign w4355 = ~w4353 & ~w4354;
assign w4356 = w4353 & w4354;
assign w4357 = ~w4355 & ~w4356;
assign w4358 = w5 & ~w4357;
assign w4359 = ~w4349 & ~w4350;
assign w4360 = ~w4358 & w4359;
assign w4361 = b[35] & w24;
assign w4362 = a[2] & ~w4361;
assign w4363 = w4360 & ~w4362;
assign w4364 = a[2] & ~w4360;
assign w4365 = ~w4363 & ~w4364;
assign w4366 = ~w4348 & ~w4365;
assign w4367 = w4348 & w4365;
assign w4368 = ~w4366 & ~w4367;
assign w4369 = w4145 & ~w4368;
assign w4370 = ~w4145 & w4368;
assign w4371 = ~w4369 & ~w4370;
assign w4372 = (~w4342 & ~w4345) | (~w4342 & w24800) | (~w4345 & w24800);
assign w4373 = b[33] & w103;
assign w4374 = b[35] & w68;
assign w4375 = b[34] & w61;
assign w4376 = w66 & w3918;
assign w4377 = ~w4374 & ~w4375;
assign w4378 = ~w4373 & w4377;
assign w4379 = ~w4376 & w4378;
assign w4380 = a[5] & ~w4379;
assign w4381 = ~a[5] & w4379;
assign w4382 = ~w4380 & ~w4381;
assign w4383 = b[31] & w183;
assign w4384 = b[30] & ~w237;
assign w4385 = b[32] & w185;
assign w4386 = w179 & w3304;
assign w4387 = ~w4383 & ~w4384;
assign w4388 = ~w4385 & w4387;
assign w4389 = ~w4386 & w4388;
assign w4390 = a[8] & ~w4389;
assign w4391 = ~a[8] & w4389;
assign w4392 = ~w4390 & ~w4391;
assign w4393 = ~w4330 & ~w4333;
assign w4394 = b[27] & ~w419;
assign w4395 = b[28] & w358;
assign w4396 = b[29] & w360;
assign w4397 = w354 & w2734;
assign w4398 = ~w4394 & ~w4395;
assign w4399 = ~w4396 & w4398;
assign w4400 = ~w4397 & w4399;
assign w4401 = a[11] & ~w4400;
assign w4402 = ~a[11] & w4400;
assign w4403 = ~w4401 & ~w4402;
assign w4404 = b[25] & w573;
assign w4405 = b[26] & w575;
assign w4406 = b[24] & ~w649;
assign w4407 = w569 & w2219;
assign w4408 = ~w4404 & ~w4405;
assign w4409 = ~w4406 & w4408;
assign w4410 = ~w4407 & w4409;
assign w4411 = a[14] & ~w4410;
assign w4412 = ~a[14] & w4410;
assign w4413 = ~w4411 & ~w4412;
assign w4414 = (~w4308 & w4178) | (~w4308 & w24956) | (w4178 & w24956);
assign w4415 = b[19] & w1154;
assign w4416 = b[20] & w1156;
assign w4417 = b[18] & ~w1272;
assign w4418 = w1150 & w1347;
assign w4419 = ~w4415 & ~w4416;
assign w4420 = ~w4417 & w4419;
assign w4421 = ~w4418 & w4420;
assign w4422 = a[20] & ~w4421;
assign w4423 = ~a[20] & w4421;
assign w4424 = ~w4422 & ~w4423;
assign w4425 = (~w4285 & ~w4288) | (~w4285 & w25119) | (~w4288 & w25119);
assign w4426 = b[12] & ~w2114;
assign w4427 = b[13] & w1955;
assign w4428 = b[14] & w1957;
assign w4429 = w714 & w1951;
assign w4430 = ~w4426 & ~w4427;
assign w4431 = ~w4428 & w4430;
assign w4432 = ~w4429 & w4431;
assign w4433 = a[26] & ~w4432;
assign w4434 = ~a[26] & w4432;
assign w4435 = ~w4433 & ~w4434;
assign w4436 = ~w4273 & ~w4276;
assign w4437 = (~w4251 & ~w4252) | (~w4251 & w24801) | (~w4252 & w24801);
assign w4438 = w3784 & w24957;
assign w4439 = b[5] & w3580;
assign w4440 = b[4] & w3578;
assign w4441 = w116 & w3573;
assign w4442 = ~w4439 & ~w4440;
assign w4443 = (a[35] & w4441) | (a[35] & w24802) | (w4441 & w24802);
assign w4444 = ~w4441 & w24803;
assign w4445 = ~w4443 & ~w4444;
assign w4446 = (a[38] & w3989) | (a[38] & w24958) | (w3989 & w24958);
assign w4447 = w4245 & w24804;
assign w4448 = a[38] & ~w4447;
assign w4449 = b[2] & w4243;
assign w4450 = b[1] & w4241;
assign w4451 = w22 & w4236;
assign w4452 = w3989 & ~w4235;
assign w4453 = w4240 & w4452;
assign w4454 = b[0] & w4453;
assign w4455 = ~w4449 & ~w4450;
assign w4456 = ~w4451 & w4455;
assign w4457 = ~w4454 & w4456;
assign w4458 = ~w4448 & w4457;
assign w4459 = w4448 & ~w4457;
assign w4460 = ~w4458 & ~w4459;
assign w4461 = w4445 & w4460;
assign w4462 = ~w4445 & ~w4460;
assign w4463 = ~w4461 & ~w4462;
assign w4464 = ~w4437 & w4463;
assign w4465 = w4437 & ~w4463;
assign w4466 = ~w4464 & ~w4465;
assign w4467 = b[6] & w3177;
assign w4468 = b[7] & w2973;
assign w4469 = b[8] & w2978;
assign w4470 = w270 & w2980;
assign w4471 = ~w4468 & ~w4469;
assign w4472 = ~w4467 & w4471;
assign w4473 = ~w4470 & w4472;
assign w4474 = a[32] & ~w4473;
assign w4475 = ~a[32] & w4473;
assign w4476 = ~w4474 & ~w4475;
assign w4477 = w4466 & w4476;
assign w4478 = ~w4466 & ~w4476;
assign w4479 = ~w4477 & ~w4478;
assign w4480 = ~w4267 & ~w4270;
assign w4481 = ~w4479 & w4480;
assign w4482 = w4479 & ~w4480;
assign w4483 = ~w4481 & ~w4482;
assign w4484 = b[10] & w2436;
assign w4485 = b[9] & ~w2622;
assign w4486 = b[11] & w2438;
assign w4487 = w469 & w2432;
assign w4488 = ~w4484 & ~w4485;
assign w4489 = ~w4486 & w4488;
assign w4490 = ~w4487 & w4489;
assign w4491 = a[29] & ~w4490;
assign w4492 = ~a[29] & w4490;
assign w4493 = ~w4491 & ~w4492;
assign w4494 = ~w4483 & ~w4493;
assign w4495 = w4483 & w4493;
assign w4496 = ~w4494 & ~w4495;
assign w4497 = w4436 & ~w4496;
assign w4498 = ~w4436 & w4496;
assign w4499 = ~w4497 & ~w4498;
assign w4500 = ~w4435 & ~w4499;
assign w4501 = w4435 & w4499;
assign w4502 = ~w4500 & ~w4501;
assign w4503 = (~w4279 & ~w4199) | (~w4279 & w24959) | (~w4199 & w24959);
assign w4504 = w4502 & w4503;
assign w4505 = ~w4502 & ~w4503;
assign w4506 = ~w4504 & ~w4505;
assign w4507 = b[16] & w1517;
assign w4508 = b[15] & ~w1676;
assign w4509 = b[17] & w1519;
assign w4510 = w1008 & w1513;
assign w4511 = ~w4507 & ~w4508;
assign w4512 = ~w4509 & w4511;
assign w4513 = ~w4510 & w4512;
assign w4514 = a[23] & ~w4513;
assign w4515 = ~a[23] & w4513;
assign w4516 = ~w4514 & ~w4515;
assign w4517 = w4506 & w4516;
assign w4518 = ~w4506 & ~w4516;
assign w4519 = ~w4517 & ~w4518;
assign w4520 = ~w4425 & ~w4519;
assign w4521 = w4425 & w4519;
assign w4522 = ~w4520 & ~w4521;
assign w4523 = w4424 & ~w4522;
assign w4524 = ~w4424 & w4522;
assign w4525 = ~w4523 & ~w4524;
assign w4526 = ~w4302 & ~w4306;
assign w4527 = ~w4525 & w4526;
assign w4528 = w4525 & ~w4526;
assign w4529 = ~w4527 & ~w4528;
assign w4530 = b[22] & w838;
assign w4531 = b[23] & w834;
assign w4532 = b[21] & ~w934;
assign w4533 = ~w4530 & ~w4531;
assign w4534 = ~w4532 & w4533;
assign w4535 = w826 & w1755;
assign w4536 = ~a[17] & ~w4535;
assign w4537 = ~a[16] & w4535;
assign w4538 = ~w4536 & ~w4537;
assign w4539 = w4534 & ~w4538;
assign w4540 = a[17] & ~w4534;
assign w4541 = ~w4539 & ~w4540;
assign w4542 = ~w4529 & ~w4541;
assign w4543 = w4529 & w4541;
assign w4544 = ~w4542 & ~w4543;
assign w4545 = w4414 & w4544;
assign w4546 = ~w4414 & ~w4544;
assign w4547 = ~w4545 & ~w4546;
assign w4548 = ~w4413 & w4547;
assign w4549 = w4413 & ~w4547;
assign w4550 = ~w4548 & ~w4549;
assign w4551 = ~w4324 & ~w4326;
assign w4552 = w4550 & ~w4551;
assign w4553 = ~w4550 & w4551;
assign w4554 = ~w4552 & ~w4553;
assign w4555 = ~w4403 & ~w4554;
assign w4556 = w4403 & w4554;
assign w4557 = ~w4555 & ~w4556;
assign w4558 = w4393 & w4557;
assign w4559 = ~w4393 & ~w4557;
assign w4560 = ~w4558 & ~w4559;
assign w4561 = ~w4392 & w4560;
assign w4562 = w4392 & ~w4560;
assign w4563 = ~w4561 & ~w4562;
assign w4564 = (~w4336 & ~w4156) | (~w4336 & w25120) | (~w4156 & w25120);
assign w4565 = w4563 & w4564;
assign w4566 = ~w4563 & ~w4564;
assign w4567 = ~w4565 & ~w4566;
assign w4568 = ~w4382 & ~w4567;
assign w4569 = w4382 & w4567;
assign w4570 = ~w4568 & ~w4569;
assign w4571 = w4372 & w4570;
assign w4572 = ~w4372 & ~w4570;
assign w4573 = ~w4571 & ~w4572;
assign w4574 = b[38] & w11;
assign w4575 = b[37] & w9;
assign w4576 = ~b[37] & ~b[38];
assign w4577 = b[37] & b[38];
assign w4578 = ~w4576 & ~w4577;
assign w4579 = ~w4351 & ~w4356;
assign w4580 = w4578 & w4579;
assign w4581 = ~w4578 & ~w4579;
assign w4582 = ~w4580 & ~w4581;
assign w4583 = w5 & w4582;
assign w4584 = ~w4574 & ~w4575;
assign w4585 = ~w4583 & w4584;
assign w4586 = b[36] & w24;
assign w4587 = a[2] & ~w4586;
assign w4588 = w4585 & ~w4587;
assign w4589 = a[2] & ~w4585;
assign w4590 = ~w4588 & ~w4589;
assign w4591 = ~w4573 & w4590;
assign w4592 = w4573 & ~w4590;
assign w4593 = ~w4591 & ~w4592;
assign w4594 = (~w4367 & w4145) | (~w4367 & w24372) | (w4145 & w24372);
assign w4595 = w4593 & ~w4594;
assign w4596 = ~w4593 & w4594;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = b[34] & w103;
assign w4599 = b[36] & w68;
assign w4600 = b[35] & w61;
assign w4601 = w66 & w4129;
assign w4602 = ~w4599 & ~w4600;
assign w4603 = ~w4598 & w4602;
assign w4604 = ~w4601 & w4603;
assign w4605 = a[5] & ~w4604;
assign w4606 = ~a[5] & w4604;
assign w4607 = ~w4605 & ~w4606;
assign w4608 = ~w4562 & ~w4565;
assign w4609 = (~w4549 & w4551) | (~w4549 & w24960) | (w4551 & w24960);
assign w4610 = b[25] & ~w649;
assign w4611 = b[27] & w575;
assign w4612 = b[26] & w573;
assign w4613 = w569 & w2378;
assign w4614 = ~w4610 & ~w4611;
assign w4615 = ~w4612 & w4614;
assign w4616 = ~w4613 & w4615;
assign w4617 = a[14] & ~w4616;
assign w4618 = ~a[14] & w4616;
assign w4619 = ~w4617 & ~w4618;
assign w4620 = (~w4542 & ~w4414) | (~w4542 & w25121) | (~w4414 & w25121);
assign w4621 = b[22] & ~w934;
assign w4622 = b[23] & w838;
assign w4623 = b[24] & w834;
assign w4624 = w832 & w1895;
assign w4625 = ~w4621 & ~w4622;
assign w4626 = ~w4623 & w4625;
assign w4627 = ~w4624 & w4626;
assign w4628 = a[17] & ~w4627;
assign w4629 = ~a[17] & w4627;
assign w4630 = ~w4628 & ~w4629;
assign w4631 = (~w4523 & w4526) | (~w4523 & w24373) | (w4526 & w24373);
assign w4632 = b[17] & w1517;
assign w4633 = b[16] & ~w1676;
assign w4634 = b[18] & w1519;
assign w4635 = ~w1108 & w1513;
assign w4636 = ~w4632 & ~w4633;
assign w4637 = ~w4634 & w4636;
assign w4638 = ~w4635 & w4637;
assign w4639 = a[23] & ~w4638;
assign w4640 = ~a[23] & w4638;
assign w4641 = ~w4639 & ~w4640;
assign w4642 = ~w4501 & ~w4504;
assign w4643 = a[38] & ~a[39];
assign w4644 = ~a[38] & a[39];
assign w4645 = ~w4643 & ~w4644;
assign w4646 = b[0] & ~w4645;
assign w4647 = w4447 & w4457;
assign w4648 = w4452 & w24646;
assign w4649 = b[2] & w4241;
assign w4650 = b[3] & w4243;
assign w4651 = ~w4649 & ~w4650;
assign w4652 = ~w4648 & w4651;
assign w4653 = (a[38] & ~w4652) | (a[38] & w24647) | (~w4652 & w24647);
assign w4654 = w4652 & w24648;
assign w4655 = ~w4653 & ~w4654;
assign w4656 = w4647 & w4655;
assign w4657 = ~w4647 & ~w4655;
assign w4658 = ~w4656 & ~w4657;
assign w4659 = w4646 & w4658;
assign w4660 = ~w4646 & ~w4658;
assign w4661 = ~w4659 & ~w4660;
assign w4662 = b[4] & w3785;
assign w4663 = b[5] & w3578;
assign w4664 = b[6] & w3580;
assign w4665 = w157 & w3573;
assign w4666 = ~w4663 & ~w4664;
assign w4667 = ~w4662 & w4666;
assign w4668 = ~w4665 & w4667;
assign w4669 = a[35] & ~w4668;
assign w4670 = ~a[35] & w4668;
assign w4671 = ~w4669 & ~w4670;
assign w4672 = w4661 & w4671;
assign w4673 = ~w4661 & ~w4671;
assign w4674 = ~w4672 & ~w4673;
assign w4675 = (~w4461 & w4437) | (~w4461 & w24649) | (w4437 & w24649);
assign w4676 = ~w4674 & w4675;
assign w4677 = w4674 & ~w4675;
assign w4678 = ~w4676 & ~w4677;
assign w4679 = b[7] & w3177;
assign w4680 = b[8] & w2973;
assign w4681 = b[9] & w2978;
assign w4682 = w322 & w2980;
assign w4683 = ~w4680 & ~w4681;
assign w4684 = ~w4679 & w4683;
assign w4685 = ~w4682 & w4684;
assign w4686 = a[32] & ~w4685;
assign w4687 = ~a[32] & w4685;
assign w4688 = ~w4686 & ~w4687;
assign w4689 = w4678 & w4688;
assign w4690 = ~w4678 & ~w4688;
assign w4691 = ~w4689 & ~w4690;
assign w4692 = (~w4477 & w4480) | (~w4477 & w24650) | (w4480 & w24650);
assign w4693 = w4691 & ~w4692;
assign w4694 = ~w4691 & w4692;
assign w4695 = ~w4693 & ~w4694;
assign w4696 = b[12] & w2438;
assign w4697 = b[10] & ~w2622;
assign w4698 = b[11] & w2436;
assign w4699 = w536 & w2432;
assign w4700 = ~w4696 & ~w4697;
assign w4701 = ~w4698 & w4700;
assign w4702 = ~w4699 & w4701;
assign w4703 = a[29] & ~w4702;
assign w4704 = ~a[29] & w4702;
assign w4705 = ~w4703 & ~w4704;
assign w4706 = ~w4695 & ~w4705;
assign w4707 = w4695 & w4705;
assign w4708 = ~w4706 & ~w4707;
assign w4709 = ~w4495 & ~w4498;
assign w4710 = w4708 & ~w4709;
assign w4711 = ~w4708 & w4709;
assign w4712 = ~w4710 & ~w4711;
assign w4713 = b[13] & ~w2114;
assign w4714 = b[15] & w1957;
assign w4715 = b[14] & w1955;
assign w4716 = ~w799 & w1951;
assign w4717 = ~w4713 & ~w4714;
assign w4718 = ~w4715 & w4717;
assign w4719 = ~w4716 & w4718;
assign w4720 = a[26] & ~w4719;
assign w4721 = ~a[26] & w4719;
assign w4722 = ~w4720 & ~w4721;
assign w4723 = w4712 & w4722;
assign w4724 = ~w4712 & ~w4722;
assign w4725 = ~w4723 & ~w4724;
assign w4726 = w4642 & w4725;
assign w4727 = ~w4642 & ~w4725;
assign w4728 = ~w4726 & ~w4727;
assign w4729 = w4641 & ~w4728;
assign w4730 = ~w4641 & w4728;
assign w4731 = ~w4729 & ~w4730;
assign w4732 = (~w4518 & ~w4425) | (~w4518 & w24651) | (~w4425 & w24651);
assign w4733 = ~w4731 & ~w4732;
assign w4734 = w4731 & w4732;
assign w4735 = ~w4733 & ~w4734;
assign w4736 = b[20] & w1154;
assign w4737 = b[19] & ~w1272;
assign w4738 = b[21] & w1156;
assign w4739 = w1150 & w1467;
assign w4740 = ~w4736 & ~w4737;
assign w4741 = ~w4738 & w4740;
assign w4742 = ~w4739 & w4741;
assign w4743 = a[20] & ~w4742;
assign w4744 = ~a[20] & w4742;
assign w4745 = ~w4743 & ~w4744;
assign w4746 = w4735 & w4745;
assign w4747 = ~w4735 & ~w4745;
assign w4748 = ~w4746 & ~w4747;
assign w4749 = ~w4631 & ~w4748;
assign w4750 = w4631 & w4748;
assign w4751 = ~w4749 & ~w4750;
assign w4752 = ~w4630 & w4751;
assign w4753 = w4630 & ~w4751;
assign w4754 = ~w4752 & ~w4753;
assign w4755 = w4620 & w4754;
assign w4756 = ~w4620 & ~w4754;
assign w4757 = ~w4755 & ~w4756;
assign w4758 = w4619 & w4757;
assign w4759 = ~w4619 & ~w4757;
assign w4760 = ~w4758 & ~w4759;
assign w4761 = ~w4609 & w4760;
assign w4762 = w4609 & ~w4760;
assign w4763 = ~w4761 & ~w4762;
assign w4764 = b[29] & w358;
assign w4765 = b[30] & w360;
assign w4766 = b[28] & ~w419;
assign w4767 = w354 & ~w2908;
assign w4768 = ~w4764 & ~w4765;
assign w4769 = ~w4766 & w4768;
assign w4770 = ~w4767 & w4769;
assign w4771 = a[11] & ~w4770;
assign w4772 = ~a[11] & w4770;
assign w4773 = ~w4771 & ~w4772;
assign w4774 = w4763 & w4773;
assign w4775 = ~w4763 & ~w4773;
assign w4776 = ~w4774 & ~w4775;
assign w4777 = ~w4555 & ~w4558;
assign w4778 = w4776 & w4777;
assign w4779 = ~w4776 & ~w4777;
assign w4780 = ~w4778 & ~w4779;
assign w4781 = b[33] & w185;
assign w4782 = b[31] & ~w237;
assign w4783 = b[32] & w183;
assign w4784 = w179 & w3499;
assign w4785 = ~w4781 & ~w4782;
assign w4786 = ~w4783 & w4785;
assign w4787 = ~w4784 & w4786;
assign w4788 = a[8] & ~w4787;
assign w4789 = ~a[8] & w4787;
assign w4790 = ~w4788 & ~w4789;
assign w4791 = w4780 & w4790;
assign w4792 = ~w4780 & ~w4790;
assign w4793 = ~w4791 & ~w4792;
assign w4794 = w4608 & w4793;
assign w4795 = ~w4608 & ~w4793;
assign w4796 = ~w4794 & ~w4795;
assign w4797 = ~w4607 & w4796;
assign w4798 = w4607 & ~w4796;
assign w4799 = ~w4797 & ~w4798;
assign w4800 = (~w4568 & ~w4372) | (~w4568 & w25122) | (~w4372 & w25122);
assign w4801 = w4799 & w4800;
assign w4802 = ~w4799 & ~w4800;
assign w4803 = ~w4801 & ~w4802;
assign w4804 = b[39] & w11;
assign w4805 = b[38] & w9;
assign w4806 = (~w4577 & ~w4579) | (~w4577 & w24652) | (~w4579 & w24652);
assign w4807 = ~b[38] & ~b[39];
assign w4808 = b[38] & b[39];
assign w4809 = ~w4807 & ~w4808;
assign w4810 = ~w4806 & ~w4809;
assign w4811 = w4806 & w4809;
assign w4812 = ~w4810 & ~w4811;
assign w4813 = w5 & ~w4812;
assign w4814 = ~w4804 & ~w4805;
assign w4815 = ~w4813 & w4814;
assign w4816 = b[37] & w24;
assign w4817 = a[2] & ~w4816;
assign w4818 = w4815 & ~w4817;
assign w4819 = a[2] & ~w4815;
assign w4820 = ~w4818 & ~w4819;
assign w4821 = w4803 & w4820;
assign w4822 = ~w4803 & ~w4820;
assign w4823 = ~w4821 & ~w4822;
assign w4824 = (~w4591 & w4594) | (~w4591 & w24805) | (w4594 & w24805);
assign w4825 = w4823 & w4824;
assign w4826 = ~w4823 & ~w4824;
assign w4827 = ~w4825 & ~w4826;
assign w4828 = ~w4798 & ~w4801;
assign w4829 = b[33] & w183;
assign w4830 = b[34] & w185;
assign w4831 = b[32] & ~w237;
assign w4832 = w179 & ~w3710;
assign w4833 = ~w4829 & ~w4830;
assign w4834 = ~w4831 & w4833;
assign w4835 = ~w4832 & w4834;
assign w4836 = a[8] & ~w4835;
assign w4837 = ~a[8] & w4835;
assign w4838 = ~w4836 & ~w4837;
assign w4839 = (~w4774 & ~w4777) | (~w4774 & w24961) | (~w4777 & w24961);
assign w4840 = b[29] & ~w419;
assign w4841 = b[30] & w358;
assign w4842 = b[31] & w360;
assign w4843 = w354 & ~w3112;
assign w4844 = ~w4840 & ~w4841;
assign w4845 = ~w4842 & w4844;
assign w4846 = ~w4843 & w4845;
assign w4847 = a[11] & ~w4846;
assign w4848 = ~a[11] & w4846;
assign w4849 = ~w4847 & ~w4848;
assign w4850 = (~w4758 & w4609) | (~w4758 & w25123) | (w4609 & w25123);
assign w4851 = b[28] & w575;
assign w4852 = b[26] & ~w649;
assign w4853 = b[27] & w573;
assign w4854 = w569 & w2559;
assign w4855 = ~w4851 & ~w4852;
assign w4856 = ~w4853 & w4855;
assign w4857 = ~w4854 & w4856;
assign w4858 = a[14] & ~w4857;
assign w4859 = ~a[14] & w4857;
assign w4860 = ~w4858 & ~w4859;
assign w4861 = (~w4753 & ~w4620) | (~w4753 & w24374) | (~w4620 & w24374);
assign w4862 = b[22] & w1156;
assign w4863 = b[21] & w1154;
assign w4864 = b[20] & ~w1272;
assign w4865 = w1150 & w1615;
assign w4866 = ~w4862 & ~w4863;
assign w4867 = ~w4864 & w4866;
assign w4868 = ~w4865 & w4867;
assign w4869 = a[20] & ~w4868;
assign w4870 = ~a[20] & w4868;
assign w4871 = ~w4869 & ~w4870;
assign w4872 = b[18] & w1517;
assign w4873 = b[17] & ~w1676;
assign w4874 = b[19] & w1519;
assign w4875 = ~w1231 & w1513;
assign w4876 = ~w4872 & ~w4873;
assign w4877 = ~w4874 & w4876;
assign w4878 = ~w4875 & w4877;
assign w4879 = a[23] & ~w4878;
assign w4880 = ~a[23] & w4878;
assign w4881 = ~w4879 & ~w4880;
assign w4882 = (~w4707 & w4709) | (~w4707 & w24653) | (w4709 & w24653);
assign w4883 = b[11] & ~w2622;
assign w4884 = b[12] & w2436;
assign w4885 = b[13] & w2438;
assign w4886 = w628 & w2432;
assign w4887 = ~w4883 & ~w4884;
assign w4888 = ~w4885 & w4887;
assign w4889 = ~w4886 & w4888;
assign w4890 = a[29] & ~w4889;
assign w4891 = ~a[29] & w4889;
assign w4892 = ~w4890 & ~w4891;
assign w4893 = ~w4689 & ~w4693;
assign w4894 = b[8] & w3177;
assign w4895 = b[9] & w2973;
assign w4896 = b[10] & w2978;
assign w4897 = w397 & w2980;
assign w4898 = ~w4895 & ~w4896;
assign w4899 = ~w4894 & w4898;
assign w4900 = ~w4897 & w4899;
assign w4901 = a[32] & ~w4900;
assign w4902 = ~a[32] & w4900;
assign w4903 = ~w4901 & ~w4902;
assign w4904 = w4452 & w24806;
assign w4905 = b[3] & w4241;
assign w4906 = b[4] & w4243;
assign w4907 = w84 & w4236;
assign w4908 = ~w4905 & ~w4906;
assign w4909 = ~w4904 & w4908;
assign w4910 = ~w4907 & w4909;
assign w4911 = a[38] & ~w4910;
assign w4912 = ~a[38] & w4910;
assign w4913 = ~w4911 & ~w4912;
assign w4914 = a[41] & w4646;
assign w4915 = a[39] & ~a[40];
assign w4916 = ~a[39] & a[40];
assign w4917 = ~w4915 & ~w4916;
assign w4918 = w4645 & ~w4917;
assign w4919 = b[0] & w4918;
assign w4920 = a[40] & ~a[41];
assign w4921 = ~a[40] & a[41];
assign w4922 = ~w4920 & ~w4921;
assign w4923 = ~w4645 & ~w4922;
assign w4924 = ~w8 & w4923;
assign w4925 = ~w4645 & w4922;
assign w4926 = b[1] & w4925;
assign w4927 = ~w4919 & ~w4924;
assign w4928 = ~w4926 & w4927;
assign w4929 = w4914 & ~w4928;
assign w4930 = ~w4914 & w4928;
assign w4931 = ~w4929 & ~w4930;
assign w4932 = ~w4913 & ~w4931;
assign w4933 = w4913 & w4931;
assign w4934 = ~w4932 & ~w4933;
assign w4935 = (~w4656 & ~w4658) | (~w4656 & w24654) | (~w4658 & w24654);
assign w4936 = w4934 & ~w4935;
assign w4937 = ~w4934 & w4935;
assign w4938 = ~w4936 & ~w4937;
assign w4939 = b[5] & w3785;
assign w4940 = b[6] & w3578;
assign w4941 = b[7] & w3580;
assign w4942 = w216 & w3573;
assign w4943 = ~w4940 & ~w4941;
assign w4944 = ~w4939 & w4943;
assign w4945 = ~w4942 & w4944;
assign w4946 = a[35] & ~w4945;
assign w4947 = ~a[35] & w4945;
assign w4948 = ~w4946 & ~w4947;
assign w4949 = w4938 & w4948;
assign w4950 = ~w4938 & ~w4948;
assign w4951 = ~w4949 & ~w4950;
assign w4952 = (~w4672 & ~w4674) | (~w4672 & w24807) | (~w4674 & w24807);
assign w4953 = w4951 & w4952;
assign w4954 = ~w4951 & ~w4952;
assign w4955 = ~w4953 & ~w4954;
assign w4956 = w4903 & ~w4955;
assign w4957 = ~w4903 & w4955;
assign w4958 = ~w4956 & ~w4957;
assign w4959 = ~w4893 & w4958;
assign w4960 = w4893 & ~w4958;
assign w4961 = ~w4959 & ~w4960;
assign w4962 = w4892 & w4961;
assign w4963 = ~w4892 & ~w4961;
assign w4964 = ~w4962 & ~w4963;
assign w4965 = ~w4882 & w4964;
assign w4966 = w4882 & ~w4964;
assign w4967 = ~w4965 & ~w4966;
assign w4968 = b[14] & ~w2114;
assign w4969 = b[16] & w1957;
assign w4970 = b[15] & w1955;
assign w4971 = w905 & w1951;
assign w4972 = ~w4968 & ~w4969;
assign w4973 = ~w4970 & w4972;
assign w4974 = ~w4971 & w4973;
assign w4975 = a[26] & ~w4974;
assign w4976 = ~a[26] & w4974;
assign w4977 = ~w4975 & ~w4976;
assign w4978 = w4967 & w4977;
assign w4979 = ~w4967 & ~w4977;
assign w4980 = ~w4978 & ~w4979;
assign w4981 = (~w4724 & ~w4642) | (~w4724 & w24655) | (~w4642 & w24655);
assign w4982 = w4980 & w4981;
assign w4983 = ~w4980 & ~w4981;
assign w4984 = ~w4982 & ~w4983;
assign w4985 = w4881 & w4984;
assign w4986 = ~w4881 & ~w4984;
assign w4987 = ~w4985 & ~w4986;
assign w4988 = ~w4729 & ~w4734;
assign w4989 = w4987 & w4988;
assign w4990 = ~w4987 & ~w4988;
assign w4991 = ~w4989 & ~w4990;
assign w4992 = w4871 & ~w4991;
assign w4993 = ~w4871 & w4991;
assign w4994 = ~w4992 & ~w4993;
assign w4995 = (~w4747 & ~w4631) | (~w4747 & w24656) | (~w4631 & w24656);
assign w4996 = ~w4994 & ~w4995;
assign w4997 = w4994 & w4995;
assign w4998 = ~w4996 & ~w4997;
assign w4999 = b[25] & w834;
assign w5000 = b[23] & ~w934;
assign w5001 = b[24] & w838;
assign w5002 = w832 & w2061;
assign w5003 = ~w4999 & ~w5000;
assign w5004 = ~w5001 & w5003;
assign w5005 = ~w5002 & w5004;
assign w5006 = a[17] & ~w5005;
assign w5007 = ~a[17] & w5005;
assign w5008 = ~w5006 & ~w5007;
assign w5009 = w4998 & w5008;
assign w5010 = ~w4998 & ~w5008;
assign w5011 = ~w5009 & ~w5010;
assign w5012 = w4861 & w5011;
assign w5013 = ~w4861 & ~w5011;
assign w5014 = ~w5012 & ~w5013;
assign w5015 = ~w4860 & w5014;
assign w5016 = w4860 & ~w5014;
assign w5017 = ~w5015 & ~w5016;
assign w5018 = ~w4850 & w5017;
assign w5019 = w4850 & ~w5017;
assign w5020 = ~w5018 & ~w5019;
assign w5021 = ~w4849 & ~w5020;
assign w5022 = w4849 & w5020;
assign w5023 = ~w5021 & ~w5022;
assign w5024 = ~w4839 & ~w5023;
assign w5025 = w4839 & w5023;
assign w5026 = ~w5024 & ~w5025;
assign w5027 = ~w4838 & w5026;
assign w5028 = w4838 & ~w5026;
assign w5029 = ~w5027 & ~w5028;
assign w5030 = ~w4792 & ~w4794;
assign w5031 = w5029 & w5030;
assign w5032 = ~w5029 & ~w5030;
assign w5033 = ~w5031 & ~w5032;
assign w5034 = b[35] & w103;
assign w5035 = b[37] & w68;
assign w5036 = b[36] & w61;
assign w5037 = w66 & ~w4357;
assign w5038 = ~w5035 & ~w5036;
assign w5039 = ~w5034 & w5038;
assign w5040 = ~w5037 & w5039;
assign w5041 = a[5] & ~w5040;
assign w5042 = ~a[5] & w5040;
assign w5043 = ~w5041 & ~w5042;
assign w5044 = w5033 & w5043;
assign w5045 = ~w5033 & ~w5043;
assign w5046 = ~w5044 & ~w5045;
assign w5047 = ~w4828 & ~w5046;
assign w5048 = w4828 & w5046;
assign w5049 = ~w5047 & ~w5048;
assign w5050 = b[40] & w11;
assign w5051 = b[39] & w9;
assign w5052 = ~b[39] & ~b[40];
assign w5053 = b[39] & b[40];
assign w5054 = ~w5052 & ~w5053;
assign w5055 = ~w4807 & ~w4811;
assign w5056 = w5054 & ~w5055;
assign w5057 = ~w5054 & w5055;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = w5 & ~w5058;
assign w5060 = ~w5050 & ~w5051;
assign w5061 = ~w5059 & w5060;
assign w5062 = b[38] & w24;
assign w5063 = a[2] & ~w5062;
assign w5064 = w5061 & ~w5063;
assign w5065 = a[2] & ~w5061;
assign w5066 = ~w5064 & ~w5065;
assign w5067 = ~w5049 & w5066;
assign w5068 = w5049 & ~w5066;
assign w5069 = ~w5067 & ~w5068;
assign w5070 = (~w4822 & ~w4824) | (~w4822 & w25124) | (~w4824 & w25124);
assign w5071 = w5069 & w5070;
assign w5072 = ~w5069 & ~w5070;
assign w5073 = ~w5071 & ~w5072;
assign w5074 = ~w5067 & ~w5071;
assign w5075 = b[36] & w103;
assign w5076 = b[37] & w61;
assign w5077 = b[38] & w68;
assign w5078 = w66 & w4582;
assign w5079 = ~w5076 & ~w5077;
assign w5080 = ~w5075 & w5079;
assign w5081 = ~w5078 & w5080;
assign w5082 = a[5] & ~w5081;
assign w5083 = ~a[5] & w5081;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = (~w5028 & ~w5030) | (~w5028 & w24962) | (~w5030 & w24962);
assign w5086 = b[30] & ~w419;
assign w5087 = b[32] & w360;
assign w5088 = b[31] & w358;
assign w5089 = w354 & w3304;
assign w5090 = ~w5086 & ~w5087;
assign w5091 = ~w5088 & w5090;
assign w5092 = ~w5089 & w5091;
assign w5093 = a[11] & ~w5092;
assign w5094 = ~a[11] & w5092;
assign w5095 = ~w5093 & ~w5094;
assign w5096 = (~w5016 & w4850) | (~w5016 & w24375) | (w4850 & w24375);
assign w5097 = b[28] & w573;
assign w5098 = b[27] & ~w649;
assign w5099 = b[29] & w575;
assign w5100 = w569 & w2734;
assign w5101 = ~w5097 & ~w5098;
assign w5102 = ~w5099 & w5101;
assign w5103 = ~w5100 & w5102;
assign w5104 = a[14] & ~w5103;
assign w5105 = ~a[14] & w5103;
assign w5106 = ~w5104 & ~w5105;
assign w5107 = b[24] & ~w934;
assign w5108 = b[25] & w838;
assign w5109 = b[26] & w834;
assign w5110 = w832 & w2219;
assign w5111 = ~w5107 & ~w5108;
assign w5112 = ~w5109 & w5111;
assign w5113 = ~w5110 & w5112;
assign w5114 = a[17] & ~w5113;
assign w5115 = ~a[17] & w5113;
assign w5116 = ~w5114 & ~w5115;
assign w5117 = ~w4992 & ~w4997;
assign w5118 = b[20] & w1519;
assign w5119 = b[19] & w1517;
assign w5120 = b[18] & ~w1676;
assign w5121 = w1347 & w1513;
assign w5122 = ~w5118 & ~w5119;
assign w5123 = ~w5120 & w5122;
assign w5124 = ~w5121 & w5123;
assign w5125 = a[23] & ~w5124;
assign w5126 = ~a[23] & w5124;
assign w5127 = ~w5125 & ~w5126;
assign w5128 = (~w4978 & ~w4981) | (~w4978 & w24963) | (~w4981 & w24963);
assign w5129 = b[16] & w1955;
assign w5130 = b[17] & w1957;
assign w5131 = b[15] & ~w2114;
assign w5132 = w1008 & w1951;
assign w5133 = ~w5129 & ~w5130;
assign w5134 = ~w5131 & w5133;
assign w5135 = ~w5132 & w5134;
assign w5136 = a[26] & ~w5135;
assign w5137 = ~a[26] & w5135;
assign w5138 = ~w5136 & ~w5137;
assign w5139 = ~w4962 & ~w4965;
assign w5140 = b[14] & w2438;
assign w5141 = b[12] & ~w2622;
assign w5142 = b[13] & w2436;
assign w5143 = w714 & w2432;
assign w5144 = ~w5140 & ~w5141;
assign w5145 = ~w5142 & w5144;
assign w5146 = ~w5143 & w5145;
assign w5147 = a[29] & ~w5146;
assign w5148 = ~a[29] & w5146;
assign w5149 = ~w5147 & ~w5148;
assign w5150 = (~w4956 & w4893) | (~w4956 & w24964) | (w4893 & w24964);
assign w5151 = ~w4933 & ~w4936;
assign w5152 = w4452 & w25125;
assign w5153 = b[5] & w4243;
assign w5154 = b[4] & w4241;
assign w5155 = w116 & w4236;
assign w5156 = ~w5153 & ~w5154;
assign w5157 = (a[38] & w5155) | (a[38] & w24965) | (w5155 & w24965);
assign w5158 = ~w5155 & w24966;
assign w5159 = ~w5157 & ~w5158;
assign w5160 = (a[41] & w4645) | (a[41] & w25126) | (w4645 & w25126);
assign w5161 = w4927 & w24967;
assign w5162 = a[41] & ~w5161;
assign w5163 = w22 & w4923;
assign w5164 = b[1] & w4918;
assign w5165 = b[2] & w4925;
assign w5166 = w4645 & w4917;
assign w5167 = ~w4922 & w5166;
assign w5168 = b[0] & w5167;
assign w5169 = ~w5163 & ~w5164;
assign w5170 = ~w5165 & w5169;
assign w5171 = ~w5168 & w5170;
assign w5172 = ~w5162 & w5171;
assign w5173 = w5162 & ~w5171;
assign w5174 = ~w5172 & ~w5173;
assign w5175 = w5159 & w5174;
assign w5176 = ~w5159 & ~w5174;
assign w5177 = ~w5175 & ~w5176;
assign w5178 = ~w4936 & w24968;
assign w5179 = (w5177 & w4936) | (w5177 & w24969) | (w4936 & w24969);
assign w5180 = ~w5178 & ~w5179;
assign w5181 = b[6] & w3785;
assign w5182 = b[8] & w3580;
assign w5183 = b[7] & w3578;
assign w5184 = w270 & w3573;
assign w5185 = ~w5182 & ~w5183;
assign w5186 = ~w5181 & w5185;
assign w5187 = ~w5184 & w5186;
assign w5188 = a[35] & ~w5187;
assign w5189 = ~a[35] & w5187;
assign w5190 = ~w5188 & ~w5189;
assign w5191 = ~w5180 & ~w5190;
assign w5192 = w5180 & w5190;
assign w5193 = ~w5191 & ~w5192;
assign w5194 = ~w4950 & ~w4953;
assign w5195 = w5193 & w5194;
assign w5196 = ~w5193 & ~w5194;
assign w5197 = ~w5195 & ~w5196;
assign w5198 = b[9] & w3177;
assign w5199 = b[10] & w2973;
assign w5200 = b[11] & w2978;
assign w5201 = w469 & w2980;
assign w5202 = ~w5199 & ~w5200;
assign w5203 = ~w5198 & w5202;
assign w5204 = ~w5201 & w5203;
assign w5205 = a[32] & ~w5204;
assign w5206 = ~a[32] & w5204;
assign w5207 = ~w5205 & ~w5206;
assign w5208 = ~w5197 & ~w5207;
assign w5209 = w5197 & w5207;
assign w5210 = ~w5208 & ~w5209;
assign w5211 = w5150 & w5210;
assign w5212 = ~w5150 & ~w5210;
assign w5213 = ~w5211 & ~w5212;
assign w5214 = w5149 & ~w5213;
assign w5215 = ~w5149 & w5213;
assign w5216 = ~w5214 & ~w5215;
assign w5217 = ~w5139 & w5216;
assign w5218 = w5139 & ~w5216;
assign w5219 = ~w5217 & ~w5218;
assign w5220 = ~w5138 & ~w5219;
assign w5221 = w5138 & w5219;
assign w5222 = ~w5220 & ~w5221;
assign w5223 = ~w5128 & w5222;
assign w5224 = w5128 & ~w5222;
assign w5225 = ~w5223 & ~w5224;
assign w5226 = w5127 & w5225;
assign w5227 = ~w5127 & ~w5225;
assign w5228 = ~w5226 & ~w5227;
assign w5229 = ~w4986 & ~w4989;
assign w5230 = ~w5228 & ~w5229;
assign w5231 = w5228 & w5229;
assign w5232 = ~w5230 & ~w5231;
assign w5233 = b[21] & ~w1272;
assign w5234 = b[22] & w1154;
assign w5235 = b[23] & w1156;
assign w5236 = ~w5233 & ~w5234;
assign w5237 = ~w5235 & w5236;
assign w5238 = w1144 & w1755;
assign w5239 = ~a[20] & ~w5238;
assign w5240 = ~a[19] & w5238;
assign w5241 = ~w5239 & ~w5240;
assign w5242 = w5237 & ~w5241;
assign w5243 = a[20] & ~w5237;
assign w5244 = ~w5242 & ~w5243;
assign w5245 = ~w5232 & ~w5244;
assign w5246 = w5232 & w5244;
assign w5247 = ~w5245 & ~w5246;
assign w5248 = w5117 & w5247;
assign w5249 = ~w5117 & ~w5247;
assign w5250 = ~w5248 & ~w5249;
assign w5251 = ~w5116 & w5250;
assign w5252 = w5116 & ~w5250;
assign w5253 = ~w5251 & ~w5252;
assign w5254 = (~w5010 & ~w4861) | (~w5010 & w24657) | (~w4861 & w24657);
assign w5255 = w5253 & w5254;
assign w5256 = ~w5253 & ~w5254;
assign w5257 = ~w5255 & ~w5256;
assign w5258 = w5106 & w5257;
assign w5259 = ~w5106 & ~w5257;
assign w5260 = ~w5258 & ~w5259;
assign w5261 = w5096 & ~w5260;
assign w5262 = ~w5096 & w5260;
assign w5263 = ~w5261 & ~w5262;
assign w5264 = ~w5095 & ~w5263;
assign w5265 = w5095 & w5263;
assign w5266 = ~w5264 & ~w5265;
assign w5267 = (~w5021 & ~w4839) | (~w5021 & w25127) | (~w4839 & w25127);
assign w5268 = w5266 & w5267;
assign w5269 = ~w5266 & ~w5267;
assign w5270 = ~w5268 & ~w5269;
assign w5271 = b[35] & w185;
assign w5272 = b[33] & ~w237;
assign w5273 = b[34] & w183;
assign w5274 = w179 & w3918;
assign w5275 = ~w5271 & ~w5272;
assign w5276 = ~w5273 & w5275;
assign w5277 = ~w5274 & w5276;
assign w5278 = a[8] & ~w5277;
assign w5279 = ~a[8] & w5277;
assign w5280 = ~w5278 & ~w5279;
assign w5281 = w5270 & w5280;
assign w5282 = ~w5270 & ~w5280;
assign w5283 = ~w5281 & ~w5282;
assign w5284 = ~w5085 & ~w5283;
assign w5285 = w5085 & w5283;
assign w5286 = ~w5284 & ~w5285;
assign w5287 = w5084 & ~w5286;
assign w5288 = ~w5084 & w5286;
assign w5289 = ~w5287 & ~w5288;
assign w5290 = ~w5045 & ~w5048;
assign w5291 = ~w5289 & ~w5290;
assign w5292 = w5289 & w5290;
assign w5293 = ~w5291 & ~w5292;
assign w5294 = b[41] & w11;
assign w5295 = b[40] & w9;
assign w5296 = ~b[40] & ~b[41];
assign w5297 = b[40] & b[41];
assign w5298 = ~w5296 & ~w5297;
assign w5299 = ~w5052 & ~w5056;
assign w5300 = ~w5298 & ~w5299;
assign w5301 = w5298 & w5299;
assign w5302 = ~w5300 & ~w5301;
assign w5303 = w5 & w5302;
assign w5304 = ~w5294 & ~w5295;
assign w5305 = ~w5303 & w5304;
assign w5306 = b[39] & w24;
assign w5307 = a[2] & ~w5306;
assign w5308 = w5305 & ~w5307;
assign w5309 = a[2] & ~w5305;
assign w5310 = ~w5308 & ~w5309;
assign w5311 = ~w5293 & ~w5310;
assign w5312 = w5293 & w5310;
assign w5313 = ~w5311 & ~w5312;
assign w5314 = w5074 & ~w5313;
assign w5315 = ~w5074 & w5313;
assign w5316 = ~w5314 & ~w5315;
assign w5317 = (~w5287 & ~w5290) | (~w5287 & w24970) | (~w5290 & w24970);
assign w5318 = b[37] & w103;
assign w5319 = b[39] & w68;
assign w5320 = b[38] & w61;
assign w5321 = w66 & ~w4812;
assign w5322 = ~w5319 & ~w5320;
assign w5323 = ~w5318 & w5322;
assign w5324 = ~w5321 & w5323;
assign w5325 = a[5] & ~w5324;
assign w5326 = ~a[5] & w5324;
assign w5327 = ~w5325 & ~w5326;
assign w5328 = b[34] & ~w237;
assign w5329 = b[35] & w183;
assign w5330 = b[36] & w185;
assign w5331 = w179 & w4129;
assign w5332 = ~w5328 & ~w5329;
assign w5333 = ~w5330 & w5332;
assign w5334 = ~w5331 & w5333;
assign w5335 = a[8] & ~w5334;
assign w5336 = ~a[8] & w5334;
assign w5337 = ~w5335 & ~w5336;
assign w5338 = (~w5265 & ~w5267) | (~w5265 & w24376) | (~w5267 & w24376);
assign w5339 = (~w5258 & w5096) | (~w5258 & w24658) | (w5096 & w24658);
assign w5340 = b[30] & w575;
assign w5341 = b[29] & w573;
assign w5342 = b[28] & ~w649;
assign w5343 = w569 & ~w2908;
assign w5344 = ~w5340 & ~w5341;
assign w5345 = ~w5342 & w5344;
assign w5346 = ~w5343 & w5345;
assign w5347 = a[14] & ~w5346;
assign w5348 = ~a[14] & w5346;
assign w5349 = ~w5347 & ~w5348;
assign w5350 = ~w5252 & ~w5255;
assign w5351 = b[24] & w1156;
assign w5352 = b[22] & ~w1272;
assign w5353 = b[23] & w1154;
assign w5354 = w1150 & w1895;
assign w5355 = ~w5351 & ~w5352;
assign w5356 = ~w5353 & w5355;
assign w5357 = ~w5354 & w5356;
assign w5358 = a[20] & ~w5357;
assign w5359 = ~a[20] & w5357;
assign w5360 = ~w5358 & ~w5359;
assign w5361 = (~w5226 & ~w5229) | (~w5226 & w25259) | (~w5229 & w25259);
assign w5362 = b[21] & w1519;
assign w5363 = b[20] & w1517;
assign w5364 = b[19] & ~w1676;
assign w5365 = w1467 & w1513;
assign w5366 = ~w5362 & ~w5363;
assign w5367 = ~w5364 & w5366;
assign w5368 = ~w5365 & w5367;
assign w5369 = a[23] & ~w5368;
assign w5370 = ~a[23] & w5368;
assign w5371 = ~w5369 & ~w5370;
assign w5372 = ~w5221 & ~w5223;
assign w5373 = b[17] & w1955;
assign w5374 = b[18] & w1957;
assign w5375 = b[16] & ~w2114;
assign w5376 = ~w1108 & w1951;
assign w5377 = ~w5373 & ~w5374;
assign w5378 = ~w5375 & w5377;
assign w5379 = ~w5376 & w5378;
assign w5380 = a[26] & ~w5379;
assign w5381 = ~a[26] & w5379;
assign w5382 = ~w5380 & ~w5381;
assign w5383 = (~w5214 & w5139) | (~w5214 & w24971) | (w5139 & w24971);
assign w5384 = b[13] & ~w2622;
assign w5385 = b[14] & w2436;
assign w5386 = b[15] & w2438;
assign w5387 = ~w799 & w2432;
assign w5388 = ~w5384 & ~w5385;
assign w5389 = ~w5386 & w5388;
assign w5390 = ~w5387 & w5389;
assign w5391 = a[29] & ~w5390;
assign w5392 = ~a[29] & w5390;
assign w5393 = ~w5391 & ~w5392;
assign w5394 = (~w5192 & ~w5194) | (~w5192 & w24972) | (~w5194 & w24972);
assign w5395 = a[41] & ~a[42];
assign w5396 = ~a[41] & a[42];
assign w5397 = ~w5395 & ~w5396;
assign w5398 = b[0] & ~w5397;
assign w5399 = w5161 & w5171;
assign w5400 = w5166 & w24808;
assign w5401 = b[2] & w4918;
assign w5402 = b[3] & w4925;
assign w5403 = ~w5401 & ~w5402;
assign w5404 = ~w5400 & w5403;
assign w5405 = (a[41] & ~w5404) | (a[41] & w24809) | (~w5404 & w24809);
assign w5406 = w5404 & w24810;
assign w5407 = ~w5405 & ~w5406;
assign w5408 = w5399 & w5407;
assign w5409 = ~w5399 & ~w5407;
assign w5410 = ~w5408 & ~w5409;
assign w5411 = ~w5398 & ~w5410;
assign w5412 = w5398 & w5410;
assign w5413 = ~w5411 & ~w5412;
assign w5414 = b[4] & w4453;
assign w5415 = b[5] & w4241;
assign w5416 = b[6] & w4243;
assign w5417 = w157 & w4236;
assign w5418 = ~w5415 & ~w5416;
assign w5419 = ~w5414 & w5418;
assign w5420 = ~w5417 & w5419;
assign w5421 = a[38] & ~w5420;
assign w5422 = ~a[38] & w5420;
assign w5423 = ~w5421 & ~w5422;
assign w5424 = w5413 & w5423;
assign w5425 = ~w5413 & ~w5423;
assign w5426 = ~w5424 & ~w5425;
assign w5427 = (~w5175 & w5151) | (~w5175 & w24811) | (w5151 & w24811);
assign w5428 = ~w5426 & w5427;
assign w5429 = w5426 & ~w5427;
assign w5430 = ~w5428 & ~w5429;
assign w5431 = b[7] & w3785;
assign w5432 = b[8] & w3578;
assign w5433 = b[9] & w3580;
assign w5434 = w322 & w3573;
assign w5435 = ~w5432 & ~w5433;
assign w5436 = ~w5431 & w5435;
assign w5437 = ~w5434 & w5436;
assign w5438 = a[35] & ~w5437;
assign w5439 = ~a[35] & w5437;
assign w5440 = ~w5438 & ~w5439;
assign w5441 = ~w5430 & ~w5440;
assign w5442 = w5430 & w5440;
assign w5443 = ~w5441 & ~w5442;
assign w5444 = w5394 & w5443;
assign w5445 = ~w5394 & ~w5443;
assign w5446 = ~w5444 & ~w5445;
assign w5447 = b[10] & w3177;
assign w5448 = b[11] & w2973;
assign w5449 = b[12] & w2978;
assign w5450 = w536 & w2980;
assign w5451 = ~w5448 & ~w5449;
assign w5452 = ~w5447 & w5451;
assign w5453 = ~w5450 & w5452;
assign w5454 = a[32] & ~w5453;
assign w5455 = ~a[32] & w5453;
assign w5456 = ~w5454 & ~w5455;
assign w5457 = w5446 & ~w5456;
assign w5458 = ~w5446 & w5456;
assign w5459 = ~w5457 & ~w5458;
assign w5460 = ~w5208 & ~w5211;
assign w5461 = w5459 & w5460;
assign w5462 = ~w5459 & ~w5460;
assign w5463 = ~w5461 & ~w5462;
assign w5464 = w5393 & w5463;
assign w5465 = ~w5393 & ~w5463;
assign w5466 = ~w5464 & ~w5465;
assign w5467 = ~w5383 & ~w5466;
assign w5468 = w5383 & w5466;
assign w5469 = ~w5467 & ~w5468;
assign w5470 = ~w5382 & w5469;
assign w5471 = w5382 & ~w5469;
assign w5472 = ~w5470 & ~w5471;
assign w5473 = ~w5372 & w5472;
assign w5474 = w5372 & ~w5472;
assign w5475 = ~w5473 & ~w5474;
assign w5476 = w5371 & w5475;
assign w5477 = ~w5371 & ~w5475;
assign w5478 = ~w5476 & ~w5477;
assign w5479 = ~w5361 & w5478;
assign w5480 = w5361 & ~w5478;
assign w5481 = ~w5479 & ~w5480;
assign w5482 = ~w5360 & ~w5481;
assign w5483 = w5360 & w5481;
assign w5484 = ~w5482 & ~w5483;
assign w5485 = ~w5245 & ~w5248;
assign w5486 = w5484 & w5485;
assign w5487 = ~w5484 & ~w5485;
assign w5488 = ~w5486 & ~w5487;
assign w5489 = b[25] & ~w934;
assign w5490 = b[26] & w838;
assign w5491 = b[27] & w834;
assign w5492 = w832 & w2378;
assign w5493 = ~w5489 & ~w5490;
assign w5494 = ~w5491 & w5493;
assign w5495 = ~w5492 & w5494;
assign w5496 = a[17] & ~w5495;
assign w5497 = ~a[17] & w5495;
assign w5498 = ~w5496 & ~w5497;
assign w5499 = w5488 & w5498;
assign w5500 = ~w5488 & ~w5498;
assign w5501 = ~w5499 & ~w5500;
assign w5502 = w5350 & ~w5501;
assign w5503 = ~w5350 & w5501;
assign w5504 = ~w5502 & ~w5503;
assign w5505 = ~w5349 & ~w5504;
assign w5506 = w5349 & w5504;
assign w5507 = ~w5505 & ~w5506;
assign w5508 = ~w5339 & w5507;
assign w5509 = w5339 & ~w5507;
assign w5510 = ~w5508 & ~w5509;
assign w5511 = b[32] & w358;
assign w5512 = b[31] & ~w419;
assign w5513 = b[33] & w360;
assign w5514 = w354 & w3499;
assign w5515 = ~w5511 & ~w5512;
assign w5516 = ~w5513 & w5515;
assign w5517 = ~w5514 & w5516;
assign w5518 = a[11] & ~w5517;
assign w5519 = ~a[11] & w5517;
assign w5520 = ~w5518 & ~w5519;
assign w5521 = w5510 & w5520;
assign w5522 = ~w5510 & ~w5520;
assign w5523 = ~w5521 & ~w5522;
assign w5524 = w5338 & w5523;
assign w5525 = ~w5338 & ~w5523;
assign w5526 = ~w5524 & ~w5525;
assign w5527 = ~w5337 & w5526;
assign w5528 = w5337 & ~w5526;
assign w5529 = ~w5527 & ~w5528;
assign w5530 = (~w5282 & ~w5085) | (~w5282 & w25128) | (~w5085 & w25128);
assign w5531 = w5529 & w5530;
assign w5532 = ~w5529 & ~w5530;
assign w5533 = ~w5531 & ~w5532;
assign w5534 = ~w5327 & ~w5533;
assign w5535 = w5327 & w5533;
assign w5536 = ~w5534 & ~w5535;
assign w5537 = w5317 & w5536;
assign w5538 = ~w5317 & ~w5536;
assign w5539 = ~w5537 & ~w5538;
assign w5540 = b[42] & w11;
assign w5541 = b[41] & w9;
assign w5542 = ~w5297 & ~w5301;
assign w5543 = ~b[41] & ~b[42];
assign w5544 = b[41] & b[42];
assign w5545 = ~w5543 & ~w5544;
assign w5546 = w5542 & ~w5545;
assign w5547 = ~w5542 & w5545;
assign w5548 = ~w5546 & ~w5547;
assign w5549 = w5 & w5548;
assign w5550 = ~w5540 & ~w5541;
assign w5551 = ~w5549 & w5550;
assign w5552 = b[40] & w24;
assign w5553 = a[2] & ~w5552;
assign w5554 = w5551 & ~w5553;
assign w5555 = a[2] & ~w5551;
assign w5556 = ~w5554 & ~w5555;
assign w5557 = ~w5539 & w5556;
assign w5558 = w5539 & ~w5556;
assign w5559 = ~w5557 & ~w5558;
assign w5560 = ~w5312 & ~w5315;
assign w5561 = w5559 & ~w5560;
assign w5562 = ~w5559 & w5560;
assign w5563 = ~w5561 & ~w5562;
assign w5564 = b[38] & w103;
assign w5565 = b[39] & w61;
assign w5566 = b[40] & w68;
assign w5567 = w66 & ~w5058;
assign w5568 = ~w5565 & ~w5566;
assign w5569 = ~w5564 & w5568;
assign w5570 = ~w5567 & w5569;
assign w5571 = a[5] & ~w5570;
assign w5572 = ~a[5] & w5570;
assign w5573 = ~w5571 & ~w5572;
assign w5574 = b[34] & w360;
assign w5575 = b[33] & w358;
assign w5576 = b[32] & ~w419;
assign w5577 = w354 & ~w3710;
assign w5578 = ~w5574 & ~w5575;
assign w5579 = ~w5576 & w5578;
assign w5580 = ~w5577 & w5579;
assign w5581 = a[11] & ~w5580;
assign w5582 = ~a[11] & w5580;
assign w5583 = ~w5581 & ~w5582;
assign w5584 = ~w5506 & ~w5508;
assign w5585 = b[31] & w575;
assign w5586 = b[30] & w573;
assign w5587 = b[29] & ~w649;
assign w5588 = w569 & ~w3112;
assign w5589 = ~w5585 & ~w5586;
assign w5590 = ~w5587 & w5589;
assign w5591 = ~w5588 & w5590;
assign w5592 = a[14] & ~w5591;
assign w5593 = ~a[14] & w5591;
assign w5594 = ~w5592 & ~w5593;
assign w5595 = b[28] & w834;
assign w5596 = b[27] & w838;
assign w5597 = b[26] & ~w934;
assign w5598 = w832 & w2559;
assign w5599 = ~w5595 & ~w5596;
assign w5600 = ~w5597 & w5599;
assign w5601 = ~w5598 & w5600;
assign w5602 = a[17] & ~w5601;
assign w5603 = ~a[17] & w5601;
assign w5604 = ~w5602 & ~w5603;
assign w5605 = (~w5483 & ~w5485) | (~w5483 & w25260) | (~w5485 & w25260);
assign w5606 = ~w5476 & ~w5479;
assign w5607 = b[22] & w1519;
assign w5608 = b[21] & w1517;
assign w5609 = b[20] & ~w1676;
assign w5610 = w1513 & w1615;
assign w5611 = ~w5607 & ~w5608;
assign w5612 = ~w5609 & w5611;
assign w5613 = ~w5610 & w5612;
assign w5614 = a[23] & ~w5613;
assign w5615 = ~a[23] & w5613;
assign w5616 = ~w5614 & ~w5615;
assign w5617 = (~w5471 & w5372) | (~w5471 & w25129) | (w5372 & w25129);
assign w5618 = b[14] & ~w2622;
assign w5619 = b[15] & w2436;
assign w5620 = b[16] & w2438;
assign w5621 = w905 & w2432;
assign w5622 = ~w5618 & ~w5619;
assign w5623 = ~w5620 & w5622;
assign w5624 = ~w5621 & w5623;
assign w5625 = a[29] & ~w5624;
assign w5626 = ~a[29] & w5624;
assign w5627 = ~w5625 & ~w5626;
assign w5628 = (~w5458 & ~w5460) | (~w5458 & w25130) | (~w5460 & w25130);
assign w5629 = b[11] & w3177;
assign w5630 = b[12] & w2973;
assign w5631 = b[13] & w2978;
assign w5632 = w628 & w2980;
assign w5633 = ~w5630 & ~w5631;
assign w5634 = ~w5629 & w5633;
assign w5635 = ~w5632 & w5634;
assign w5636 = a[32] & ~w5635;
assign w5637 = ~a[32] & w5635;
assign w5638 = ~w5636 & ~w5637;
assign w5639 = b[8] & w3785;
assign w5640 = b[9] & w3578;
assign w5641 = b[10] & w3580;
assign w5642 = w397 & w3573;
assign w5643 = ~w5640 & ~w5641;
assign w5644 = ~w5639 & w5643;
assign w5645 = ~w5642 & w5644;
assign w5646 = a[35] & ~w5645;
assign w5647 = ~a[35] & w5645;
assign w5648 = ~w5646 & ~w5647;
assign w5649 = w5166 & w25131;
assign w5650 = b[4] & w4925;
assign w5651 = b[3] & w4918;
assign w5652 = w84 & w4923;
assign w5653 = ~w5650 & ~w5651;
assign w5654 = ~w5649 & w5653;
assign w5655 = ~w5652 & w5654;
assign w5656 = a[41] & ~w5655;
assign w5657 = ~a[41] & w5655;
assign w5658 = ~w5656 & ~w5657;
assign w5659 = a[44] & w5398;
assign w5660 = a[43] & ~a[44];
assign w5661 = ~a[43] & a[44];
assign w5662 = ~w5660 & ~w5661;
assign w5663 = ~w5397 & ~w5662;
assign w5664 = ~w8 & w5663;
assign w5665 = ~w5397 & w5662;
assign w5666 = b[1] & w5665;
assign w5667 = a[42] & ~a[43];
assign w5668 = ~a[42] & a[43];
assign w5669 = ~w5667 & ~w5668;
assign w5670 = w5397 & ~w5669;
assign w5671 = b[0] & w5670;
assign w5672 = ~w5664 & ~w5666;
assign w5673 = ~w5671 & w5672;
assign w5674 = ~w5659 & w5673;
assign w5675 = w5659 & ~w5673;
assign w5676 = ~w5674 & ~w5675;
assign w5677 = ~w5658 & ~w5676;
assign w5678 = w5658 & w5676;
assign w5679 = ~w5677 & ~w5678;
assign w5680 = (~w5408 & ~w5410) | (~w5408 & w24973) | (~w5410 & w24973);
assign w5681 = w5679 & ~w5680;
assign w5682 = ~w5679 & w5680;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = b[5] & w4453;
assign w5685 = b[7] & w4243;
assign w5686 = b[6] & w4241;
assign w5687 = w216 & w4236;
assign w5688 = ~w5685 & ~w5686;
assign w5689 = ~w5684 & w5688;
assign w5690 = ~w5687 & w5689;
assign w5691 = a[38] & ~w5690;
assign w5692 = ~a[38] & w5690;
assign w5693 = ~w5691 & ~w5692;
assign w5694 = w5683 & w5693;
assign w5695 = ~w5683 & ~w5693;
assign w5696 = ~w5694 & ~w5695;
assign w5697 = ~w5424 & ~w5429;
assign w5698 = w5696 & w5697;
assign w5699 = ~w5696 & ~w5697;
assign w5700 = ~w5698 & ~w5699;
assign w5701 = w5648 & ~w5700;
assign w5702 = ~w5648 & w5700;
assign w5703 = ~w5701 & ~w5702;
assign w5704 = ~w5441 & ~w5444;
assign w5705 = w5703 & w5704;
assign w5706 = ~w5703 & ~w5704;
assign w5707 = ~w5705 & ~w5706;
assign w5708 = ~w5638 & ~w5707;
assign w5709 = w5638 & w5707;
assign w5710 = ~w5708 & ~w5709;
assign w5711 = ~w5628 & ~w5710;
assign w5712 = w5628 & w5710;
assign w5713 = ~w5711 & ~w5712;
assign w5714 = w5627 & ~w5713;
assign w5715 = ~w5627 & w5713;
assign w5716 = ~w5714 & ~w5715;
assign w5717 = ~w5465 & ~w5468;
assign w5718 = ~w5716 & ~w5717;
assign w5719 = w5716 & w5717;
assign w5720 = ~w5718 & ~w5719;
assign w5721 = b[17] & ~w2114;
assign w5722 = b[19] & w1957;
assign w5723 = b[18] & w1955;
assign w5724 = ~w1231 & w1951;
assign w5725 = ~w5721 & ~w5722;
assign w5726 = ~w5723 & w5725;
assign w5727 = ~w5724 & w5726;
assign w5728 = a[26] & ~w5727;
assign w5729 = ~a[26] & w5727;
assign w5730 = ~w5728 & ~w5729;
assign w5731 = w5720 & w5730;
assign w5732 = ~w5720 & ~w5730;
assign w5733 = ~w5731 & ~w5732;
assign w5734 = ~w5617 & ~w5733;
assign w5735 = w5617 & w5733;
assign w5736 = ~w5734 & ~w5735;
assign w5737 = ~w5616 & w5736;
assign w5738 = w5616 & ~w5736;
assign w5739 = ~w5737 & ~w5738;
assign w5740 = w5606 & ~w5739;
assign w5741 = ~w5606 & w5739;
assign w5742 = ~w5740 & ~w5741;
assign w5743 = b[24] & w1154;
assign w5744 = b[25] & w1156;
assign w5745 = b[23] & ~w1272;
assign w5746 = w1150 & w2061;
assign w5747 = ~w5743 & ~w5744;
assign w5748 = ~w5745 & w5747;
assign w5749 = ~w5746 & w5748;
assign w5750 = a[20] & ~w5749;
assign w5751 = ~a[20] & w5749;
assign w5752 = ~w5750 & ~w5751;
assign w5753 = w5742 & w5752;
assign w5754 = ~w5742 & ~w5752;
assign w5755 = ~w5753 & ~w5754;
assign w5756 = ~w5605 & ~w5755;
assign w5757 = w5605 & w5755;
assign w5758 = ~w5756 & ~w5757;
assign w5759 = ~w5604 & w5758;
assign w5760 = w5604 & ~w5758;
assign w5761 = ~w5759 & ~w5760;
assign w5762 = ~w5499 & ~w5503;
assign w5763 = w5761 & ~w5762;
assign w5764 = ~w5761 & w5762;
assign w5765 = ~w5763 & ~w5764;
assign w5766 = w5594 & w5765;
assign w5767 = ~w5594 & ~w5765;
assign w5768 = ~w5766 & ~w5767;
assign w5769 = w5584 & ~w5768;
assign w5770 = ~w5584 & w5768;
assign w5771 = ~w5769 & ~w5770;
assign w5772 = w5583 & w5771;
assign w5773 = ~w5583 & ~w5771;
assign w5774 = ~w5772 & ~w5773;
assign w5775 = (~w5522 & ~w5338) | (~w5522 & w24659) | (~w5338 & w24659);
assign w5776 = ~w5774 & ~w5775;
assign w5777 = w5774 & w5775;
assign w5778 = ~w5776 & ~w5777;
assign w5779 = b[37] & w185;
assign w5780 = b[35] & ~w237;
assign w5781 = b[36] & w183;
assign w5782 = w179 & ~w4357;
assign w5783 = ~w5779 & ~w5780;
assign w5784 = ~w5781 & w5783;
assign w5785 = ~w5782 & w5784;
assign w5786 = a[8] & ~w5785;
assign w5787 = ~a[8] & w5785;
assign w5788 = ~w5786 & ~w5787;
assign w5789 = w5778 & w5788;
assign w5790 = ~w5778 & ~w5788;
assign w5791 = ~w5789 & ~w5790;
assign w5792 = (~w5528 & ~w5530) | (~w5528 & w24377) | (~w5530 & w24377);
assign w5793 = w5791 & w5792;
assign w5794 = ~w5791 & ~w5792;
assign w5795 = ~w5793 & ~w5794;
assign w5796 = w5573 & ~w5795;
assign w5797 = ~w5573 & w5795;
assign w5798 = ~w5796 & ~w5797;
assign w5799 = (~w5534 & ~w5317) | (~w5534 & w25132) | (~w5317 & w25132);
assign w5800 = w5798 & w5799;
assign w5801 = ~w5798 & ~w5799;
assign w5802 = ~w5800 & ~w5801;
assign w5803 = b[43] & w11;
assign w5804 = b[42] & w9;
assign w5805 = ~b[42] & ~b[43];
assign w5806 = b[42] & b[43];
assign w5807 = ~w5805 & ~w5806;
assign w5808 = ~w5544 & ~w5547;
assign w5809 = w5807 & ~w5808;
assign w5810 = ~w5807 & w5808;
assign w5811 = ~w5809 & ~w5810;
assign w5812 = w5 & w5811;
assign w5813 = ~w5803 & ~w5804;
assign w5814 = ~w5812 & w5813;
assign w5815 = b[41] & w24;
assign w5816 = a[2] & ~w5815;
assign w5817 = w5814 & ~w5816;
assign w5818 = a[2] & ~w5814;
assign w5819 = ~w5817 & ~w5818;
assign w5820 = w5802 & w5819;
assign w5821 = ~w5802 & ~w5819;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = (~w5557 & w5560) | (~w5557 & w24974) | (w5560 & w24974);
assign w5824 = ~w5822 & ~w5823;
assign w5825 = w5822 & w5823;
assign w5826 = ~w5824 & ~w5825;
assign w5827 = (~w5796 & ~w5799) | (~w5796 & w24378) | (~w5799 & w24378);
assign w5828 = b[39] & w103;
assign w5829 = b[40] & w61;
assign w5830 = b[41] & w68;
assign w5831 = w66 & w5302;
assign w5832 = ~w5829 & ~w5830;
assign w5833 = ~w5828 & w5832;
assign w5834 = ~w5831 & w5833;
assign w5835 = a[5] & ~w5834;
assign w5836 = ~a[5] & w5834;
assign w5837 = ~w5835 & ~w5836;
assign w5838 = b[36] & ~w237;
assign w5839 = b[38] & w185;
assign w5840 = b[37] & w183;
assign w5841 = w179 & w4582;
assign w5842 = ~w5838 & ~w5839;
assign w5843 = ~w5840 & w5842;
assign w5844 = ~w5841 & w5843;
assign w5845 = a[8] & ~w5844;
assign w5846 = ~a[8] & w5844;
assign w5847 = ~w5845 & ~w5846;
assign w5848 = ~w5766 & ~w5770;
assign w5849 = b[30] & ~w649;
assign w5850 = b[31] & w573;
assign w5851 = b[32] & w575;
assign w5852 = w569 & w3304;
assign w5853 = ~w5849 & ~w5850;
assign w5854 = ~w5851 & w5853;
assign w5855 = ~w5852 & w5854;
assign w5856 = a[14] & ~w5855;
assign w5857 = ~a[14] & w5855;
assign w5858 = ~w5856 & ~w5857;
assign w5859 = (~w5760 & w5762) | (~w5760 & w25261) | (w5762 & w25261);
assign w5860 = b[27] & ~w934;
assign w5861 = b[29] & w834;
assign w5862 = b[28] & w838;
assign w5863 = w832 & w2734;
assign w5864 = ~w5860 & ~w5861;
assign w5865 = ~w5862 & w5864;
assign w5866 = ~w5863 & w5865;
assign w5867 = a[17] & ~w5866;
assign w5868 = ~a[17] & w5866;
assign w5869 = ~w5867 & ~w5868;
assign w5870 = b[24] & ~w1272;
assign w5871 = b[25] & w1154;
assign w5872 = b[26] & w1156;
assign w5873 = w1150 & w2219;
assign w5874 = ~w5870 & ~w5871;
assign w5875 = ~w5872 & w5874;
assign w5876 = ~w5873 & w5875;
assign w5877 = a[20] & ~w5876;
assign w5878 = ~a[20] & w5876;
assign w5879 = ~w5877 & ~w5878;
assign w5880 = ~w5738 & ~w5741;
assign w5881 = b[18] & ~w2114;
assign w5882 = b[20] & w1957;
assign w5883 = b[19] & w1955;
assign w5884 = w1347 & w1951;
assign w5885 = ~w5881 & ~w5882;
assign w5886 = ~w5883 & w5885;
assign w5887 = ~w5884 & w5886;
assign w5888 = a[26] & ~w5887;
assign w5889 = ~a[26] & w5887;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = (~w5714 & ~w5717) | (~w5714 & w25133) | (~w5717 & w25133);
assign w5892 = b[16] & w2436;
assign w5893 = b[17] & w2438;
assign w5894 = b[15] & ~w2622;
assign w5895 = w1008 & w2432;
assign w5896 = ~w5892 & ~w5893;
assign w5897 = ~w5894 & w5896;
assign w5898 = ~w5895 & w5897;
assign w5899 = a[29] & ~w5898;
assign w5900 = ~a[29] & w5898;
assign w5901 = ~w5899 & ~w5900;
assign w5902 = b[12] & w3177;
assign w5903 = b[13] & w2973;
assign w5904 = b[14] & w2978;
assign w5905 = w714 & w2980;
assign w5906 = ~w5903 & ~w5904;
assign w5907 = ~w5902 & w5906;
assign w5908 = ~w5905 & w5907;
assign w5909 = a[32] & ~w5908;
assign w5910 = ~a[32] & w5908;
assign w5911 = ~w5909 & ~w5910;
assign w5912 = ~w5701 & ~w5705;
assign w5913 = b[9] & w3785;
assign w5914 = b[10] & w3578;
assign w5915 = b[11] & w3580;
assign w5916 = w469 & w3573;
assign w5917 = ~w5914 & ~w5915;
assign w5918 = ~w5913 & w5917;
assign w5919 = ~w5916 & w5918;
assign w5920 = a[35] & ~w5919;
assign w5921 = ~a[35] & w5919;
assign w5922 = ~w5920 & ~w5921;
assign w5923 = ~w5678 & ~w5681;
assign w5924 = w5166 & w25418;
assign w5925 = b[5] & w4925;
assign w5926 = b[4] & w4918;
assign w5927 = w116 & w4923;
assign w5928 = ~w5925 & ~w5926;
assign w5929 = (a[41] & w5927) | (a[41] & w25134) | (w5927 & w25134);
assign w5930 = ~w5927 & w25135;
assign w5931 = ~w5929 & ~w5930;
assign w5932 = (a[44] & w5397) | (a[44] & w25419) | (w5397 & w25419);
assign w5933 = w5672 & w24975;
assign w5934 = a[44] & ~w5933;
assign w5935 = w22 & w5663;
assign w5936 = b[2] & w5665;
assign w5937 = b[1] & w5670;
assign w5938 = w5397 & ~w5662;
assign w5939 = w5669 & w5938;
assign w5940 = b[0] & w5939;
assign w5941 = ~w5935 & ~w5936;
assign w5942 = ~w5937 & w5941;
assign w5943 = ~w5940 & w5942;
assign w5944 = ~w5934 & w5943;
assign w5945 = w5934 & ~w5943;
assign w5946 = ~w5944 & ~w5945;
assign w5947 = w5931 & w5946;
assign w5948 = ~w5931 & ~w5946;
assign w5949 = ~w5947 & ~w5948;
assign w5950 = ~w5681 & w25136;
assign w5951 = (~w5949 & w5681) | (~w5949 & w25137) | (w5681 & w25137);
assign w5952 = ~w5950 & ~w5951;
assign w5953 = b[6] & w4453;
assign w5954 = b[7] & w4241;
assign w5955 = b[8] & w4243;
assign w5956 = w270 & w4236;
assign w5957 = ~w5954 & ~w5955;
assign w5958 = ~w5953 & w5957;
assign w5959 = ~w5956 & w5958;
assign w5960 = a[38] & ~w5959;
assign w5961 = ~a[38] & w5959;
assign w5962 = ~w5960 & ~w5961;
assign w5963 = w5952 & ~w5962;
assign w5964 = ~w5952 & w5962;
assign w5965 = ~w5963 & ~w5964;
assign w5966 = (~w5695 & ~w5697) | (~w5695 & w24976) | (~w5697 & w24976);
assign w5967 = w5965 & w5966;
assign w5968 = ~w5965 & ~w5966;
assign w5969 = ~w5967 & ~w5968;
assign w5970 = ~w5922 & ~w5969;
assign w5971 = w5922 & w5969;
assign w5972 = ~w5970 & ~w5971;
assign w5973 = w5912 & ~w5972;
assign w5974 = ~w5912 & w5972;
assign w5975 = ~w5973 & ~w5974;
assign w5976 = ~w5911 & ~w5975;
assign w5977 = w5911 & w5975;
assign w5978 = ~w5976 & ~w5977;
assign w5979 = ~w5708 & ~w5712;
assign w5980 = w5978 & w5979;
assign w5981 = ~w5978 & ~w5979;
assign w5982 = ~w5980 & ~w5981;
assign w5983 = ~w5901 & ~w5982;
assign w5984 = w5901 & w5982;
assign w5985 = ~w5983 & ~w5984;
assign w5986 = ~w5891 & ~w5985;
assign w5987 = w5891 & w5985;
assign w5988 = ~w5986 & ~w5987;
assign w5989 = ~w5890 & w5988;
assign w5990 = w5890 & ~w5988;
assign w5991 = ~w5989 & ~w5990;
assign w5992 = ~w5732 & ~w5735;
assign w5993 = ~w5991 & ~w5992;
assign w5994 = w5991 & w5992;
assign w5995 = ~w5993 & ~w5994;
assign w5996 = b[23] & w1519;
assign w5997 = b[22] & w1517;
assign w5998 = b[21] & ~w1676;
assign w5999 = w1513 & w1755;
assign w6000 = ~w5996 & ~w5997;
assign w6001 = ~w5998 & w6000;
assign w6002 = ~w5999 & w6001;
assign w6003 = a[23] & ~w6002;
assign w6004 = ~a[23] & w6002;
assign w6005 = ~w6003 & ~w6004;
assign w6006 = ~w5995 & ~w6005;
assign w6007 = w5995 & w6005;
assign w6008 = ~w6006 & ~w6007;
assign w6009 = w5880 & w6008;
assign w6010 = ~w5880 & ~w6008;
assign w6011 = ~w6009 & ~w6010;
assign w6012 = ~w5879 & w6011;
assign w6013 = w5879 & ~w6011;
assign w6014 = ~w6012 & ~w6013;
assign w6015 = ~w5754 & ~w5757;
assign w6016 = w6014 & w6015;
assign w6017 = ~w6014 & ~w6015;
assign w6018 = ~w6016 & ~w6017;
assign w6019 = ~w5869 & ~w6018;
assign w6020 = w5869 & w6018;
assign w6021 = ~w6019 & ~w6020;
assign w6022 = w5859 & ~w6021;
assign w6023 = ~w5859 & w6021;
assign w6024 = ~w6022 & ~w6023;
assign w6025 = ~w5858 & ~w6024;
assign w6026 = w5858 & w6024;
assign w6027 = ~w6025 & ~w6026;
assign w6028 = ~w5848 & w6027;
assign w6029 = w5848 & ~w6027;
assign w6030 = ~w6028 & ~w6029;
assign w6031 = b[35] & w360;
assign w6032 = b[33] & ~w419;
assign w6033 = b[34] & w358;
assign w6034 = w354 & w3918;
assign w6035 = ~w6031 & ~w6032;
assign w6036 = ~w6033 & w6035;
assign w6037 = ~w6034 & w6036;
assign w6038 = a[11] & ~w6037;
assign w6039 = ~a[11] & w6037;
assign w6040 = ~w6038 & ~w6039;
assign w6041 = w6030 & w6040;
assign w6042 = ~w6030 & ~w6040;
assign w6043 = ~w6041 & ~w6042;
assign w6044 = ~w5772 & ~w5777;
assign w6045 = w6043 & w6044;
assign w6046 = ~w6043 & ~w6044;
assign w6047 = ~w6045 & ~w6046;
assign w6048 = w5847 & ~w6047;
assign w6049 = ~w5847 & w6047;
assign w6050 = ~w6048 & ~w6049;
assign w6051 = (~w5790 & ~w5792) | (~w5790 & w24660) | (~w5792 & w24660);
assign w6052 = w6050 & w6051;
assign w6053 = ~w6050 & ~w6051;
assign w6054 = ~w6052 & ~w6053;
assign w6055 = ~w5837 & ~w6054;
assign w6056 = w5837 & w6054;
assign w6057 = ~w6055 & ~w6056;
assign w6058 = ~w5827 & ~w6057;
assign w6059 = w5827 & w6057;
assign w6060 = ~w6058 & ~w6059;
assign w6061 = b[44] & w11;
assign w6062 = b[43] & w9;
assign w6063 = ~b[43] & ~b[44];
assign w6064 = b[43] & b[44];
assign w6065 = ~w6063 & ~w6064;
assign w6066 = ~w5806 & ~w5809;
assign w6067 = w6065 & ~w6066;
assign w6068 = ~w6065 & w6066;
assign w6069 = ~w6067 & ~w6068;
assign w6070 = w5 & w6069;
assign w6071 = ~w6061 & ~w6062;
assign w6072 = ~w6070 & w6071;
assign w6073 = b[42] & w24;
assign w6074 = a[2] & ~w6073;
assign w6075 = w6072 & ~w6074;
assign w6076 = a[2] & ~w6072;
assign w6077 = ~w6075 & ~w6076;
assign w6078 = ~w6060 & w6077;
assign w6079 = w6060 & ~w6077;
assign w6080 = ~w6078 & ~w6079;
assign w6081 = (~w5821 & ~w5823) | (~w5821 & w25138) | (~w5823 & w25138);
assign w6082 = w6080 & w6081;
assign w6083 = ~w6080 & ~w6081;
assign w6084 = ~w6082 & ~w6083;
assign w6085 = (~w6078 & ~w6081) | (~w6078 & w24379) | (~w6081 & w24379);
assign w6086 = b[40] & w103;
assign w6087 = b[42] & w68;
assign w6088 = b[41] & w61;
assign w6089 = w66 & w5548;
assign w6090 = ~w6087 & ~w6088;
assign w6091 = ~w6086 & w6090;
assign w6092 = ~w6089 & w6091;
assign w6093 = a[5] & ~w6092;
assign w6094 = ~a[5] & w6092;
assign w6095 = ~w6093 & ~w6094;
assign w6096 = b[36] & w360;
assign w6097 = b[35] & w358;
assign w6098 = b[34] & ~w419;
assign w6099 = w354 & w4129;
assign w6100 = ~w6096 & ~w6097;
assign w6101 = ~w6098 & w6100;
assign w6102 = ~w6099 & w6101;
assign w6103 = a[11] & ~w6102;
assign w6104 = ~a[11] & w6102;
assign w6105 = ~w6103 & ~w6104;
assign w6106 = (~w6026 & w5848) | (~w6026 & w25262) | (w5848 & w25262);
assign w6107 = b[33] & w575;
assign w6108 = b[32] & w573;
assign w6109 = b[31] & ~w649;
assign w6110 = w569 & w3499;
assign w6111 = ~w6107 & ~w6108;
assign w6112 = ~w6109 & w6111;
assign w6113 = ~w6110 & w6112;
assign w6114 = a[14] & ~w6113;
assign w6115 = ~a[14] & w6113;
assign w6116 = ~w6114 & ~w6115;
assign w6117 = b[30] & w834;
assign w6118 = b[28] & ~w934;
assign w6119 = b[29] & w838;
assign w6120 = w832 & ~w2908;
assign w6121 = ~w6117 & ~w6118;
assign w6122 = ~w6119 & w6121;
assign w6123 = ~w6120 & w6122;
assign w6124 = a[17] & ~w6123;
assign w6125 = ~a[17] & w6123;
assign w6126 = ~w6124 & ~w6125;
assign w6127 = ~w6013 & ~w6016;
assign w6128 = b[23] & w1517;
assign w6129 = b[24] & w1519;
assign w6130 = b[22] & ~w1676;
assign w6131 = w1513 & w1895;
assign w6132 = ~w6128 & ~w6129;
assign w6133 = ~w6130 & w6132;
assign w6134 = ~w6131 & w6133;
assign w6135 = a[23] & ~w6134;
assign w6136 = ~a[23] & w6134;
assign w6137 = ~w6135 & ~w6136;
assign w6138 = (~w5990 & ~w5992) | (~w5990 & w25263) | (~w5992 & w25263);
assign w6139 = b[17] & w2436;
assign w6140 = b[18] & w2438;
assign w6141 = b[16] & ~w2622;
assign w6142 = ~w1108 & w2432;
assign w6143 = ~w6139 & ~w6140;
assign w6144 = ~w6141 & w6143;
assign w6145 = ~w6142 & w6144;
assign w6146 = a[29] & ~w6145;
assign w6147 = ~a[29] & w6145;
assign w6148 = ~w6146 & ~w6147;
assign w6149 = b[13] & w3177;
assign w6150 = b[15] & w2978;
assign w6151 = b[14] & w2973;
assign w6152 = ~w799 & w2980;
assign w6153 = ~w6150 & ~w6151;
assign w6154 = ~w6149 & w6153;
assign w6155 = ~w6152 & w6154;
assign w6156 = a[32] & ~w6155;
assign w6157 = ~a[32] & w6155;
assign w6158 = ~w6156 & ~w6157;
assign w6159 = (~w5964 & ~w5966) | (~w5964 & w25139) | (~w5966 & w25139);
assign w6160 = a[44] & ~a[45];
assign w6161 = ~a[44] & a[45];
assign w6162 = ~w6160 & ~w6161;
assign w6163 = b[0] & ~w6162;
assign w6164 = w5933 & w5943;
assign w6165 = w46 & w5663;
assign w6166 = b[2] & w5670;
assign w6167 = b[3] & w5665;
assign w6168 = w5938 & w24977;
assign w6169 = ~w6166 & ~w6167;
assign w6170 = ~w6165 & w6169;
assign w6171 = (a[44] & ~w6170) | (a[44] & w24812) | (~w6170 & w24812);
assign w6172 = w6170 & w24813;
assign w6173 = ~w6171 & ~w6172;
assign w6174 = w6164 & w6173;
assign w6175 = ~w6164 & ~w6173;
assign w6176 = ~w6174 & ~w6175;
assign w6177 = ~w6163 & ~w6176;
assign w6178 = w6163 & w6176;
assign w6179 = ~w6177 & ~w6178;
assign w6180 = b[4] & w5167;
assign w6181 = b[6] & w4925;
assign w6182 = b[5] & w4918;
assign w6183 = w157 & w4923;
assign w6184 = ~w6181 & ~w6182;
assign w6185 = ~w6180 & w6184;
assign w6186 = ~w6183 & w6185;
assign w6187 = a[41] & ~w6186;
assign w6188 = ~a[41] & w6186;
assign w6189 = ~w6187 & ~w6188;
assign w6190 = w6179 & w6189;
assign w6191 = ~w6179 & ~w6189;
assign w6192 = ~w6190 & ~w6191;
assign w6193 = (~w5948 & ~w5923) | (~w5948 & w24814) | (~w5923 & w24814);
assign w6194 = ~w6192 & ~w6193;
assign w6195 = w6192 & w6193;
assign w6196 = ~w6194 & ~w6195;
assign w6197 = b[7] & w4453;
assign w6198 = b[8] & w4241;
assign w6199 = b[9] & w4243;
assign w6200 = w322 & w4236;
assign w6201 = ~w6198 & ~w6199;
assign w6202 = ~w6197 & w6201;
assign w6203 = ~w6200 & w6202;
assign w6204 = a[38] & ~w6203;
assign w6205 = ~a[38] & w6203;
assign w6206 = ~w6204 & ~w6205;
assign w6207 = ~w6196 & ~w6206;
assign w6208 = w6196 & w6206;
assign w6209 = ~w6207 & ~w6208;
assign w6210 = w6159 & ~w6209;
assign w6211 = ~w6159 & w6209;
assign w6212 = ~w6210 & ~w6211;
assign w6213 = b[10] & w3785;
assign w6214 = b[12] & w3580;
assign w6215 = b[11] & w3578;
assign w6216 = w536 & w3573;
assign w6217 = ~w6214 & ~w6215;
assign w6218 = ~w6213 & w6217;
assign w6219 = ~w6216 & w6218;
assign w6220 = a[35] & ~w6219;
assign w6221 = ~a[35] & w6219;
assign w6222 = ~w6220 & ~w6221;
assign w6223 = ~w6212 & ~w6222;
assign w6224 = w6212 & w6222;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = (~w5971 & w5912) | (~w5971 & w24815) | (w5912 & w24815);
assign w6227 = w6225 & ~w6226;
assign w6228 = ~w6225 & w6226;
assign w6229 = ~w6227 & ~w6228;
assign w6230 = w6158 & w6229;
assign w6231 = ~w6158 & ~w6229;
assign w6232 = ~w6230 & ~w6231;
assign w6233 = (~w6232 & w5980) | (~w6232 & w24816) | (w5980 & w24816);
assign w6234 = ~w5980 & w24817;
assign w6235 = ~w6233 & ~w6234;
assign w6236 = w6148 & ~w6235;
assign w6237 = ~w6148 & w6235;
assign w6238 = ~w6236 & ~w6237;
assign w6239 = ~w5983 & ~w5987;
assign w6240 = w6238 & w6239;
assign w6241 = ~w6238 & ~w6239;
assign w6242 = ~w6240 & ~w6241;
assign w6243 = b[20] & w1955;
assign w6244 = b[19] & ~w2114;
assign w6245 = b[21] & w1957;
assign w6246 = w1467 & w1951;
assign w6247 = ~w6243 & ~w6244;
assign w6248 = ~w6245 & w6247;
assign w6249 = ~w6246 & w6248;
assign w6250 = a[26] & ~w6249;
assign w6251 = ~a[26] & w6249;
assign w6252 = ~w6250 & ~w6251;
assign w6253 = w6242 & w6252;
assign w6254 = ~w6242 & ~w6252;
assign w6255 = ~w6253 & ~w6254;
assign w6256 = w6138 & w6255;
assign w6257 = ~w6138 & ~w6255;
assign w6258 = ~w6256 & ~w6257;
assign w6259 = w6137 & ~w6258;
assign w6260 = ~w6137 & w6258;
assign w6261 = ~w6259 & ~w6260;
assign w6262 = (~w6006 & ~w5880) | (~w6006 & w24380) | (~w5880 & w24380);
assign w6263 = w6261 & w6262;
assign w6264 = ~w6261 & ~w6262;
assign w6265 = ~w6263 & ~w6264;
assign w6266 = b[27] & w1156;
assign w6267 = b[26] & w1154;
assign w6268 = b[25] & ~w1272;
assign w6269 = w1150 & w2378;
assign w6270 = ~w6266 & ~w6267;
assign w6271 = ~w6268 & w6270;
assign w6272 = ~w6269 & w6271;
assign w6273 = a[20] & ~w6272;
assign w6274 = ~a[20] & w6272;
assign w6275 = ~w6273 & ~w6274;
assign w6276 = w6265 & w6275;
assign w6277 = ~w6265 & ~w6275;
assign w6278 = ~w6276 & ~w6277;
assign w6279 = w6127 & ~w6278;
assign w6280 = ~w6127 & w6278;
assign w6281 = ~w6279 & ~w6280;
assign w6282 = ~w6126 & ~w6281;
assign w6283 = w6126 & w6281;
assign w6284 = ~w6282 & ~w6283;
assign w6285 = ~w6020 & ~w6023;
assign w6286 = w6284 & ~w6285;
assign w6287 = ~w6284 & w6285;
assign w6288 = ~w6286 & ~w6287;
assign w6289 = w6116 & w6288;
assign w6290 = ~w6116 & ~w6288;
assign w6291 = ~w6289 & ~w6290;
assign w6292 = ~w6106 & w6291;
assign w6293 = w6106 & ~w6291;
assign w6294 = ~w6292 & ~w6293;
assign w6295 = w6105 & w6294;
assign w6296 = ~w6105 & ~w6294;
assign w6297 = ~w6295 & ~w6296;
assign w6298 = ~w6042 & ~w6045;
assign w6299 = ~w6297 & ~w6298;
assign w6300 = w6297 & w6298;
assign w6301 = ~w6299 & ~w6300;
assign w6302 = b[37] & ~w237;
assign w6303 = b[38] & w183;
assign w6304 = b[39] & w185;
assign w6305 = w179 & ~w4812;
assign w6306 = ~w6302 & ~w6303;
assign w6307 = ~w6304 & w6306;
assign w6308 = ~w6305 & w6307;
assign w6309 = a[8] & ~w6308;
assign w6310 = ~a[8] & w6308;
assign w6311 = ~w6309 & ~w6310;
assign w6312 = w6301 & w6311;
assign w6313 = ~w6301 & ~w6311;
assign w6314 = ~w6312 & ~w6313;
assign w6315 = ~w6048 & ~w6052;
assign w6316 = w6314 & w6315;
assign w6317 = ~w6314 & ~w6315;
assign w6318 = ~w6316 & ~w6317;
assign w6319 = w6095 & ~w6318;
assign w6320 = ~w6095 & w6318;
assign w6321 = ~w6319 & ~w6320;
assign w6322 = (~w6055 & ~w5827) | (~w6055 & w24661) | (~w5827 & w24661);
assign w6323 = ~w6321 & ~w6322;
assign w6324 = w6321 & w6322;
assign w6325 = ~w6323 & ~w6324;
assign w6326 = b[45] & w11;
assign w6327 = b[44] & w9;
assign w6328 = (~w6064 & w6066) | (~w6064 & w24818) | (w6066 & w24818);
assign w6329 = ~b[44] & ~b[45];
assign w6330 = b[44] & b[45];
assign w6331 = ~w6329 & ~w6330;
assign w6332 = w6328 & ~w6331;
assign w6333 = ~w6328 & w6331;
assign w6334 = ~w6332 & ~w6333;
assign w6335 = w5 & w6334;
assign w6336 = ~w6326 & ~w6327;
assign w6337 = ~w6335 & w6336;
assign w6338 = b[43] & w24;
assign w6339 = a[2] & ~w6338;
assign w6340 = w6337 & ~w6339;
assign w6341 = a[2] & ~w6337;
assign w6342 = ~w6340 & ~w6341;
assign w6343 = ~w6325 & ~w6342;
assign w6344 = w6325 & w6342;
assign w6345 = ~w6343 & ~w6344;
assign w6346 = w6085 & ~w6345;
assign w6347 = ~w6085 & w6345;
assign w6348 = ~w6346 & ~w6347;
assign w6349 = ~w6319 & ~w6324;
assign w6350 = b[41] & w103;
assign w6351 = b[42] & w61;
assign w6352 = b[43] & w68;
assign w6353 = w66 & w5811;
assign w6354 = ~w6351 & ~w6352;
assign w6355 = ~w6350 & w6354;
assign w6356 = ~w6353 & w6355;
assign w6357 = a[5] & ~w6356;
assign w6358 = ~a[5] & w6356;
assign w6359 = ~w6357 & ~w6358;
assign w6360 = b[38] & ~w237;
assign w6361 = b[40] & w185;
assign w6362 = b[39] & w183;
assign w6363 = w179 & ~w5058;
assign w6364 = ~w6360 & ~w6361;
assign w6365 = ~w6362 & w6364;
assign w6366 = ~w6363 & w6365;
assign w6367 = a[8] & ~w6366;
assign w6368 = ~a[8] & w6366;
assign w6369 = ~w6367 & ~w6368;
assign w6370 = ~w6289 & ~w6292;
assign w6371 = b[34] & w575;
assign w6372 = b[32] & ~w649;
assign w6373 = b[33] & w573;
assign w6374 = w569 & ~w3710;
assign w6375 = ~w6371 & ~w6372;
assign w6376 = ~w6373 & w6375;
assign w6377 = ~w6374 & w6376;
assign w6378 = a[14] & ~w6377;
assign w6379 = ~a[14] & w6377;
assign w6380 = ~w6378 & ~w6379;
assign w6381 = ~w6283 & ~w6286;
assign w6382 = b[30] & w838;
assign w6383 = b[31] & w834;
assign w6384 = b[29] & ~w934;
assign w6385 = w832 & ~w3112;
assign w6386 = ~w6382 & ~w6383;
assign w6387 = ~w6384 & w6386;
assign w6388 = ~w6385 & w6387;
assign w6389 = a[17] & ~w6388;
assign w6390 = ~a[17] & w6388;
assign w6391 = ~w6389 & ~w6390;
assign w6392 = b[28] & w1156;
assign w6393 = b[27] & w1154;
assign w6394 = b[26] & ~w1272;
assign w6395 = w1150 & w2559;
assign w6396 = ~w6392 & ~w6393;
assign w6397 = ~w6394 & w6396;
assign w6398 = ~w6395 & w6397;
assign w6399 = a[20] & ~w6398;
assign w6400 = ~a[20] & w6398;
assign w6401 = ~w6399 & ~w6400;
assign w6402 = (~w6259 & ~w6262) | (~w6259 & w24819) | (~w6262 & w24819);
assign w6403 = b[23] & ~w1676;
assign w6404 = b[24] & w1517;
assign w6405 = b[25] & w1519;
assign w6406 = w1513 & w2061;
assign w6407 = ~w6403 & ~w6404;
assign w6408 = ~w6405 & w6407;
assign w6409 = ~w6406 & w6408;
assign w6410 = a[23] & ~w6409;
assign w6411 = ~a[23] & w6409;
assign w6412 = ~w6410 & ~w6411;
assign w6413 = b[20] & ~w2114;
assign w6414 = b[22] & w1957;
assign w6415 = b[21] & w1955;
assign w6416 = w1615 & w1951;
assign w6417 = ~w6413 & ~w6414;
assign w6418 = ~w6415 & w6417;
assign w6419 = ~w6416 & w6418;
assign w6420 = a[26] & ~w6419;
assign w6421 = ~a[26] & w6419;
assign w6422 = ~w6420 & ~w6421;
assign w6423 = (~w6236 & ~w6239) | (~w6236 & w24820) | (~w6239 & w24820);
assign w6424 = b[14] & w3177;
assign w6425 = b[16] & w2978;
assign w6426 = b[15] & w2973;
assign w6427 = w905 & w2980;
assign w6428 = ~w6425 & ~w6426;
assign w6429 = ~w6424 & w6428;
assign w6430 = ~w6427 & w6429;
assign w6431 = a[32] & ~w6430;
assign w6432 = ~a[32] & w6430;
assign w6433 = ~w6431 & ~w6432;
assign w6434 = (~w6224 & w6226) | (~w6224 & w25140) | (w6226 & w25140);
assign w6435 = b[11] & w3785;
assign w6436 = b[12] & w3578;
assign w6437 = b[13] & w3580;
assign w6438 = w628 & w3573;
assign w6439 = ~w6436 & ~w6437;
assign w6440 = ~w6435 & w6439;
assign w6441 = ~w6438 & w6440;
assign w6442 = a[35] & ~w6441;
assign w6443 = ~a[35] & w6441;
assign w6444 = ~w6442 & ~w6443;
assign w6445 = b[8] & w4453;
assign w6446 = b[9] & w4241;
assign w6447 = b[10] & w4243;
assign w6448 = w397 & w4236;
assign w6449 = ~w6446 & ~w6447;
assign w6450 = ~w6445 & w6449;
assign w6451 = ~w6448 & w6450;
assign w6452 = a[38] & ~w6451;
assign w6453 = ~a[38] & w6451;
assign w6454 = ~w6452 & ~w6453;
assign w6455 = w5938 & w24978;
assign w6456 = b[3] & w5670;
assign w6457 = b[4] & w5665;
assign w6458 = w84 & w5663;
assign w6459 = ~w6456 & ~w6457;
assign w6460 = ~w6455 & w6459;
assign w6461 = ~w6458 & w6460;
assign w6462 = a[44] & ~w6461;
assign w6463 = ~a[44] & w6461;
assign w6464 = ~w6462 & ~w6463;
assign w6465 = a[47] & w6163;
assign w6466 = a[46] & ~a[47];
assign w6467 = ~a[46] & a[47];
assign w6468 = ~w6466 & ~w6467;
assign w6469 = ~w6162 & ~w6468;
assign w6470 = ~w8 & w6469;
assign w6471 = a[45] & ~a[46];
assign w6472 = ~a[45] & a[46];
assign w6473 = ~w6471 & ~w6472;
assign w6474 = w6162 & ~w6473;
assign w6475 = b[0] & w6474;
assign w6476 = ~w6162 & w6468;
assign w6477 = b[1] & w6476;
assign w6478 = ~w6470 & ~w6475;
assign w6479 = ~w6477 & w6478;
assign w6480 = ~w6465 & w6479;
assign w6481 = w6465 & ~w6479;
assign w6482 = ~w6480 & ~w6481;
assign w6483 = ~w6464 & ~w6482;
assign w6484 = w6464 & w6482;
assign w6485 = ~w6483 & ~w6484;
assign w6486 = (~w6174 & ~w6176) | (~w6174 & w24821) | (~w6176 & w24821);
assign w6487 = ~w6485 & w6486;
assign w6488 = w6485 & ~w6486;
assign w6489 = ~w6487 & ~w6488;
assign w6490 = b[5] & w5167;
assign w6491 = b[7] & w4925;
assign w6492 = b[6] & w4918;
assign w6493 = w216 & w4923;
assign w6494 = ~w6491 & ~w6492;
assign w6495 = ~w6490 & w6494;
assign w6496 = ~w6493 & w6495;
assign w6497 = a[41] & ~w6496;
assign w6498 = ~a[41] & w6496;
assign w6499 = ~w6497 & ~w6498;
assign w6500 = w6489 & w6499;
assign w6501 = ~w6489 & ~w6499;
assign w6502 = ~w6500 & ~w6501;
assign w6503 = ~w6190 & ~w6195;
assign w6504 = ~w6502 & w6503;
assign w6505 = w6502 & ~w6503;
assign w6506 = ~w6504 & ~w6505;
assign w6507 = w6454 & w6506;
assign w6508 = ~w6454 & ~w6506;
assign w6509 = ~w6507 & ~w6508;
assign w6510 = (~w6208 & w6159) | (~w6208 & w24822) | (w6159 & w24822);
assign w6511 = w6509 & ~w6510;
assign w6512 = ~w6509 & w6510;
assign w6513 = ~w6511 & ~w6512;
assign w6514 = ~w6444 & ~w6513;
assign w6515 = w6444 & w6513;
assign w6516 = ~w6514 & ~w6515;
assign w6517 = w6434 & ~w6516;
assign w6518 = ~w6434 & w6516;
assign w6519 = ~w6517 & ~w6518;
assign w6520 = w6433 & w6519;
assign w6521 = ~w6433 & ~w6519;
assign w6522 = ~w6520 & ~w6521;
assign w6523 = (~w6231 & ~w24817) | (~w6231 & w25141) | (~w24817 & w25141);
assign w6524 = ~w6522 & ~w6523;
assign w6525 = w6522 & w6523;
assign w6526 = ~w6524 & ~w6525;
assign w6527 = b[17] & ~w2622;
assign w6528 = b[18] & w2436;
assign w6529 = b[19] & w2438;
assign w6530 = ~w1231 & w2432;
assign w6531 = ~w6527 & ~w6528;
assign w6532 = ~w6529 & w6531;
assign w6533 = ~w6530 & w6532;
assign w6534 = a[29] & ~w6533;
assign w6535 = ~a[29] & w6533;
assign w6536 = ~w6534 & ~w6535;
assign w6537 = w6526 & w6536;
assign w6538 = ~w6526 & ~w6536;
assign w6539 = ~w6537 & ~w6538;
assign w6540 = ~w6423 & ~w6539;
assign w6541 = w6423 & w6539;
assign w6542 = ~w6540 & ~w6541;
assign w6543 = ~w6422 & w6542;
assign w6544 = w6422 & ~w6542;
assign w6545 = ~w6543 & ~w6544;
assign w6546 = (~w6254 & ~w6138) | (~w6254 & w24823) | (~w6138 & w24823);
assign w6547 = w6545 & w6546;
assign w6548 = ~w6545 & ~w6546;
assign w6549 = ~w6547 & ~w6548;
assign w6550 = w6412 & w6549;
assign w6551 = ~w6412 & ~w6549;
assign w6552 = ~w6550 & ~w6551;
assign w6553 = ~w6402 & w6552;
assign w6554 = w6402 & ~w6552;
assign w6555 = ~w6553 & ~w6554;
assign w6556 = ~w6401 & ~w6555;
assign w6557 = w6401 & w6555;
assign w6558 = ~w6556 & ~w6557;
assign w6559 = (~w6276 & w6127) | (~w6276 & w24381) | (w6127 & w24381);
assign w6560 = w6558 & ~w6559;
assign w6561 = ~w6558 & w6559;
assign w6562 = ~w6560 & ~w6561;
assign w6563 = ~w6391 & ~w6562;
assign w6564 = w6391 & w6562;
assign w6565 = ~w6563 & ~w6564;
assign w6566 = ~w6381 & w6565;
assign w6567 = w6381 & ~w6565;
assign w6568 = ~w6566 & ~w6567;
assign w6569 = w6380 & w6568;
assign w6570 = ~w6380 & ~w6568;
assign w6571 = ~w6569 & ~w6570;
assign w6572 = w6370 & ~w6571;
assign w6573 = ~w6370 & w6571;
assign w6574 = ~w6572 & ~w6573;
assign w6575 = b[37] & w360;
assign w6576 = b[35] & ~w419;
assign w6577 = b[36] & w358;
assign w6578 = w354 & ~w4357;
assign w6579 = ~w6575 & ~w6576;
assign w6580 = ~w6577 & w6579;
assign w6581 = ~w6578 & w6580;
assign w6582 = a[11] & ~w6581;
assign w6583 = ~a[11] & w6581;
assign w6584 = ~w6582 & ~w6583;
assign w6585 = w6574 & w6584;
assign w6586 = ~w6574 & ~w6584;
assign w6587 = ~w6585 & ~w6586;
assign w6588 = (~w6295 & ~w6298) | (~w6295 & w25264) | (~w6298 & w25264);
assign w6589 = w6587 & w6588;
assign w6590 = ~w6587 & ~w6588;
assign w6591 = ~w6589 & ~w6590;
assign w6592 = w6369 & ~w6591;
assign w6593 = ~w6369 & w6591;
assign w6594 = ~w6592 & ~w6593;
assign w6595 = ~w6313 & ~w6316;
assign w6596 = w6594 & w6595;
assign w6597 = ~w6594 & ~w6595;
assign w6598 = ~w6596 & ~w6597;
assign w6599 = w6359 & w6598;
assign w6600 = ~w6359 & ~w6598;
assign w6601 = ~w6599 & ~w6600;
assign w6602 = w6349 & w6601;
assign w6603 = ~w6349 & ~w6601;
assign w6604 = ~w6602 & ~w6603;
assign w6605 = b[46] & w11;
assign w6606 = b[45] & w9;
assign w6607 = ~b[45] & ~b[46];
assign w6608 = b[45] & b[46];
assign w6609 = ~w6607 & ~w6608;
assign w6610 = ~w6330 & ~w6333;
assign w6611 = ~w6609 & ~w6610;
assign w6612 = w6609 & w6610;
assign w6613 = ~w6611 & ~w6612;
assign w6614 = w5 & ~w6613;
assign w6615 = ~w6605 & ~w6606;
assign w6616 = ~w6614 & w6615;
assign w6617 = b[44] & w24;
assign w6618 = a[2] & ~w6617;
assign w6619 = w6616 & ~w6618;
assign w6620 = a[2] & ~w6616;
assign w6621 = ~w6619 & ~w6620;
assign w6622 = ~w6604 & w6621;
assign w6623 = w6604 & ~w6621;
assign w6624 = ~w6622 & ~w6623;
assign w6625 = (~w6344 & w6085) | (~w6344 & w24662) | (w6085 & w24662);
assign w6626 = w6624 & ~w6625;
assign w6627 = ~w6624 & w6625;
assign w6628 = ~w6626 & ~w6627;
assign w6629 = b[42] & w103;
assign w6630 = b[43] & w61;
assign w6631 = b[44] & w68;
assign w6632 = w66 & w6069;
assign w6633 = ~w6630 & ~w6631;
assign w6634 = ~w6629 & w6633;
assign w6635 = ~w6632 & w6634;
assign w6636 = a[5] & ~w6635;
assign w6637 = ~a[5] & w6635;
assign w6638 = ~w6636 & ~w6637;
assign w6639 = (~w6592 & ~w6595) | (~w6592 & w25265) | (~w6595 & w25265);
assign w6640 = b[38] & w360;
assign w6641 = b[37] & w358;
assign w6642 = b[36] & ~w419;
assign w6643 = w354 & w4582;
assign w6644 = ~w6640 & ~w6641;
assign w6645 = ~w6642 & w6644;
assign w6646 = ~w6643 & w6645;
assign w6647 = a[11] & ~w6646;
assign w6648 = ~a[11] & w6646;
assign w6649 = ~w6647 & ~w6648;
assign w6650 = ~w6569 & ~w6573;
assign w6651 = b[34] & w573;
assign w6652 = b[33] & ~w649;
assign w6653 = b[35] & w575;
assign w6654 = w569 & w3918;
assign w6655 = ~w6651 & ~w6652;
assign w6656 = ~w6653 & w6655;
assign w6657 = ~w6654 & w6656;
assign w6658 = a[14] & ~w6657;
assign w6659 = ~a[14] & w6657;
assign w6660 = ~w6658 & ~w6659;
assign w6661 = b[32] & w834;
assign w6662 = b[31] & w838;
assign w6663 = b[30] & ~w934;
assign w6664 = w832 & w3304;
assign w6665 = ~w6661 & ~w6662;
assign w6666 = ~w6663 & w6665;
assign w6667 = ~w6664 & w6666;
assign w6668 = a[17] & ~w6667;
assign w6669 = ~a[17] & w6667;
assign w6670 = ~w6668 & ~w6669;
assign w6671 = (~w6557 & w6559) | (~w6557 & w24824) | (w6559 & w24824);
assign w6672 = b[28] & w1154;
assign w6673 = b[27] & ~w1272;
assign w6674 = b[29] & w1156;
assign w6675 = w1150 & w2734;
assign w6676 = ~w6672 & ~w6673;
assign w6677 = ~w6674 & w6676;
assign w6678 = ~w6675 & w6677;
assign w6679 = a[20] & ~w6678;
assign w6680 = ~a[20] & w6678;
assign w6681 = ~w6679 & ~w6680;
assign w6682 = b[25] & w1517;
assign w6683 = b[24] & ~w1676;
assign w6684 = b[26] & w1519;
assign w6685 = w1513 & w2219;
assign w6686 = ~w6682 & ~w6683;
assign w6687 = ~w6684 & w6686;
assign w6688 = ~w6685 & w6687;
assign w6689 = a[23] & ~w6688;
assign w6690 = ~a[23] & w6688;
assign w6691 = ~w6689 & ~w6690;
assign w6692 = (~w6544 & ~w6546) | (~w6544 & w24663) | (~w6546 & w24663);
assign w6693 = b[18] & ~w2622;
assign w6694 = b[19] & w2436;
assign w6695 = b[20] & w2438;
assign w6696 = w1347 & w2432;
assign w6697 = ~w6693 & ~w6694;
assign w6698 = ~w6695 & w6697;
assign w6699 = ~w6696 & w6698;
assign w6700 = a[29] & ~w6699;
assign w6701 = ~a[29] & w6699;
assign w6702 = ~w6700 & ~w6701;
assign w6703 = (~w6520 & ~w6523) | (~w6520 & w24664) | (~w6523 & w24664);
assign w6704 = b[12] & w3785;
assign w6705 = b[14] & w3580;
assign w6706 = b[13] & w3578;
assign w6707 = w714 & w3573;
assign w6708 = ~w6705 & ~w6706;
assign w6709 = ~w6704 & w6708;
assign w6710 = ~w6707 & w6709;
assign w6711 = a[35] & ~w6710;
assign w6712 = ~a[35] & w6710;
assign w6713 = ~w6711 & ~w6712;
assign w6714 = ~w6507 & ~w6511;
assign w6715 = ~w6484 & ~w6488;
assign w6716 = b[3] & w5939;
assign w6717 = b[5] & w5665;
assign w6718 = b[4] & w5670;
assign w6719 = w116 & w5663;
assign w6720 = ~w6717 & ~w6718;
assign w6721 = ~w6716 & w6720;
assign w6722 = (a[44] & w6719) | (a[44] & w25266) | (w6719 & w25266);
assign w6723 = ~w6719 & w25267;
assign w6724 = ~w6722 & ~w6723;
assign w6725 = a[47] & ~w6163;
assign w6726 = w6478 & w24979;
assign w6727 = a[47] & ~w6726;
assign w6728 = w22 & w6469;
assign w6729 = b[1] & w6474;
assign w6730 = b[2] & w6476;
assign w6731 = w6162 & ~w6468;
assign w6732 = w6473 & w6731;
assign w6733 = b[0] & w6732;
assign w6734 = ~w6728 & ~w6729;
assign w6735 = ~w6730 & w6734;
assign w6736 = ~w6733 & w6735;
assign w6737 = ~w6727 & w6736;
assign w6738 = w6727 & ~w6736;
assign w6739 = ~w6737 & ~w6738;
assign w6740 = w6724 & w6739;
assign w6741 = ~w6724 & ~w6739;
assign w6742 = ~w6740 & ~w6741;
assign w6743 = (w6742 & w6488) | (w6742 & w25268) | (w6488 & w25268);
assign w6744 = ~w6488 & w25269;
assign w6745 = ~w6743 & ~w6744;
assign w6746 = b[6] & w5167;
assign w6747 = b[8] & w4925;
assign w6748 = b[7] & w4918;
assign w6749 = w270 & w4923;
assign w6750 = ~w6747 & ~w6748;
assign w6751 = ~w6746 & w6750;
assign w6752 = ~w6749 & w6751;
assign w6753 = a[41] & ~w6752;
assign w6754 = ~a[41] & w6752;
assign w6755 = ~w6753 & ~w6754;
assign w6756 = ~w6745 & ~w6755;
assign w6757 = w6745 & w6755;
assign w6758 = ~w6756 & ~w6757;
assign w6759 = (~w6500 & w6503) | (~w6500 & w24665) | (w6503 & w24665);
assign w6760 = w6758 & ~w6759;
assign w6761 = ~w6758 & w6759;
assign w6762 = ~w6760 & ~w6761;
assign w6763 = b[9] & w4453;
assign w6764 = b[11] & w4243;
assign w6765 = b[10] & w4241;
assign w6766 = w469 & w4236;
assign w6767 = ~w6764 & ~w6765;
assign w6768 = ~w6763 & w6767;
assign w6769 = ~w6766 & w6768;
assign w6770 = a[38] & ~w6769;
assign w6771 = ~a[38] & w6769;
assign w6772 = ~w6770 & ~w6771;
assign w6773 = ~w6762 & ~w6772;
assign w6774 = w6762 & w6772;
assign w6775 = ~w6773 & ~w6774;
assign w6776 = w6714 & w6775;
assign w6777 = ~w6714 & ~w6775;
assign w6778 = ~w6776 & ~w6777;
assign w6779 = w6713 & ~w6778;
assign w6780 = ~w6713 & w6778;
assign w6781 = ~w6779 & ~w6780;
assign w6782 = (~w6515 & w6434) | (~w6515 & w24666) | (w6434 & w24666);
assign w6783 = w6781 & ~w6782;
assign w6784 = ~w6781 & w6782;
assign w6785 = ~w6783 & ~w6784;
assign w6786 = b[15] & w3177;
assign w6787 = b[17] & w2978;
assign w6788 = b[16] & w2973;
assign w6789 = w1008 & w2980;
assign w6790 = ~w6787 & ~w6788;
assign w6791 = ~w6786 & w6790;
assign w6792 = ~w6789 & w6791;
assign w6793 = a[32] & ~w6792;
assign w6794 = ~a[32] & w6792;
assign w6795 = ~w6793 & ~w6794;
assign w6796 = ~w6785 & ~w6795;
assign w6797 = w6785 & w6795;
assign w6798 = ~w6796 & ~w6797;
assign w6799 = w6703 & w6798;
assign w6800 = ~w6703 & ~w6798;
assign w6801 = ~w6799 & ~w6800;
assign w6802 = w6702 & ~w6801;
assign w6803 = ~w6702 & w6801;
assign w6804 = ~w6802 & ~w6803;
assign w6805 = (~w6538 & ~w6423) | (~w6538 & w25142) | (~w6423 & w25142);
assign w6806 = ~w6804 & ~w6805;
assign w6807 = w6804 & w6805;
assign w6808 = ~w6806 & ~w6807;
assign w6809 = b[23] & w1957;
assign w6810 = b[21] & ~w2114;
assign w6811 = b[22] & w1955;
assign w6812 = w1755 & w1951;
assign w6813 = ~w6809 & ~w6810;
assign w6814 = ~w6811 & w6813;
assign w6815 = ~w6812 & w6814;
assign w6816 = a[26] & ~w6815;
assign w6817 = ~a[26] & w6815;
assign w6818 = ~w6816 & ~w6817;
assign w6819 = ~w6808 & ~w6818;
assign w6820 = w6808 & w6818;
assign w6821 = ~w6819 & ~w6820;
assign w6822 = w6692 & w6821;
assign w6823 = ~w6692 & ~w6821;
assign w6824 = ~w6822 & ~w6823;
assign w6825 = ~w6691 & w6824;
assign w6826 = w6691 & ~w6824;
assign w6827 = ~w6825 & ~w6826;
assign w6828 = (~w6550 & w6402) | (~w6550 & w24667) | (w6402 & w24667);
assign w6829 = w6827 & ~w6828;
assign w6830 = ~w6827 & w6828;
assign w6831 = ~w6829 & ~w6830;
assign w6832 = ~w6681 & ~w6831;
assign w6833 = w6681 & w6831;
assign w6834 = ~w6832 & ~w6833;
assign w6835 = ~w6671 & ~w6834;
assign w6836 = w6671 & w6834;
assign w6837 = ~w6835 & ~w6836;
assign w6838 = ~w6670 & w6837;
assign w6839 = w6670 & ~w6837;
assign w6840 = ~w6838 & ~w6839;
assign w6841 = (~w6564 & w6381) | (~w6564 & w24382) | (w6381 & w24382);
assign w6842 = w6840 & ~w6841;
assign w6843 = ~w6840 & w6841;
assign w6844 = ~w6842 & ~w6843;
assign w6845 = w6660 & w6844;
assign w6846 = ~w6660 & ~w6844;
assign w6847 = ~w6845 & ~w6846;
assign w6848 = ~w6650 & w6847;
assign w6849 = w6650 & ~w6847;
assign w6850 = ~w6848 & ~w6849;
assign w6851 = w6649 & w6850;
assign w6852 = ~w6649 & ~w6850;
assign w6853 = ~w6851 & ~w6852;
assign w6854 = ~w6586 & ~w6589;
assign w6855 = ~w6853 & ~w6854;
assign w6856 = w6853 & w6854;
assign w6857 = ~w6855 & ~w6856;
assign w6858 = b[41] & w185;
assign w6859 = b[39] & ~w237;
assign w6860 = b[40] & w183;
assign w6861 = w179 & w5302;
assign w6862 = ~w6858 & ~w6859;
assign w6863 = ~w6860 & w6862;
assign w6864 = ~w6861 & w6863;
assign w6865 = a[8] & ~w6864;
assign w6866 = ~a[8] & w6864;
assign w6867 = ~w6865 & ~w6866;
assign w6868 = w6857 & w6867;
assign w6869 = ~w6857 & ~w6867;
assign w6870 = ~w6868 & ~w6869;
assign w6871 = w6639 & w6870;
assign w6872 = ~w6639 & ~w6870;
assign w6873 = ~w6871 & ~w6872;
assign w6874 = ~w6638 & w6873;
assign w6875 = w6638 & ~w6873;
assign w6876 = ~w6874 & ~w6875;
assign w6877 = ~w6600 & ~w6602;
assign w6878 = w6876 & w6877;
assign w6879 = ~w6876 & ~w6877;
assign w6880 = ~w6878 & ~w6879;
assign w6881 = b[47] & w11;
assign w6882 = b[46] & w9;
assign w6883 = ~b[46] & ~b[47];
assign w6884 = b[46] & b[47];
assign w6885 = ~w6883 & ~w6884;
assign w6886 = (~w6607 & ~w6610) | (~w6607 & w24668) | (~w6610 & w24668);
assign w6887 = ~w6885 & ~w6886;
assign w6888 = w6885 & w6886;
assign w6889 = ~w6887 & ~w6888;
assign w6890 = w5 & w6889;
assign w6891 = ~w6881 & ~w6882;
assign w6892 = ~w6890 & w6891;
assign w6893 = b[45] & w24;
assign w6894 = a[2] & ~w6893;
assign w6895 = w6892 & ~w6894;
assign w6896 = a[2] & ~w6892;
assign w6897 = ~w6895 & ~w6896;
assign w6898 = w6880 & w6897;
assign w6899 = ~w6880 & ~w6897;
assign w6900 = ~w6898 & ~w6899;
assign w6901 = ~w6622 & ~w6626;
assign w6902 = ~w6900 & ~w6901;
assign w6903 = w6900 & w6901;
assign w6904 = ~w6902 & ~w6903;
assign w6905 = (~w6875 & ~w6877) | (~w6875 & w25270) | (~w6877 & w25270);
assign w6906 = b[43] & w103;
assign w6907 = b[44] & w61;
assign w6908 = b[45] & w68;
assign w6909 = w66 & w6334;
assign w6910 = ~w6907 & ~w6908;
assign w6911 = ~w6906 & w6910;
assign w6912 = ~w6909 & w6911;
assign w6913 = a[5] & ~w6912;
assign w6914 = ~a[5] & w6912;
assign w6915 = ~w6913 & ~w6914;
assign w6916 = b[41] & w183;
assign w6917 = b[40] & ~w237;
assign w6918 = b[42] & w185;
assign w6919 = w179 & w5548;
assign w6920 = ~w6916 & ~w6917;
assign w6921 = ~w6918 & w6920;
assign w6922 = ~w6919 & w6921;
assign w6923 = a[8] & ~w6922;
assign w6924 = ~a[8] & w6922;
assign w6925 = ~w6923 & ~w6924;
assign w6926 = (~w6845 & w6650) | (~w6845 & w24383) | (w6650 & w24383);
assign w6927 = b[34] & ~w649;
assign w6928 = b[36] & w575;
assign w6929 = b[35] & w573;
assign w6930 = w569 & w4129;
assign w6931 = ~w6927 & ~w6928;
assign w6932 = ~w6929 & w6931;
assign w6933 = ~w6930 & w6932;
assign w6934 = a[14] & ~w6933;
assign w6935 = ~a[14] & w6933;
assign w6936 = ~w6934 & ~w6935;
assign w6937 = (~w6839 & w6841) | (~w6839 & w24825) | (w6841 & w24825);
assign w6938 = b[28] & ~w1272;
assign w6939 = b[30] & w1156;
assign w6940 = b[29] & w1154;
assign w6941 = w1150 & ~w2908;
assign w6942 = ~w6938 & ~w6939;
assign w6943 = ~w6940 & w6942;
assign w6944 = ~w6941 & w6943;
assign w6945 = a[20] & ~w6944;
assign w6946 = ~a[20] & w6944;
assign w6947 = ~w6945 & ~w6946;
assign w6948 = ~w6826 & ~w6829;
assign w6949 = b[25] & ~w1676;
assign w6950 = b[26] & w1517;
assign w6951 = b[27] & w1519;
assign w6952 = w1513 & w2378;
assign w6953 = ~w6949 & ~w6950;
assign w6954 = ~w6951 & w6953;
assign w6955 = ~w6952 & w6954;
assign w6956 = a[23] & ~w6955;
assign w6957 = ~a[23] & w6955;
assign w6958 = ~w6956 & ~w6957;
assign w6959 = (~w6819 & ~w6692) | (~w6819 & w25271) | (~w6692 & w25271);
assign w6960 = b[23] & w1955;
assign w6961 = b[24] & w1957;
assign w6962 = b[22] & ~w2114;
assign w6963 = w1895 & w1951;
assign w6964 = ~w6960 & ~w6961;
assign w6965 = ~w6962 & w6964;
assign w6966 = ~w6963 & w6965;
assign w6967 = a[26] & ~w6966;
assign w6968 = ~a[26] & w6966;
assign w6969 = ~w6967 & ~w6968;
assign w6970 = (~w6802 & ~w6805) | (~w6802 & w24669) | (~w6805 & w24669);
assign w6971 = b[16] & w3177;
assign w6972 = b[18] & w2978;
assign w6973 = b[17] & w2973;
assign w6974 = ~w1108 & w2980;
assign w6975 = ~w6972 & ~w6973;
assign w6976 = ~w6971 & w6975;
assign w6977 = ~w6974 & w6976;
assign w6978 = a[32] & ~w6977;
assign w6979 = ~a[32] & w6977;
assign w6980 = ~w6978 & ~w6979;
assign w6981 = ~w6779 & ~w6783;
assign w6982 = b[13] & w3785;
assign w6983 = b[14] & w3578;
assign w6984 = b[15] & w3580;
assign w6985 = ~w799 & w3573;
assign w6986 = ~w6983 & ~w6984;
assign w6987 = ~w6982 & w6986;
assign w6988 = ~w6985 & w6987;
assign w6989 = a[35] & ~w6988;
assign w6990 = ~a[35] & w6988;
assign w6991 = ~w6989 & ~w6990;
assign w6992 = (~w6757 & w6759) | (~w6757 & w25272) | (w6759 & w25272);
assign w6993 = a[47] & ~a[48];
assign w6994 = ~a[47] & a[48];
assign w6995 = ~w6993 & ~w6994;
assign w6996 = b[0] & ~w6995;
assign w6997 = w6726 & w6736;
assign w6998 = w6731 & w24826;
assign w6999 = b[3] & w6476;
assign w7000 = b[2] & w6474;
assign w7001 = ~w6999 & ~w7000;
assign w7002 = ~w6998 & w7001;
assign w7003 = (a[47] & ~w7002) | (a[47] & w24827) | (~w7002 & w24827);
assign w7004 = w7002 & w24828;
assign w7005 = ~w7003 & ~w7004;
assign w7006 = w6997 & w7005;
assign w7007 = ~w6997 & ~w7005;
assign w7008 = ~w7006 & ~w7007;
assign w7009 = w6996 & w7008;
assign w7010 = ~w6996 & ~w7008;
assign w7011 = ~w7009 & ~w7010;
assign w7012 = b[4] & w5939;
assign w7013 = b[6] & w5665;
assign w7014 = b[5] & w5670;
assign w7015 = w157 & w5663;
assign w7016 = ~w7013 & ~w7014;
assign w7017 = ~w7012 & w7016;
assign w7018 = ~w7015 & w7017;
assign w7019 = a[44] & ~w7018;
assign w7020 = ~a[44] & w7018;
assign w7021 = ~w7019 & ~w7020;
assign w7022 = w7011 & w7021;
assign w7023 = ~w7011 & ~w7021;
assign w7024 = ~w7022 & ~w7023;
assign w7025 = (~w6740 & w6715) | (~w6740 & w24980) | (w6715 & w24980);
assign w7026 = ~w7024 & w7025;
assign w7027 = w7024 & ~w7025;
assign w7028 = ~w7026 & ~w7027;
assign w7029 = b[7] & w5167;
assign w7030 = b[8] & w4918;
assign w7031 = b[9] & w4925;
assign w7032 = w322 & w4923;
assign w7033 = ~w7030 & ~w7031;
assign w7034 = ~w7029 & w7033;
assign w7035 = ~w7032 & w7034;
assign w7036 = a[41] & ~w7035;
assign w7037 = ~a[41] & w7035;
assign w7038 = ~w7036 & ~w7037;
assign w7039 = w7028 & w7038;
assign w7040 = ~w7028 & ~w7038;
assign w7041 = ~w7039 & ~w7040;
assign w7042 = w6992 & ~w7041;
assign w7043 = ~w6992 & w7041;
assign w7044 = ~w7042 & ~w7043;
assign w7045 = b[10] & w4453;
assign w7046 = b[12] & w4243;
assign w7047 = b[11] & w4241;
assign w7048 = w536 & w4236;
assign w7049 = ~w7046 & ~w7047;
assign w7050 = ~w7045 & w7049;
assign w7051 = ~w7048 & w7050;
assign w7052 = a[38] & ~w7051;
assign w7053 = ~a[38] & w7051;
assign w7054 = ~w7052 & ~w7053;
assign w7055 = ~w7044 & ~w7054;
assign w7056 = w7044 & w7054;
assign w7057 = ~w7055 & ~w7056;
assign w7058 = (~w6773 & ~w6714) | (~w6773 & w24670) | (~w6714 & w24670);
assign w7059 = w7057 & w7058;
assign w7060 = ~w7057 & ~w7058;
assign w7061 = ~w7059 & ~w7060;
assign w7062 = w6991 & w7061;
assign w7063 = ~w6991 & ~w7061;
assign w7064 = ~w7062 & ~w7063;
assign w7065 = ~w6981 & ~w7064;
assign w7066 = w6981 & w7064;
assign w7067 = ~w7065 & ~w7066;
assign w7068 = w6980 & ~w7067;
assign w7069 = ~w6980 & w7067;
assign w7070 = ~w7068 & ~w7069;
assign w7071 = ~w6796 & ~w6799;
assign w7072 = ~w7070 & ~w7071;
assign w7073 = w7070 & w7071;
assign w7074 = ~w7072 & ~w7073;
assign w7075 = b[21] & w2438;
assign w7076 = b[20] & w2436;
assign w7077 = b[19] & ~w2622;
assign w7078 = w1467 & w2432;
assign w7079 = ~w7075 & ~w7076;
assign w7080 = ~w7077 & w7079;
assign w7081 = ~w7078 & w7080;
assign w7082 = a[29] & ~w7081;
assign w7083 = ~a[29] & w7081;
assign w7084 = ~w7082 & ~w7083;
assign w7085 = w7074 & w7084;
assign w7086 = ~w7074 & ~w7084;
assign w7087 = ~w7085 & ~w7086;
assign w7088 = w6970 & w7087;
assign w7089 = ~w6970 & ~w7087;
assign w7090 = ~w7088 & ~w7089;
assign w7091 = w6969 & ~w7090;
assign w7092 = ~w6969 & w7090;
assign w7093 = ~w7091 & ~w7092;
assign w7094 = w6959 & w7093;
assign w7095 = ~w6959 & ~w7093;
assign w7096 = ~w7094 & ~w7095;
assign w7097 = w6958 & w7096;
assign w7098 = ~w6958 & ~w7096;
assign w7099 = ~w7097 & ~w7098;
assign w7100 = ~w6948 & w7099;
assign w7101 = w6948 & ~w7099;
assign w7102 = ~w7100 & ~w7101;
assign w7103 = w6947 & w7102;
assign w7104 = ~w6947 & ~w7102;
assign w7105 = ~w7103 & ~w7104;
assign w7106 = (~w6832 & ~w6671) | (~w6832 & w24671) | (~w6671 & w24671);
assign w7107 = w7105 & w7106;
assign w7108 = ~w7105 & ~w7106;
assign w7109 = ~w7107 & ~w7108;
assign w7110 = b[31] & ~w934;
assign w7111 = b[32] & w838;
assign w7112 = b[33] & w834;
assign w7113 = w832 & w3499;
assign w7114 = ~w7110 & ~w7111;
assign w7115 = ~w7112 & w7114;
assign w7116 = ~w7113 & w7115;
assign w7117 = a[17] & ~w7116;
assign w7118 = ~a[17] & w7116;
assign w7119 = ~w7117 & ~w7118;
assign w7120 = w7109 & w7119;
assign w7121 = ~w7109 & ~w7119;
assign w7122 = ~w7120 & ~w7121;
assign w7123 = w6937 & ~w7122;
assign w7124 = ~w6937 & w7122;
assign w7125 = ~w7123 & ~w7124;
assign w7126 = ~w6936 & ~w7125;
assign w7127 = w6936 & w7125;
assign w7128 = ~w7126 & ~w7127;
assign w7129 = w6926 & ~w7128;
assign w7130 = ~w6926 & w7128;
assign w7131 = ~w7129 & ~w7130;
assign w7132 = b[38] & w358;
assign w7133 = b[39] & w360;
assign w7134 = b[37] & ~w419;
assign w7135 = w354 & ~w4812;
assign w7136 = ~w7132 & ~w7133;
assign w7137 = ~w7134 & w7136;
assign w7138 = ~w7135 & w7137;
assign w7139 = a[11] & ~w7138;
assign w7140 = ~a[11] & w7138;
assign w7141 = ~w7139 & ~w7140;
assign w7142 = w7131 & w7141;
assign w7143 = ~w7131 & ~w7141;
assign w7144 = ~w7142 & ~w7143;
assign w7145 = ~w6851 & ~w6856;
assign w7146 = w7144 & w7145;
assign w7147 = ~w7144 & ~w7145;
assign w7148 = ~w7146 & ~w7147;
assign w7149 = w6925 & ~w7148;
assign w7150 = ~w6925 & w7148;
assign w7151 = ~w7149 & ~w7150;
assign w7152 = ~w6869 & ~w6871;
assign w7153 = w7151 & w7152;
assign w7154 = ~w7151 & ~w7152;
assign w7155 = ~w7153 & ~w7154;
assign w7156 = w6915 & w7155;
assign w7157 = ~w6915 & ~w7155;
assign w7158 = ~w7156 & ~w7157;
assign w7159 = w6905 & w7158;
assign w7160 = ~w6905 & ~w7158;
assign w7161 = ~w7159 & ~w7160;
assign w7162 = b[48] & w11;
assign w7163 = b[47] & w9;
assign w7164 = ~w6884 & ~w6888;
assign w7165 = ~b[47] & ~b[48];
assign w7166 = b[47] & b[48];
assign w7167 = ~w7165 & ~w7166;
assign w7168 = ~w7164 & ~w7167;
assign w7169 = w7164 & w7167;
assign w7170 = ~w7168 & ~w7169;
assign w7171 = w5 & ~w7170;
assign w7172 = ~w7162 & ~w7163;
assign w7173 = ~w7171 & w7172;
assign w7174 = b[46] & w24;
assign w7175 = a[2] & ~w7174;
assign w7176 = w7173 & ~w7175;
assign w7177 = a[2] & ~w7173;
assign w7178 = ~w7176 & ~w7177;
assign w7179 = w7161 & ~w7178;
assign w7180 = ~w7161 & w7178;
assign w7181 = ~w7179 & ~w7180;
assign w7182 = ~w6899 & ~w6903;
assign w7183 = w7181 & w7182;
assign w7184 = ~w7181 & ~w7182;
assign w7185 = ~w7183 & ~w7184;
assign w7186 = (~w7180 & ~w7182) | (~w7180 & w25273) | (~w7182 & w25273);
assign w7187 = b[44] & w103;
assign w7188 = b[46] & w68;
assign w7189 = b[45] & w61;
assign w7190 = w66 & ~w6613;
assign w7191 = ~w7188 & ~w7189;
assign w7192 = ~w7187 & w7191;
assign w7193 = ~w7190 & w7192;
assign w7194 = a[5] & ~w7193;
assign w7195 = ~a[5] & w7193;
assign w7196 = ~w7194 & ~w7195;
assign w7197 = b[38] & ~w419;
assign w7198 = b[40] & w360;
assign w7199 = b[39] & w358;
assign w7200 = w354 & ~w5058;
assign w7201 = ~w7197 & ~w7198;
assign w7202 = ~w7199 & w7201;
assign w7203 = ~w7200 & w7202;
assign w7204 = a[11] & ~w7203;
assign w7205 = ~a[11] & w7203;
assign w7206 = ~w7204 & ~w7205;
assign w7207 = (~w7127 & w6926) | (~w7127 & w24829) | (w6926 & w24829);
assign w7208 = b[36] & w573;
assign w7209 = b[35] & ~w649;
assign w7210 = b[37] & w575;
assign w7211 = w569 & ~w4357;
assign w7212 = ~w7208 & ~w7209;
assign w7213 = ~w7210 & w7212;
assign w7214 = ~w7211 & w7213;
assign w7215 = a[14] & ~w7214;
assign w7216 = ~a[14] & w7214;
assign w7217 = ~w7215 & ~w7216;
assign w7218 = b[34] & w834;
assign w7219 = b[32] & ~w934;
assign w7220 = b[33] & w838;
assign w7221 = w832 & ~w3710;
assign w7222 = ~w7218 & ~w7219;
assign w7223 = ~w7220 & w7222;
assign w7224 = ~w7221 & w7223;
assign w7225 = a[17] & ~w7224;
assign w7226 = ~a[17] & w7224;
assign w7227 = ~w7225 & ~w7226;
assign w7228 = ~w7103 & ~w7107;
assign w7229 = b[29] & ~w1272;
assign w7230 = b[31] & w1156;
assign w7231 = b[30] & w1154;
assign w7232 = w1150 & ~w3112;
assign w7233 = ~w7229 & ~w7230;
assign w7234 = ~w7231 & w7233;
assign w7235 = ~w7232 & w7234;
assign w7236 = a[20] & ~w7235;
assign w7237 = ~a[20] & w7235;
assign w7238 = ~w7236 & ~w7237;
assign w7239 = (~w7097 & w6948) | (~w7097 & w25274) | (w6948 & w25274);
assign w7240 = b[26] & ~w1676;
assign w7241 = b[28] & w1519;
assign w7242 = b[27] & w1517;
assign w7243 = w1513 & w2559;
assign w7244 = ~w7240 & ~w7241;
assign w7245 = ~w7242 & w7244;
assign w7246 = ~w7243 & w7245;
assign w7247 = a[23] & ~w7246;
assign w7248 = ~a[23] & w7246;
assign w7249 = ~w7247 & ~w7248;
assign w7250 = (~w7091 & ~w6959) | (~w7091 & w25420) | (~w6959 & w25420);
assign w7251 = b[20] & ~w2622;
assign w7252 = b[21] & w2436;
assign w7253 = b[22] & w2438;
assign w7254 = w1615 & w2432;
assign w7255 = ~w7251 & ~w7252;
assign w7256 = ~w7253 & w7255;
assign w7257 = ~w7254 & w7256;
assign w7258 = a[29] & ~w7257;
assign w7259 = ~a[29] & w7257;
assign w7260 = ~w7258 & ~w7259;
assign w7261 = b[17] & w3177;
assign w7262 = b[18] & w2973;
assign w7263 = b[19] & w2978;
assign w7264 = ~w1231 & w2980;
assign w7265 = ~w7262 & ~w7263;
assign w7266 = ~w7261 & w7265;
assign w7267 = ~w7264 & w7266;
assign w7268 = a[32] & ~w7267;
assign w7269 = ~a[32] & w7267;
assign w7270 = ~w7268 & ~w7269;
assign w7271 = (~w7056 & ~w7058) | (~w7056 & w25275) | (~w7058 & w25275);
assign w7272 = b[11] & w4453;
assign w7273 = b[13] & w4243;
assign w7274 = b[12] & w4241;
assign w7275 = w628 & w4236;
assign w7276 = ~w7273 & ~w7274;
assign w7277 = ~w7272 & w7276;
assign w7278 = ~w7275 & w7277;
assign w7279 = a[38] & ~w7278;
assign w7280 = ~a[38] & w7278;
assign w7281 = ~w7279 & ~w7280;
assign w7282 = (~w7039 & w6992) | (~w7039 & w25143) | (w6992 & w25143);
assign w7283 = b[8] & w5167;
assign w7284 = b[9] & w4918;
assign w7285 = b[10] & w4925;
assign w7286 = w397 & w4923;
assign w7287 = ~w7284 & ~w7285;
assign w7288 = ~w7283 & w7287;
assign w7289 = ~w7286 & w7288;
assign w7290 = a[41] & ~w7289;
assign w7291 = ~a[41] & w7289;
assign w7292 = ~w7290 & ~w7291;
assign w7293 = w6731 & w25276;
assign w7294 = b[4] & w6476;
assign w7295 = b[3] & w6474;
assign w7296 = w84 & w6469;
assign w7297 = ~w7294 & ~w7295;
assign w7298 = ~w7293 & w7297;
assign w7299 = ~w7296 & w7298;
assign w7300 = a[47] & ~w7299;
assign w7301 = ~a[47] & w7299;
assign w7302 = ~w7300 & ~w7301;
assign w7303 = a[50] & w6996;
assign w7304 = a[48] & ~a[49];
assign w7305 = ~a[48] & a[49];
assign w7306 = ~w7304 & ~w7305;
assign w7307 = w6995 & ~w7306;
assign w7308 = b[0] & w7307;
assign w7309 = a[49] & ~a[50];
assign w7310 = ~a[49] & a[50];
assign w7311 = ~w7309 & ~w7310;
assign w7312 = ~w6995 & ~w7311;
assign w7313 = ~w8 & w7312;
assign w7314 = ~w6995 & w7311;
assign w7315 = b[1] & w7314;
assign w7316 = ~w7308 & ~w7313;
assign w7317 = ~w7315 & w7316;
assign w7318 = w7303 & ~w7317;
assign w7319 = ~w7303 & w7317;
assign w7320 = ~w7318 & ~w7319;
assign w7321 = ~w7302 & ~w7320;
assign w7322 = w7302 & w7320;
assign w7323 = ~w7321 & ~w7322;
assign w7324 = (~w7006 & ~w7008) | (~w7006 & w24981) | (~w7008 & w24981);
assign w7325 = w7323 & ~w7324;
assign w7326 = ~w7323 & w7324;
assign w7327 = ~w7325 & ~w7326;
assign w7328 = b[5] & w5939;
assign w7329 = b[7] & w5665;
assign w7330 = b[6] & w5670;
assign w7331 = w216 & w5663;
assign w7332 = ~w7329 & ~w7330;
assign w7333 = ~w7328 & w7332;
assign w7334 = ~w7331 & w7333;
assign w7335 = a[44] & ~w7334;
assign w7336 = ~a[44] & w7334;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = w7327 & w7337;
assign w7339 = ~w7327 & ~w7337;
assign w7340 = ~w7338 & ~w7339;
assign w7341 = ~w7022 & ~w7027;
assign w7342 = w7340 & w7341;
assign w7343 = ~w7340 & ~w7341;
assign w7344 = ~w7342 & ~w7343;
assign w7345 = w7292 & ~w7344;
assign w7346 = ~w7292 & w7344;
assign w7347 = ~w7345 & ~w7346;
assign w7348 = ~w7282 & w7347;
assign w7349 = w7282 & ~w7347;
assign w7350 = ~w7348 & ~w7349;
assign w7351 = w7281 & w7350;
assign w7352 = ~w7281 & ~w7350;
assign w7353 = ~w7351 & ~w7352;
assign w7354 = ~w7271 & w7353;
assign w7355 = w7271 & ~w7353;
assign w7356 = ~w7354 & ~w7355;
assign w7357 = b[14] & w3785;
assign w7358 = b[15] & w3578;
assign w7359 = b[16] & w3580;
assign w7360 = w905 & w3573;
assign w7361 = ~w7358 & ~w7359;
assign w7362 = ~w7357 & w7361;
assign w7363 = ~w7360 & w7362;
assign w7364 = a[35] & ~w7363;
assign w7365 = ~a[35] & w7363;
assign w7366 = ~w7364 & ~w7365;
assign w7367 = w7356 & w7366;
assign w7368 = ~w7356 & ~w7366;
assign w7369 = ~w7367 & ~w7368;
assign w7370 = (~w7063 & ~w6981) | (~w7063 & w25144) | (~w6981 & w25144);
assign w7371 = w7369 & w7370;
assign w7372 = ~w7369 & ~w7370;
assign w7373 = ~w7371 & ~w7372;
assign w7374 = w7270 & w7373;
assign w7375 = ~w7270 & ~w7373;
assign w7376 = ~w7374 & ~w7375;
assign w7377 = ~w7068 & ~w7073;
assign w7378 = ~w7376 & ~w7377;
assign w7379 = w7376 & w7377;
assign w7380 = ~w7378 & ~w7379;
assign w7381 = w7260 & ~w7380;
assign w7382 = ~w7260 & w7380;
assign w7383 = ~w7381 & ~w7382;
assign w7384 = ~w7086 & ~w7088;
assign w7385 = ~w7383 & ~w7384;
assign w7386 = w7383 & w7384;
assign w7387 = ~w7385 & ~w7386;
assign w7388 = b[23] & ~w2114;
assign w7389 = b[25] & w1957;
assign w7390 = b[24] & w1955;
assign w7391 = w1951 & w2061;
assign w7392 = ~w7388 & ~w7389;
assign w7393 = ~w7390 & w7392;
assign w7394 = ~w7391 & w7393;
assign w7395 = a[26] & ~w7394;
assign w7396 = ~a[26] & w7394;
assign w7397 = ~w7395 & ~w7396;
assign w7398 = w7387 & w7397;
assign w7399 = ~w7387 & ~w7397;
assign w7400 = ~w7398 & ~w7399;
assign w7401 = w7250 & w7400;
assign w7402 = ~w7250 & ~w7400;
assign w7403 = ~w7401 & ~w7402;
assign w7404 = w7249 & ~w7403;
assign w7405 = ~w7249 & w7403;
assign w7406 = ~w7404 & ~w7405;
assign w7407 = ~w7239 & w7406;
assign w7408 = w7239 & ~w7406;
assign w7409 = ~w7407 & ~w7408;
assign w7410 = w7238 & w7409;
assign w7411 = ~w7238 & ~w7409;
assign w7412 = ~w7410 & ~w7411;
assign w7413 = ~w7228 & ~w7412;
assign w7414 = w7228 & w7412;
assign w7415 = ~w7413 & ~w7414;
assign w7416 = w7227 & ~w7415;
assign w7417 = ~w7227 & w7415;
assign w7418 = ~w7416 & ~w7417;
assign w7419 = (~w7120 & w6937) | (~w7120 & w24672) | (w6937 & w24672);
assign w7420 = w7418 & ~w7419;
assign w7421 = ~w7418 & w7419;
assign w7422 = ~w7420 & ~w7421;
assign w7423 = w7217 & w7422;
assign w7424 = ~w7217 & ~w7422;
assign w7425 = ~w7423 & ~w7424;
assign w7426 = ~w7207 & w7425;
assign w7427 = w7207 & ~w7425;
assign w7428 = ~w7426 & ~w7427;
assign w7429 = w7206 & w7428;
assign w7430 = ~w7206 & ~w7428;
assign w7431 = ~w7429 & ~w7430;
assign w7432 = (~w7143 & ~w7145) | (~w7143 & w24384) | (~w7145 & w24384);
assign w7433 = ~w7431 & ~w7432;
assign w7434 = w7431 & w7432;
assign w7435 = ~w7433 & ~w7434;
assign w7436 = b[43] & w185;
assign w7437 = b[41] & ~w237;
assign w7438 = b[42] & w183;
assign w7439 = w179 & w5811;
assign w7440 = ~w7436 & ~w7437;
assign w7441 = ~w7438 & w7440;
assign w7442 = ~w7439 & w7441;
assign w7443 = a[8] & ~w7442;
assign w7444 = ~a[8] & w7442;
assign w7445 = ~w7443 & ~w7444;
assign w7446 = w7435 & w7445;
assign w7447 = ~w7435 & ~w7445;
assign w7448 = ~w7446 & ~w7447;
assign w7449 = ~w7149 & ~w7153;
assign w7450 = w7448 & w7449;
assign w7451 = ~w7448 & ~w7449;
assign w7452 = ~w7450 & ~w7451;
assign w7453 = w7196 & ~w7452;
assign w7454 = ~w7196 & w7452;
assign w7455 = ~w7453 & ~w7454;
assign w7456 = ~w7157 & ~w7159;
assign w7457 = ~w7455 & ~w7456;
assign w7458 = w7455 & w7456;
assign w7459 = ~w7457 & ~w7458;
assign w7460 = b[49] & w11;
assign w7461 = b[48] & w9;
assign w7462 = ~b[48] & ~b[49];
assign w7463 = b[48] & b[49];
assign w7464 = ~w7462 & ~w7463;
assign w7465 = ~w7165 & ~w7169;
assign w7466 = ~w7464 & w7465;
assign w7467 = w7464 & ~w7465;
assign w7468 = ~w7466 & ~w7467;
assign w7469 = w5 & ~w7468;
assign w7470 = ~w7460 & ~w7461;
assign w7471 = ~w7469 & w7470;
assign w7472 = b[47] & w24;
assign w7473 = a[2] & ~w7472;
assign w7474 = w7471 & ~w7473;
assign w7475 = a[2] & ~w7471;
assign w7476 = ~w7474 & ~w7475;
assign w7477 = ~w7459 & ~w7476;
assign w7478 = w7459 & w7476;
assign w7479 = ~w7477 & ~w7478;
assign w7480 = w7186 & ~w7479;
assign w7481 = ~w7186 & w7479;
assign w7482 = ~w7480 & ~w7481;
assign w7483 = b[45] & w103;
assign w7484 = b[46] & w61;
assign w7485 = b[47] & w68;
assign w7486 = w66 & w6889;
assign w7487 = ~w7484 & ~w7485;
assign w7488 = ~w7483 & w7487;
assign w7489 = ~w7486 & w7488;
assign w7490 = a[5] & ~w7489;
assign w7491 = ~a[5] & w7489;
assign w7492 = ~w7490 & ~w7491;
assign w7493 = b[44] & w185;
assign w7494 = b[42] & ~w237;
assign w7495 = b[43] & w183;
assign w7496 = w179 & w6069;
assign w7497 = ~w7493 & ~w7494;
assign w7498 = ~w7495 & w7497;
assign w7499 = ~w7496 & w7498;
assign w7500 = a[8] & ~w7499;
assign w7501 = ~a[8] & w7499;
assign w7502 = ~w7500 & ~w7501;
assign w7503 = (~w7423 & w7207) | (~w7423 & w24673) | (w7207 & w24673);
assign w7504 = b[36] & ~w649;
assign w7505 = b[38] & w575;
assign w7506 = b[37] & w573;
assign w7507 = w569 & w4582;
assign w7508 = ~w7504 & ~w7505;
assign w7509 = ~w7506 & w7508;
assign w7510 = ~w7507 & w7509;
assign w7511 = a[14] & ~w7510;
assign w7512 = ~a[14] & w7510;
assign w7513 = ~w7511 & ~w7512;
assign w7514 = ~w7416 & ~w7420;
assign w7515 = b[30] & ~w1272;
assign w7516 = b[31] & w1154;
assign w7517 = b[32] & w1156;
assign w7518 = w1150 & w3304;
assign w7519 = ~w7515 & ~w7516;
assign w7520 = ~w7517 & w7519;
assign w7521 = ~w7518 & w7520;
assign w7522 = a[20] & ~w7521;
assign w7523 = ~a[20] & w7521;
assign w7524 = ~w7522 & ~w7523;
assign w7525 = (~w7404 & w7239) | (~w7404 & w25421) | (w7239 & w25421);
assign w7526 = b[28] & w1517;
assign w7527 = b[27] & ~w1676;
assign w7528 = b[29] & w1519;
assign w7529 = w1513 & w2734;
assign w7530 = ~w7526 & ~w7527;
assign w7531 = ~w7528 & w7530;
assign w7532 = ~w7529 & w7531;
assign w7533 = a[23] & ~w7532;
assign w7534 = ~a[23] & w7532;
assign w7535 = ~w7533 & ~w7534;
assign w7536 = b[24] & ~w2114;
assign w7537 = b[25] & w1955;
assign w7538 = b[26] & w1957;
assign w7539 = w1951 & w2219;
assign w7540 = ~w7536 & ~w7537;
assign w7541 = ~w7538 & w7540;
assign w7542 = ~w7539 & w7541;
assign w7543 = a[26] & ~w7542;
assign w7544 = ~a[26] & w7542;
assign w7545 = ~w7543 & ~w7544;
assign w7546 = ~w7381 & ~w7386;
assign w7547 = (~w7367 & ~w7370) | (~w7367 & w25422) | (~w7370 & w25422);
assign w7548 = b[15] & w3785;
assign w7549 = b[17] & w3580;
assign w7550 = b[16] & w3578;
assign w7551 = w1008 & w3573;
assign w7552 = ~w7549 & ~w7550;
assign w7553 = ~w7548 & w7552;
assign w7554 = ~w7551 & w7553;
assign w7555 = a[35] & ~w7554;
assign w7556 = ~a[35] & w7554;
assign w7557 = ~w7555 & ~w7556;
assign w7558 = (~w7351 & w7271) | (~w7351 & w25145) | (w7271 & w25145);
assign w7559 = b[12] & w4453;
assign w7560 = b[13] & w4241;
assign w7561 = b[14] & w4243;
assign w7562 = w714 & w4236;
assign w7563 = ~w7560 & ~w7561;
assign w7564 = ~w7559 & w7563;
assign w7565 = ~w7562 & w7564;
assign w7566 = a[38] & ~w7565;
assign w7567 = ~a[38] & w7565;
assign w7568 = ~w7566 & ~w7567;
assign w7569 = ~w7345 & ~w7348;
assign w7570 = ~w7322 & ~w7325;
assign w7571 = w6731 & w25423;
assign w7572 = b[5] & w6476;
assign w7573 = b[4] & w6474;
assign w7574 = w116 & w6469;
assign w7575 = ~w7572 & ~w7573;
assign w7576 = (a[47] & w7574) | (a[47] & w25146) | (w7574 & w25146);
assign w7577 = ~w7574 & w25147;
assign w7578 = ~w7576 & ~w7577;
assign w7579 = (a[50] & w6995) | (a[50] & w25424) | (w6995 & w25424);
assign w7580 = w7316 & w25148;
assign w7581 = a[50] & ~w7580;
assign w7582 = b[1] & w7307;
assign w7583 = b[2] & w7314;
assign w7584 = w22 & w7312;
assign w7585 = w6995 & w7306;
assign w7586 = ~w7311 & w7585;
assign w7587 = b[0] & w7586;
assign w7588 = ~w7582 & ~w7583;
assign w7589 = ~w7584 & w7588;
assign w7590 = ~w7587 & w7589;
assign w7591 = ~w7581 & w7590;
assign w7592 = w7581 & ~w7590;
assign w7593 = ~w7591 & ~w7592;
assign w7594 = w7578 & w7593;
assign w7595 = ~w7578 & ~w7593;
assign w7596 = ~w7594 & ~w7595;
assign w7597 = (w7596 & w7325) | (w7596 & w25277) | (w7325 & w25277);
assign w7598 = ~w7325 & w25278;
assign w7599 = ~w7597 & ~w7598;
assign w7600 = b[6] & w5939;
assign w7601 = b[7] & w5670;
assign w7602 = b[8] & w5665;
assign w7603 = w270 & w5663;
assign w7604 = ~w7601 & ~w7602;
assign w7605 = ~w7600 & w7604;
assign w7606 = ~w7603 & w7605;
assign w7607 = a[44] & ~w7606;
assign w7608 = ~a[44] & w7606;
assign w7609 = ~w7607 & ~w7608;
assign w7610 = ~w7599 & ~w7609;
assign w7611 = w7599 & w7609;
assign w7612 = ~w7610 & ~w7611;
assign w7613 = (~w7339 & ~w7341) | (~w7339 & w25149) | (~w7341 & w25149);
assign w7614 = w7612 & w7613;
assign w7615 = ~w7612 & ~w7613;
assign w7616 = ~w7614 & ~w7615;
assign w7617 = b[9] & w5167;
assign w7618 = b[10] & w4918;
assign w7619 = b[11] & w4925;
assign w7620 = w469 & w4923;
assign w7621 = ~w7618 & ~w7619;
assign w7622 = ~w7617 & w7621;
assign w7623 = ~w7620 & w7622;
assign w7624 = a[41] & ~w7623;
assign w7625 = ~a[41] & w7623;
assign w7626 = ~w7624 & ~w7625;
assign w7627 = ~w7616 & ~w7626;
assign w7628 = w7616 & w7626;
assign w7629 = ~w7627 & ~w7628;
assign w7630 = w7569 & w7629;
assign w7631 = ~w7569 & ~w7629;
assign w7632 = ~w7630 & ~w7631;
assign w7633 = w7568 & ~w7632;
assign w7634 = ~w7568 & w7632;
assign w7635 = ~w7633 & ~w7634;
assign w7636 = ~w7558 & w7635;
assign w7637 = w7558 & ~w7635;
assign w7638 = ~w7636 & ~w7637;
assign w7639 = w7557 & w7638;
assign w7640 = ~w7557 & ~w7638;
assign w7641 = ~w7639 & ~w7640;
assign w7642 = ~w7547 & w7641;
assign w7643 = w7547 & ~w7641;
assign w7644 = ~w7642 & ~w7643;
assign w7645 = b[18] & w3177;
assign w7646 = b[20] & w2978;
assign w7647 = b[19] & w2973;
assign w7648 = w1347 & w2980;
assign w7649 = ~w7646 & ~w7647;
assign w7650 = ~w7645 & w7649;
assign w7651 = ~w7648 & w7650;
assign w7652 = a[32] & ~w7651;
assign w7653 = ~a[32] & w7651;
assign w7654 = ~w7652 & ~w7653;
assign w7655 = ~w7644 & ~w7654;
assign w7656 = w7644 & w7654;
assign w7657 = ~w7655 & ~w7656;
assign w7658 = (~w7375 & ~w7377) | (~w7375 & w25150) | (~w7377 & w25150);
assign w7659 = ~w7657 & ~w7658;
assign w7660 = w7657 & w7658;
assign w7661 = ~w7659 & ~w7660;
assign w7662 = b[22] & w2436;
assign w7663 = b[21] & ~w2622;
assign w7664 = b[23] & w2438;
assign w7665 = w1755 & w2432;
assign w7666 = ~w7662 & ~w7663;
assign w7667 = ~w7664 & w7666;
assign w7668 = ~w7665 & w7667;
assign w7669 = a[29] & ~w7668;
assign w7670 = ~a[29] & w7668;
assign w7671 = ~w7669 & ~w7670;
assign w7672 = ~w7661 & ~w7671;
assign w7673 = w7661 & w7671;
assign w7674 = ~w7672 & ~w7673;
assign w7675 = w7546 & w7674;
assign w7676 = ~w7546 & ~w7674;
assign w7677 = ~w7675 & ~w7676;
assign w7678 = ~w7545 & w7677;
assign w7679 = w7545 & ~w7677;
assign w7680 = ~w7678 & ~w7679;
assign w7681 = (~w7399 & ~w7250) | (~w7399 & w25151) | (~w7250 & w25151);
assign w7682 = w7680 & w7681;
assign w7683 = ~w7680 & ~w7681;
assign w7684 = ~w7682 & ~w7683;
assign w7685 = w7535 & w7684;
assign w7686 = ~w7535 & ~w7684;
assign w7687 = ~w7685 & ~w7686;
assign w7688 = ~w7525 & w7687;
assign w7689 = w7525 & ~w7687;
assign w7690 = ~w7688 & ~w7689;
assign w7691 = ~w7524 & ~w7690;
assign w7692 = w7524 & w7690;
assign w7693 = ~w7691 & ~w7692;
assign w7694 = (~w7411 & ~w7228) | (~w7411 & w25279) | (~w7228 & w25279);
assign w7695 = w7693 & w7694;
assign w7696 = ~w7693 & ~w7694;
assign w7697 = ~w7695 & ~w7696;
assign w7698 = b[33] & ~w934;
assign w7699 = b[34] & w838;
assign w7700 = b[35] & w834;
assign w7701 = w832 & w3918;
assign w7702 = ~w7698 & ~w7699;
assign w7703 = ~w7700 & w7702;
assign w7704 = ~w7701 & w7703;
assign w7705 = a[17] & ~w7704;
assign w7706 = ~a[17] & w7704;
assign w7707 = ~w7705 & ~w7706;
assign w7708 = w7697 & w7707;
assign w7709 = ~w7697 & ~w7707;
assign w7710 = ~w7708 & ~w7709;
assign w7711 = w7514 & w7710;
assign w7712 = ~w7514 & ~w7710;
assign w7713 = ~w7711 & ~w7712;
assign w7714 = ~w7513 & w7713;
assign w7715 = w7513 & ~w7713;
assign w7716 = ~w7714 & ~w7715;
assign w7717 = w7503 & ~w7716;
assign w7718 = ~w7503 & w7716;
assign w7719 = ~w7717 & ~w7718;
assign w7720 = b[39] & ~w419;
assign w7721 = b[40] & w358;
assign w7722 = b[41] & w360;
assign w7723 = w354 & w5302;
assign w7724 = ~w7720 & ~w7721;
assign w7725 = ~w7722 & w7724;
assign w7726 = ~w7723 & w7725;
assign w7727 = a[11] & ~w7726;
assign w7728 = ~a[11] & w7726;
assign w7729 = ~w7727 & ~w7728;
assign w7730 = w7719 & w7729;
assign w7731 = ~w7719 & ~w7729;
assign w7732 = ~w7730 & ~w7731;
assign w7733 = (~w7429 & ~w7432) | (~w7429 & w24830) | (~w7432 & w24830);
assign w7734 = w7732 & w7733;
assign w7735 = ~w7732 & ~w7733;
assign w7736 = ~w7734 & ~w7735;
assign w7737 = w7502 & ~w7736;
assign w7738 = ~w7502 & w7736;
assign w7739 = ~w7737 & ~w7738;
assign w7740 = (~w7447 & ~w7449) | (~w7447 & w24385) | (~w7449 & w24385);
assign w7741 = w7739 & w7740;
assign w7742 = ~w7739 & ~w7740;
assign w7743 = ~w7741 & ~w7742;
assign w7744 = w7492 & w7743;
assign w7745 = ~w7492 & ~w7743;
assign w7746 = ~w7744 & ~w7745;
assign w7747 = ~w7453 & ~w7458;
assign w7748 = w7746 & w7747;
assign w7749 = ~w7746 & ~w7747;
assign w7750 = ~w7748 & ~w7749;
assign w7751 = b[50] & w11;
assign w7752 = b[49] & w9;
assign w7753 = ~b[49] & ~b[50];
assign w7754 = b[49] & b[50];
assign w7755 = ~w7753 & ~w7754;
assign w7756 = (~w7462 & w7465) | (~w7462 & w25152) | (w7465 & w25152);
assign w7757 = w7755 & w7756;
assign w7758 = ~w7755 & ~w7756;
assign w7759 = ~w7757 & ~w7758;
assign w7760 = w5 & w7759;
assign w7761 = ~w7751 & ~w7752;
assign w7762 = ~w7760 & w7761;
assign w7763 = b[48] & w24;
assign w7764 = a[2] & ~w7763;
assign w7765 = w7762 & ~w7764;
assign w7766 = a[2] & ~w7762;
assign w7767 = ~w7765 & ~w7766;
assign w7768 = ~w7750 & w7767;
assign w7769 = w7750 & ~w7767;
assign w7770 = ~w7768 & ~w7769;
assign w7771 = ~w7478 & ~w7481;
assign w7772 = w7770 & ~w7771;
assign w7773 = ~w7770 & w7771;
assign w7774 = ~w7772 & ~w7773;
assign w7775 = ~w7768 & ~w7772;
assign w7776 = b[46] & w103;
assign w7777 = b[48] & w68;
assign w7778 = b[47] & w61;
assign w7779 = w66 & ~w7170;
assign w7780 = ~w7777 & ~w7778;
assign w7781 = ~w7776 & w7780;
assign w7782 = ~w7779 & w7781;
assign w7783 = a[5] & ~w7782;
assign w7784 = ~a[5] & w7782;
assign w7785 = ~w7783 & ~w7784;
assign w7786 = (~w7737 & ~w7740) | (~w7737 & w24831) | (~w7740 & w24831);
assign w7787 = b[40] & ~w419;
assign w7788 = b[42] & w360;
assign w7789 = b[41] & w358;
assign w7790 = w354 & w5548;
assign w7791 = ~w7787 & ~w7788;
assign w7792 = ~w7789 & w7791;
assign w7793 = ~w7790 & w7792;
assign w7794 = a[11] & ~w7793;
assign w7795 = ~a[11] & w7793;
assign w7796 = ~w7794 & ~w7795;
assign w7797 = ~w7715 & ~w7718;
assign w7798 = b[38] & w573;
assign w7799 = b[37] & ~w649;
assign w7800 = b[39] & w575;
assign w7801 = w569 & ~w4812;
assign w7802 = ~w7798 & ~w7799;
assign w7803 = ~w7800 & w7802;
assign w7804 = ~w7801 & w7803;
assign w7805 = a[14] & ~w7804;
assign w7806 = ~a[14] & w7804;
assign w7807 = ~w7805 & ~w7806;
assign w7808 = b[35] & w838;
assign w7809 = b[36] & w834;
assign w7810 = b[34] & ~w934;
assign w7811 = w832 & w4129;
assign w7812 = ~w7808 & ~w7809;
assign w7813 = ~w7810 & w7812;
assign w7814 = ~w7811 & w7813;
assign w7815 = a[17] & ~w7814;
assign w7816 = ~a[17] & w7814;
assign w7817 = ~w7815 & ~w7816;
assign w7818 = (~w7692 & ~w7694) | (~w7692 & w25425) | (~w7694 & w25425);
assign w7819 = (~w7685 & w7525) | (~w7685 & w25153) | (w7525 & w25153);
assign w7820 = b[28] & ~w1676;
assign w7821 = b[29] & w1517;
assign w7822 = b[30] & w1519;
assign w7823 = w1513 & ~w2908;
assign w7824 = ~w7820 & ~w7821;
assign w7825 = ~w7822 & w7824;
assign w7826 = ~w7823 & w7825;
assign w7827 = a[23] & ~w7826;
assign w7828 = ~a[23] & w7826;
assign w7829 = ~w7827 & ~w7828;
assign w7830 = ~w7679 & ~w7682;
assign w7831 = b[24] & w2438;
assign w7832 = b[23] & w2436;
assign w7833 = b[22] & ~w2622;
assign w7834 = w1895 & w2432;
assign w7835 = ~w7831 & ~w7832;
assign w7836 = ~w7833 & w7835;
assign w7837 = ~w7834 & w7836;
assign w7838 = a[29] & ~w7837;
assign w7839 = ~a[29] & w7837;
assign w7840 = ~w7838 & ~w7839;
assign w7841 = (~w7656 & ~w7658) | (~w7656 & w25426) | (~w7658 & w25426);
assign w7842 = (~w7639 & w7547) | (~w7639 & w25154) | (w7547 & w25154);
assign w7843 = b[16] & w3785;
assign w7844 = b[17] & w3578;
assign w7845 = b[18] & w3580;
assign w7846 = ~w1108 & w3573;
assign w7847 = ~w7844 & ~w7845;
assign w7848 = ~w7843 & w7847;
assign w7849 = ~w7846 & w7848;
assign w7850 = a[35] & ~w7849;
assign w7851 = ~a[35] & w7849;
assign w7852 = ~w7850 & ~w7851;
assign w7853 = ~w7633 & ~w7636;
assign w7854 = b[13] & w4453;
assign w7855 = b[14] & w4241;
assign w7856 = b[15] & w4243;
assign w7857 = ~w799 & w4236;
assign w7858 = ~w7855 & ~w7856;
assign w7859 = ~w7854 & w7858;
assign w7860 = ~w7857 & w7859;
assign w7861 = a[38] & ~w7860;
assign w7862 = ~a[38] & w7860;
assign w7863 = ~w7861 & ~w7862;
assign w7864 = (~w7611 & ~w7613) | (~w7611 & w25280) | (~w7613 & w25280);
assign w7865 = a[50] & ~a[51];
assign w7866 = ~a[50] & a[51];
assign w7867 = ~w7865 & ~w7866;
assign w7868 = b[0] & ~w7867;
assign w7869 = w7580 & w7590;
assign w7870 = w46 & w7312;
assign w7871 = b[2] & w7307;
assign w7872 = b[3] & w7314;
assign w7873 = w7585 & w25155;
assign w7874 = ~w7871 & ~w7872;
assign w7875 = ~w7870 & w7874;
assign w7876 = (a[50] & ~w7875) | (a[50] & w24982) | (~w7875 & w24982);
assign w7877 = w7875 & w24983;
assign w7878 = ~w7876 & ~w7877;
assign w7879 = w7869 & w7878;
assign w7880 = ~w7869 & ~w7878;
assign w7881 = ~w7879 & ~w7880;
assign w7882 = w7868 & w7881;
assign w7883 = ~w7868 & ~w7881;
assign w7884 = ~w7882 & ~w7883;
assign w7885 = b[4] & w6732;
assign w7886 = b[5] & w6474;
assign w7887 = b[6] & w6476;
assign w7888 = w157 & w6469;
assign w7889 = ~w7886 & ~w7887;
assign w7890 = ~w7885 & w7889;
assign w7891 = ~w7888 & w7890;
assign w7892 = a[47] & ~w7891;
assign w7893 = ~a[47] & w7891;
assign w7894 = ~w7892 & ~w7893;
assign w7895 = w7884 & w7894;
assign w7896 = ~w7884 & ~w7894;
assign w7897 = ~w7895 & ~w7896;
assign w7898 = (~w7594 & w7570) | (~w7594 & w24984) | (w7570 & w24984);
assign w7899 = ~w7897 & w7898;
assign w7900 = w7897 & ~w7898;
assign w7901 = ~w7899 & ~w7900;
assign w7902 = b[7] & w5939;
assign w7903 = b[9] & w5665;
assign w7904 = b[8] & w5670;
assign w7905 = w322 & w5663;
assign w7906 = ~w7903 & ~w7904;
assign w7907 = ~w7902 & w7906;
assign w7908 = ~w7905 & w7907;
assign w7909 = a[44] & ~w7908;
assign w7910 = ~a[44] & w7908;
assign w7911 = ~w7909 & ~w7910;
assign w7912 = ~w7901 & ~w7911;
assign w7913 = w7901 & w7911;
assign w7914 = ~w7912 & ~w7913;
assign w7915 = ~w7614 & w24985;
assign w7916 = ~w7864 & ~w7914;
assign w7917 = b[10] & w5167;
assign w7918 = b[11] & w4918;
assign w7919 = b[12] & w4925;
assign w7920 = w536 & w4923;
assign w7921 = ~w7918 & ~w7919;
assign w7922 = ~w7917 & w7921;
assign w7923 = ~w7920 & w7922;
assign w7924 = a[41] & ~w7923;
assign w7925 = ~a[41] & w7923;
assign w7926 = ~w7924 & ~w7925;
assign w7927 = ~w7915 & w25281;
assign w7928 = (w7926 & w7915) | (w7926 & w25282) | (w7915 & w25282);
assign w7929 = ~w7927 & ~w7928;
assign w7930 = (~w7627 & ~w7569) | (~w7627 & w24986) | (~w7569 & w24986);
assign w7931 = w7929 & w7930;
assign w7932 = ~w7929 & ~w7930;
assign w7933 = ~w7931 & ~w7932;
assign w7934 = w7863 & w7933;
assign w7935 = ~w7863 & ~w7933;
assign w7936 = ~w7934 & ~w7935;
assign w7937 = w7853 & w7936;
assign w7938 = ~w7853 & ~w7936;
assign w7939 = ~w7937 & ~w7938;
assign w7940 = w7852 & ~w7939;
assign w7941 = ~w7852 & w7939;
assign w7942 = ~w7940 & ~w7941;
assign w7943 = ~w7842 & w7942;
assign w7944 = w7842 & ~w7942;
assign w7945 = ~w7943 & ~w7944;
assign w7946 = b[19] & w3177;
assign w7947 = b[21] & w2978;
assign w7948 = b[20] & w2973;
assign w7949 = w1467 & w2980;
assign w7950 = ~w7947 & ~w7948;
assign w7951 = ~w7946 & w7950;
assign w7952 = ~w7949 & w7951;
assign w7953 = a[32] & ~w7952;
assign w7954 = ~a[32] & w7952;
assign w7955 = ~w7953 & ~w7954;
assign w7956 = w7945 & w7955;
assign w7957 = ~w7945 & ~w7955;
assign w7958 = ~w7956 & ~w7957;
assign w7959 = ~w7841 & w7958;
assign w7960 = w7841 & ~w7958;
assign w7961 = ~w7959 & ~w7960;
assign w7962 = ~w7840 & ~w7961;
assign w7963 = w7840 & w7961;
assign w7964 = ~w7962 & ~w7963;
assign w7965 = (~w7672 & ~w7546) | (~w7672 & w25156) | (~w7546 & w25156);
assign w7966 = w7964 & w7965;
assign w7967 = ~w7964 & ~w7965;
assign w7968 = ~w7966 & ~w7967;
assign w7969 = b[26] & w1955;
assign w7970 = b[25] & ~w2114;
assign w7971 = b[27] & w1957;
assign w7972 = w1951 & w2378;
assign w7973 = ~w7969 & ~w7970;
assign w7974 = ~w7971 & w7973;
assign w7975 = ~w7972 & w7974;
assign w7976 = a[26] & ~w7975;
assign w7977 = ~a[26] & w7975;
assign w7978 = ~w7976 & ~w7977;
assign w7979 = w7968 & w7978;
assign w7980 = ~w7968 & ~w7978;
assign w7981 = ~w7979 & ~w7980;
assign w7982 = w7830 & w7981;
assign w7983 = ~w7830 & ~w7981;
assign w7984 = ~w7982 & ~w7983;
assign w7985 = w7829 & ~w7984;
assign w7986 = ~w7829 & w7984;
assign w7987 = ~w7985 & ~w7986;
assign w7988 = ~w7819 & w7987;
assign w7989 = w7819 & ~w7987;
assign w7990 = ~w7988 & ~w7989;
assign w7991 = b[31] & ~w1272;
assign w7992 = b[33] & w1156;
assign w7993 = b[32] & w1154;
assign w7994 = w1150 & w3499;
assign w7995 = ~w7991 & ~w7992;
assign w7996 = ~w7993 & w7995;
assign w7997 = ~w7994 & w7996;
assign w7998 = a[20] & ~w7997;
assign w7999 = ~a[20] & w7997;
assign w8000 = ~w7998 & ~w7999;
assign w8001 = w7990 & w8000;
assign w8002 = ~w7990 & ~w8000;
assign w8003 = ~w8001 & ~w8002;
assign w8004 = w7818 & ~w8003;
assign w8005 = ~w7818 & w8003;
assign w8006 = ~w8004 & ~w8005;
assign w8007 = w7817 & w8006;
assign w8008 = ~w7817 & ~w8006;
assign w8009 = ~w8007 & ~w8008;
assign w8010 = (~w7709 & ~w7514) | (~w7709 & w25283) | (~w7514 & w25283);
assign w8011 = w8009 & w8010;
assign w8012 = ~w8009 & ~w8010;
assign w8013 = ~w8011 & ~w8012;
assign w8014 = w7807 & w8013;
assign w8015 = ~w7807 & ~w8013;
assign w8016 = ~w8014 & ~w8015;
assign w8017 = ~w7797 & w8016;
assign w8018 = w7797 & ~w8016;
assign w8019 = ~w8017 & ~w8018;
assign w8020 = ~w7796 & ~w8019;
assign w8021 = w7796 & w8019;
assign w8022 = ~w8020 & ~w8021;
assign w8023 = (~w7731 & ~w7733) | (~w7731 & w24674) | (~w7733 & w24674);
assign w8024 = w8022 & w8023;
assign w8025 = ~w8022 & ~w8023;
assign w8026 = ~w8024 & ~w8025;
assign w8027 = b[44] & w183;
assign w8028 = b[43] & ~w237;
assign w8029 = b[45] & w185;
assign w8030 = w179 & w6334;
assign w8031 = ~w8027 & ~w8028;
assign w8032 = ~w8029 & w8031;
assign w8033 = ~w8030 & w8032;
assign w8034 = a[8] & ~w8033;
assign w8035 = ~a[8] & w8033;
assign w8036 = ~w8034 & ~w8035;
assign w8037 = w8026 & w8036;
assign w8038 = ~w8026 & ~w8036;
assign w8039 = ~w8037 & ~w8038;
assign w8040 = w7786 & w8039;
assign w8041 = ~w7786 & ~w8039;
assign w8042 = ~w8040 & ~w8041;
assign w8043 = ~w7785 & w8042;
assign w8044 = w7785 & ~w8042;
assign w8045 = ~w8043 & ~w8044;
assign w8046 = (~w7745 & ~w7747) | (~w7745 & w24386) | (~w7747 & w24386);
assign w8047 = w8045 & w8046;
assign w8048 = ~w8045 & ~w8046;
assign w8049 = ~w8047 & ~w8048;
assign w8050 = b[51] & w11;
assign w8051 = b[50] & w9;
assign w8052 = (~w7754 & ~w7756) | (~w7754 & w24987) | (~w7756 & w24987);
assign w8053 = ~b[50] & ~b[51];
assign w8054 = b[50] & b[51];
assign w8055 = ~w8053 & ~w8054;
assign w8056 = ~w8052 & ~w8055;
assign w8057 = w8052 & w8055;
assign w8058 = ~w8056 & ~w8057;
assign w8059 = w5 & ~w8058;
assign w8060 = ~w8050 & ~w8051;
assign w8061 = ~w8059 & w8060;
assign w8062 = b[49] & w24;
assign w8063 = a[2] & ~w8062;
assign w8064 = w8061 & ~w8063;
assign w8065 = a[2] & ~w8061;
assign w8066 = ~w8064 & ~w8065;
assign w8067 = w8049 & w8066;
assign w8068 = ~w8049 & ~w8066;
assign w8069 = ~w8067 & ~w8068;
assign w8070 = ~w7775 & w8069;
assign w8071 = w7775 & ~w8069;
assign w8072 = ~w8070 & ~w8071;
assign w8073 = (~w8044 & ~w8046) | (~w8044 & w24832) | (~w8046 & w24832);
assign w8074 = b[44] & ~w237;
assign w8075 = b[45] & w183;
assign w8076 = b[46] & w185;
assign w8077 = w179 & ~w6613;
assign w8078 = ~w8074 & ~w8075;
assign w8079 = ~w8076 & w8078;
assign w8080 = ~w8077 & w8079;
assign w8081 = a[8] & ~w8080;
assign w8082 = ~a[8] & w8080;
assign w8083 = ~w8081 & ~w8082;
assign w8084 = (~w8014 & w7797) | (~w8014 & w25284) | (w7797 & w25284);
assign w8085 = b[38] & ~w649;
assign w8086 = b[39] & w573;
assign w8087 = b[40] & w575;
assign w8088 = w569 & ~w5058;
assign w8089 = ~w8085 & ~w8086;
assign w8090 = ~w8087 & w8089;
assign w8091 = ~w8088 & w8090;
assign w8092 = a[14] & ~w8091;
assign w8093 = ~a[14] & w8091;
assign w8094 = ~w8092 & ~w8093;
assign w8095 = (~w8007 & ~w8010) | (~w8007 & w25427) | (~w8010 & w25427);
assign w8096 = b[34] & w1156;
assign w8097 = b[33] & w1154;
assign w8098 = b[32] & ~w1272;
assign w8099 = w1150 & ~w3710;
assign w8100 = ~w8096 & ~w8097;
assign w8101 = ~w8098 & w8100;
assign w8102 = ~w8099 & w8101;
assign w8103 = a[20] & ~w8102;
assign w8104 = ~a[20] & w8102;
assign w8105 = ~w8103 & ~w8104;
assign w8106 = (~w7985 & w7819) | (~w7985 & w24988) | (w7819 & w24988);
assign w8107 = b[31] & w1519;
assign w8108 = b[29] & ~w1676;
assign w8109 = b[30] & w1517;
assign w8110 = w1513 & ~w3112;
assign w8111 = ~w8107 & ~w8108;
assign w8112 = ~w8109 & w8111;
assign w8113 = ~w8110 & w8112;
assign w8114 = a[23] & ~w8113;
assign w8115 = ~a[23] & w8113;
assign w8116 = ~w8114 & ~w8115;
assign w8117 = b[26] & ~w2114;
assign w8118 = b[27] & w1955;
assign w8119 = b[28] & w1957;
assign w8120 = w1951 & w2559;
assign w8121 = ~w8117 & ~w8118;
assign w8122 = ~w8119 & w8121;
assign w8123 = ~w8120 & w8122;
assign w8124 = a[26] & ~w8123;
assign w8125 = ~a[26] & w8123;
assign w8126 = ~w8124 & ~w8125;
assign w8127 = (~w7963 & ~w7965) | (~w7963 & w25428) | (~w7965 & w25428);
assign w8128 = (~w7956 & w7841) | (~w7956 & w24989) | (w7841 & w24989);
assign w8129 = b[20] & w3177;
assign w8130 = b[21] & w2973;
assign w8131 = b[22] & w2978;
assign w8132 = w1615 & w2980;
assign w8133 = ~w8130 & ~w8131;
assign w8134 = ~w8129 & w8133;
assign w8135 = ~w8132 & w8134;
assign w8136 = a[32] & ~w8135;
assign w8137 = ~a[32] & w8135;
assign w8138 = ~w8136 & ~w8137;
assign w8139 = (~w7940 & w7842) | (~w7940 & w24990) | (w7842 & w24990);
assign w8140 = b[17] & w3785;
assign w8141 = b[19] & w3580;
assign w8142 = b[18] & w3578;
assign w8143 = ~w1231 & w3573;
assign w8144 = ~w8141 & ~w8142;
assign w8145 = ~w8140 & w8144;
assign w8146 = ~w8143 & w8145;
assign w8147 = a[35] & ~w8146;
assign w8148 = ~a[35] & w8146;
assign w8149 = ~w8147 & ~w8148;
assign w8150 = b[14] & w4453;
assign w8151 = b[15] & w4241;
assign w8152 = b[16] & w4243;
assign w8153 = w905 & w4236;
assign w8154 = ~w8151 & ~w8152;
assign w8155 = ~w8150 & w8154;
assign w8156 = ~w8153 & w8155;
assign w8157 = a[38] & ~w8156;
assign w8158 = ~a[38] & w8156;
assign w8159 = ~w8157 & ~w8158;
assign w8160 = (~w7928 & ~w7930) | (~w7928 & w25285) | (~w7930 & w25285);
assign w8161 = b[11] & w5167;
assign w8162 = b[13] & w4925;
assign w8163 = b[12] & w4918;
assign w8164 = w628 & w4923;
assign w8165 = ~w8162 & ~w8163;
assign w8166 = ~w8161 & w8165;
assign w8167 = ~w8164 & w8166;
assign w8168 = a[41] & ~w8167;
assign w8169 = ~a[41] & w8167;
assign w8170 = ~w8168 & ~w8169;
assign w8171 = b[8] & w5939;
assign w8172 = b[9] & w5670;
assign w8173 = b[10] & w5665;
assign w8174 = w397 & w5663;
assign w8175 = ~w8172 & ~w8173;
assign w8176 = ~w8171 & w8175;
assign w8177 = ~w8174 & w8176;
assign w8178 = a[44] & ~w8177;
assign w8179 = ~a[44] & w8177;
assign w8180 = ~w8178 & ~w8179;
assign w8181 = w7585 & w25157;
assign w8182 = b[3] & w7307;
assign w8183 = b[4] & w7314;
assign w8184 = w84 & w7312;
assign w8185 = ~w8182 & ~w8183;
assign w8186 = ~w8181 & w8185;
assign w8187 = ~w8184 & w8186;
assign w8188 = a[50] & ~w8187;
assign w8189 = ~a[50] & w8187;
assign w8190 = ~w8188 & ~w8189;
assign w8191 = a[53] & w7868;
assign w8192 = a[52] & ~a[53];
assign w8193 = ~a[52] & a[53];
assign w8194 = ~w8192 & ~w8193;
assign w8195 = ~w7867 & ~w8194;
assign w8196 = ~w8 & w8195;
assign w8197 = a[51] & ~a[52];
assign w8198 = ~a[51] & a[52];
assign w8199 = ~w8197 & ~w8198;
assign w8200 = w7867 & ~w8199;
assign w8201 = b[0] & w8200;
assign w8202 = ~w7867 & w8194;
assign w8203 = b[1] & w8202;
assign w8204 = ~w8196 & ~w8201;
assign w8205 = ~w8203 & w8204;
assign w8206 = ~w8191 & w8205;
assign w8207 = w8191 & ~w8205;
assign w8208 = ~w8206 & ~w8207;
assign w8209 = ~w8190 & ~w8208;
assign w8210 = w8190 & w8208;
assign w8211 = ~w8209 & ~w8210;
assign w8212 = (~w7879 & ~w7881) | (~w7879 & w24991) | (~w7881 & w24991);
assign w8213 = w8211 & ~w8212;
assign w8214 = ~w8211 & w8212;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = b[5] & w6732;
assign w8217 = b[6] & w6474;
assign w8218 = b[7] & w6476;
assign w8219 = w216 & w6469;
assign w8220 = ~w8217 & ~w8218;
assign w8221 = ~w8216 & w8220;
assign w8222 = ~w8219 & w8221;
assign w8223 = a[47] & ~w8222;
assign w8224 = ~a[47] & w8222;
assign w8225 = ~w8223 & ~w8224;
assign w8226 = w8215 & w8225;
assign w8227 = ~w8215 & ~w8225;
assign w8228 = ~w8226 & ~w8227;
assign w8229 = ~w7895 & ~w7900;
assign w8230 = w8228 & w8229;
assign w8231 = ~w8228 & ~w8229;
assign w8232 = ~w8230 & ~w8231;
assign w8233 = w8180 & ~w8232;
assign w8234 = ~w8180 & w8232;
assign w8235 = ~w8233 & ~w8234;
assign w8236 = (~w7912 & ~w24985) | (~w7912 & w25158) | (~w24985 & w25158);
assign w8237 = w8235 & w8236;
assign w8238 = ~w8235 & ~w8236;
assign w8239 = ~w8237 & ~w8238;
assign w8240 = ~w8170 & ~w8239;
assign w8241 = w8170 & w8239;
assign w8242 = ~w8240 & ~w8241;
assign w8243 = ~w8160 & ~w8242;
assign w8244 = w8160 & w8242;
assign w8245 = ~w8243 & ~w8244;
assign w8246 = w8159 & ~w8245;
assign w8247 = ~w8159 & w8245;
assign w8248 = ~w8246 & ~w8247;
assign w8249 = (~w7935 & ~w7853) | (~w7935 & w24992) | (~w7853 & w24992);
assign w8250 = ~w8248 & ~w8249;
assign w8251 = w8248 & w8249;
assign w8252 = ~w8250 & ~w8251;
assign w8253 = ~w8149 & ~w8252;
assign w8254 = w8149 & w8252;
assign w8255 = ~w8253 & ~w8254;
assign w8256 = ~w8139 & ~w8255;
assign w8257 = w8139 & w8255;
assign w8258 = ~w8256 & ~w8257;
assign w8259 = w8138 & ~w8258;
assign w8260 = ~w8138 & w8258;
assign w8261 = ~w8259 & ~w8260;
assign w8262 = w8128 & ~w8261;
assign w8263 = ~w8128 & w8261;
assign w8264 = ~w8262 & ~w8263;
assign w8265 = b[25] & w2438;
assign w8266 = b[23] & ~w2622;
assign w8267 = b[24] & w2436;
assign w8268 = w2061 & w2432;
assign w8269 = ~w8265 & ~w8266;
assign w8270 = ~w8267 & w8269;
assign w8271 = ~w8268 & w8270;
assign w8272 = a[29] & ~w8271;
assign w8273 = ~a[29] & w8271;
assign w8274 = ~w8272 & ~w8273;
assign w8275 = w8264 & w8274;
assign w8276 = ~w8264 & ~w8274;
assign w8277 = ~w8275 & ~w8276;
assign w8278 = ~w8127 & ~w8277;
assign w8279 = w8127 & w8277;
assign w8280 = ~w8278 & ~w8279;
assign w8281 = ~w8126 & w8280;
assign w8282 = w8126 & ~w8280;
assign w8283 = ~w8281 & ~w8282;
assign w8284 = (~w7980 & ~w7830) | (~w7980 & w24993) | (~w7830 & w24993);
assign w8285 = w8283 & w8284;
assign w8286 = ~w8283 & ~w8284;
assign w8287 = ~w8285 & ~w8286;
assign w8288 = w8116 & w8287;
assign w8289 = ~w8116 & ~w8287;
assign w8290 = ~w8288 & ~w8289;
assign w8291 = ~w8106 & w8290;
assign w8292 = w8106 & ~w8290;
assign w8293 = ~w8291 & ~w8292;
assign w8294 = w8105 & w8293;
assign w8295 = ~w8105 & ~w8293;
assign w8296 = ~w8294 & ~w8295;
assign w8297 = (~w8001 & w7818) | (~w8001 & w25159) | (w7818 & w25159);
assign w8298 = ~w8296 & w8297;
assign w8299 = w8296 & ~w8297;
assign w8300 = ~w8298 & ~w8299;
assign w8301 = b[35] & ~w934;
assign w8302 = b[36] & w838;
assign w8303 = b[37] & w834;
assign w8304 = w832 & ~w4357;
assign w8305 = ~w8301 & ~w8302;
assign w8306 = ~w8303 & w8305;
assign w8307 = ~w8304 & w8306;
assign w8308 = a[17] & ~w8307;
assign w8309 = ~a[17] & w8307;
assign w8310 = ~w8308 & ~w8309;
assign w8311 = w8300 & w8310;
assign w8312 = ~w8300 & ~w8310;
assign w8313 = ~w8311 & ~w8312;
assign w8314 = w8095 & w8313;
assign w8315 = ~w8095 & ~w8313;
assign w8316 = ~w8314 & ~w8315;
assign w8317 = ~w8094 & w8316;
assign w8318 = w8094 & ~w8316;
assign w8319 = ~w8317 & ~w8318;
assign w8320 = w8084 & ~w8319;
assign w8321 = ~w8084 & w8319;
assign w8322 = ~w8320 & ~w8321;
assign w8323 = b[41] & ~w419;
assign w8324 = b[43] & w360;
assign w8325 = b[42] & w358;
assign w8326 = w354 & w5811;
assign w8327 = ~w8323 & ~w8324;
assign w8328 = ~w8325 & w8327;
assign w8329 = ~w8326 & w8328;
assign w8330 = a[11] & ~w8329;
assign w8331 = ~a[11] & w8329;
assign w8332 = ~w8330 & ~w8331;
assign w8333 = w8322 & w8332;
assign w8334 = ~w8322 & ~w8332;
assign w8335 = ~w8333 & ~w8334;
assign w8336 = ~w8021 & ~w8024;
assign w8337 = w8335 & w8336;
assign w8338 = ~w8335 & ~w8336;
assign w8339 = ~w8337 & ~w8338;
assign w8340 = w8083 & ~w8339;
assign w8341 = ~w8083 & w8339;
assign w8342 = ~w8340 & ~w8341;
assign w8343 = (~w8038 & ~w7786) | (~w8038 & w24675) | (~w7786 & w24675);
assign w8344 = ~w8342 & ~w8343;
assign w8345 = w8342 & w8343;
assign w8346 = ~w8344 & ~w8345;
assign w8347 = b[47] & w103;
assign w8348 = b[48] & w61;
assign w8349 = b[49] & w68;
assign w8350 = w66 & ~w7468;
assign w8351 = ~w8348 & ~w8349;
assign w8352 = ~w8347 & w8351;
assign w8353 = ~w8350 & w8352;
assign w8354 = a[5] & ~w8353;
assign w8355 = ~a[5] & w8353;
assign w8356 = ~w8354 & ~w8355;
assign w8357 = w8346 & w8356;
assign w8358 = ~w8346 & ~w8356;
assign w8359 = ~w8357 & ~w8358;
assign w8360 = ~w8073 & ~w8359;
assign w8361 = w8073 & w8359;
assign w8362 = ~w8360 & ~w8361;
assign w8363 = b[52] & w11;
assign w8364 = b[51] & w9;
assign w8365 = ~b[51] & ~b[52];
assign w8366 = b[51] & b[52];
assign w8367 = ~w8365 & ~w8366;
assign w8368 = ~w8053 & ~w8057;
assign w8369 = ~w8367 & w8368;
assign w8370 = w8367 & ~w8368;
assign w8371 = ~w8369 & ~w8370;
assign w8372 = w5 & ~w8371;
assign w8373 = ~w8363 & ~w8364;
assign w8374 = ~w8372 & w8373;
assign w8375 = b[50] & w24;
assign w8376 = a[2] & ~w8375;
assign w8377 = w8374 & ~w8376;
assign w8378 = a[2] & ~w8374;
assign w8379 = ~w8377 & ~w8378;
assign w8380 = ~w8362 & w8379;
assign w8381 = w8362 & ~w8379;
assign w8382 = ~w8380 & ~w8381;
assign w8383 = (~w8067 & w7775) | (~w8067 & w24387) | (w7775 & w24387);
assign w8384 = w8382 & ~w8383;
assign w8385 = ~w8382 & w8383;
assign w8386 = ~w8384 & ~w8385;
assign w8387 = (~w8380 & w8383) | (~w8380 & w24833) | (w8383 & w24833);
assign w8388 = b[48] & w103;
assign w8389 = b[49] & w61;
assign w8390 = b[50] & w68;
assign w8391 = w66 & w7759;
assign w8392 = ~w8389 & ~w8390;
assign w8393 = ~w8388 & w8392;
assign w8394 = ~w8391 & w8393;
assign w8395 = a[5] & ~w8394;
assign w8396 = ~a[5] & w8394;
assign w8397 = ~w8395 & ~w8396;
assign w8398 = ~w8340 & ~w8345;
assign w8399 = b[46] & w183;
assign w8400 = b[47] & w185;
assign w8401 = b[45] & ~w237;
assign w8402 = w179 & w6889;
assign w8403 = ~w8399 & ~w8400;
assign w8404 = ~w8401 & w8403;
assign w8405 = ~w8402 & w8404;
assign w8406 = a[8] & ~w8405;
assign w8407 = ~a[8] & w8405;
assign w8408 = ~w8406 & ~w8407;
assign w8409 = b[43] & w358;
assign w8410 = b[42] & ~w419;
assign w8411 = b[44] & w360;
assign w8412 = w354 & w6069;
assign w8413 = ~w8409 & ~w8410;
assign w8414 = ~w8411 & w8413;
assign w8415 = ~w8412 & w8414;
assign w8416 = a[11] & ~w8415;
assign w8417 = ~a[11] & w8415;
assign w8418 = ~w8416 & ~w8417;
assign w8419 = (~w8318 & w8084) | (~w8318 & w25429) | (w8084 & w25429);
assign w8420 = b[40] & w573;
assign w8421 = b[39] & ~w649;
assign w8422 = b[41] & w575;
assign w8423 = w569 & w5302;
assign w8424 = ~w8420 & ~w8421;
assign w8425 = ~w8422 & w8424;
assign w8426 = ~w8423 & w8425;
assign w8427 = a[14] & ~w8426;
assign w8428 = ~a[14] & w8426;
assign w8429 = ~w8427 & ~w8428;
assign w8430 = b[38] & w834;
assign w8431 = b[37] & w838;
assign w8432 = b[36] & ~w934;
assign w8433 = w832 & w4582;
assign w8434 = ~w8430 & ~w8431;
assign w8435 = ~w8432 & w8434;
assign w8436 = ~w8433 & w8435;
assign w8437 = a[17] & ~w8436;
assign w8438 = ~a[17] & w8436;
assign w8439 = ~w8437 & ~w8438;
assign w8440 = (~w8294 & w8297) | (~w8294 & w24994) | (w8297 & w24994);
assign w8441 = (~w8288 & w8106) | (~w8288 & w24388) | (w8106 & w24388);
assign w8442 = b[31] & w1517;
assign w8443 = b[30] & ~w1676;
assign w8444 = b[32] & w1519;
assign w8445 = w1513 & w3304;
assign w8446 = ~w8442 & ~w8443;
assign w8447 = ~w8444 & w8446;
assign w8448 = ~w8445 & w8447;
assign w8449 = a[23] & ~w8448;
assign w8450 = ~a[23] & w8448;
assign w8451 = ~w8449 & ~w8450;
assign w8452 = (~w8282 & ~w8284) | (~w8282 & w24834) | (~w8284 & w24834);
assign w8453 = b[25] & w2436;
assign w8454 = b[26] & w2438;
assign w8455 = b[24] & ~w2622;
assign w8456 = w2219 & w2432;
assign w8457 = ~w8453 & ~w8454;
assign w8458 = ~w8455 & w8457;
assign w8459 = ~w8456 & w8458;
assign w8460 = a[29] & ~w8459;
assign w8461 = ~a[29] & w8459;
assign w8462 = ~w8460 & ~w8461;
assign w8463 = (~w8259 & w8128) | (~w8259 & w24835) | (w8128 & w24835);
assign w8464 = (~w8253 & ~w8139) | (~w8253 & w24836) | (~w8139 & w24836);
assign w8465 = b[18] & w3785;
assign w8466 = b[20] & w3580;
assign w8467 = b[19] & w3578;
assign w8468 = w1347 & w3573;
assign w8469 = ~w8466 & ~w8467;
assign w8470 = ~w8465 & w8469;
assign w8471 = ~w8468 & w8470;
assign w8472 = a[35] & ~w8471;
assign w8473 = ~a[35] & w8471;
assign w8474 = ~w8472 & ~w8473;
assign w8475 = (~w8246 & ~w8249) | (~w8246 & w25286) | (~w8249 & w25286);
assign w8476 = b[12] & w5167;
assign w8477 = b[13] & w4918;
assign w8478 = b[14] & w4925;
assign w8479 = w714 & w4923;
assign w8480 = ~w8477 & ~w8478;
assign w8481 = ~w8476 & w8480;
assign w8482 = ~w8479 & w8481;
assign w8483 = a[41] & ~w8482;
assign w8484 = ~a[41] & w8482;
assign w8485 = ~w8483 & ~w8484;
assign w8486 = (~w8233 & ~w8236) | (~w8233 & w24837) | (~w8236 & w24837);
assign w8487 = b[9] & w5939;
assign w8488 = b[10] & w5670;
assign w8489 = b[11] & w5665;
assign w8490 = w469 & w5663;
assign w8491 = ~w8488 & ~w8489;
assign w8492 = ~w8487 & w8491;
assign w8493 = ~w8490 & w8492;
assign w8494 = a[44] & ~w8493;
assign w8495 = ~a[44] & w8493;
assign w8496 = ~w8494 & ~w8495;
assign w8497 = ~w8210 & ~w8213;
assign w8498 = b[3] & w7586;
assign w8499 = b[5] & w7314;
assign w8500 = b[4] & w7307;
assign w8501 = w116 & w7312;
assign w8502 = ~w8499 & ~w8500;
assign w8503 = ~w8498 & w8502;
assign w8504 = ~w8501 & w8503;
assign w8505 = a[50] & ~w8504;
assign w8506 = ~a[50] & w8504;
assign w8507 = ~w8505 & ~w8506;
assign w8508 = a[53] & ~w7868;
assign w8509 = w8204 & w25160;
assign w8510 = a[53] & ~w8509;
assign w8511 = b[1] & w8200;
assign w8512 = b[2] & w8202;
assign w8513 = w22 & w8195;
assign w8514 = w7867 & ~w8194;
assign w8515 = w8199 & w8514;
assign w8516 = b[0] & w8515;
assign w8517 = ~w8511 & ~w8512;
assign w8518 = ~w8513 & w8517;
assign w8519 = ~w8516 & w8518;
assign w8520 = ~w8510 & w8519;
assign w8521 = w8510 & ~w8519;
assign w8522 = ~w8520 & ~w8521;
assign w8523 = w8507 & w8522;
assign w8524 = ~w8507 & ~w8522;
assign w8525 = ~w8523 & ~w8524;
assign w8526 = w8497 & w8525;
assign w8527 = ~w8497 & ~w8525;
assign w8528 = ~w8526 & ~w8527;
assign w8529 = b[6] & w6732;
assign w8530 = b[7] & w6474;
assign w8531 = b[8] & w6476;
assign w8532 = w270 & w6469;
assign w8533 = ~w8530 & ~w8531;
assign w8534 = ~w8529 & w8533;
assign w8535 = ~w8532 & w8534;
assign w8536 = a[47] & ~w8535;
assign w8537 = ~a[47] & w8535;
assign w8538 = ~w8536 & ~w8537;
assign w8539 = w8528 & ~w8538;
assign w8540 = ~w8528 & w8538;
assign w8541 = ~w8539 & ~w8540;
assign w8542 = (~w8227 & ~w8229) | (~w8227 & w24838) | (~w8229 & w24838);
assign w8543 = w8541 & w8542;
assign w8544 = ~w8541 & ~w8542;
assign w8545 = ~w8543 & ~w8544;
assign w8546 = ~w8496 & ~w8545;
assign w8547 = w8496 & w8545;
assign w8548 = ~w8546 & ~w8547;
assign w8549 = w8486 & w8548;
assign w8550 = ~w8486 & ~w8548;
assign w8551 = ~w8549 & ~w8550;
assign w8552 = w8485 & ~w8551;
assign w8553 = ~w8485 & w8551;
assign w8554 = ~w8552 & ~w8553;
assign w8555 = (~w8240 & ~w8160) | (~w8240 & w24839) | (~w8160 & w24839);
assign w8556 = w8554 & w8555;
assign w8557 = ~w8554 & ~w8555;
assign w8558 = ~w8556 & ~w8557;
assign w8559 = b[15] & w4453;
assign w8560 = b[16] & w4241;
assign w8561 = b[17] & w4243;
assign w8562 = w1008 & w4236;
assign w8563 = ~w8560 & ~w8561;
assign w8564 = ~w8559 & w8563;
assign w8565 = ~w8562 & w8564;
assign w8566 = a[38] & ~w8565;
assign w8567 = ~a[38] & w8565;
assign w8568 = ~w8566 & ~w8567;
assign w8569 = ~w8558 & ~w8568;
assign w8570 = w8558 & w8568;
assign w8571 = ~w8569 & ~w8570;
assign w8572 = ~w8475 & ~w8571;
assign w8573 = w8475 & w8571;
assign w8574 = ~w8572 & ~w8573;
assign w8575 = w8474 & ~w8574;
assign w8576 = ~w8474 & w8574;
assign w8577 = ~w8575 & ~w8576;
assign w8578 = w8464 & w8577;
assign w8579 = ~w8464 & ~w8577;
assign w8580 = ~w8578 & ~w8579;
assign w8581 = b[21] & w3177;
assign w8582 = b[23] & w2978;
assign w8583 = b[22] & w2973;
assign w8584 = w1755 & w2980;
assign w8585 = ~w8582 & ~w8583;
assign w8586 = ~w8581 & w8585;
assign w8587 = ~w8584 & w8586;
assign w8588 = a[32] & ~w8587;
assign w8589 = ~a[32] & w8587;
assign w8590 = ~w8588 & ~w8589;
assign w8591 = w8580 & w8590;
assign w8592 = ~w8580 & ~w8590;
assign w8593 = ~w8591 & ~w8592;
assign w8594 = ~w8463 & w8593;
assign w8595 = w8463 & ~w8593;
assign w8596 = ~w8594 & ~w8595;
assign w8597 = ~w8462 & ~w8596;
assign w8598 = w8462 & w8596;
assign w8599 = ~w8597 & ~w8598;
assign w8600 = (~w8276 & ~w8127) | (~w8276 & w24995) | (~w8127 & w24995);
assign w8601 = w8599 & w8600;
assign w8602 = ~w8599 & ~w8600;
assign w8603 = ~w8601 & ~w8602;
assign w8604 = b[29] & w1957;
assign w8605 = b[27] & ~w2114;
assign w8606 = b[28] & w1955;
assign w8607 = w1951 & w2734;
assign w8608 = ~w8604 & ~w8605;
assign w8609 = ~w8606 & w8608;
assign w8610 = ~w8607 & w8609;
assign w8611 = a[26] & ~w8610;
assign w8612 = ~a[26] & w8610;
assign w8613 = ~w8611 & ~w8612;
assign w8614 = ~w8603 & ~w8613;
assign w8615 = w8603 & w8613;
assign w8616 = ~w8614 & ~w8615;
assign w8617 = ~w8452 & ~w8616;
assign w8618 = w8452 & w8616;
assign w8619 = ~w8617 & ~w8618;
assign w8620 = w8451 & ~w8619;
assign w8621 = ~w8451 & w8619;
assign w8622 = ~w8620 & ~w8621;
assign w8623 = ~w8441 & w8622;
assign w8624 = w8441 & ~w8622;
assign w8625 = ~w8623 & ~w8624;
assign w8626 = b[33] & ~w1272;
assign w8627 = b[35] & w1156;
assign w8628 = b[34] & w1154;
assign w8629 = w1150 & w3918;
assign w8630 = ~w8626 & ~w8627;
assign w8631 = ~w8628 & w8630;
assign w8632 = ~w8629 & w8631;
assign w8633 = a[20] & ~w8632;
assign w8634 = ~a[20] & w8632;
assign w8635 = ~w8633 & ~w8634;
assign w8636 = w8625 & w8635;
assign w8637 = ~w8625 & ~w8635;
assign w8638 = ~w8636 & ~w8637;
assign w8639 = ~w8440 & ~w8638;
assign w8640 = w8440 & w8638;
assign w8641 = ~w8639 & ~w8640;
assign w8642 = ~w8439 & w8641;
assign w8643 = w8439 & ~w8641;
assign w8644 = ~w8642 & ~w8643;
assign w8645 = (~w8312 & ~w8095) | (~w8312 & w25161) | (~w8095 & w25161);
assign w8646 = w8644 & w8645;
assign w8647 = ~w8644 & ~w8645;
assign w8648 = ~w8646 & ~w8647;
assign w8649 = w8429 & w8648;
assign w8650 = ~w8429 & ~w8648;
assign w8651 = ~w8649 & ~w8650;
assign w8652 = ~w8419 & w8651;
assign w8653 = w8419 & ~w8651;
assign w8654 = ~w8652 & ~w8653;
assign w8655 = w8418 & w8654;
assign w8656 = ~w8418 & ~w8654;
assign w8657 = ~w8655 & ~w8656;
assign w8658 = (~w8334 & ~w8336) | (~w8334 & w25287) | (~w8336 & w25287);
assign w8659 = w8657 & w8658;
assign w8660 = ~w8657 & ~w8658;
assign w8661 = ~w8659 & ~w8660;
assign w8662 = w8408 & w8661;
assign w8663 = ~w8408 & ~w8661;
assign w8664 = ~w8662 & ~w8663;
assign w8665 = w8398 & w8664;
assign w8666 = ~w8398 & ~w8664;
assign w8667 = ~w8665 & ~w8666;
assign w8668 = w8397 & ~w8667;
assign w8669 = ~w8397 & w8667;
assign w8670 = ~w8668 & ~w8669;
assign w8671 = (~w8358 & ~w8073) | (~w8358 & w24676) | (~w8073 & w24676);
assign w8672 = w8670 & w8671;
assign w8673 = ~w8670 & ~w8671;
assign w8674 = ~w8672 & ~w8673;
assign w8675 = b[53] & w11;
assign w8676 = b[52] & w9;
assign w8677 = ~b[52] & ~b[53];
assign w8678 = b[52] & b[53];
assign w8679 = ~w8677 & ~w8678;
assign w8680 = (~w8365 & w8368) | (~w8365 & w24840) | (w8368 & w24840);
assign w8681 = w8679 & w8680;
assign w8682 = ~w8679 & ~w8680;
assign w8683 = ~w8681 & ~w8682;
assign w8684 = w5 & w8683;
assign w8685 = ~w8675 & ~w8676;
assign w8686 = ~w8684 & w8685;
assign w8687 = b[51] & w24;
assign w8688 = a[2] & ~w8687;
assign w8689 = w8686 & ~w8688;
assign w8690 = a[2] & ~w8686;
assign w8691 = ~w8689 & ~w8690;
assign w8692 = w8674 & w8691;
assign w8693 = ~w8674 & ~w8691;
assign w8694 = ~w8692 & ~w8693;
assign w8695 = w8387 & ~w8694;
assign w8696 = ~w8387 & w8694;
assign w8697 = ~w8695 & ~w8696;
assign w8698 = ~w8668 & ~w8672;
assign w8699 = b[48] & w185;
assign w8700 = b[46] & ~w237;
assign w8701 = b[47] & w183;
assign w8702 = w179 & ~w7170;
assign w8703 = ~w8699 & ~w8700;
assign w8704 = ~w8701 & w8703;
assign w8705 = ~w8702 & w8704;
assign w8706 = a[8] & ~w8705;
assign w8707 = ~a[8] & w8705;
assign w8708 = ~w8706 & ~w8707;
assign w8709 = (~w8655 & ~w8658) | (~w8655 & w25430) | (~w8658 & w25430);
assign w8710 = b[45] & w360;
assign w8711 = b[44] & w358;
assign w8712 = b[43] & ~w419;
assign w8713 = w354 & w6334;
assign w8714 = ~w8710 & ~w8711;
assign w8715 = ~w8712 & w8714;
assign w8716 = ~w8713 & w8715;
assign w8717 = a[11] & ~w8716;
assign w8718 = ~a[11] & w8716;
assign w8719 = ~w8717 & ~w8718;
assign w8720 = (~w8649 & w8419) | (~w8649 & w25162) | (w8419 & w25162);
assign w8721 = b[41] & w573;
assign w8722 = b[42] & w575;
assign w8723 = b[40] & ~w649;
assign w8724 = w569 & w5548;
assign w8725 = ~w8721 & ~w8722;
assign w8726 = ~w8723 & w8725;
assign w8727 = ~w8724 & w8726;
assign w8728 = a[14] & ~w8727;
assign w8729 = ~a[14] & w8727;
assign w8730 = ~w8728 & ~w8729;
assign w8731 = (~w8643 & ~w8645) | (~w8643 & w24996) | (~w8645 & w24996);
assign w8732 = b[34] & ~w1272;
assign w8733 = b[36] & w1156;
assign w8734 = b[35] & w1154;
assign w8735 = w1150 & w4129;
assign w8736 = ~w8732 & ~w8733;
assign w8737 = ~w8734 & w8736;
assign w8738 = ~w8735 & w8737;
assign w8739 = a[20] & ~w8738;
assign w8740 = ~a[20] & w8738;
assign w8741 = ~w8739 & ~w8740;
assign w8742 = (~w8620 & w8441) | (~w8620 & w24841) | (w8441 & w24841);
assign w8743 = b[32] & w1517;
assign w8744 = b[33] & w1519;
assign w8745 = b[31] & ~w1676;
assign w8746 = w1513 & w3499;
assign w8747 = ~w8743 & ~w8744;
assign w8748 = ~w8745 & w8747;
assign w8749 = ~w8746 & w8748;
assign w8750 = a[23] & ~w8749;
assign w8751 = ~a[23] & w8749;
assign w8752 = ~w8750 & ~w8751;
assign w8753 = b[30] & w1957;
assign w8754 = b[29] & w1955;
assign w8755 = b[28] & ~w2114;
assign w8756 = w1951 & ~w2908;
assign w8757 = ~w8753 & ~w8754;
assign w8758 = ~w8755 & w8757;
assign w8759 = ~w8756 & w8758;
assign w8760 = a[26] & ~w8759;
assign w8761 = ~a[26] & w8759;
assign w8762 = ~w8760 & ~w8761;
assign w8763 = (~w8598 & ~w8600) | (~w8598 & w24842) | (~w8600 & w24842);
assign w8764 = b[25] & ~w2622;
assign w8765 = b[27] & w2438;
assign w8766 = b[26] & w2436;
assign w8767 = w2378 & w2432;
assign w8768 = ~w8764 & ~w8765;
assign w8769 = ~w8766 & w8768;
assign w8770 = ~w8767 & w8769;
assign w8771 = a[29] & ~w8770;
assign w8772 = ~a[29] & w8770;
assign w8773 = ~w8771 & ~w8772;
assign w8774 = (~w8591 & w8463) | (~w8591 & w25163) | (w8463 & w25163);
assign w8775 = b[22] & w3177;
assign w8776 = b[23] & w2973;
assign w8777 = b[24] & w2978;
assign w8778 = w1895 & w2980;
assign w8779 = ~w8776 & ~w8777;
assign w8780 = ~w8775 & w8779;
assign w8781 = ~w8778 & w8780;
assign w8782 = a[32] & ~w8781;
assign w8783 = ~a[32] & w8781;
assign w8784 = ~w8782 & ~w8783;
assign w8785 = (~w8575 & ~w8464) | (~w8575 & w25288) | (~w8464 & w25288);
assign w8786 = b[16] & w4453;
assign w8787 = b[18] & w4243;
assign w8788 = b[17] & w4241;
assign w8789 = ~w1108 & w4236;
assign w8790 = ~w8787 & ~w8788;
assign w8791 = ~w8786 & w8790;
assign w8792 = ~w8789 & w8791;
assign w8793 = a[38] & ~w8792;
assign w8794 = ~a[38] & w8792;
assign w8795 = ~w8793 & ~w8794;
assign w8796 = ~w8552 & ~w8556;
assign w8797 = b[13] & w5167;
assign w8798 = b[15] & w4925;
assign w8799 = b[14] & w4918;
assign w8800 = ~w799 & w4923;
assign w8801 = ~w8798 & ~w8799;
assign w8802 = ~w8797 & w8801;
assign w8803 = ~w8800 & w8802;
assign w8804 = a[41] & ~w8803;
assign w8805 = ~a[41] & w8803;
assign w8806 = ~w8804 & ~w8805;
assign w8807 = b[10] & w5939;
assign w8808 = b[11] & w5670;
assign w8809 = b[12] & w5665;
assign w8810 = w536 & w5663;
assign w8811 = ~w8808 & ~w8809;
assign w8812 = ~w8807 & w8811;
assign w8813 = ~w8810 & w8812;
assign w8814 = a[44] & ~w8813;
assign w8815 = ~a[44] & w8813;
assign w8816 = ~w8814 & ~w8815;
assign w8817 = ~w8540 & ~w8543;
assign w8818 = b[7] & w6732;
assign w8819 = b[9] & w6476;
assign w8820 = b[8] & w6474;
assign w8821 = w322 & w6469;
assign w8822 = ~w8819 & ~w8820;
assign w8823 = ~w8818 & w8822;
assign w8824 = ~w8821 & w8823;
assign w8825 = a[47] & ~w8824;
assign w8826 = ~a[47] & w8824;
assign w8827 = ~w8825 & ~w8826;
assign w8828 = a[53] & ~a[54];
assign w8829 = ~a[53] & a[54];
assign w8830 = ~w8828 & ~w8829;
assign w8831 = b[0] & ~w8830;
assign w8832 = w8509 & w8519;
assign w8833 = w8514 & w24997;
assign w8834 = b[3] & w8202;
assign w8835 = b[2] & w8200;
assign w8836 = w46 & w8195;
assign w8837 = ~w8834 & ~w8835;
assign w8838 = ~w8833 & w8837;
assign w8839 = (a[53] & ~w8838) | (a[53] & w24998) | (~w8838 & w24998);
assign w8840 = w8838 & w24999;
assign w8841 = ~w8839 & ~w8840;
assign w8842 = w8832 & w8841;
assign w8843 = ~w8832 & ~w8841;
assign w8844 = ~w8842 & ~w8843;
assign w8845 = w8831 & w8844;
assign w8846 = ~w8831 & ~w8844;
assign w8847 = ~w8845 & ~w8846;
assign w8848 = b[4] & w7586;
assign w8849 = b[6] & w7314;
assign w8850 = b[5] & w7307;
assign w8851 = w157 & w7312;
assign w8852 = ~w8849 & ~w8850;
assign w8853 = ~w8848 & w8852;
assign w8854 = ~w8851 & w8853;
assign w8855 = a[50] & ~w8854;
assign w8856 = ~a[50] & w8854;
assign w8857 = ~w8855 & ~w8856;
assign w8858 = w8847 & w8857;
assign w8859 = ~w8847 & ~w8857;
assign w8860 = ~w8858 & ~w8859;
assign w8861 = (~w8524 & ~w8497) | (~w8524 & w25164) | (~w8497 & w25164);
assign w8862 = w8860 & w8861;
assign w8863 = ~w8860 & ~w8861;
assign w8864 = ~w8862 & ~w8863;
assign w8865 = ~w8827 & ~w8864;
assign w8866 = w8827 & w8864;
assign w8867 = ~w8865 & ~w8866;
assign w8868 = w8817 & w8867;
assign w8869 = ~w8817 & ~w8867;
assign w8870 = ~w8868 & ~w8869;
assign w8871 = ~w8816 & w8870;
assign w8872 = w8816 & ~w8870;
assign w8873 = ~w8871 & ~w8872;
assign w8874 = (~w8546 & ~w8486) | (~w8546 & w25165) | (~w8486 & w25165);
assign w8875 = w8873 & w8874;
assign w8876 = ~w8873 & ~w8874;
assign w8877 = ~w8875 & ~w8876;
assign w8878 = w8806 & w8877;
assign w8879 = ~w8806 & ~w8877;
assign w8880 = ~w8878 & ~w8879;
assign w8881 = w8796 & w8880;
assign w8882 = ~w8796 & ~w8880;
assign w8883 = ~w8881 & ~w8882;
assign w8884 = ~w8795 & w8883;
assign w8885 = w8795 & ~w8883;
assign w8886 = ~w8884 & ~w8885;
assign w8887 = (~w8569 & ~w8475) | (~w8569 & w24843) | (~w8475 & w24843);
assign w8888 = w8886 & w8887;
assign w8889 = ~w8886 & ~w8887;
assign w8890 = ~w8888 & ~w8889;
assign w8891 = b[19] & w3785;
assign w8892 = b[20] & w3578;
assign w8893 = b[21] & w3580;
assign w8894 = w1467 & w3573;
assign w8895 = ~w8892 & ~w8893;
assign w8896 = ~w8891 & w8895;
assign w8897 = ~w8894 & w8896;
assign w8898 = a[35] & ~w8897;
assign w8899 = ~a[35] & w8897;
assign w8900 = ~w8898 & ~w8899;
assign w8901 = w8890 & w8900;
assign w8902 = ~w8890 & ~w8900;
assign w8903 = ~w8901 & ~w8902;
assign w8904 = ~w8785 & ~w8903;
assign w8905 = w8785 & w8903;
assign w8906 = ~w8904 & ~w8905;
assign w8907 = w8784 & ~w8906;
assign w8908 = ~w8784 & w8906;
assign w8909 = ~w8907 & ~w8908;
assign w8910 = ~w8774 & w8909;
assign w8911 = w8774 & ~w8909;
assign w8912 = ~w8910 & ~w8911;
assign w8913 = w8773 & w8912;
assign w8914 = ~w8773 & ~w8912;
assign w8915 = ~w8913 & ~w8914;
assign w8916 = w8763 & w8915;
assign w8917 = ~w8763 & ~w8915;
assign w8918 = ~w8916 & ~w8917;
assign w8919 = w8762 & ~w8918;
assign w8920 = ~w8762 & w8918;
assign w8921 = ~w8919 & ~w8920;
assign w8922 = (~w8614 & ~w8452) | (~w8614 & w25000) | (~w8452 & w25000);
assign w8923 = w8921 & w8922;
assign w8924 = ~w8921 & ~w8922;
assign w8925 = ~w8923 & ~w8924;
assign w8926 = w8752 & w8925;
assign w8927 = ~w8752 & ~w8925;
assign w8928 = ~w8926 & ~w8927;
assign w8929 = ~w8742 & w8928;
assign w8930 = w8742 & ~w8928;
assign w8931 = ~w8929 & ~w8930;
assign w8932 = w8741 & w8931;
assign w8933 = ~w8741 & ~w8931;
assign w8934 = ~w8932 & ~w8933;
assign w8935 = (~w8637 & ~w8440) | (~w8637 & w24389) | (~w8440 & w24389);
assign w8936 = ~w8934 & ~w8935;
assign w8937 = w8934 & w8935;
assign w8938 = ~w8936 & ~w8937;
assign w8939 = b[39] & w834;
assign w8940 = b[37] & ~w934;
assign w8941 = b[38] & w838;
assign w8942 = w832 & ~w4812;
assign w8943 = ~w8939 & ~w8940;
assign w8944 = ~w8941 & w8943;
assign w8945 = ~w8942 & w8944;
assign w8946 = a[17] & ~w8945;
assign w8947 = ~a[17] & w8945;
assign w8948 = ~w8946 & ~w8947;
assign w8949 = w8938 & w8948;
assign w8950 = ~w8938 & ~w8948;
assign w8951 = ~w8949 & ~w8950;
assign w8952 = w8731 & ~w8951;
assign w8953 = ~w8731 & w8951;
assign w8954 = ~w8952 & ~w8953;
assign w8955 = ~w8730 & ~w8954;
assign w8956 = w8730 & w8954;
assign w8957 = ~w8955 & ~w8956;
assign w8958 = ~w8720 & w8957;
assign w8959 = w8720 & ~w8957;
assign w8960 = ~w8958 & ~w8959;
assign w8961 = ~w8719 & ~w8960;
assign w8962 = w8719 & w8960;
assign w8963 = ~w8961 & ~w8962;
assign w8964 = ~w8709 & ~w8963;
assign w8965 = w8709 & w8963;
assign w8966 = ~w8964 & ~w8965;
assign w8967 = w8708 & ~w8966;
assign w8968 = ~w8708 & w8966;
assign w8969 = ~w8967 & ~w8968;
assign w8970 = (~w8663 & ~w8398) | (~w8663 & w25289) | (~w8398 & w25289);
assign w8971 = ~w8969 & ~w8970;
assign w8972 = w8969 & w8970;
assign w8973 = ~w8971 & ~w8972;
assign w8974 = b[49] & w103;
assign w8975 = b[51] & w68;
assign w8976 = b[50] & w61;
assign w8977 = w66 & ~w8058;
assign w8978 = ~w8975 & ~w8976;
assign w8979 = ~w8974 & w8978;
assign w8980 = ~w8977 & w8979;
assign w8981 = a[5] & ~w8980;
assign w8982 = ~a[5] & w8980;
assign w8983 = ~w8981 & ~w8982;
assign w8984 = ~w8973 & ~w8983;
assign w8985 = w8973 & w8983;
assign w8986 = ~w8984 & ~w8985;
assign w8987 = w8698 & w8986;
assign w8988 = ~w8698 & ~w8986;
assign w8989 = ~w8987 & ~w8988;
assign w8990 = b[54] & w11;
assign w8991 = b[53] & w9;
assign w8992 = ~w8678 & ~w8681;
assign w8993 = ~b[53] & ~b[54];
assign w8994 = b[53] & b[54];
assign w8995 = ~w8993 & ~w8994;
assign w8996 = ~w8992 & ~w8995;
assign w8997 = w8992 & w8995;
assign w8998 = ~w8996 & ~w8997;
assign w8999 = w5 & ~w8998;
assign w9000 = ~w8990 & ~w8991;
assign w9001 = ~w8999 & w9000;
assign w9002 = b[52] & w24;
assign w9003 = a[2] & ~w9002;
assign w9004 = w9001 & ~w9003;
assign w9005 = a[2] & ~w9001;
assign w9006 = ~w9004 & ~w9005;
assign w9007 = ~w8989 & w9006;
assign w9008 = w8989 & ~w9006;
assign w9009 = ~w9007 & ~w9008;
assign w9010 = (~w8692 & w8387) | (~w8692 & w24677) | (w8387 & w24677);
assign w9011 = w9009 & ~w9010;
assign w9012 = ~w9009 & w9010;
assign w9013 = ~w9011 & ~w9012;
assign w9014 = ~w9007 & ~w9011;
assign w9015 = b[50] & w103;
assign w9016 = b[51] & w61;
assign w9017 = b[52] & w68;
assign w9018 = w66 & ~w8371;
assign w9019 = ~w9016 & ~w9017;
assign w9020 = ~w9015 & w9019;
assign w9021 = ~w9018 & w9020;
assign w9022 = a[5] & ~w9021;
assign w9023 = ~a[5] & w9021;
assign w9024 = ~w9022 & ~w9023;
assign w9025 = (~w8967 & ~w8970) | (~w8967 & w25431) | (~w8970 & w25431);
assign w9026 = b[49] & w185;
assign w9027 = b[47] & ~w237;
assign w9028 = b[48] & w183;
assign w9029 = w179 & ~w7468;
assign w9030 = ~w9026 & ~w9027;
assign w9031 = ~w9028 & w9030;
assign w9032 = ~w9029 & w9031;
assign w9033 = a[8] & ~w9032;
assign w9034 = ~a[8] & w9032;
assign w9035 = ~w9033 & ~w9034;
assign w9036 = b[44] & ~w419;
assign w9037 = b[46] & w360;
assign w9038 = b[45] & w358;
assign w9039 = w354 & ~w6613;
assign w9040 = ~w9036 & ~w9037;
assign w9041 = ~w9038 & w9040;
assign w9042 = ~w9039 & w9041;
assign w9043 = a[11] & ~w9042;
assign w9044 = ~a[11] & w9042;
assign w9045 = ~w9043 & ~w9044;
assign w9046 = (~w8956 & w8720) | (~w8956 & w25001) | (w8720 & w25001);
assign w9047 = b[38] & ~w934;
assign w9048 = b[39] & w838;
assign w9049 = b[40] & w834;
assign w9050 = w832 & ~w5058;
assign w9051 = ~w9047 & ~w9048;
assign w9052 = ~w9049 & w9051;
assign w9053 = ~w9050 & w9052;
assign w9054 = a[17] & ~w9053;
assign w9055 = ~a[17] & w9053;
assign w9056 = ~w9054 & ~w9055;
assign w9057 = (~w8932 & ~w8935) | (~w8932 & w24844) | (~w8935 & w24844);
assign w9058 = (~w8926 & w8742) | (~w8926 & w25002) | (w8742 & w25002);
assign w9059 = b[34] & w1519;
assign w9060 = b[32] & ~w1676;
assign w9061 = b[33] & w1517;
assign w9062 = w1513 & ~w3710;
assign w9063 = ~w9059 & ~w9060;
assign w9064 = ~w9061 & w9063;
assign w9065 = ~w9062 & w9064;
assign w9066 = a[23] & ~w9065;
assign w9067 = ~a[23] & w9065;
assign w9068 = ~w9066 & ~w9067;
assign w9069 = (~w8919 & ~w8922) | (~w8919 & w24678) | (~w8922 & w24678);
assign w9070 = b[26] & ~w2622;
assign w9071 = b[27] & w2436;
assign w9072 = b[28] & w2438;
assign w9073 = w2432 & w2559;
assign w9074 = ~w9070 & ~w9071;
assign w9075 = ~w9072 & w9074;
assign w9076 = ~w9073 & w9075;
assign w9077 = a[29] & ~w9076;
assign w9078 = ~a[29] & w9076;
assign w9079 = ~w9077 & ~w9078;
assign w9080 = (~w8907 & w8774) | (~w8907 & w24679) | (w8774 & w24679);
assign w9081 = b[23] & w3177;
assign w9082 = b[24] & w2973;
assign w9083 = b[25] & w2978;
assign w9084 = w2061 & w2980;
assign w9085 = ~w9082 & ~w9083;
assign w9086 = ~w9081 & w9085;
assign w9087 = ~w9084 & w9086;
assign w9088 = a[32] & ~w9087;
assign w9089 = ~a[32] & w9087;
assign w9090 = ~w9088 & ~w9089;
assign w9091 = b[20] & w3785;
assign w9092 = b[21] & w3578;
assign w9093 = b[22] & w3580;
assign w9094 = w1615 & w3573;
assign w9095 = ~w9092 & ~w9093;
assign w9096 = ~w9091 & w9095;
assign w9097 = ~w9094 & w9096;
assign w9098 = a[35] & ~w9097;
assign w9099 = ~a[35] & w9097;
assign w9100 = ~w9098 & ~w9099;
assign w9101 = ~w8885 & ~w8888;
assign w9102 = b[17] & w4453;
assign w9103 = b[19] & w4243;
assign w9104 = b[18] & w4241;
assign w9105 = ~w1231 & w4236;
assign w9106 = ~w9103 & ~w9104;
assign w9107 = ~w9102 & w9106;
assign w9108 = ~w9105 & w9107;
assign w9109 = a[38] & ~w9108;
assign w9110 = ~a[38] & w9108;
assign w9111 = ~w9109 & ~w9110;
assign w9112 = b[14] & w5167;
assign w9113 = b[16] & w4925;
assign w9114 = b[15] & w4918;
assign w9115 = w905 & w4923;
assign w9116 = ~w9113 & ~w9114;
assign w9117 = ~w9112 & w9116;
assign w9118 = ~w9115 & w9117;
assign w9119 = a[41] & ~w9118;
assign w9120 = ~a[41] & w9118;
assign w9121 = ~w9119 & ~w9120;
assign w9122 = ~w8872 & ~w8875;
assign w9123 = b[11] & w5939;
assign w9124 = b[12] & w5670;
assign w9125 = b[13] & w5665;
assign w9126 = w628 & w5663;
assign w9127 = ~w9124 & ~w9125;
assign w9128 = ~w9123 & w9127;
assign w9129 = ~w9126 & w9128;
assign w9130 = a[44] & ~w9129;
assign w9131 = ~a[44] & w9129;
assign w9132 = ~w9130 & ~w9131;
assign w9133 = b[8] & w6732;
assign w9134 = b[10] & w6476;
assign w9135 = b[9] & w6474;
assign w9136 = w397 & w6469;
assign w9137 = ~w9134 & ~w9135;
assign w9138 = ~w9133 & w9137;
assign w9139 = ~w9136 & w9138;
assign w9140 = a[47] & ~w9139;
assign w9141 = ~a[47] & w9139;
assign w9142 = ~w9140 & ~w9141;
assign w9143 = ~w8858 & ~w8862;
assign w9144 = b[2] & w8515;
assign w9145 = b[3] & w8200;
assign w9146 = b[4] & w8202;
assign w9147 = w84 & w8195;
assign w9148 = ~w9145 & ~w9146;
assign w9149 = ~w9144 & w9148;
assign w9150 = ~w9147 & w9149;
assign w9151 = a[53] & ~w9150;
assign w9152 = ~a[53] & w9150;
assign w9153 = ~w9151 & ~w9152;
assign w9154 = a[56] & w8831;
assign w9155 = a[55] & ~a[56];
assign w9156 = ~a[55] & a[56];
assign w9157 = ~w9155 & ~w9156;
assign w9158 = ~w8830 & ~w9157;
assign w9159 = ~w8 & w9158;
assign w9160 = ~w8830 & w9157;
assign w9161 = b[1] & w9160;
assign w9162 = a[54] & ~a[55];
assign w9163 = ~a[54] & a[55];
assign w9164 = ~w9162 & ~w9163;
assign w9165 = w8830 & ~w9164;
assign w9166 = b[0] & w9165;
assign w9167 = ~w9159 & ~w9161;
assign w9168 = ~w9166 & w9167;
assign w9169 = ~w9154 & w9168;
assign w9170 = w9154 & ~w9168;
assign w9171 = ~w9169 & ~w9170;
assign w9172 = ~w9153 & ~w9171;
assign w9173 = w9153 & w9171;
assign w9174 = ~w9172 & ~w9173;
assign w9175 = (~w8842 & ~w8844) | (~w8842 & w25166) | (~w8844 & w25166);
assign w9176 = w9174 & ~w9175;
assign w9177 = ~w9174 & w9175;
assign w9178 = ~w9176 & ~w9177;
assign w9179 = b[5] & w7586;
assign w9180 = b[6] & w7307;
assign w9181 = b[7] & w7314;
assign w9182 = w216 & w7312;
assign w9183 = ~w9180 & ~w9181;
assign w9184 = ~w9179 & w9183;
assign w9185 = ~w9182 & w9184;
assign w9186 = a[50] & ~w9185;
assign w9187 = ~a[50] & w9185;
assign w9188 = ~w9186 & ~w9187;
assign w9189 = ~w9178 & ~w9188;
assign w9190 = w9178 & w9188;
assign w9191 = ~w9189 & ~w9190;
assign w9192 = w9143 & w9191;
assign w9193 = ~w9143 & ~w9191;
assign w9194 = ~w9192 & ~w9193;
assign w9195 = ~w9142 & w9194;
assign w9196 = w9142 & ~w9194;
assign w9197 = ~w9195 & ~w9196;
assign w9198 = (~w8865 & ~w8817) | (~w8865 & w25167) | (~w8817 & w25167);
assign w9199 = w9197 & w9198;
assign w9200 = ~w9197 & ~w9198;
assign w9201 = ~w9199 & ~w9200;
assign w9202 = ~w9132 & ~w9201;
assign w9203 = w9132 & w9201;
assign w9204 = ~w9202 & ~w9203;
assign w9205 = ~w9122 & ~w9204;
assign w9206 = w9122 & w9204;
assign w9207 = ~w9205 & ~w9206;
assign w9208 = ~w9121 & w9207;
assign w9209 = w9121 & ~w9207;
assign w9210 = ~w9208 & ~w9209;
assign w9211 = (~w8879 & ~w8796) | (~w8879 & w24680) | (~w8796 & w24680);
assign w9212 = ~w9210 & ~w9211;
assign w9213 = w9210 & w9211;
assign w9214 = ~w9212 & ~w9213;
assign w9215 = ~w9111 & ~w9214;
assign w9216 = w9111 & w9214;
assign w9217 = ~w9215 & ~w9216;
assign w9218 = ~w9101 & ~w9217;
assign w9219 = w9101 & w9217;
assign w9220 = ~w9218 & ~w9219;
assign w9221 = w9100 & ~w9220;
assign w9222 = ~w9100 & w9220;
assign w9223 = ~w9221 & ~w9222;
assign w9224 = (~w8902 & ~w8785) | (~w8902 & w24681) | (~w8785 & w24681);
assign w9225 = w9223 & w9224;
assign w9226 = ~w9223 & ~w9224;
assign w9227 = ~w9225 & ~w9226;
assign w9228 = w9090 & w9227;
assign w9229 = ~w9090 & ~w9227;
assign w9230 = ~w9228 & ~w9229;
assign w9231 = ~w9080 & w9230;
assign w9232 = w9080 & ~w9230;
assign w9233 = ~w9231 & ~w9232;
assign w9234 = w9079 & w9233;
assign w9235 = ~w9079 & ~w9233;
assign w9236 = ~w9234 & ~w9235;
assign w9237 = (~w8914 & ~w8763) | (~w8914 & w25168) | (~w8763 & w25168);
assign w9238 = ~w9236 & ~w9237;
assign w9239 = w9236 & w9237;
assign w9240 = ~w9238 & ~w9239;
assign w9241 = b[29] & ~w2114;
assign w9242 = b[31] & w1957;
assign w9243 = b[30] & w1955;
assign w9244 = w1951 & ~w3112;
assign w9245 = ~w9241 & ~w9242;
assign w9246 = ~w9243 & w9245;
assign w9247 = ~w9244 & w9246;
assign w9248 = a[26] & ~w9247;
assign w9249 = ~a[26] & w9247;
assign w9250 = ~w9248 & ~w9249;
assign w9251 = w9240 & w9250;
assign w9252 = ~w9240 & ~w9250;
assign w9253 = ~w9251 & ~w9252;
assign w9254 = w9069 & ~w9253;
assign w9255 = ~w9069 & w9253;
assign w9256 = ~w9254 & ~w9255;
assign w9257 = ~w9068 & ~w9256;
assign w9258 = w9068 & w9256;
assign w9259 = ~w9257 & ~w9258;
assign w9260 = w9058 & ~w9259;
assign w9261 = ~w9058 & w9259;
assign w9262 = ~w9260 & ~w9261;
assign w9263 = b[35] & ~w1272;
assign w9264 = b[37] & w1156;
assign w9265 = b[36] & w1154;
assign w9266 = w1150 & ~w4357;
assign w9267 = ~w9263 & ~w9264;
assign w9268 = ~w9265 & w9267;
assign w9269 = ~w9266 & w9268;
assign w9270 = a[20] & ~w9269;
assign w9271 = ~a[20] & w9269;
assign w9272 = ~w9270 & ~w9271;
assign w9273 = w9262 & w9272;
assign w9274 = ~w9262 & ~w9272;
assign w9275 = ~w9273 & ~w9274;
assign w9276 = ~w9057 & ~w9275;
assign w9277 = w9057 & w9275;
assign w9278 = ~w9276 & ~w9277;
assign w9279 = ~w9056 & w9278;
assign w9280 = w9056 & ~w9278;
assign w9281 = ~w9279 & ~w9280;
assign w9282 = (~w8949 & w8731) | (~w8949 & w24390) | (w8731 & w24390);
assign w9283 = ~w9281 & w9282;
assign w9284 = w9281 & ~w9282;
assign w9285 = ~w9283 & ~w9284;
assign w9286 = b[41] & ~w649;
assign w9287 = b[42] & w573;
assign w9288 = b[43] & w575;
assign w9289 = w569 & w5811;
assign w9290 = ~w9286 & ~w9287;
assign w9291 = ~w9288 & w9290;
assign w9292 = ~w9289 & w9291;
assign w9293 = a[14] & ~w9292;
assign w9294 = ~a[14] & w9292;
assign w9295 = ~w9293 & ~w9294;
assign w9296 = ~w9285 & ~w9295;
assign w9297 = w9285 & w9295;
assign w9298 = ~w9296 & ~w9297;
assign w9299 = w9046 & ~w9298;
assign w9300 = ~w9046 & w9298;
assign w9301 = ~w9299 & ~w9300;
assign w9302 = w9045 & w9301;
assign w9303 = ~w9045 & ~w9301;
assign w9304 = ~w9302 & ~w9303;
assign w9305 = (~w8961 & ~w8709) | (~w8961 & w25169) | (~w8709 & w25169);
assign w9306 = w9304 & w9305;
assign w9307 = ~w9304 & ~w9305;
assign w9308 = ~w9306 & ~w9307;
assign w9309 = ~w9035 & ~w9308;
assign w9310 = w9035 & w9308;
assign w9311 = ~w9309 & ~w9310;
assign w9312 = w9025 & w9311;
assign w9313 = ~w9025 & ~w9311;
assign w9314 = ~w9312 & ~w9313;
assign w9315 = w9024 & ~w9314;
assign w9316 = ~w9024 & w9314;
assign w9317 = ~w9315 & ~w9316;
assign w9318 = (~w8984 & ~w8698) | (~w8984 & w25290) | (~w8698 & w25290);
assign w9319 = w9317 & w9318;
assign w9320 = ~w9317 & ~w9318;
assign w9321 = ~w9319 & ~w9320;
assign w9322 = b[55] & w11;
assign w9323 = b[54] & w9;
assign w9324 = ~b[54] & ~b[55];
assign w9325 = b[54] & b[55];
assign w9326 = ~w9324 & ~w9325;
assign w9327 = (~w8993 & ~w8992) | (~w8993 & w24682) | (~w8992 & w24682);
assign w9328 = ~w9326 & w9327;
assign w9329 = w9326 & ~w9327;
assign w9330 = ~w9328 & ~w9329;
assign w9331 = w5 & ~w9330;
assign w9332 = ~w9322 & ~w9323;
assign w9333 = ~w9331 & w9332;
assign w9334 = b[53] & w24;
assign w9335 = a[2] & ~w9334;
assign w9336 = w9333 & ~w9335;
assign w9337 = a[2] & ~w9333;
assign w9338 = ~w9336 & ~w9337;
assign w9339 = w9321 & w9338;
assign w9340 = ~w9321 & ~w9338;
assign w9341 = ~w9339 & ~w9340;
assign w9342 = w9014 & ~w9341;
assign w9343 = ~w9014 & w9341;
assign w9344 = ~w9342 & ~w9343;
assign w9345 = (~w9315 & ~w9318) | (~w9315 & w25432) | (~w9318 & w25432);
assign w9346 = b[51] & w103;
assign w9347 = b[52] & w61;
assign w9348 = b[53] & w68;
assign w9349 = w66 & w8683;
assign w9350 = ~w9347 & ~w9348;
assign w9351 = ~w9346 & w9350;
assign w9352 = ~w9349 & w9351;
assign w9353 = a[5] & ~w9352;
assign w9354 = ~a[5] & w9352;
assign w9355 = ~w9353 & ~w9354;
assign w9356 = b[48] & ~w237;
assign w9357 = b[50] & w185;
assign w9358 = b[49] & w183;
assign w9359 = w179 & w7759;
assign w9360 = ~w9356 & ~w9357;
assign w9361 = ~w9358 & w9360;
assign w9362 = ~w9359 & w9361;
assign w9363 = a[8] & ~w9362;
assign w9364 = ~a[8] & w9362;
assign w9365 = ~w9363 & ~w9364;
assign w9366 = (~w9302 & ~w9305) | (~w9302 & w25003) | (~w9305 & w25003);
assign w9367 = b[46] & w358;
assign w9368 = b[45] & ~w419;
assign w9369 = b[47] & w360;
assign w9370 = w354 & w6889;
assign w9371 = ~w9367 & ~w9368;
assign w9372 = ~w9369 & w9371;
assign w9373 = ~w9370 & w9372;
assign w9374 = a[11] & ~w9373;
assign w9375 = ~a[11] & w9373;
assign w9376 = ~w9374 & ~w9375;
assign w9377 = b[42] & ~w649;
assign w9378 = b[43] & w573;
assign w9379 = b[44] & w575;
assign w9380 = w569 & w6069;
assign w9381 = ~w9377 & ~w9378;
assign w9382 = ~w9379 & w9381;
assign w9383 = ~w9380 & w9382;
assign w9384 = a[14] & ~w9383;
assign w9385 = ~a[14] & w9383;
assign w9386 = ~w9384 & ~w9385;
assign w9387 = (~w9280 & w9282) | (~w9280 & w24845) | (w9282 & w24845);
assign w9388 = b[37] & w1154;
assign w9389 = b[38] & w1156;
assign w9390 = b[36] & ~w1272;
assign w9391 = w1150 & w4582;
assign w9392 = ~w9388 & ~w9389;
assign w9393 = ~w9390 & w9392;
assign w9394 = ~w9391 & w9393;
assign w9395 = a[20] & ~w9394;
assign w9396 = ~a[20] & w9394;
assign w9397 = ~w9395 & ~w9396;
assign w9398 = (~w9258 & w9058) | (~w9258 & w24683) | (w9058 & w24683);
assign w9399 = b[35] & w1519;
assign w9400 = b[33] & ~w1676;
assign w9401 = b[34] & w1517;
assign w9402 = w1513 & w3918;
assign w9403 = ~w9399 & ~w9400;
assign w9404 = ~w9401 & w9403;
assign w9405 = ~w9402 & w9404;
assign w9406 = a[23] & ~w9405;
assign w9407 = ~a[23] & w9405;
assign w9408 = ~w9406 & ~w9407;
assign w9409 = b[31] & w1955;
assign w9410 = b[32] & w1957;
assign w9411 = b[30] & ~w2114;
assign w9412 = w1951 & w3304;
assign w9413 = ~w9409 & ~w9410;
assign w9414 = ~w9411 & w9413;
assign w9415 = ~w9412 & w9414;
assign w9416 = a[26] & ~w9415;
assign w9417 = ~a[26] & w9415;
assign w9418 = ~w9416 & ~w9417;
assign w9419 = (~w9234 & ~w9237) | (~w9234 & w24684) | (~w9237 & w24684);
assign w9420 = ~w9228 & ~w9231;
assign w9421 = b[24] & w3177;
assign w9422 = b[25] & w2973;
assign w9423 = b[26] & w2978;
assign w9424 = w2219 & w2980;
assign w9425 = ~w9422 & ~w9423;
assign w9426 = ~w9421 & w9425;
assign w9427 = ~w9424 & w9426;
assign w9428 = a[32] & ~w9427;
assign w9429 = ~a[32] & w9427;
assign w9430 = ~w9428 & ~w9429;
assign w9431 = ~w9221 & ~w9225;
assign w9432 = b[18] & w4453;
assign w9433 = b[20] & w4243;
assign w9434 = b[19] & w4241;
assign w9435 = w1347 & w4236;
assign w9436 = ~w9433 & ~w9434;
assign w9437 = ~w9432 & w9436;
assign w9438 = ~w9435 & w9437;
assign w9439 = a[38] & ~w9438;
assign w9440 = ~a[38] & w9438;
assign w9441 = ~w9439 & ~w9440;
assign w9442 = ~w9209 & ~w9213;
assign w9443 = b[15] & w5167;
assign w9444 = b[17] & w4925;
assign w9445 = b[16] & w4918;
assign w9446 = w1008 & w4923;
assign w9447 = ~w9444 & ~w9445;
assign w9448 = ~w9443 & w9447;
assign w9449 = ~w9446 & w9448;
assign w9450 = a[41] & ~w9449;
assign w9451 = ~a[41] & w9449;
assign w9452 = ~w9450 & ~w9451;
assign w9453 = b[12] & w5939;
assign w9454 = b[14] & w5665;
assign w9455 = b[13] & w5670;
assign w9456 = w714 & w5663;
assign w9457 = ~w9454 & ~w9455;
assign w9458 = ~w9453 & w9457;
assign w9459 = ~w9456 & w9458;
assign w9460 = a[44] & ~w9459;
assign w9461 = ~a[44] & w9459;
assign w9462 = ~w9460 & ~w9461;
assign w9463 = ~w9196 & ~w9199;
assign w9464 = ~w9173 & ~w9176;
assign w9465 = b[3] & w8515;
assign w9466 = b[5] & w8202;
assign w9467 = b[4] & w8200;
assign w9468 = w116 & w8195;
assign w9469 = ~w9466 & ~w9467;
assign w9470 = ~w9465 & w9469;
assign w9471 = ~w9468 & w9470;
assign w9472 = a[53] & ~w9471;
assign w9473 = ~a[53] & w9471;
assign w9474 = ~w9472 & ~w9473;
assign w9475 = a[56] & ~w8831;
assign w9476 = w9168 & w9475;
assign w9477 = a[56] & ~w9476;
assign w9478 = b[1] & w9165;
assign w9479 = b[2] & w9160;
assign w9480 = w22 & w9158;
assign w9481 = w8830 & ~w9157;
assign w9482 = w9164 & w9481;
assign w9483 = b[0] & w9482;
assign w9484 = ~w9478 & ~w9479;
assign w9485 = ~w9480 & w9484;
assign w9486 = ~w9483 & w9485;
assign w9487 = ~w9477 & w9486;
assign w9488 = w9477 & ~w9486;
assign w9489 = ~w9487 & ~w9488;
assign w9490 = w9474 & w9489;
assign w9491 = ~w9474 & ~w9489;
assign w9492 = ~w9490 & ~w9491;
assign w9493 = w9464 & w9492;
assign w9494 = ~w9464 & ~w9492;
assign w9495 = ~w9493 & ~w9494;
assign w9496 = b[6] & w7586;
assign w9497 = b[7] & w7307;
assign w9498 = b[8] & w7314;
assign w9499 = w270 & w7312;
assign w9500 = ~w9497 & ~w9498;
assign w9501 = ~w9496 & w9500;
assign w9502 = ~w9499 & w9501;
assign w9503 = a[50] & ~w9502;
assign w9504 = ~a[50] & w9502;
assign w9505 = ~w9503 & ~w9504;
assign w9506 = w9495 & ~w9505;
assign w9507 = ~w9495 & w9505;
assign w9508 = ~w9506 & ~w9507;
assign w9509 = ~w9189 & ~w9192;
assign w9510 = w9508 & w9509;
assign w9511 = ~w9508 & ~w9509;
assign w9512 = ~w9510 & ~w9511;
assign w9513 = b[9] & w6732;
assign w9514 = b[11] & w6476;
assign w9515 = b[10] & w6474;
assign w9516 = w469 & w6469;
assign w9517 = ~w9514 & ~w9515;
assign w9518 = ~w9513 & w9517;
assign w9519 = ~w9516 & w9518;
assign w9520 = a[47] & ~w9519;
assign w9521 = ~a[47] & w9519;
assign w9522 = ~w9520 & ~w9521;
assign w9523 = ~w9512 & ~w9522;
assign w9524 = w9512 & w9522;
assign w9525 = ~w9523 & ~w9524;
assign w9526 = w9463 & w9525;
assign w9527 = ~w9463 & ~w9525;
assign w9528 = ~w9526 & ~w9527;
assign w9529 = w9462 & ~w9528;
assign w9530 = ~w9462 & w9528;
assign w9531 = ~w9529 & ~w9530;
assign w9532 = (~w9202 & ~w9122) | (~w9202 & w25548) | (~w9122 & w25548);
assign w9533 = w9531 & w9532;
assign w9534 = ~w9531 & ~w9532;
assign w9535 = ~w9533 & ~w9534;
assign w9536 = ~w9452 & ~w9535;
assign w9537 = w9452 & w9535;
assign w9538 = ~w9536 & ~w9537;
assign w9539 = ~w9442 & ~w9538;
assign w9540 = w9442 & w9538;
assign w9541 = ~w9539 & ~w9540;
assign w9542 = w9441 & ~w9541;
assign w9543 = ~w9441 & w9541;
assign w9544 = ~w9542 & ~w9543;
assign w9545 = (~w9215 & ~w9101) | (~w9215 & w24685) | (~w9101 & w24685);
assign w9546 = w9544 & w9545;
assign w9547 = ~w9544 & ~w9545;
assign w9548 = ~w9546 & ~w9547;
assign w9549 = b[21] & w3785;
assign w9550 = b[22] & w3578;
assign w9551 = b[23] & w3580;
assign w9552 = w1755 & w3573;
assign w9553 = ~w9550 & ~w9551;
assign w9554 = ~w9549 & w9553;
assign w9555 = ~w9552 & w9554;
assign w9556 = a[35] & ~w9555;
assign w9557 = ~a[35] & w9555;
assign w9558 = ~w9556 & ~w9557;
assign w9559 = w9548 & w9558;
assign w9560 = ~w9548 & ~w9558;
assign w9561 = ~w9559 & ~w9560;
assign w9562 = w9431 & ~w9561;
assign w9563 = ~w9431 & w9561;
assign w9564 = ~w9562 & ~w9563;
assign w9565 = w9430 & w9564;
assign w9566 = ~w9430 & ~w9564;
assign w9567 = ~w9565 & ~w9566;
assign w9568 = ~w9420 & w9567;
assign w9569 = w9420 & ~w9567;
assign w9570 = ~w9568 & ~w9569;
assign w9571 = b[28] & w2436;
assign w9572 = b[29] & w2438;
assign w9573 = b[27] & ~w2622;
assign w9574 = w2432 & w2734;
assign w9575 = ~w9571 & ~w9572;
assign w9576 = ~w9573 & w9575;
assign w9577 = ~w9574 & w9576;
assign w9578 = a[29] & ~w9577;
assign w9579 = ~a[29] & w9577;
assign w9580 = ~w9578 & ~w9579;
assign w9581 = ~w9570 & ~w9580;
assign w9582 = w9570 & w9580;
assign w9583 = ~w9581 & ~w9582;
assign w9584 = w9419 & w9583;
assign w9585 = ~w9419 & ~w9583;
assign w9586 = ~w9584 & ~w9585;
assign w9587 = w9418 & ~w9586;
assign w9588 = ~w9418 & w9586;
assign w9589 = ~w9587 & ~w9588;
assign w9590 = (~w9251 & w9069) | (~w9251 & w25170) | (w9069 & w25170);
assign w9591 = w9589 & ~w9590;
assign w9592 = ~w9589 & w9590;
assign w9593 = ~w9591 & ~w9592;
assign w9594 = w9408 & w9593;
assign w9595 = ~w9408 & ~w9593;
assign w9596 = ~w9594 & ~w9595;
assign w9597 = ~w9398 & w9596;
assign w9598 = w9398 & ~w9596;
assign w9599 = ~w9597 & ~w9598;
assign w9600 = w9397 & w9599;
assign w9601 = ~w9397 & ~w9599;
assign w9602 = ~w9600 & ~w9601;
assign w9603 = (~w9274 & ~w9057) | (~w9274 & w25004) | (~w9057 & w25004);
assign w9604 = ~w9602 & ~w9603;
assign w9605 = w9602 & w9603;
assign w9606 = ~w9604 & ~w9605;
assign w9607 = b[39] & ~w934;
assign w9608 = b[41] & w834;
assign w9609 = b[40] & w838;
assign w9610 = w832 & w5302;
assign w9611 = ~w9607 & ~w9608;
assign w9612 = ~w9609 & w9611;
assign w9613 = ~w9610 & w9612;
assign w9614 = a[17] & ~w9613;
assign w9615 = ~a[17] & w9613;
assign w9616 = ~w9614 & ~w9615;
assign w9617 = w9606 & w9616;
assign w9618 = ~w9606 & ~w9616;
assign w9619 = ~w9617 & ~w9618;
assign w9620 = ~w9387 & ~w9619;
assign w9621 = w9387 & w9619;
assign w9622 = ~w9620 & ~w9621;
assign w9623 = ~w9386 & w9622;
assign w9624 = w9386 & ~w9622;
assign w9625 = ~w9623 & ~w9624;
assign w9626 = (~w9297 & w9046) | (~w9297 & w24391) | (w9046 & w24391);
assign w9627 = w9625 & ~w9626;
assign w9628 = ~w9625 & w9626;
assign w9629 = ~w9627 & ~w9628;
assign w9630 = w9376 & w9629;
assign w9631 = ~w9376 & ~w9629;
assign w9632 = ~w9630 & ~w9631;
assign w9633 = ~w9366 & ~w9632;
assign w9634 = w9366 & w9632;
assign w9635 = ~w9633 & ~w9634;
assign w9636 = ~w9365 & w9635;
assign w9637 = w9365 & ~w9635;
assign w9638 = ~w9636 & ~w9637;
assign w9639 = (~w9309 & ~w9025) | (~w9309 & w25171) | (~w9025 & w25171);
assign w9640 = w9638 & w9639;
assign w9641 = ~w9638 & ~w9639;
assign w9642 = ~w9640 & ~w9641;
assign w9643 = ~w9355 & ~w9642;
assign w9644 = w9355 & w9642;
assign w9645 = ~w9643 & ~w9644;
assign w9646 = w9345 & w9645;
assign w9647 = ~w9345 & ~w9645;
assign w9648 = ~w9646 & ~w9647;
assign w9649 = b[56] & w11;
assign w9650 = b[55] & w9;
assign w9651 = ~b[55] & ~b[56];
assign w9652 = b[55] & b[56];
assign w9653 = ~w9651 & ~w9652;
assign w9654 = ~w9324 & ~w9329;
assign w9655 = ~w9653 & ~w9654;
assign w9656 = w9653 & w9654;
assign w9657 = ~w9655 & ~w9656;
assign w9658 = w5 & w9657;
assign w9659 = ~w9649 & ~w9650;
assign w9660 = ~w9658 & w9659;
assign w9661 = b[54] & w24;
assign w9662 = a[2] & ~w9661;
assign w9663 = w9660 & ~w9662;
assign w9664 = a[2] & ~w9660;
assign w9665 = ~w9663 & ~w9664;
assign w9666 = ~w9648 & w9665;
assign w9667 = w9648 & ~w9665;
assign w9668 = ~w9666 & ~w9667;
assign w9669 = (~w9339 & w9014) | (~w9339 & w25291) | (w9014 & w25291);
assign w9670 = w9668 & ~w9669;
assign w9671 = ~w9668 & w9669;
assign w9672 = ~w9670 & ~w9671;
assign w9673 = (~w9666 & w9669) | (~w9666 & w25433) | (w9669 & w25433);
assign w9674 = b[52] & w103;
assign w9675 = b[54] & w68;
assign w9676 = b[53] & w61;
assign w9677 = w66 & ~w8998;
assign w9678 = ~w9675 & ~w9676;
assign w9679 = ~w9674 & w9678;
assign w9680 = ~w9677 & w9679;
assign w9681 = a[5] & ~w9680;
assign w9682 = ~a[5] & w9680;
assign w9683 = ~w9681 & ~w9682;
assign w9684 = (~w9637 & ~w9639) | (~w9637 & w25005) | (~w9639 & w25005);
assign w9685 = b[51] & w185;
assign w9686 = b[49] & ~w237;
assign w9687 = b[50] & w183;
assign w9688 = w179 & ~w8058;
assign w9689 = ~w9685 & ~w9686;
assign w9690 = ~w9687 & w9689;
assign w9691 = ~w9688 & w9690;
assign w9692 = a[8] & ~w9691;
assign w9693 = ~a[8] & w9691;
assign w9694 = ~w9692 & ~w9693;
assign w9695 = b[46] & ~w419;
assign w9696 = b[48] & w360;
assign w9697 = b[47] & w358;
assign w9698 = w354 & ~w7170;
assign w9699 = ~w9695 & ~w9696;
assign w9700 = ~w9697 & w9699;
assign w9701 = ~w9698 & w9700;
assign w9702 = a[11] & ~w9701;
assign w9703 = ~a[11] & w9701;
assign w9704 = ~w9702 & ~w9703;
assign w9705 = (~w9624 & w9626) | (~w9624 & w24846) | (w9626 & w24846);
assign w9706 = b[43] & ~w649;
assign w9707 = b[45] & w575;
assign w9708 = b[44] & w573;
assign w9709 = w569 & w6334;
assign w9710 = ~w9706 & ~w9707;
assign w9711 = ~w9708 & w9710;
assign w9712 = ~w9709 & w9711;
assign w9713 = a[14] & ~w9712;
assign w9714 = ~a[14] & w9712;
assign w9715 = ~w9713 & ~w9714;
assign w9716 = b[41] & w838;
assign w9717 = b[40] & ~w934;
assign w9718 = b[42] & w834;
assign w9719 = w832 & w5548;
assign w9720 = ~w9716 & ~w9717;
assign w9721 = ~w9718 & w9720;
assign w9722 = ~w9719 & w9721;
assign w9723 = a[17] & ~w9722;
assign w9724 = ~a[17] & w9722;
assign w9725 = ~w9723 & ~w9724;
assign w9726 = b[35] & w1517;
assign w9727 = b[34] & ~w1676;
assign w9728 = b[36] & w1519;
assign w9729 = w1513 & w4129;
assign w9730 = ~w9726 & ~w9727;
assign w9731 = ~w9728 & w9730;
assign w9732 = ~w9729 & w9731;
assign w9733 = a[23] & ~w9732;
assign w9734 = ~a[23] & w9732;
assign w9735 = ~w9733 & ~w9734;
assign w9736 = (~w9587 & w9590) | (~w9587 & w25292) | (w9590 & w25292);
assign w9737 = ~w9565 & ~w9568;
assign w9738 = b[25] & w3177;
assign w9739 = b[27] & w2978;
assign w9740 = b[26] & w2973;
assign w9741 = w2378 & w2980;
assign w9742 = ~w9739 & ~w9740;
assign w9743 = ~w9738 & w9742;
assign w9744 = ~w9741 & w9743;
assign w9745 = a[32] & ~w9744;
assign w9746 = ~a[32] & w9744;
assign w9747 = ~w9745 & ~w9746;
assign w9748 = b[22] & w3785;
assign w9749 = b[23] & w3578;
assign w9750 = b[24] & w3580;
assign w9751 = w1895 & w3573;
assign w9752 = ~w9749 & ~w9750;
assign w9753 = ~w9748 & w9752;
assign w9754 = ~w9751 & w9753;
assign w9755 = a[35] & ~w9754;
assign w9756 = ~a[35] & w9754;
assign w9757 = ~w9755 & ~w9756;
assign w9758 = ~w9542 & ~w9546;
assign w9759 = b[16] & w5167;
assign w9760 = b[17] & w4918;
assign w9761 = b[18] & w4925;
assign w9762 = ~w1108 & w4923;
assign w9763 = ~w9760 & ~w9761;
assign w9764 = ~w9759 & w9763;
assign w9765 = ~w9762 & w9764;
assign w9766 = a[41] & ~w9765;
assign w9767 = ~a[41] & w9765;
assign w9768 = ~w9766 & ~w9767;
assign w9769 = ~w9529 & ~w9533;
assign w9770 = b[13] & w5939;
assign w9771 = b[14] & w5670;
assign w9772 = b[15] & w5665;
assign w9773 = ~w799 & w5663;
assign w9774 = ~w9771 & ~w9772;
assign w9775 = ~w9770 & w9774;
assign w9776 = ~w9773 & w9775;
assign w9777 = a[44] & ~w9776;
assign w9778 = ~a[44] & w9776;
assign w9779 = ~w9777 & ~w9778;
assign w9780 = b[10] & w6732;
assign w9781 = b[12] & w6476;
assign w9782 = b[11] & w6474;
assign w9783 = w536 & w6469;
assign w9784 = ~w9781 & ~w9782;
assign w9785 = ~w9780 & w9784;
assign w9786 = ~w9783 & w9785;
assign w9787 = a[47] & ~w9786;
assign w9788 = ~a[47] & w9786;
assign w9789 = ~w9787 & ~w9788;
assign w9790 = ~w9507 & ~w9510;
assign w9791 = b[7] & w7586;
assign w9792 = b[8] & w7307;
assign w9793 = b[9] & w7314;
assign w9794 = w322 & w7312;
assign w9795 = ~w9792 & ~w9793;
assign w9796 = ~w9791 & w9795;
assign w9797 = ~w9794 & w9796;
assign w9798 = a[50] & ~w9797;
assign w9799 = ~a[50] & w9797;
assign w9800 = ~w9798 & ~w9799;
assign w9801 = b[1] & w9482;
assign w9802 = b[2] & w9165;
assign w9803 = b[3] & w9160;
assign w9804 = w46 & w9158;
assign w9805 = ~w9802 & ~w9803;
assign w9806 = ~w9801 & w9805;
assign w9807 = ~w9804 & w9806;
assign w9808 = a[56] & ~w9807;
assign w9809 = ~a[56] & w9807;
assign w9810 = ~w9808 & ~w9809;
assign w9811 = w9476 & w9486;
assign w9812 = a[56] & ~a[57];
assign w9813 = ~a[56] & a[57];
assign w9814 = ~w9812 & ~w9813;
assign w9815 = b[0] & ~w9814;
assign w9816 = w9811 & w9815;
assign w9817 = ~w9811 & ~w9815;
assign w9818 = ~w9816 & ~w9817;
assign w9819 = w9810 & w9818;
assign w9820 = ~w9810 & ~w9818;
assign w9821 = ~w9819 & ~w9820;
assign w9822 = b[4] & w8515;
assign w9823 = b[5] & w8200;
assign w9824 = b[6] & w8202;
assign w9825 = w157 & w8195;
assign w9826 = ~w9823 & ~w9824;
assign w9827 = ~w9822 & w9826;
assign w9828 = ~w9825 & w9827;
assign w9829 = a[53] & ~w9828;
assign w9830 = ~a[53] & w9828;
assign w9831 = ~w9829 & ~w9830;
assign w9832 = w9821 & w9831;
assign w9833 = ~w9821 & ~w9831;
assign w9834 = ~w9832 & ~w9833;
assign w9835 = ~w9491 & ~w9493;
assign w9836 = w9834 & w9835;
assign w9837 = ~w9834 & ~w9835;
assign w9838 = ~w9836 & ~w9837;
assign w9839 = w9800 & w9838;
assign w9840 = ~w9800 & ~w9838;
assign w9841 = ~w9839 & ~w9840;
assign w9842 = w9790 & ~w9841;
assign w9843 = ~w9790 & w9841;
assign w9844 = ~w9842 & ~w9843;
assign w9845 = ~w9789 & ~w9844;
assign w9846 = w9789 & w9844;
assign w9847 = ~w9845 & ~w9846;
assign w9848 = ~w9523 & ~w9526;
assign w9849 = w9847 & w9848;
assign w9850 = ~w9847 & ~w9848;
assign w9851 = ~w9849 & ~w9850;
assign w9852 = w9779 & w9851;
assign w9853 = ~w9779 & ~w9851;
assign w9854 = ~w9852 & ~w9853;
assign w9855 = w9769 & ~w9854;
assign w9856 = ~w9769 & w9854;
assign w9857 = ~w9855 & ~w9856;
assign w9858 = ~w9768 & ~w9857;
assign w9859 = w9768 & w9857;
assign w9860 = ~w9858 & ~w9859;
assign w9861 = (~w9536 & ~w9442) | (~w9536 & w25549) | (~w9442 & w25549);
assign w9862 = w9860 & w9861;
assign w9863 = ~w9860 & ~w9861;
assign w9864 = ~w9862 & ~w9863;
assign w9865 = b[19] & w4453;
assign w9866 = b[21] & w4243;
assign w9867 = b[20] & w4241;
assign w9868 = w1467 & w4236;
assign w9869 = ~w9866 & ~w9867;
assign w9870 = ~w9865 & w9869;
assign w9871 = ~w9868 & w9870;
assign w9872 = a[38] & ~w9871;
assign w9873 = ~a[38] & w9871;
assign w9874 = ~w9872 & ~w9873;
assign w9875 = w9864 & w9874;
assign w9876 = ~w9864 & ~w9874;
assign w9877 = ~w9875 & ~w9876;
assign w9878 = w9758 & w9877;
assign w9879 = ~w9758 & ~w9877;
assign w9880 = ~w9878 & ~w9879;
assign w9881 = ~w9757 & w9880;
assign w9882 = w9757 & ~w9880;
assign w9883 = ~w9881 & ~w9882;
assign w9884 = (~w9559 & w9431) | (~w9559 & w25434) | (w9431 & w25434);
assign w9885 = w9883 & ~w9884;
assign w9886 = ~w9883 & w9884;
assign w9887 = ~w9885 & ~w9886;
assign w9888 = w9747 & w9887;
assign w9889 = ~w9747 & ~w9887;
assign w9890 = ~w9888 & ~w9889;
assign w9891 = ~w9737 & w9890;
assign w9892 = w9737 & ~w9890;
assign w9893 = ~w9891 & ~w9892;
assign w9894 = b[28] & ~w2622;
assign w9895 = b[29] & w2436;
assign w9896 = b[30] & w2438;
assign w9897 = w2432 & ~w2908;
assign w9898 = ~w9894 & ~w9895;
assign w9899 = ~w9896 & w9898;
assign w9900 = ~w9897 & w9899;
assign w9901 = a[29] & ~w9900;
assign w9902 = ~a[29] & w9900;
assign w9903 = ~w9901 & ~w9902;
assign w9904 = w9893 & w9903;
assign w9905 = ~w9893 & ~w9903;
assign w9906 = ~w9904 & ~w9905;
assign w9907 = ~w9581 & ~w9584;
assign w9908 = w9906 & w9907;
assign w9909 = ~w9906 & ~w9907;
assign w9910 = ~w9908 & ~w9909;
assign w9911 = b[32] & w1955;
assign w9912 = b[31] & ~w2114;
assign w9913 = b[33] & w1957;
assign w9914 = w1951 & w3499;
assign w9915 = ~w9911 & ~w9912;
assign w9916 = ~w9913 & w9915;
assign w9917 = ~w9914 & w9916;
assign w9918 = a[26] & ~w9917;
assign w9919 = ~a[26] & w9917;
assign w9920 = ~w9918 & ~w9919;
assign w9921 = w9910 & w9920;
assign w9922 = ~w9910 & ~w9920;
assign w9923 = ~w9921 & ~w9922;
assign w9924 = ~w9736 & ~w9923;
assign w9925 = w9736 & w9923;
assign w9926 = ~w9924 & ~w9925;
assign w9927 = ~w9735 & w9926;
assign w9928 = w9735 & ~w9926;
assign w9929 = ~w9927 & ~w9928;
assign w9930 = (~w9594 & w9398) | (~w9594 & w25172) | (w9398 & w25172);
assign w9931 = ~w9929 & w9930;
assign w9932 = w9929 & ~w9930;
assign w9933 = ~w9931 & ~w9932;
assign w9934 = b[37] & ~w1272;
assign w9935 = b[38] & w1154;
assign w9936 = b[39] & w1156;
assign w9937 = w1150 & ~w4812;
assign w9938 = ~w9934 & ~w9935;
assign w9939 = ~w9936 & w9938;
assign w9940 = ~w9937 & w9939;
assign w9941 = a[20] & ~w9940;
assign w9942 = ~a[20] & w9940;
assign w9943 = ~w9941 & ~w9942;
assign w9944 = w9933 & w9943;
assign w9945 = ~w9933 & ~w9943;
assign w9946 = ~w9944 & ~w9945;
assign w9947 = (~w9600 & ~w9603) | (~w9600 & w24686) | (~w9603 & w24686);
assign w9948 = w9946 & w9947;
assign w9949 = ~w9946 & ~w9947;
assign w9950 = ~w9948 & ~w9949;
assign w9951 = ~w9725 & w9950;
assign w9952 = w9725 & ~w9950;
assign w9953 = ~w9951 & ~w9952;
assign w9954 = (~w9618 & ~w9387) | (~w9618 & w25006) | (~w9387 & w25006);
assign w9955 = w9953 & w9954;
assign w9956 = ~w9953 & ~w9954;
assign w9957 = ~w9955 & ~w9956;
assign w9958 = ~w9715 & ~w9957;
assign w9959 = w9715 & w9957;
assign w9960 = ~w9958 & ~w9959;
assign w9961 = ~w9705 & w9960;
assign w9962 = w9705 & ~w9960;
assign w9963 = ~w9961 & ~w9962;
assign w9964 = ~w9704 & ~w9963;
assign w9965 = w9704 & w9963;
assign w9966 = ~w9964 & ~w9965;
assign w9967 = (~w9631 & ~w9366) | (~w9631 & w24392) | (~w9366 & w24392);
assign w9968 = w9966 & w9967;
assign w9969 = ~w9966 & ~w9967;
assign w9970 = ~w9968 & ~w9969;
assign w9971 = ~w9694 & ~w9970;
assign w9972 = w9694 & w9970;
assign w9973 = ~w9971 & ~w9972;
assign w9974 = ~w9684 & ~w9973;
assign w9975 = w9684 & w9973;
assign w9976 = ~w9974 & ~w9975;
assign w9977 = ~w9683 & w9976;
assign w9978 = w9683 & ~w9976;
assign w9979 = ~w9977 & ~w9978;
assign w9980 = (~w9643 & ~w9345) | (~w9643 & w25173) | (~w9345 & w25173);
assign w9981 = w9979 & w9980;
assign w9982 = ~w9979 & ~w9980;
assign w9983 = ~w9981 & ~w9982;
assign w9984 = b[57] & w11;
assign w9985 = b[56] & w9;
assign w9986 = ~w9652 & ~w9656;
assign w9987 = ~b[56] & ~b[57];
assign w9988 = b[56] & b[57];
assign w9989 = ~w9987 & ~w9988;
assign w9990 = ~w9986 & ~w9989;
assign w9991 = w9986 & w9989;
assign w9992 = ~w9990 & ~w9991;
assign w9993 = w5 & ~w9992;
assign w9994 = ~w9984 & ~w9985;
assign w9995 = ~w9993 & w9994;
assign w9996 = b[55] & w24;
assign w9997 = a[2] & ~w9996;
assign w9998 = w9995 & ~w9997;
assign w9999 = a[2] & ~w9995;
assign w10000 = ~w9998 & ~w9999;
assign w10001 = w9983 & w10000;
assign w10002 = ~w9983 & ~w10000;
assign w10003 = ~w10001 & ~w10002;
assign w10004 = ~w9673 & w10003;
assign w10005 = w9673 & ~w10003;
assign w10006 = ~w10004 & ~w10005;
assign w10007 = (~w9978 & ~w9980) | (~w9978 & w25007) | (~w9980 & w25007);
assign w10008 = b[53] & w103;
assign w10009 = b[55] & w68;
assign w10010 = b[54] & w61;
assign w10011 = w66 & ~w9330;
assign w10012 = ~w10009 & ~w10010;
assign w10013 = ~w10008 & w10012;
assign w10014 = ~w10011 & w10013;
assign w10015 = a[5] & ~w10014;
assign w10016 = ~a[5] & w10014;
assign w10017 = ~w10015 & ~w10016;
assign w10018 = b[50] & ~w237;
assign w10019 = b[51] & w183;
assign w10020 = b[52] & w185;
assign w10021 = w179 & ~w8371;
assign w10022 = ~w10018 & ~w10019;
assign w10023 = ~w10020 & w10022;
assign w10024 = ~w10021 & w10023;
assign w10025 = a[8] & ~w10024;
assign w10026 = ~a[8] & w10024;
assign w10027 = ~w10025 & ~w10026;
assign w10028 = (~w9965 & ~w9967) | (~w9965 & w24847) | (~w9967 & w24847);
assign w10029 = b[47] & ~w419;
assign w10030 = b[48] & w358;
assign w10031 = b[49] & w360;
assign w10032 = w354 & ~w7468;
assign w10033 = ~w10029 & ~w10030;
assign w10034 = ~w10031 & w10033;
assign w10035 = ~w10032 & w10034;
assign w10036 = a[11] & ~w10035;
assign w10037 = ~a[11] & w10035;
assign w10038 = ~w10036 & ~w10037;
assign w10039 = (~w9959 & w9705) | (~w9959 & w25008) | (w9705 & w25008);
assign w10040 = b[44] & ~w649;
assign w10041 = b[46] & w575;
assign w10042 = b[45] & w573;
assign w10043 = w569 & ~w6613;
assign w10044 = ~w10040 & ~w10041;
assign w10045 = ~w10042 & w10044;
assign w10046 = ~w10043 & w10045;
assign w10047 = a[14] & ~w10046;
assign w10048 = ~a[14] & w10046;
assign w10049 = ~w10047 & ~w10048;
assign w10050 = (~w9952 & ~w9954) | (~w9952 & w24687) | (~w9954 & w24687);
assign w10051 = b[39] & w1154;
assign w10052 = b[40] & w1156;
assign w10053 = b[38] & ~w1272;
assign w10054 = w1150 & ~w5058;
assign w10055 = ~w10051 & ~w10052;
assign w10056 = ~w10053 & w10055;
assign w10057 = ~w10054 & w10056;
assign w10058 = a[20] & ~w10057;
assign w10059 = ~a[20] & w10057;
assign w10060 = ~w10058 & ~w10059;
assign w10061 = (~w9928 & w9930) | (~w9928 & w25293) | (w9930 & w25293);
assign w10062 = b[35] & ~w1676;
assign w10063 = b[36] & w1517;
assign w10064 = b[37] & w1519;
assign w10065 = w1513 & ~w4357;
assign w10066 = ~w10062 & ~w10063;
assign w10067 = ~w10064 & w10066;
assign w10068 = ~w10065 & w10067;
assign w10069 = a[23] & ~w10068;
assign w10070 = ~a[23] & w10068;
assign w10071 = ~w10069 & ~w10070;
assign w10072 = b[32] & ~w2114;
assign w10073 = b[34] & w1957;
assign w10074 = b[33] & w1955;
assign w10075 = w1951 & ~w3710;
assign w10076 = ~w10072 & ~w10073;
assign w10077 = ~w10074 & w10076;
assign w10078 = ~w10075 & w10077;
assign w10079 = a[26] & ~w10078;
assign w10080 = ~a[26] & w10078;
assign w10081 = ~w10079 & ~w10080;
assign w10082 = ~w9904 & ~w9908;
assign w10083 = b[30] & w2436;
assign w10084 = b[31] & w2438;
assign w10085 = b[29] & ~w2622;
assign w10086 = w2432 & ~w3112;
assign w10087 = ~w10083 & ~w10084;
assign w10088 = ~w10085 & w10087;
assign w10089 = ~w10086 & w10088;
assign w10090 = a[29] & ~w10089;
assign w10091 = ~a[29] & w10089;
assign w10092 = ~w10090 & ~w10091;
assign w10093 = (~w9888 & w9737) | (~w9888 & w25435) | (w9737 & w25435);
assign w10094 = b[26] & w3177;
assign w10095 = b[28] & w2978;
assign w10096 = b[27] & w2973;
assign w10097 = w2559 & w2980;
assign w10098 = ~w10095 & ~w10096;
assign w10099 = ~w10094 & w10098;
assign w10100 = ~w10097 & w10099;
assign w10101 = a[32] & ~w10100;
assign w10102 = ~a[32] & w10100;
assign w10103 = ~w10101 & ~w10102;
assign w10104 = ~w9882 & ~w9885;
assign w10105 = b[20] & w4453;
assign w10106 = b[22] & w4243;
assign w10107 = b[21] & w4241;
assign w10108 = w1615 & w4236;
assign w10109 = ~w10106 & ~w10107;
assign w10110 = ~w10105 & w10109;
assign w10111 = ~w10108 & w10110;
assign w10112 = a[38] & ~w10111;
assign w10113 = ~a[38] & w10111;
assign w10114 = ~w10112 & ~w10113;
assign w10115 = b[14] & w5939;
assign w10116 = b[16] & w5665;
assign w10117 = b[15] & w5670;
assign w10118 = w905 & w5663;
assign w10119 = ~w10116 & ~w10117;
assign w10120 = ~w10115 & w10119;
assign w10121 = ~w10118 & w10120;
assign w10122 = a[44] & ~w10121;
assign w10123 = ~a[44] & w10121;
assign w10124 = ~w10122 & ~w10123;
assign w10125 = ~w9832 & ~w9836;
assign w10126 = ~w9816 & ~w9819;
assign w10127 = b[2] & w9482;
assign w10128 = b[3] & w9165;
assign w10129 = b[4] & w9160;
assign w10130 = w84 & w9158;
assign w10131 = ~w10128 & ~w10129;
assign w10132 = ~w10127 & w10131;
assign w10133 = ~w10130 & w10132;
assign w10134 = a[56] & ~w10133;
assign w10135 = ~a[56] & w10133;
assign w10136 = ~w10134 & ~w10135;
assign w10137 = a[59] & w9815;
assign w10138 = a[58] & ~a[59];
assign w10139 = ~a[58] & a[59];
assign w10140 = ~w10138 & ~w10139;
assign w10141 = ~w9814 & ~w10140;
assign w10142 = ~w8 & w10141;
assign w10143 = a[57] & ~a[58];
assign w10144 = ~a[57] & a[58];
assign w10145 = ~w10143 & ~w10144;
assign w10146 = w9814 & ~w10145;
assign w10147 = b[0] & w10146;
assign w10148 = ~w9814 & w10140;
assign w10149 = b[1] & w10148;
assign w10150 = ~w10142 & ~w10147;
assign w10151 = ~w10149 & w10150;
assign w10152 = ~w10137 & w10151;
assign w10153 = w10137 & ~w10151;
assign w10154 = ~w10152 & ~w10153;
assign w10155 = ~w10136 & ~w10154;
assign w10156 = w10136 & w10154;
assign w10157 = ~w10155 & ~w10156;
assign w10158 = ~w10126 & w10157;
assign w10159 = w10126 & ~w10157;
assign w10160 = ~w10158 & ~w10159;
assign w10161 = b[5] & w8515;
assign w10162 = b[7] & w8202;
assign w10163 = b[6] & w8200;
assign w10164 = w216 & w8195;
assign w10165 = ~w10162 & ~w10163;
assign w10166 = ~w10161 & w10165;
assign w10167 = ~w10164 & w10166;
assign w10168 = a[53] & ~w10167;
assign w10169 = ~a[53] & w10167;
assign w10170 = ~w10168 & ~w10169;
assign w10171 = ~w10160 & ~w10170;
assign w10172 = w10160 & w10170;
assign w10173 = ~w10171 & ~w10172;
assign w10174 = w10125 & ~w10173;
assign w10175 = ~w10125 & w10173;
assign w10176 = ~w10174 & ~w10175;
assign w10177 = b[8] & w7586;
assign w10178 = b[9] & w7307;
assign w10179 = b[10] & w7314;
assign w10180 = w397 & w7312;
assign w10181 = ~w10178 & ~w10179;
assign w10182 = ~w10177 & w10181;
assign w10183 = ~w10180 & w10182;
assign w10184 = a[50] & ~w10183;
assign w10185 = ~a[50] & w10183;
assign w10186 = ~w10184 & ~w10185;
assign w10187 = w10176 & w10186;
assign w10188 = ~w10176 & ~w10186;
assign w10189 = ~w10187 & ~w10188;
assign w10190 = ~w9839 & ~w9843;
assign w10191 = ~w10189 & w10190;
assign w10192 = w10189 & ~w10190;
assign w10193 = ~w10191 & ~w10192;
assign w10194 = b[11] & w6732;
assign w10195 = b[12] & w6474;
assign w10196 = b[13] & w6476;
assign w10197 = w628 & w6469;
assign w10198 = ~w10195 & ~w10196;
assign w10199 = ~w10194 & w10198;
assign w10200 = ~w10197 & w10199;
assign w10201 = a[47] & ~w10200;
assign w10202 = ~a[47] & w10200;
assign w10203 = ~w10201 & ~w10202;
assign w10204 = w10193 & w10203;
assign w10205 = ~w10193 & ~w10203;
assign w10206 = ~w10204 & ~w10205;
assign w10207 = ~w9846 & ~w9849;
assign w10208 = w10206 & w10207;
assign w10209 = ~w10206 & ~w10207;
assign w10210 = ~w10208 & ~w10209;
assign w10211 = w10124 & ~w10210;
assign w10212 = ~w10124 & w10210;
assign w10213 = ~w10211 & ~w10212;
assign w10214 = ~w9852 & ~w9856;
assign w10215 = ~w10213 & w10214;
assign w10216 = w10213 & ~w10214;
assign w10217 = ~w10215 & ~w10216;
assign w10218 = b[17] & w5167;
assign w10219 = b[18] & w4918;
assign w10220 = b[19] & w4925;
assign w10221 = ~w1231 & w4923;
assign w10222 = ~w10219 & ~w10220;
assign w10223 = ~w10218 & w10222;
assign w10224 = ~w10221 & w10223;
assign w10225 = a[41] & ~w10224;
assign w10226 = ~a[41] & w10224;
assign w10227 = ~w10225 & ~w10226;
assign w10228 = w10217 & w10227;
assign w10229 = ~w10217 & ~w10227;
assign w10230 = ~w10228 & ~w10229;
assign w10231 = ~w9859 & ~w9862;
assign w10232 = ~w10230 & w10231;
assign w10233 = w10230 & ~w10231;
assign w10234 = ~w10232 & ~w10233;
assign w10235 = w10114 & w10234;
assign w10236 = ~w10114 & ~w10234;
assign w10237 = ~w10235 & ~w10236;
assign w10238 = (~w9876 & ~w9758) | (~w9876 & w25550) | (~w9758 & w25550);
assign w10239 = ~w10237 & ~w10238;
assign w10240 = w10237 & w10238;
assign w10241 = ~w10239 & ~w10240;
assign w10242 = b[23] & w3785;
assign w10243 = b[25] & w3580;
assign w10244 = b[24] & w3578;
assign w10245 = w2061 & w3573;
assign w10246 = ~w10243 & ~w10244;
assign w10247 = ~w10242 & w10246;
assign w10248 = ~w10245 & w10247;
assign w10249 = a[35] & ~w10248;
assign w10250 = ~a[35] & w10248;
assign w10251 = ~w10249 & ~w10250;
assign w10252 = w10241 & w10251;
assign w10253 = ~w10241 & ~w10251;
assign w10254 = ~w10252 & ~w10253;
assign w10255 = w10104 & ~w10254;
assign w10256 = ~w10104 & w10254;
assign w10257 = ~w10255 & ~w10256;
assign w10258 = w10103 & w10257;
assign w10259 = ~w10103 & ~w10257;
assign w10260 = ~w10258 & ~w10259;
assign w10261 = ~w10093 & w10260;
assign w10262 = w10093 & ~w10260;
assign w10263 = ~w10261 & ~w10262;
assign w10264 = w10092 & w10263;
assign w10265 = ~w10092 & ~w10263;
assign w10266 = ~w10264 & ~w10265;
assign w10267 = ~w10082 & ~w10266;
assign w10268 = w10082 & w10266;
assign w10269 = ~w10267 & ~w10268;
assign w10270 = ~w10081 & w10269;
assign w10271 = w10081 & ~w10269;
assign w10272 = ~w10270 & ~w10271;
assign w10273 = ~w9922 & ~w9925;
assign w10274 = w10272 & w10273;
assign w10275 = ~w10272 & ~w10273;
assign w10276 = ~w10274 & ~w10275;
assign w10277 = w10071 & w10276;
assign w10278 = ~w10071 & ~w10276;
assign w10279 = ~w10277 & ~w10278;
assign w10280 = ~w10061 & w10279;
assign w10281 = w10061 & ~w10279;
assign w10282 = ~w10280 & ~w10281;
assign w10283 = w10060 & w10282;
assign w10284 = ~w10060 & ~w10282;
assign w10285 = ~w10283 & ~w10284;
assign w10286 = (~w9945 & ~w9947) | (~w9945 & w25174) | (~w9947 & w25174);
assign w10287 = ~w10285 & ~w10286;
assign w10288 = w10285 & w10286;
assign w10289 = ~w10287 & ~w10288;
assign w10290 = b[41] & ~w934;
assign w10291 = b[43] & w834;
assign w10292 = b[42] & w838;
assign w10293 = w832 & w5811;
assign w10294 = ~w10290 & ~w10291;
assign w10295 = ~w10292 & w10294;
assign w10296 = ~w10293 & w10295;
assign w10297 = a[17] & ~w10296;
assign w10298 = ~a[17] & w10296;
assign w10299 = ~w10297 & ~w10298;
assign w10300 = ~w10289 & ~w10299;
assign w10301 = w10289 & w10299;
assign w10302 = ~w10300 & ~w10301;
assign w10303 = w10050 & w10302;
assign w10304 = ~w10050 & ~w10302;
assign w10305 = ~w10303 & ~w10304;
assign w10306 = ~w10049 & w10305;
assign w10307 = w10049 & ~w10305;
assign w10308 = ~w10306 & ~w10307;
assign w10309 = ~w10039 & w10308;
assign w10310 = w10039 & ~w10308;
assign w10311 = ~w10309 & ~w10310;
assign w10312 = w10038 & w10311;
assign w10313 = ~w10038 & ~w10311;
assign w10314 = ~w10312 & ~w10313;
assign w10315 = w10028 & ~w10314;
assign w10316 = ~w10028 & w10314;
assign w10317 = ~w10315 & ~w10316;
assign w10318 = ~w10027 & ~w10317;
assign w10319 = w10027 & w10317;
assign w10320 = ~w10318 & ~w10319;
assign w10321 = (~w9971 & ~w9684) | (~w9971 & w24393) | (~w9684 & w24393);
assign w10322 = w10320 & w10321;
assign w10323 = ~w10320 & ~w10321;
assign w10324 = ~w10322 & ~w10323;
assign w10325 = ~w10017 & ~w10324;
assign w10326 = w10017 & w10324;
assign w10327 = ~w10325 & ~w10326;
assign w10328 = w10007 & w10327;
assign w10329 = ~w10007 & ~w10327;
assign w10330 = ~w10328 & ~w10329;
assign w10331 = b[58] & w11;
assign w10332 = b[57] & w9;
assign w10333 = ~b[57] & ~b[58];
assign w10334 = b[57] & b[58];
assign w10335 = ~w10333 & ~w10334;
assign w10336 = ~w9987 & ~w9991;
assign w10337 = ~w10335 & w10336;
assign w10338 = w10335 & ~w10336;
assign w10339 = ~w10337 & ~w10338;
assign w10340 = w5 & ~w10339;
assign w10341 = ~w10331 & ~w10332;
assign w10342 = ~w10340 & w10341;
assign w10343 = b[56] & w24;
assign w10344 = a[2] & ~w10343;
assign w10345 = w10342 & ~w10344;
assign w10346 = a[2] & ~w10342;
assign w10347 = ~w10345 & ~w10346;
assign w10348 = w10330 & ~w10347;
assign w10349 = ~w10330 & w10347;
assign w10350 = ~w10348 & ~w10349;
assign w10351 = (~w10001 & w9673) | (~w10001 & w25175) | (w9673 & w25175);
assign w10352 = w10350 & w10351;
assign w10353 = ~w10350 & ~w10351;
assign w10354 = ~w10352 & ~w10353;
assign w10355 = b[54] & w103;
assign w10356 = b[56] & w68;
assign w10357 = b[55] & w61;
assign w10358 = w66 & w9657;
assign w10359 = ~w10356 & ~w10357;
assign w10360 = ~w10355 & w10359;
assign w10361 = ~w10358 & w10360;
assign w10362 = a[5] & ~w10361;
assign w10363 = ~a[5] & w10361;
assign w10364 = ~w10362 & ~w10363;
assign w10365 = ~b[58] & ~b[59];
assign w10366 = b[58] & b[59];
assign w10367 = ~w10365 & ~w10366;
assign w10368 = ~w10333 & ~w10338;
assign w10369 = w10367 & w10368;
assign w10370 = ~w10367 & ~w10368;
assign w10371 = ~w10369 & ~w10370;
assign w10372 = w117 & w10371;
assign w10373 = b[59] & w11;
assign w10374 = b[58] & w9;
assign w10375 = ~w10373 & ~w10374;
assign w10376 = ~a[2] & ~w10375;
assign w10377 = ~a[2] & ~w10371;
assign w10378 = ~a[2] & ~w5;
assign w10379 = b[57] & w25;
assign w10380 = ~w10378 & ~w10379;
assign w10381 = w10375 & w10380;
assign w10382 = ~w10377 & w10381;
assign w10383 = ~w10376 & ~w10382;
assign w10384 = ~w10372 & ~w10383;
assign w10385 = w10364 & w10384;
assign w10386 = ~w10364 & ~w10384;
assign w10387 = ~w10385 & ~w10386;
assign w10388 = b[53] & w185;
assign w10389 = b[51] & ~w237;
assign w10390 = b[52] & w183;
assign w10391 = w179 & w8683;
assign w10392 = ~w10388 & ~w10389;
assign w10393 = ~w10390 & w10392;
assign w10394 = ~w10391 & w10393;
assign w10395 = a[8] & ~w10394;
assign w10396 = ~a[8] & w10394;
assign w10397 = ~w10395 & ~w10396;
assign w10398 = b[48] & ~w419;
assign w10399 = b[50] & w360;
assign w10400 = b[49] & w358;
assign w10401 = w354 & w7759;
assign w10402 = ~w10398 & ~w10399;
assign w10403 = ~w10400 & w10402;
assign w10404 = ~w10401 & w10403;
assign w10405 = a[11] & ~w10404;
assign w10406 = ~a[11] & w10404;
assign w10407 = ~w10405 & ~w10406;
assign w10408 = (~w10307 & w10039) | (~w10307 & w24688) | (w10039 & w24688);
assign w10409 = b[45] & ~w649;
assign w10410 = b[47] & w575;
assign w10411 = b[46] & w573;
assign w10412 = w569 & w6889;
assign w10413 = ~w10409 & ~w10410;
assign w10414 = ~w10411 & w10413;
assign w10415 = ~w10412 & w10414;
assign w10416 = a[14] & ~w10415;
assign w10417 = ~a[14] & w10415;
assign w10418 = ~w10416 & ~w10417;
assign w10419 = (~w10300 & ~w10050) | (~w10300 & w25176) | (~w10050 & w25176);
assign w10420 = b[44] & w834;
assign w10421 = b[42] & ~w934;
assign w10422 = b[43] & w838;
assign w10423 = w832 & w6069;
assign w10424 = ~w10420 & ~w10421;
assign w10425 = ~w10422 & w10424;
assign w10426 = ~w10423 & w10425;
assign w10427 = a[17] & ~w10426;
assign w10428 = ~a[17] & w10426;
assign w10429 = ~w10427 & ~w10428;
assign w10430 = (~w10283 & ~w10286) | (~w10283 & w25294) | (~w10286 & w25294);
assign w10431 = ~w10277 & ~w10280;
assign w10432 = b[36] & ~w1676;
assign w10433 = b[38] & w1519;
assign w10434 = b[37] & w1517;
assign w10435 = w1513 & w4582;
assign w10436 = ~w10432 & ~w10433;
assign w10437 = ~w10434 & w10436;
assign w10438 = ~w10435 & w10437;
assign w10439 = a[23] & ~w10438;
assign w10440 = ~a[23] & w10438;
assign w10441 = ~w10439 & ~w10440;
assign w10442 = ~w10271 & ~w10274;
assign w10443 = b[31] & w2436;
assign w10444 = b[32] & w2438;
assign w10445 = b[30] & ~w2622;
assign w10446 = w2432 & w3304;
assign w10447 = ~w10443 & ~w10444;
assign w10448 = ~w10445 & w10447;
assign w10449 = ~w10446 & w10448;
assign w10450 = a[29] & ~w10449;
assign w10451 = ~a[29] & w10449;
assign w10452 = ~w10450 & ~w10451;
assign w10453 = ~w10258 & ~w10261;
assign w10454 = b[24] & w3785;
assign w10455 = b[25] & w3578;
assign w10456 = b[26] & w3580;
assign w10457 = w2219 & w3573;
assign w10458 = ~w10455 & ~w10456;
assign w10459 = ~w10454 & w10458;
assign w10460 = ~w10457 & w10459;
assign w10461 = a[35] & ~w10460;
assign w10462 = ~a[35] & w10460;
assign w10463 = ~w10461 & ~w10462;
assign w10464 = ~w10235 & ~w10240;
assign w10465 = b[21] & w4453;
assign w10466 = b[22] & w4241;
assign w10467 = b[23] & w4243;
assign w10468 = w1755 & w4236;
assign w10469 = ~w10466 & ~w10467;
assign w10470 = ~w10465 & w10469;
assign w10471 = ~w10468 & w10470;
assign w10472 = a[38] & ~w10471;
assign w10473 = ~a[38] & w10471;
assign w10474 = ~w10472 & ~w10473;
assign w10475 = ~w10211 & ~w10216;
assign w10476 = ~w10187 & ~w10192;
assign w10477 = ~w10172 & ~w10175;
assign w10478 = ~w10156 & ~w10158;
assign w10479 = b[3] & w9482;
assign w10480 = b[4] & w9165;
assign w10481 = b[5] & w9160;
assign w10482 = w116 & w9158;
assign w10483 = ~w10480 & ~w10481;
assign w10484 = ~w10479 & w10483;
assign w10485 = ~w10482 & w10484;
assign w10486 = a[56] & ~w10485;
assign w10487 = ~a[56] & w10485;
assign w10488 = ~w10486 & ~w10487;
assign w10489 = a[59] & ~w9815;
assign w10490 = w10151 & w10489;
assign w10491 = a[59] & ~w10490;
assign w10492 = b[1] & w10146;
assign w10493 = b[2] & w10148;
assign w10494 = w22 & w10141;
assign w10495 = w9814 & ~w10140;
assign w10496 = w10145 & w10495;
assign w10497 = b[0] & w10496;
assign w10498 = ~w10492 & ~w10493;
assign w10499 = ~w10494 & w10498;
assign w10500 = ~w10497 & w10499;
assign w10501 = ~w10491 & w10500;
assign w10502 = w10491 & ~w10500;
assign w10503 = ~w10501 & ~w10502;
assign w10504 = w10488 & w10503;
assign w10505 = ~w10488 & ~w10503;
assign w10506 = ~w10504 & ~w10505;
assign w10507 = w10478 & w10506;
assign w10508 = ~w10478 & ~w10506;
assign w10509 = ~w10507 & ~w10508;
assign w10510 = b[6] & w8515;
assign w10511 = b[7] & w8200;
assign w10512 = b[8] & w8202;
assign w10513 = w270 & w8195;
assign w10514 = ~w10511 & ~w10512;
assign w10515 = ~w10510 & w10514;
assign w10516 = ~w10513 & w10515;
assign w10517 = a[53] & ~w10516;
assign w10518 = ~a[53] & w10516;
assign w10519 = ~w10517 & ~w10518;
assign w10520 = w10509 & ~w10519;
assign w10521 = ~w10509 & w10519;
assign w10522 = ~w10520 & ~w10521;
assign w10523 = ~w10477 & w10522;
assign w10524 = w10477 & ~w10522;
assign w10525 = ~w10523 & ~w10524;
assign w10526 = b[9] & w7586;
assign w10527 = b[10] & w7307;
assign w10528 = b[11] & w7314;
assign w10529 = w469 & w7312;
assign w10530 = ~w10527 & ~w10528;
assign w10531 = ~w10526 & w10530;
assign w10532 = ~w10529 & w10531;
assign w10533 = a[50] & ~w10532;
assign w10534 = ~a[50] & w10532;
assign w10535 = ~w10533 & ~w10534;
assign w10536 = ~w10525 & ~w10535;
assign w10537 = w10525 & w10535;
assign w10538 = ~w10536 & ~w10537;
assign w10539 = w10476 & ~w10538;
assign w10540 = ~w10476 & w10538;
assign w10541 = ~w10539 & ~w10540;
assign w10542 = b[12] & w6732;
assign w10543 = b[13] & w6474;
assign w10544 = b[14] & w6476;
assign w10545 = w714 & w6469;
assign w10546 = ~w10543 & ~w10544;
assign w10547 = ~w10542 & w10546;
assign w10548 = ~w10545 & w10547;
assign w10549 = a[47] & ~w10548;
assign w10550 = ~a[47] & w10548;
assign w10551 = ~w10549 & ~w10550;
assign w10552 = w10541 & w10551;
assign w10553 = ~w10541 & ~w10551;
assign w10554 = ~w10552 & ~w10553;
assign w10555 = ~w10205 & ~w10208;
assign w10556 = w10554 & w10555;
assign w10557 = ~w10554 & ~w10555;
assign w10558 = ~w10556 & ~w10557;
assign w10559 = b[15] & w5939;
assign w10560 = b[17] & w5665;
assign w10561 = b[16] & w5670;
assign w10562 = w1008 & w5663;
assign w10563 = ~w10560 & ~w10561;
assign w10564 = ~w10559 & w10563;
assign w10565 = ~w10562 & w10564;
assign w10566 = a[44] & ~w10565;
assign w10567 = ~a[44] & w10565;
assign w10568 = ~w10566 & ~w10567;
assign w10569 = ~w10558 & ~w10568;
assign w10570 = w10558 & w10568;
assign w10571 = ~w10569 & ~w10570;
assign w10572 = w10475 & ~w10571;
assign w10573 = ~w10475 & w10571;
assign w10574 = ~w10572 & ~w10573;
assign w10575 = b[18] & w5167;
assign w10576 = b[20] & w4925;
assign w10577 = b[19] & w4918;
assign w10578 = w1347 & w4923;
assign w10579 = ~w10576 & ~w10577;
assign w10580 = ~w10575 & w10579;
assign w10581 = ~w10578 & w10580;
assign w10582 = a[41] & ~w10581;
assign w10583 = ~a[41] & w10581;
assign w10584 = ~w10582 & ~w10583;
assign w10585 = w10574 & w10584;
assign w10586 = ~w10574 & ~w10584;
assign w10587 = ~w10585 & ~w10586;
assign w10588 = ~w10228 & ~w10233;
assign w10589 = w10587 & ~w10588;
assign w10590 = ~w10587 & w10588;
assign w10591 = ~w10589 & ~w10590;
assign w10592 = w10474 & w10591;
assign w10593 = ~w10474 & ~w10591;
assign w10594 = ~w10592 & ~w10593;
assign w10595 = w10464 & ~w10594;
assign w10596 = ~w10464 & w10594;
assign w10597 = ~w10595 & ~w10596;
assign w10598 = w10463 & w10597;
assign w10599 = ~w10463 & ~w10597;
assign w10600 = ~w10598 & ~w10599;
assign w10601 = (~w10252 & w10104) | (~w10252 & w25551) | (w10104 & w25551);
assign w10602 = ~w10600 & w10601;
assign w10603 = w10600 & ~w10601;
assign w10604 = ~w10602 & ~w10603;
assign w10605 = b[27] & w3177;
assign w10606 = b[28] & w2973;
assign w10607 = b[29] & w2978;
assign w10608 = w2734 & w2980;
assign w10609 = ~w10606 & ~w10607;
assign w10610 = ~w10605 & w10609;
assign w10611 = ~w10608 & w10610;
assign w10612 = a[32] & ~w10611;
assign w10613 = ~a[32] & w10611;
assign w10614 = ~w10612 & ~w10613;
assign w10615 = ~w10604 & ~w10614;
assign w10616 = w10604 & w10614;
assign w10617 = ~w10615 & ~w10616;
assign w10618 = w10453 & ~w10617;
assign w10619 = ~w10453 & w10617;
assign w10620 = ~w10618 & ~w10619;
assign w10621 = w10452 & w10620;
assign w10622 = ~w10452 & ~w10620;
assign w10623 = ~w10621 & ~w10622;
assign w10624 = (~w10265 & ~w10082) | (~w10265 & w25436) | (~w10082 & w25436);
assign w10625 = w10623 & w10624;
assign w10626 = ~w10623 & ~w10624;
assign w10627 = ~w10625 & ~w10626;
assign w10628 = b[34] & w1955;
assign w10629 = b[33] & ~w2114;
assign w10630 = b[35] & w1957;
assign w10631 = w1951 & w3918;
assign w10632 = ~w10628 & ~w10629;
assign w10633 = ~w10630 & w10632;
assign w10634 = ~w10631 & w10633;
assign w10635 = a[26] & ~w10634;
assign w10636 = ~a[26] & w10634;
assign w10637 = ~w10635 & ~w10636;
assign w10638 = w10627 & w10637;
assign w10639 = ~w10627 & ~w10637;
assign w10640 = ~w10638 & ~w10639;
assign w10641 = ~w10442 & ~w10640;
assign w10642 = w10442 & w10640;
assign w10643 = ~w10641 & ~w10642;
assign w10644 = ~w10441 & w10643;
assign w10645 = w10441 & ~w10643;
assign w10646 = ~w10644 & ~w10645;
assign w10647 = w10431 & ~w10646;
assign w10648 = ~w10431 & w10646;
assign w10649 = ~w10647 & ~w10648;
assign w10650 = b[41] & w1156;
assign w10651 = b[40] & w1154;
assign w10652 = b[39] & ~w1272;
assign w10653 = w1150 & w5302;
assign w10654 = ~w10650 & ~w10651;
assign w10655 = ~w10652 & w10654;
assign w10656 = ~w10653 & w10655;
assign w10657 = a[20] & ~w10656;
assign w10658 = ~a[20] & w10656;
assign w10659 = ~w10657 & ~w10658;
assign w10660 = ~w10649 & ~w10659;
assign w10661 = w10649 & w10659;
assign w10662 = ~w10660 & ~w10661;
assign w10663 = ~w10430 & ~w10662;
assign w10664 = w10430 & w10662;
assign w10665 = ~w10663 & ~w10664;
assign w10666 = w10429 & ~w10665;
assign w10667 = ~w10429 & w10665;
assign w10668 = ~w10666 & ~w10667;
assign w10669 = w10419 & w10668;
assign w10670 = ~w10419 & ~w10668;
assign w10671 = ~w10669 & ~w10670;
assign w10672 = w10418 & w10671;
assign w10673 = ~w10418 & ~w10671;
assign w10674 = ~w10672 & ~w10673;
assign w10675 = ~w10408 & ~w10674;
assign w10676 = w10408 & w10674;
assign w10677 = ~w10675 & ~w10676;
assign w10678 = ~w10407 & w10677;
assign w10679 = w10407 & ~w10677;
assign w10680 = ~w10678 & ~w10679;
assign w10681 = (~w10312 & w10028) | (~w10312 & w25009) | (w10028 & w25009);
assign w10682 = w10680 & ~w10681;
assign w10683 = ~w10680 & w10681;
assign w10684 = ~w10682 & ~w10683;
assign w10685 = ~w10397 & ~w10684;
assign w10686 = w10397 & w10684;
assign w10687 = ~w10685 & ~w10686;
assign w10688 = (~w10319 & ~w10321) | (~w10319 & w24848) | (~w10321 & w24848);
assign w10689 = w10687 & w10688;
assign w10690 = ~w10687 & ~w10688;
assign w10691 = ~w10689 & ~w10690;
assign w10692 = w10387 & ~w10691;
assign w10693 = ~w10387 & w10691;
assign w10694 = ~w10692 & ~w10693;
assign w10695 = (~w10325 & ~w10007) | (~w10325 & w24689) | (~w10007 & w24689);
assign w10696 = w10694 & w10695;
assign w10697 = ~w10694 & ~w10695;
assign w10698 = ~w10696 & ~w10697;
assign w10699 = ~w10348 & ~w10352;
assign w10700 = ~w10352 & w24394;
assign w10701 = ~w10698 & ~w10699;
assign w10702 = ~w10700 & ~w10701;
assign w10703 = (~w10696 & w10352) | (~w10696 & w24690) | (w10352 & w24690);
assign w10704 = b[55] & w103;
assign w10705 = b[56] & w61;
assign w10706 = b[57] & w68;
assign w10707 = w66 & ~w9992;
assign w10708 = ~w10705 & ~w10706;
assign w10709 = ~w10704 & w10708;
assign w10710 = ~w10707 & w10709;
assign w10711 = a[5] & ~w10710;
assign w10712 = ~a[5] & w10710;
assign w10713 = ~w10711 & ~w10712;
assign w10714 = b[52] & ~w237;
assign w10715 = b[53] & w183;
assign w10716 = b[54] & w185;
assign w10717 = w179 & ~w8998;
assign w10718 = ~w10714 & ~w10715;
assign w10719 = ~w10716 & w10718;
assign w10720 = ~w10717 & w10719;
assign w10721 = a[8] & ~w10720;
assign w10722 = ~a[8] & w10720;
assign w10723 = ~w10721 & ~w10722;
assign w10724 = (~w10679 & w10681) | (~w10679 & w24691) | (w10681 & w24691);
assign w10725 = b[48] & w575;
assign w10726 = b[47] & w573;
assign w10727 = b[46] & ~w649;
assign w10728 = w569 & ~w7170;
assign w10729 = ~w10725 & ~w10726;
assign w10730 = ~w10727 & w10729;
assign w10731 = ~w10728 & w10730;
assign w10732 = a[14] & ~w10731;
assign w10733 = ~a[14] & w10731;
assign w10734 = ~w10732 & ~w10733;
assign w10735 = (~w10666 & ~w10419) | (~w10666 & w25295) | (~w10419 & w25295);
assign w10736 = b[45] & w834;
assign w10737 = b[44] & w838;
assign w10738 = b[43] & ~w934;
assign w10739 = w832 & w6334;
assign w10740 = ~w10736 & ~w10737;
assign w10741 = ~w10738 & w10740;
assign w10742 = ~w10739 & w10741;
assign w10743 = a[17] & ~w10742;
assign w10744 = ~a[17] & w10742;
assign w10745 = ~w10743 & ~w10744;
assign w10746 = b[42] & w1156;
assign w10747 = b[41] & w1154;
assign w10748 = b[40] & ~w1272;
assign w10749 = w1150 & w5548;
assign w10750 = ~w10746 & ~w10747;
assign w10751 = ~w10748 & w10750;
assign w10752 = ~w10749 & w10751;
assign w10753 = a[20] & ~w10752;
assign w10754 = ~a[20] & w10752;
assign w10755 = ~w10753 & ~w10754;
assign w10756 = ~w10645 & ~w10648;
assign w10757 = b[36] & w1957;
assign w10758 = b[34] & ~w2114;
assign w10759 = b[35] & w1955;
assign w10760 = w1951 & w4129;
assign w10761 = ~w10757 & ~w10758;
assign w10762 = ~w10759 & w10761;
assign w10763 = ~w10760 & w10762;
assign w10764 = a[26] & ~w10763;
assign w10765 = ~a[26] & w10763;
assign w10766 = ~w10764 & ~w10765;
assign w10767 = ~w10621 & ~w10625;
assign w10768 = b[28] & w3177;
assign w10769 = b[30] & w2978;
assign w10770 = b[29] & w2973;
assign w10771 = ~w2908 & w2980;
assign w10772 = ~w10769 & ~w10770;
assign w10773 = ~w10768 & w10772;
assign w10774 = ~w10771 & w10773;
assign w10775 = a[32] & ~w10774;
assign w10776 = ~a[32] & w10774;
assign w10777 = ~w10775 & ~w10776;
assign w10778 = ~w10598 & ~w10603;
assign w10779 = b[25] & w3785;
assign w10780 = b[26] & w3578;
assign w10781 = b[27] & w3580;
assign w10782 = w2378 & w3573;
assign w10783 = ~w10780 & ~w10781;
assign w10784 = ~w10779 & w10783;
assign w10785 = ~w10782 & w10784;
assign w10786 = a[35] & ~w10785;
assign w10787 = ~a[35] & w10785;
assign w10788 = ~w10786 & ~w10787;
assign w10789 = b[22] & w4453;
assign w10790 = b[24] & w4243;
assign w10791 = b[23] & w4241;
assign w10792 = w1895 & w4236;
assign w10793 = ~w10790 & ~w10791;
assign w10794 = ~w10789 & w10793;
assign w10795 = ~w10792 & w10794;
assign w10796 = a[38] & ~w10795;
assign w10797 = ~a[38] & w10795;
assign w10798 = ~w10796 & ~w10797;
assign w10799 = ~w10585 & ~w10589;
assign w10800 = b[19] & w5167;
assign w10801 = b[21] & w4925;
assign w10802 = b[20] & w4918;
assign w10803 = w1467 & w4923;
assign w10804 = ~w10801 & ~w10802;
assign w10805 = ~w10800 & w10804;
assign w10806 = ~w10803 & w10805;
assign w10807 = a[41] & ~w10806;
assign w10808 = ~a[41] & w10806;
assign w10809 = ~w10807 & ~w10808;
assign w10810 = b[16] & w5939;
assign w10811 = b[17] & w5670;
assign w10812 = b[18] & w5665;
assign w10813 = ~w1108 & w5663;
assign w10814 = ~w10811 & ~w10812;
assign w10815 = ~w10810 & w10814;
assign w10816 = ~w10813 & w10815;
assign w10817 = a[44] & ~w10816;
assign w10818 = ~a[44] & w10816;
assign w10819 = ~w10817 & ~w10818;
assign w10820 = ~w10552 & ~w10556;
assign w10821 = b[13] & w6732;
assign w10822 = b[15] & w6476;
assign w10823 = b[14] & w6474;
assign w10824 = ~w799 & w6469;
assign w10825 = ~w10822 & ~w10823;
assign w10826 = ~w10821 & w10825;
assign w10827 = ~w10824 & w10826;
assign w10828 = a[47] & ~w10827;
assign w10829 = ~a[47] & w10827;
assign w10830 = ~w10828 & ~w10829;
assign w10831 = ~w10537 & ~w10540;
assign w10832 = ~w10521 & ~w10523;
assign w10833 = b[7] & w8515;
assign w10834 = b[8] & w8200;
assign w10835 = b[9] & w8202;
assign w10836 = w322 & w8195;
assign w10837 = ~w10834 & ~w10835;
assign w10838 = ~w10833 & w10837;
assign w10839 = ~w10836 & w10838;
assign w10840 = a[53] & ~w10839;
assign w10841 = ~a[53] & w10839;
assign w10842 = ~w10840 & ~w10841;
assign w10843 = b[1] & w10496;
assign w10844 = b[2] & w10146;
assign w10845 = b[3] & w10148;
assign w10846 = w46 & w10141;
assign w10847 = ~w10844 & ~w10845;
assign w10848 = ~w10843 & w10847;
assign w10849 = ~w10846 & w10848;
assign w10850 = a[59] & ~w10849;
assign w10851 = ~a[59] & w10849;
assign w10852 = ~w10850 & ~w10851;
assign w10853 = w10490 & w10500;
assign w10854 = a[59] & ~a[60];
assign w10855 = ~a[59] & a[60];
assign w10856 = ~w10854 & ~w10855;
assign w10857 = b[0] & ~w10856;
assign w10858 = w10853 & w10857;
assign w10859 = ~w10853 & ~w10857;
assign w10860 = ~w10858 & ~w10859;
assign w10861 = w10852 & w10860;
assign w10862 = ~w10852 & ~w10860;
assign w10863 = ~w10861 & ~w10862;
assign w10864 = b[4] & w9482;
assign w10865 = b[5] & w9165;
assign w10866 = b[6] & w9160;
assign w10867 = w157 & w9158;
assign w10868 = ~w10865 & ~w10866;
assign w10869 = ~w10864 & w10868;
assign w10870 = ~w10867 & w10869;
assign w10871 = a[56] & ~w10870;
assign w10872 = ~a[56] & w10870;
assign w10873 = ~w10871 & ~w10872;
assign w10874 = w10863 & w10873;
assign w10875 = ~w10863 & ~w10873;
assign w10876 = ~w10874 & ~w10875;
assign w10877 = ~w10505 & ~w10507;
assign w10878 = w10876 & w10877;
assign w10879 = ~w10876 & ~w10877;
assign w10880 = ~w10878 & ~w10879;
assign w10881 = w10842 & w10880;
assign w10882 = ~w10842 & ~w10880;
assign w10883 = ~w10881 & ~w10882;
assign w10884 = w10832 & ~w10883;
assign w10885 = ~w10832 & w10883;
assign w10886 = ~w10884 & ~w10885;
assign w10887 = b[10] & w7586;
assign w10888 = b[11] & w7307;
assign w10889 = b[12] & w7314;
assign w10890 = w536 & w7312;
assign w10891 = ~w10888 & ~w10889;
assign w10892 = ~w10887 & w10891;
assign w10893 = ~w10890 & w10892;
assign w10894 = a[50] & ~w10893;
assign w10895 = ~a[50] & w10893;
assign w10896 = ~w10894 & ~w10895;
assign w10897 = ~w10886 & ~w10896;
assign w10898 = w10886 & w10896;
assign w10899 = ~w10897 & ~w10898;
assign w10900 = ~w10831 & w10899;
assign w10901 = w10831 & ~w10899;
assign w10902 = ~w10900 & ~w10901;
assign w10903 = w10830 & w10902;
assign w10904 = ~w10830 & ~w10902;
assign w10905 = ~w10903 & ~w10904;
assign w10906 = w10820 & ~w10905;
assign w10907 = ~w10820 & w10905;
assign w10908 = ~w10906 & ~w10907;
assign w10909 = ~w10819 & ~w10908;
assign w10910 = w10819 & w10908;
assign w10911 = ~w10909 & ~w10910;
assign w10912 = ~w10570 & ~w10573;
assign w10913 = w10911 & ~w10912;
assign w10914 = ~w10911 & w10912;
assign w10915 = ~w10913 & ~w10914;
assign w10916 = w10809 & w10915;
assign w10917 = ~w10809 & ~w10915;
assign w10918 = ~w10916 & ~w10917;
assign w10919 = w10799 & ~w10918;
assign w10920 = ~w10799 & w10918;
assign w10921 = ~w10919 & ~w10920;
assign w10922 = w10798 & w10921;
assign w10923 = ~w10798 & ~w10921;
assign w10924 = ~w10922 & ~w10923;
assign w10925 = ~w10592 & ~w10596;
assign w10926 = w10924 & ~w10925;
assign w10927 = ~w10924 & w10925;
assign w10928 = ~w10926 & ~w10927;
assign w10929 = w10788 & w10928;
assign w10930 = ~w10788 & ~w10928;
assign w10931 = ~w10929 & ~w10930;
assign w10932 = w10778 & ~w10931;
assign w10933 = ~w10778 & w10931;
assign w10934 = ~w10932 & ~w10933;
assign w10935 = w10777 & w10934;
assign w10936 = ~w10777 & ~w10934;
assign w10937 = ~w10935 & ~w10936;
assign w10938 = (~w10616 & w10453) | (~w10616 & w25552) | (w10453 & w25552);
assign w10939 = w10937 & ~w10938;
assign w10940 = ~w10937 & w10938;
assign w10941 = ~w10939 & ~w10940;
assign w10942 = b[33] & w2438;
assign w10943 = b[32] & w2436;
assign w10944 = b[31] & ~w2622;
assign w10945 = w2432 & w3499;
assign w10946 = ~w10942 & ~w10943;
assign w10947 = ~w10944 & w10946;
assign w10948 = ~w10945 & w10947;
assign w10949 = a[29] & ~w10948;
assign w10950 = ~a[29] & w10948;
assign w10951 = ~w10949 & ~w10950;
assign w10952 = w10941 & w10951;
assign w10953 = ~w10941 & ~w10951;
assign w10954 = ~w10952 & ~w10953;
assign w10955 = w10767 & ~w10954;
assign w10956 = ~w10767 & w10954;
assign w10957 = ~w10955 & ~w10956;
assign w10958 = w10766 & w10957;
assign w10959 = ~w10766 & ~w10957;
assign w10960 = ~w10958 & ~w10959;
assign w10961 = (~w10639 & ~w10442) | (~w10639 & w24395) | (~w10442 & w24395);
assign w10962 = ~w10960 & ~w10961;
assign w10963 = w10960 & w10961;
assign w10964 = ~w10962 & ~w10963;
assign w10965 = b[37] & ~w1676;
assign w10966 = b[39] & w1519;
assign w10967 = b[38] & w1517;
assign w10968 = w1513 & ~w4812;
assign w10969 = ~w10965 & ~w10966;
assign w10970 = ~w10967 & w10969;
assign w10971 = ~w10968 & w10970;
assign w10972 = a[23] & ~w10971;
assign w10973 = ~a[23] & w10971;
assign w10974 = ~w10972 & ~w10973;
assign w10975 = w10964 & w10974;
assign w10976 = ~w10964 & ~w10974;
assign w10977 = ~w10975 & ~w10976;
assign w10978 = ~w10756 & ~w10977;
assign w10979 = w10756 & w10977;
assign w10980 = ~w10978 & ~w10979;
assign w10981 = ~w10755 & w10980;
assign w10982 = w10755 & ~w10980;
assign w10983 = ~w10981 & ~w10982;
assign w10984 = ~w10660 & ~w10664;
assign w10985 = w10983 & w10984;
assign w10986 = ~w10983 & ~w10984;
assign w10987 = ~w10985 & ~w10986;
assign w10988 = ~w10745 & ~w10987;
assign w10989 = w10745 & w10987;
assign w10990 = ~w10988 & ~w10989;
assign w10991 = w10735 & w10990;
assign w10992 = ~w10735 & ~w10990;
assign w10993 = ~w10991 & ~w10992;
assign w10994 = w10734 & ~w10993;
assign w10995 = ~w10734 & w10993;
assign w10996 = ~w10994 & ~w10995;
assign w10997 = (~w10673 & ~w10408) | (~w10673 & w25177) | (~w10408 & w25177);
assign w10998 = w10996 & w10997;
assign w10999 = ~w10996 & ~w10997;
assign w11000 = ~w10998 & ~w10999;
assign w11001 = b[49] & ~w419;
assign w11002 = b[50] & w358;
assign w11003 = b[51] & w360;
assign w11004 = w354 & ~w8058;
assign w11005 = ~w11001 & ~w11002;
assign w11006 = ~w11003 & w11005;
assign w11007 = ~w11004 & w11006;
assign w11008 = a[11] & ~w11007;
assign w11009 = ~a[11] & w11007;
assign w11010 = ~w11008 & ~w11009;
assign w11011 = w11000 & w11010;
assign w11012 = ~w11000 & ~w11010;
assign w11013 = ~w11011 & ~w11012;
assign w11014 = ~w10724 & w11013;
assign w11015 = w10724 & ~w11013;
assign w11016 = ~w11014 & ~w11015;
assign w11017 = w10723 & w11016;
assign w11018 = ~w10723 & ~w11016;
assign w11019 = ~w11017 & ~w11018;
assign w11020 = ~w10685 & ~w10689;
assign w11021 = w11019 & w11020;
assign w11022 = ~w11019 & ~w11020;
assign w11023 = ~w11021 & ~w11022;
assign w11024 = ~w10713 & ~w11023;
assign w11025 = w10713 & w11023;
assign w11026 = ~w11024 & ~w11025;
assign w11027 = b[60] & w11;
assign w11028 = b[59] & w9;
assign w11029 = ~w10366 & ~w10369;
assign w11030 = ~b[59] & ~b[60];
assign w11031 = b[59] & b[60];
assign w11032 = ~w11030 & ~w11031;
assign w11033 = ~w11029 & w11032;
assign w11034 = w11029 & ~w11032;
assign w11035 = ~w11033 & ~w11034;
assign w11036 = w5 & w11035;
assign w11037 = ~w11027 & ~w11028;
assign w11038 = ~w11036 & w11037;
assign w11039 = b[58] & w24;
assign w11040 = a[2] & ~w11039;
assign w11041 = w11038 & ~w11040;
assign w11042 = a[2] & ~w11038;
assign w11043 = ~w11041 & ~w11042;
assign w11044 = w11026 & w11043;
assign w11045 = ~w11026 & ~w11043;
assign w11046 = ~w11044 & ~w11045;
assign w11047 = ~w10385 & ~w10692;
assign w11048 = w11046 & ~w11047;
assign w11049 = ~w11046 & w11047;
assign w11050 = ~w11048 & ~w11049;
assign w11051 = w10703 & ~w11050;
assign w11052 = ~w10703 & w11050;
assign w11053 = ~w11051 & ~w11052;
assign w11054 = ~w11025 & ~w11044;
assign w11055 = b[56] & w103;
assign w11056 = b[58] & w68;
assign w11057 = b[57] & w61;
assign w11058 = w66 & ~w10339;
assign w11059 = ~w11056 & ~w11057;
assign w11060 = ~w11055 & w11059;
assign w11061 = ~w11058 & w11060;
assign w11062 = a[5] & ~w11061;
assign w11063 = ~a[5] & w11061;
assign w11064 = ~w11062 & ~w11063;
assign w11065 = (~w11011 & w10724) | (~w11011 & w25178) | (w10724 & w25178);
assign w11066 = b[51] & w358;
assign w11067 = b[50] & ~w419;
assign w11068 = b[52] & w360;
assign w11069 = w354 & ~w8371;
assign w11070 = ~w11066 & ~w11067;
assign w11071 = ~w11068 & w11070;
assign w11072 = ~w11069 & w11071;
assign w11073 = a[11] & ~w11072;
assign w11074 = ~a[11] & w11072;
assign w11075 = ~w11073 & ~w11074;
assign w11076 = (~w10994 & ~w10997) | (~w10994 & w25296) | (~w10997 & w25296);
assign w11077 = b[49] & w575;
assign w11078 = b[47] & ~w649;
assign w11079 = b[48] & w573;
assign w11080 = w569 & ~w7468;
assign w11081 = ~w11077 & ~w11078;
assign w11082 = ~w11079 & w11081;
assign w11083 = ~w11080 & w11082;
assign w11084 = a[14] & ~w11083;
assign w11085 = ~a[14] & w11083;
assign w11086 = ~w11084 & ~w11085;
assign w11087 = b[44] & ~w934;
assign w11088 = b[46] & w834;
assign w11089 = b[45] & w838;
assign w11090 = w832 & ~w6613;
assign w11091 = ~w11087 & ~w11088;
assign w11092 = ~w11089 & w11091;
assign w11093 = ~w11090 & w11092;
assign w11094 = a[17] & ~w11093;
assign w11095 = ~a[17] & w11093;
assign w11096 = ~w11094 & ~w11095;
assign w11097 = ~w10982 & ~w10985;
assign w11098 = b[38] & ~w1676;
assign w11099 = b[40] & w1519;
assign w11100 = b[39] & w1517;
assign w11101 = w1513 & ~w5058;
assign w11102 = ~w11098 & ~w11099;
assign w11103 = ~w11100 & w11102;
assign w11104 = ~w11101 & w11103;
assign w11105 = a[23] & ~w11104;
assign w11106 = ~a[23] & w11104;
assign w11107 = ~w11105 & ~w11106;
assign w11108 = b[32] & ~w2622;
assign w11109 = b[34] & w2438;
assign w11110 = b[33] & w2436;
assign w11111 = w2432 & ~w3710;
assign w11112 = ~w11108 & ~w11109;
assign w11113 = ~w11110 & w11112;
assign w11114 = ~w11111 & w11113;
assign w11115 = a[29] & ~w11114;
assign w11116 = ~a[29] & w11114;
assign w11117 = ~w11115 & ~w11116;
assign w11118 = (~w10935 & w10938) | (~w10935 & w25179) | (w10938 & w25179);
assign w11119 = b[29] & w3177;
assign w11120 = b[31] & w2978;
assign w11121 = b[30] & w2973;
assign w11122 = w2980 & ~w3112;
assign w11123 = ~w11120 & ~w11121;
assign w11124 = ~w11119 & w11123;
assign w11125 = ~w11122 & w11124;
assign w11126 = a[32] & ~w11125;
assign w11127 = ~a[32] & w11125;
assign w11128 = ~w11126 & ~w11127;
assign w11129 = b[26] & w3785;
assign w11130 = b[27] & w3578;
assign w11131 = b[28] & w3580;
assign w11132 = w2559 & w3573;
assign w11133 = ~w11130 & ~w11131;
assign w11134 = ~w11129 & w11133;
assign w11135 = ~w11132 & w11134;
assign w11136 = a[35] & ~w11135;
assign w11137 = ~a[35] & w11135;
assign w11138 = ~w11136 & ~w11137;
assign w11139 = ~w10922 & ~w10926;
assign w11140 = b[23] & w4453;
assign w11141 = b[25] & w4243;
assign w11142 = b[24] & w4241;
assign w11143 = w2061 & w4236;
assign w11144 = ~w11141 & ~w11142;
assign w11145 = ~w11140 & w11144;
assign w11146 = ~w11143 & w11145;
assign w11147 = a[38] & ~w11146;
assign w11148 = ~a[38] & w11146;
assign w11149 = ~w11147 & ~w11148;
assign w11150 = b[20] & w5167;
assign w11151 = b[22] & w4925;
assign w11152 = b[21] & w4918;
assign w11153 = w1615 & w4923;
assign w11154 = ~w11151 & ~w11152;
assign w11155 = ~w11150 & w11154;
assign w11156 = ~w11153 & w11155;
assign w11157 = a[41] & ~w11156;
assign w11158 = ~a[41] & w11156;
assign w11159 = ~w11157 & ~w11158;
assign w11160 = (~w10910 & w10912) | (~w10910 & w25180) | (w10912 & w25180);
assign w11161 = ~w10903 & ~w10907;
assign w11162 = b[14] & w6732;
assign w11163 = b[16] & w6476;
assign w11164 = b[15] & w6474;
assign w11165 = w905 & w6469;
assign w11166 = ~w11163 & ~w11164;
assign w11167 = ~w11162 & w11166;
assign w11168 = ~w11165 & w11167;
assign w11169 = a[47] & ~w11168;
assign w11170 = ~a[47] & w11168;
assign w11171 = ~w11169 & ~w11170;
assign w11172 = (~w10898 & w10831) | (~w10898 & w25181) | (w10831 & w25181);
assign w11173 = (~w10874 & ~w10877) | (~w10874 & w25182) | (~w10877 & w25182);
assign w11174 = ~w10858 & ~w10861;
assign w11175 = b[2] & w10496;
assign w11176 = b[4] & w10148;
assign w11177 = b[3] & w10146;
assign w11178 = w84 & w10141;
assign w11179 = ~w11176 & ~w11177;
assign w11180 = ~w11175 & w11179;
assign w11181 = ~w11178 & w11180;
assign w11182 = a[59] & ~w11181;
assign w11183 = ~a[59] & w11181;
assign w11184 = ~w11182 & ~w11183;
assign w11185 = a[62] & w10857;
assign w11186 = a[61] & ~a[62];
assign w11187 = ~a[61] & a[62];
assign w11188 = ~w11186 & ~w11187;
assign w11189 = ~w10856 & ~w11188;
assign w11190 = ~w8 & w11189;
assign w11191 = a[60] & ~a[61];
assign w11192 = ~a[60] & a[61];
assign w11193 = ~w11191 & ~w11192;
assign w11194 = w10856 & ~w11193;
assign w11195 = b[0] & w11194;
assign w11196 = ~w10856 & w11188;
assign w11197 = b[1] & w11196;
assign w11198 = ~w11190 & ~w11195;
assign w11199 = ~w11197 & w11198;
assign w11200 = ~w11185 & w11199;
assign w11201 = w11185 & ~w11199;
assign w11202 = ~w11200 & ~w11201;
assign w11203 = ~w11184 & ~w11202;
assign w11204 = w11184 & w11202;
assign w11205 = ~w11203 & ~w11204;
assign w11206 = ~w11174 & w11205;
assign w11207 = w11174 & ~w11205;
assign w11208 = ~w11206 & ~w11207;
assign w11209 = b[5] & w9482;
assign w11210 = b[7] & w9160;
assign w11211 = b[6] & w9165;
assign w11212 = w216 & w9158;
assign w11213 = ~w11210 & ~w11211;
assign w11214 = ~w11209 & w11213;
assign w11215 = ~w11212 & w11214;
assign w11216 = a[56] & ~w11215;
assign w11217 = ~a[56] & w11215;
assign w11218 = ~w11216 & ~w11217;
assign w11219 = ~w11208 & ~w11218;
assign w11220 = w11208 & w11218;
assign w11221 = ~w11219 & ~w11220;
assign w11222 = ~w11173 & w11221;
assign w11223 = w11173 & ~w11221;
assign w11224 = ~w11222 & ~w11223;
assign w11225 = b[8] & w8515;
assign w11226 = b[9] & w8200;
assign w11227 = b[10] & w8202;
assign w11228 = w397 & w8195;
assign w11229 = ~w11226 & ~w11227;
assign w11230 = ~w11225 & w11229;
assign w11231 = ~w11228 & w11230;
assign w11232 = a[53] & ~w11231;
assign w11233 = ~a[53] & w11231;
assign w11234 = ~w11232 & ~w11233;
assign w11235 = w11224 & w11234;
assign w11236 = ~w11224 & ~w11234;
assign w11237 = ~w11235 & ~w11236;
assign w11238 = (~w10881 & w10832) | (~w10881 & w25183) | (w10832 & w25183);
assign w11239 = ~w11237 & w11238;
assign w11240 = w11237 & ~w11238;
assign w11241 = ~w11239 & ~w11240;
assign w11242 = b[11] & w7586;
assign w11243 = b[12] & w7307;
assign w11244 = b[13] & w7314;
assign w11245 = w628 & w7312;
assign w11246 = ~w11243 & ~w11244;
assign w11247 = ~w11242 & w11246;
assign w11248 = ~w11245 & w11247;
assign w11249 = a[50] & ~w11248;
assign w11250 = ~a[50] & w11248;
assign w11251 = ~w11249 & ~w11250;
assign w11252 = w11241 & w11251;
assign w11253 = ~w11241 & ~w11251;
assign w11254 = ~w11252 & ~w11253;
assign w11255 = w11172 & w11254;
assign w11256 = ~w11172 & ~w11254;
assign w11257 = ~w11255 & ~w11256;
assign w11258 = w11171 & ~w11257;
assign w11259 = ~w11171 & w11257;
assign w11260 = ~w11258 & ~w11259;
assign w11261 = w11161 & ~w11260;
assign w11262 = ~w11161 & w11260;
assign w11263 = ~w11261 & ~w11262;
assign w11264 = b[17] & w5939;
assign w11265 = b[18] & w5670;
assign w11266 = b[19] & w5665;
assign w11267 = ~w1231 & w5663;
assign w11268 = ~w11265 & ~w11266;
assign w11269 = ~w11264 & w11268;
assign w11270 = ~w11267 & w11269;
assign w11271 = a[44] & ~w11270;
assign w11272 = ~a[44] & w11270;
assign w11273 = ~w11271 & ~w11272;
assign w11274 = w11263 & w11273;
assign w11275 = ~w11263 & ~w11273;
assign w11276 = ~w11274 & ~w11275;
assign w11277 = w11160 & w11276;
assign w11278 = ~w11160 & ~w11276;
assign w11279 = ~w11277 & ~w11278;
assign w11280 = w11159 & ~w11279;
assign w11281 = ~w11159 & w11279;
assign w11282 = ~w11280 & ~w11281;
assign w11283 = ~w10916 & ~w10920;
assign w11284 = w11282 & ~w11283;
assign w11285 = ~w11282 & w11283;
assign w11286 = ~w11284 & ~w11285;
assign w11287 = w11149 & w11286;
assign w11288 = ~w11149 & ~w11286;
assign w11289 = ~w11287 & ~w11288;
assign w11290 = w11139 & ~w11289;
assign w11291 = ~w11139 & w11289;
assign w11292 = ~w11290 & ~w11291;
assign w11293 = w11138 & w11292;
assign w11294 = ~w11138 & ~w11292;
assign w11295 = ~w11293 & ~w11294;
assign w11296 = (~w10929 & w10778) | (~w10929 & w25184) | (w10778 & w25184);
assign w11297 = w11295 & w11296;
assign w11298 = ~w11295 & ~w11296;
assign w11299 = ~w11297 & ~w11298;
assign w11300 = w11128 & ~w11299;
assign w11301 = ~w11128 & w11299;
assign w11302 = ~w11300 & ~w11301;
assign w11303 = ~w11118 & w11302;
assign w11304 = w11118 & ~w11302;
assign w11305 = ~w11303 & ~w11304;
assign w11306 = w11117 & w11305;
assign w11307 = ~w11117 & ~w11305;
assign w11308 = ~w11306 & ~w11307;
assign w11309 = (~w10952 & w10767) | (~w10952 & w25553) | (w10767 & w25553);
assign w11310 = ~w11308 & w11309;
assign w11311 = w11308 & ~w11309;
assign w11312 = ~w11310 & ~w11311;
assign w11313 = b[37] & w1957;
assign w11314 = b[36] & w1955;
assign w11315 = b[35] & ~w2114;
assign w11316 = w1951 & ~w4357;
assign w11317 = ~w11313 & ~w11314;
assign w11318 = ~w11315 & w11317;
assign w11319 = ~w11316 & w11318;
assign w11320 = a[26] & ~w11319;
assign w11321 = ~a[26] & w11319;
assign w11322 = ~w11320 & ~w11321;
assign w11323 = w11312 & w11322;
assign w11324 = ~w11312 & ~w11322;
assign w11325 = ~w11323 & ~w11324;
assign w11326 = ~w10958 & ~w10963;
assign w11327 = ~w11325 & w11326;
assign w11328 = w11325 & ~w11326;
assign w11329 = ~w11327 & ~w11328;
assign w11330 = w11107 & w11329;
assign w11331 = ~w11107 & ~w11329;
assign w11332 = ~w11330 & ~w11331;
assign w11333 = (~w10976 & ~w10756) | (~w10976 & w24396) | (~w10756 & w24396);
assign w11334 = ~w11332 & ~w11333;
assign w11335 = w11332 & w11333;
assign w11336 = ~w11334 & ~w11335;
assign w11337 = b[43] & w1156;
assign w11338 = b[41] & ~w1272;
assign w11339 = b[42] & w1154;
assign w11340 = w1150 & w5811;
assign w11341 = ~w11337 & ~w11338;
assign w11342 = ~w11339 & w11341;
assign w11343 = ~w11340 & w11342;
assign w11344 = a[20] & ~w11343;
assign w11345 = ~a[20] & w11343;
assign w11346 = ~w11344 & ~w11345;
assign w11347 = w11336 & w11346;
assign w11348 = ~w11336 & ~w11346;
assign w11349 = ~w11347 & ~w11348;
assign w11350 = w11097 & ~w11349;
assign w11351 = ~w11097 & w11349;
assign w11352 = ~w11350 & ~w11351;
assign w11353 = w11096 & w11352;
assign w11354 = ~w11096 & ~w11352;
assign w11355 = ~w11353 & ~w11354;
assign w11356 = ~w10988 & ~w10991;
assign w11357 = w11355 & w11356;
assign w11358 = ~w11355 & ~w11356;
assign w11359 = ~w11357 & ~w11358;
assign w11360 = ~w11086 & ~w11359;
assign w11361 = w11086 & w11359;
assign w11362 = ~w11360 & ~w11361;
assign w11363 = w11076 & w11362;
assign w11364 = ~w11076 & ~w11362;
assign w11365 = ~w11363 & ~w11364;
assign w11366 = w11075 & ~w11365;
assign w11367 = ~w11075 & w11365;
assign w11368 = ~w11366 & ~w11367;
assign w11369 = ~w11065 & w11368;
assign w11370 = w11065 & ~w11368;
assign w11371 = ~w11369 & ~w11370;
assign w11372 = b[53] & ~w237;
assign w11373 = b[55] & w185;
assign w11374 = b[54] & w183;
assign w11375 = w179 & ~w9330;
assign w11376 = ~w11372 & ~w11373;
assign w11377 = ~w11374 & w11376;
assign w11378 = ~w11375 & w11377;
assign w11379 = a[8] & ~w11378;
assign w11380 = ~a[8] & w11378;
assign w11381 = ~w11379 & ~w11380;
assign w11382 = w11371 & w11381;
assign w11383 = ~w11371 & ~w11381;
assign w11384 = ~w11382 & ~w11383;
assign w11385 = (~w11017 & ~w11020) | (~w11017 & w24692) | (~w11020 & w24692);
assign w11386 = w11384 & w11385;
assign w11387 = ~w11384 & ~w11385;
assign w11388 = ~w11386 & ~w11387;
assign w11389 = w11064 & ~w11388;
assign w11390 = ~w11064 & w11388;
assign w11391 = ~w11389 & ~w11390;
assign w11392 = b[61] & w11;
assign w11393 = b[60] & w9;
assign w11394 = (~w11031 & w11029) | (~w11031 & w25185) | (w11029 & w25185);
assign w11395 = ~b[60] & ~b[61];
assign w11396 = b[60] & b[61];
assign w11397 = ~w11395 & ~w11396;
assign w11398 = ~w11394 & w11397;
assign w11399 = w11394 & ~w11397;
assign w11400 = ~w11398 & ~w11399;
assign w11401 = w5 & w11400;
assign w11402 = ~w11392 & ~w11393;
assign w11403 = ~w11401 & w11402;
assign w11404 = b[59] & w24;
assign w11405 = a[2] & ~w11404;
assign w11406 = w11403 & ~w11405;
assign w11407 = a[2] & ~w11403;
assign w11408 = ~w11406 & ~w11407;
assign w11409 = w11391 & w11408;
assign w11410 = ~w11391 & ~w11408;
assign w11411 = ~w11409 & ~w11410;
assign w11412 = w11054 & ~w11411;
assign w11413 = ~w11054 & w11411;
assign w11414 = ~w11412 & ~w11413;
assign w11415 = (~w11048 & ~w11050) | (~w11048 & w24693) | (~w11050 & w24693);
assign w11416 = w11414 & w11415;
assign w11417 = ~w11414 & ~w11415;
assign w11418 = ~w11416 & ~w11417;
assign w11419 = b[56] & w185;
assign w11420 = b[55] & w183;
assign w11421 = b[54] & ~w237;
assign w11422 = w179 & w9657;
assign w11423 = ~w11419 & ~w11420;
assign w11424 = ~w11421 & w11423;
assign w11425 = ~w11422 & w11424;
assign w11426 = a[8] & ~w11425;
assign w11427 = ~a[8] & w11425;
assign w11428 = ~w11426 & ~w11427;
assign w11429 = w66 & w10371;
assign w11430 = b[58] & w61;
assign w11431 = b[59] & w68;
assign w11432 = b[57] & w103;
assign w11433 = ~w11430 & ~w11431;
assign w11434 = ~w11432 & w11433;
assign w11435 = ~w11429 & w11434;
assign w11436 = ~a[5] & ~w11435;
assign w11437 = w246 & w10371;
assign w11438 = a[5] & w11434;
assign w11439 = ~w11437 & w11438;
assign w11440 = ~w11436 & ~w11439;
assign w11441 = w11428 & ~w11440;
assign w11442 = ~w11428 & w11440;
assign w11443 = ~w11441 & ~w11442;
assign w11444 = (~w11366 & w11065) | (~w11366 & w25297) | (w11065 & w25297);
assign w11445 = b[52] & w358;
assign w11446 = b[51] & ~w419;
assign w11447 = b[53] & w360;
assign w11448 = w354 & w8683;
assign w11449 = ~w11445 & ~w11446;
assign w11450 = ~w11447 & w11449;
assign w11451 = ~w11448 & w11450;
assign w11452 = a[11] & ~w11451;
assign w11453 = ~a[11] & w11451;
assign w11454 = ~w11452 & ~w11453;
assign w11455 = b[48] & ~w649;
assign w11456 = b[49] & w573;
assign w11457 = b[50] & w575;
assign w11458 = w569 & w7759;
assign w11459 = ~w11455 & ~w11456;
assign w11460 = ~w11457 & w11459;
assign w11461 = ~w11458 & w11460;
assign w11462 = a[14] & ~w11461;
assign w11463 = ~a[14] & w11461;
assign w11464 = ~w11462 & ~w11463;
assign w11465 = ~w11353 & ~w11357;
assign w11466 = b[42] & ~w1272;
assign w11467 = b[44] & w1156;
assign w11468 = b[43] & w1154;
assign w11469 = w1150 & w6069;
assign w11470 = ~w11466 & ~w11467;
assign w11471 = ~w11468 & w11470;
assign w11472 = ~w11469 & w11471;
assign w11473 = a[20] & ~w11472;
assign w11474 = ~a[20] & w11472;
assign w11475 = ~w11473 & ~w11474;
assign w11476 = ~w11330 & ~w11335;
assign w11477 = b[40] & w1517;
assign w11478 = b[39] & ~w1676;
assign w11479 = b[41] & w1519;
assign w11480 = w1513 & w5302;
assign w11481 = ~w11477 & ~w11478;
assign w11482 = ~w11479 & w11481;
assign w11483 = ~w11480 & w11482;
assign w11484 = a[23] & ~w11483;
assign w11485 = ~a[23] & w11483;
assign w11486 = ~w11484 & ~w11485;
assign w11487 = (~w11323 & w11326) | (~w11323 & w25554) | (w11326 & w25554);
assign w11488 = b[38] & w1957;
assign w11489 = b[36] & ~w2114;
assign w11490 = b[37] & w1955;
assign w11491 = w1951 & w4582;
assign w11492 = ~w11488 & ~w11489;
assign w11493 = ~w11490 & w11492;
assign w11494 = ~w11491 & w11493;
assign w11495 = a[26] & ~w11494;
assign w11496 = ~a[26] & w11494;
assign w11497 = ~w11495 & ~w11496;
assign w11498 = b[34] & w2436;
assign w11499 = b[35] & w2438;
assign w11500 = b[33] & ~w2622;
assign w11501 = w2432 & w3918;
assign w11502 = ~w11498 & ~w11499;
assign w11503 = ~w11500 & w11502;
assign w11504 = ~w11501 & w11503;
assign w11505 = a[29] & ~w11504;
assign w11506 = ~a[29] & w11504;
assign w11507 = ~w11505 & ~w11506;
assign w11508 = b[30] & w3177;
assign w11509 = b[31] & w2973;
assign w11510 = b[32] & w2978;
assign w11511 = w2980 & w3304;
assign w11512 = ~w11509 & ~w11510;
assign w11513 = ~w11508 & w11512;
assign w11514 = ~w11511 & w11513;
assign w11515 = a[32] & ~w11514;
assign w11516 = ~a[32] & w11514;
assign w11517 = ~w11515 & ~w11516;
assign w11518 = (~w11294 & ~w11296) | (~w11294 & w24694) | (~w11296 & w24694);
assign w11519 = b[27] & w3785;
assign w11520 = b[28] & w3578;
assign w11521 = b[29] & w3580;
assign w11522 = w2734 & w3573;
assign w11523 = ~w11520 & ~w11521;
assign w11524 = ~w11519 & w11523;
assign w11525 = ~w11522 & w11524;
assign w11526 = a[35] & ~w11525;
assign w11527 = ~a[35] & w11525;
assign w11528 = ~w11526 & ~w11527;
assign w11529 = (~w11280 & w11283) | (~w11280 & w25186) | (w11283 & w25186);
assign w11530 = b[18] & w5939;
assign w11531 = b[19] & w5670;
assign w11532 = b[20] & w5665;
assign w11533 = w1347 & w5663;
assign w11534 = ~w11531 & ~w11532;
assign w11535 = ~w11530 & w11534;
assign w11536 = ~w11533 & w11535;
assign w11537 = a[44] & ~w11536;
assign w11538 = ~a[44] & w11536;
assign w11539 = ~w11537 & ~w11538;
assign w11540 = (~w11258 & w11161) | (~w11258 & w25187) | (w11161 & w25187);
assign w11541 = (~w11235 & w11238) | (~w11235 & w25298) | (w11238 & w25298);
assign w11542 = (~w11220 & w11173) | (~w11220 & w25299) | (w11173 & w25299);
assign w11543 = ~w11204 & ~w11206;
assign w11544 = b[3] & w10496;
assign w11545 = b[5] & w10148;
assign w11546 = b[4] & w10146;
assign w11547 = w116 & w10141;
assign w11548 = ~w11545 & ~w11546;
assign w11549 = ~w11544 & w11548;
assign w11550 = ~w11547 & w11549;
assign w11551 = a[59] & ~w11550;
assign w11552 = ~a[59] & w11550;
assign w11553 = ~w11551 & ~w11552;
assign w11554 = a[62] & ~w10857;
assign w11555 = w11199 & w11554;
assign w11556 = a[62] & ~w11555;
assign w11557 = w22 & w11189;
assign w11558 = b[2] & w11196;
assign w11559 = b[1] & w11194;
assign w11560 = w10856 & ~w11188;
assign w11561 = w11193 & w11560;
assign w11562 = b[0] & w11561;
assign w11563 = ~w11557 & ~w11558;
assign w11564 = ~w11559 & w11563;
assign w11565 = ~w11562 & w11564;
assign w11566 = ~w11556 & w11565;
assign w11567 = w11556 & ~w11565;
assign w11568 = ~w11566 & ~w11567;
assign w11569 = ~w11553 & ~w11568;
assign w11570 = w11553 & w11568;
assign w11571 = ~w11569 & ~w11570;
assign w11572 = w11543 & w11571;
assign w11573 = ~w11543 & ~w11571;
assign w11574 = ~w11572 & ~w11573;
assign w11575 = b[6] & w9482;
assign w11576 = b[7] & w9165;
assign w11577 = b[8] & w9160;
assign w11578 = w270 & w9158;
assign w11579 = ~w11576 & ~w11577;
assign w11580 = ~w11575 & w11579;
assign w11581 = ~w11578 & w11580;
assign w11582 = a[56] & ~w11581;
assign w11583 = ~a[56] & w11581;
assign w11584 = ~w11582 & ~w11583;
assign w11585 = ~w11574 & w11584;
assign w11586 = w11574 & ~w11584;
assign w11587 = ~w11585 & ~w11586;
assign w11588 = ~w11542 & w11587;
assign w11589 = w11542 & ~w11587;
assign w11590 = ~w11588 & ~w11589;
assign w11591 = b[9] & w8515;
assign w11592 = b[10] & w8200;
assign w11593 = b[11] & w8202;
assign w11594 = w469 & w8195;
assign w11595 = ~w11592 & ~w11593;
assign w11596 = ~w11591 & w11595;
assign w11597 = ~w11594 & w11596;
assign w11598 = a[53] & ~w11597;
assign w11599 = ~a[53] & w11597;
assign w11600 = ~w11598 & ~w11599;
assign w11601 = ~w11590 & ~w11600;
assign w11602 = w11590 & w11600;
assign w11603 = ~w11601 & ~w11602;
assign w11604 = ~w11541 & w11603;
assign w11605 = w11541 & ~w11603;
assign w11606 = ~w11604 & ~w11605;
assign w11607 = b[12] & w7586;
assign w11608 = b[14] & w7314;
assign w11609 = b[13] & w7307;
assign w11610 = w714 & w7312;
assign w11611 = ~w11608 & ~w11609;
assign w11612 = ~w11607 & w11611;
assign w11613 = ~w11610 & w11612;
assign w11614 = a[50] & ~w11613;
assign w11615 = ~a[50] & w11613;
assign w11616 = ~w11614 & ~w11615;
assign w11617 = w11606 & w11616;
assign w11618 = ~w11606 & ~w11616;
assign w11619 = ~w11617 & ~w11618;
assign w11620 = (~w11253 & ~w11172) | (~w11253 & w25300) | (~w11172 & w25300);
assign w11621 = w11619 & w11620;
assign w11622 = ~w11619 & ~w11620;
assign w11623 = ~w11621 & ~w11622;
assign w11624 = b[15] & w6732;
assign w11625 = b[17] & w6476;
assign w11626 = b[16] & w6474;
assign w11627 = w1008 & w6469;
assign w11628 = ~w11625 & ~w11626;
assign w11629 = ~w11624 & w11628;
assign w11630 = ~w11627 & w11629;
assign w11631 = a[47] & ~w11630;
assign w11632 = ~a[47] & w11630;
assign w11633 = ~w11631 & ~w11632;
assign w11634 = ~w11623 & ~w11633;
assign w11635 = w11623 & w11633;
assign w11636 = ~w11634 & ~w11635;
assign w11637 = ~w11540 & w11636;
assign w11638 = w11540 & ~w11636;
assign w11639 = ~w11637 & ~w11638;
assign w11640 = w11539 & w11639;
assign w11641 = ~w11539 & ~w11639;
assign w11642 = ~w11640 & ~w11641;
assign w11643 = (~w11275 & ~w11160) | (~w11275 & w24695) | (~w11160 & w24695);
assign w11644 = w11642 & w11643;
assign w11645 = ~w11642 & ~w11643;
assign w11646 = ~w11644 & ~w11645;
assign w11647 = b[21] & w5167;
assign w11648 = b[22] & w4918;
assign w11649 = b[23] & w4925;
assign w11650 = w1755 & w4923;
assign w11651 = ~w11648 & ~w11649;
assign w11652 = ~w11647 & w11651;
assign w11653 = ~w11650 & w11652;
assign w11654 = a[41] & ~w11653;
assign w11655 = ~a[41] & w11653;
assign w11656 = ~w11654 & ~w11655;
assign w11657 = w11646 & w11656;
assign w11658 = ~w11646 & ~w11656;
assign w11659 = ~w11657 & ~w11658;
assign w11660 = w11529 & ~w11659;
assign w11661 = ~w11529 & w11659;
assign w11662 = ~w11660 & ~w11661;
assign w11663 = b[24] & w4453;
assign w11664 = b[26] & w4243;
assign w11665 = b[25] & w4241;
assign w11666 = w2219 & w4236;
assign w11667 = ~w11664 & ~w11665;
assign w11668 = ~w11663 & w11667;
assign w11669 = ~w11666 & w11668;
assign w11670 = a[38] & ~w11669;
assign w11671 = ~a[38] & w11669;
assign w11672 = ~w11670 & ~w11671;
assign w11673 = w11662 & w11672;
assign w11674 = ~w11662 & ~w11672;
assign w11675 = ~w11673 & ~w11674;
assign w11676 = ~w11287 & ~w11291;
assign w11677 = w11675 & w11676;
assign w11678 = ~w11675 & ~w11676;
assign w11679 = ~w11677 & ~w11678;
assign w11680 = w11528 & ~w11679;
assign w11681 = ~w11528 & w11679;
assign w11682 = ~w11680 & ~w11681;
assign w11683 = w11518 & w11682;
assign w11684 = ~w11518 & ~w11682;
assign w11685 = ~w11683 & ~w11684;
assign w11686 = w11517 & w11685;
assign w11687 = ~w11517 & ~w11685;
assign w11688 = ~w11686 & ~w11687;
assign w11689 = (~w11300 & w11118) | (~w11300 & w24696) | (w11118 & w24696);
assign w11690 = ~w11688 & w11689;
assign w11691 = w11688 & ~w11689;
assign w11692 = ~w11690 & ~w11691;
assign w11693 = w11507 & w11692;
assign w11694 = ~w11507 & ~w11692;
assign w11695 = ~w11693 & ~w11694;
assign w11696 = (~w11306 & w11309) | (~w11306 & w25188) | (w11309 & w25188);
assign w11697 = w11695 & w11696;
assign w11698 = ~w11695 & ~w11696;
assign w11699 = ~w11697 & ~w11698;
assign w11700 = w11497 & ~w11699;
assign w11701 = ~w11497 & w11699;
assign w11702 = ~w11700 & ~w11701;
assign w11703 = w11487 & ~w11702;
assign w11704 = ~w11487 & w11702;
assign w11705 = ~w11703 & ~w11704;
assign w11706 = ~w11486 & ~w11705;
assign w11707 = w11486 & w11705;
assign w11708 = ~w11706 & ~w11707;
assign w11709 = w11476 & w11708;
assign w11710 = ~w11476 & ~w11708;
assign w11711 = ~w11709 & ~w11710;
assign w11712 = w11475 & ~w11711;
assign w11713 = ~w11475 & w11711;
assign w11714 = ~w11712 & ~w11713;
assign w11715 = (~w11347 & w11097) | (~w11347 & w24397) | (w11097 & w24397);
assign w11716 = w11714 & ~w11715;
assign w11717 = ~w11714 & w11715;
assign w11718 = ~w11716 & ~w11717;
assign w11719 = b[45] & ~w934;
assign w11720 = b[46] & w838;
assign w11721 = b[47] & w834;
assign w11722 = w832 & w6889;
assign w11723 = ~w11719 & ~w11720;
assign w11724 = ~w11721 & w11723;
assign w11725 = ~w11722 & w11724;
assign w11726 = a[17] & ~w11725;
assign w11727 = ~a[17] & w11725;
assign w11728 = ~w11726 & ~w11727;
assign w11729 = w11718 & w11728;
assign w11730 = ~w11718 & ~w11728;
assign w11731 = ~w11729 & ~w11730;
assign w11732 = w11465 & w11731;
assign w11733 = ~w11465 & ~w11731;
assign w11734 = ~w11732 & ~w11733;
assign w11735 = w11464 & ~w11734;
assign w11736 = ~w11464 & w11734;
assign w11737 = ~w11735 & ~w11736;
assign w11738 = ~w11360 & ~w11363;
assign w11739 = w11737 & w11738;
assign w11740 = ~w11737 & ~w11738;
assign w11741 = ~w11739 & ~w11740;
assign w11742 = w11454 & w11741;
assign w11743 = ~w11454 & ~w11741;
assign w11744 = ~w11742 & ~w11743;
assign w11745 = ~w11444 & w11744;
assign w11746 = w11444 & ~w11744;
assign w11747 = ~w11745 & ~w11746;
assign w11748 = ~w11443 & ~w11747;
assign w11749 = w11443 & w11747;
assign w11750 = ~w11748 & ~w11749;
assign w11751 = (~w11383 & ~w11385) | (~w11383 & w25301) | (~w11385 & w25301);
assign w11752 = w11750 & w11751;
assign w11753 = ~w11750 & ~w11751;
assign w11754 = ~w11752 & ~w11753;
assign w11755 = b[62] & w11;
assign w11756 = b[61] & w9;
assign w11757 = (w11029 & w25302) | (w11029 & w25303) | (w25302 & w25303);
assign w11758 = ~b[61] & ~b[62];
assign w11759 = b[61] & b[62];
assign w11760 = ~w11758 & ~w11759;
assign w11761 = ~w11757 & w11760;
assign w11762 = w11757 & ~w11760;
assign w11763 = ~w11761 & ~w11762;
assign w11764 = w5 & w11763;
assign w11765 = ~w11755 & ~w11756;
assign w11766 = ~w11764 & w11765;
assign w11767 = b[60] & w24;
assign w11768 = a[2] & ~w11767;
assign w11769 = w11766 & ~w11768;
assign w11770 = a[2] & ~w11766;
assign w11771 = ~w11769 & ~w11770;
assign w11772 = ~w11754 & ~w11771;
assign w11773 = w11754 & w11771;
assign w11774 = ~w11772 & ~w11773;
assign w11775 = (~w11389 & ~w11391) | (~w11389 & w24698) | (~w11391 & w24698);
assign w11776 = w11774 & ~w11775;
assign w11777 = ~w11774 & w11775;
assign w11778 = ~w11776 & ~w11777;
assign w11779 = ~w11412 & ~w11416;
assign w11780 = ~w11416 & w24398;
assign w11781 = ~w11778 & ~w11779;
assign w11782 = ~w11780 & ~w11781;
assign w11783 = (~w11776 & w11416) | (~w11776 & w24849) | (w11416 & w24849);
assign w11784 = b[58] & w103;
assign w11785 = b[59] & w61;
assign w11786 = b[60] & w68;
assign w11787 = w66 & w11035;
assign w11788 = ~w11785 & ~w11786;
assign w11789 = ~w11784 & w11788;
assign w11790 = ~w11787 & w11789;
assign w11791 = a[5] & ~w11790;
assign w11792 = ~a[5] & w11790;
assign w11793 = ~w11791 & ~w11792;
assign w11794 = b[56] & w183;
assign w11795 = b[55] & ~w237;
assign w11796 = b[57] & w185;
assign w11797 = w179 & ~w9992;
assign w11798 = ~w11794 & ~w11795;
assign w11799 = ~w11796 & w11798;
assign w11800 = ~w11797 & w11799;
assign w11801 = a[8] & ~w11800;
assign w11802 = ~a[8] & w11800;
assign w11803 = ~w11801 & ~w11802;
assign w11804 = b[52] & ~w419;
assign w11805 = b[53] & w358;
assign w11806 = b[54] & w360;
assign w11807 = w354 & ~w8998;
assign w11808 = ~w11804 & ~w11805;
assign w11809 = ~w11806 & w11808;
assign w11810 = ~w11807 & w11809;
assign w11811 = a[11] & ~w11810;
assign w11812 = ~a[11] & w11810;
assign w11813 = ~w11811 & ~w11812;
assign w11814 = b[46] & ~w934;
assign w11815 = b[47] & w838;
assign w11816 = b[48] & w834;
assign w11817 = w832 & ~w7170;
assign w11818 = ~w11814 & ~w11815;
assign w11819 = ~w11816 & w11818;
assign w11820 = ~w11817 & w11819;
assign w11821 = a[17] & ~w11820;
assign w11822 = ~a[17] & w11820;
assign w11823 = ~w11821 & ~w11822;
assign w11824 = ~w11712 & ~w11716;
assign w11825 = b[43] & ~w1272;
assign w11826 = b[44] & w1154;
assign w11827 = b[45] & w1156;
assign w11828 = w1150 & w6334;
assign w11829 = ~w11825 & ~w11826;
assign w11830 = ~w11827 & w11829;
assign w11831 = ~w11828 & w11830;
assign w11832 = a[20] & ~w11831;
assign w11833 = ~a[20] & w11831;
assign w11834 = ~w11832 & ~w11833;
assign w11835 = b[41] & w1517;
assign w11836 = b[42] & w1519;
assign w11837 = b[40] & ~w1676;
assign w11838 = w1513 & w5548;
assign w11839 = ~w11835 & ~w11836;
assign w11840 = ~w11837 & w11839;
assign w11841 = ~w11838 & w11840;
assign w11842 = a[23] & ~w11841;
assign w11843 = ~a[23] & w11841;
assign w11844 = ~w11842 & ~w11843;
assign w11845 = (~w11700 & w11487) | (~w11700 & w25189) | (w11487 & w25189);
assign w11846 = b[35] & w2436;
assign w11847 = b[36] & w2438;
assign w11848 = b[34] & ~w2622;
assign w11849 = w2432 & w4129;
assign w11850 = ~w11846 & ~w11847;
assign w11851 = ~w11848 & w11850;
assign w11852 = ~w11849 & w11851;
assign w11853 = a[29] & ~w11852;
assign w11854 = ~a[29] & w11852;
assign w11855 = ~w11853 & ~w11854;
assign w11856 = b[28] & w3785;
assign w11857 = b[29] & w3578;
assign w11858 = b[30] & w3580;
assign w11859 = ~w2908 & w3573;
assign w11860 = ~w11857 & ~w11858;
assign w11861 = ~w11856 & w11860;
assign w11862 = ~w11859 & w11861;
assign w11863 = a[35] & ~w11862;
assign w11864 = ~a[35] & w11862;
assign w11865 = ~w11863 & ~w11864;
assign w11866 = b[25] & w4453;
assign w11867 = b[27] & w4243;
assign w11868 = b[26] & w4241;
assign w11869 = w2378 & w4236;
assign w11870 = ~w11867 & ~w11868;
assign w11871 = ~w11866 & w11870;
assign w11872 = ~w11869 & w11871;
assign w11873 = a[38] & ~w11872;
assign w11874 = ~a[38] & w11872;
assign w11875 = ~w11873 & ~w11874;
assign w11876 = (~w11640 & ~w11643) | (~w11640 & w25190) | (~w11643 & w25190);
assign w11877 = b[19] & w5939;
assign w11878 = b[20] & w5670;
assign w11879 = b[21] & w5665;
assign w11880 = w1467 & w5663;
assign w11881 = ~w11878 & ~w11879;
assign w11882 = ~w11877 & w11881;
assign w11883 = ~w11880 & w11882;
assign w11884 = a[44] & ~w11883;
assign w11885 = ~a[44] & w11883;
assign w11886 = ~w11884 & ~w11885;
assign w11887 = (~w11635 & w11540) | (~w11635 & w25304) | (w11540 & w25304);
assign w11888 = b[16] & w6732;
assign w11889 = b[17] & w6474;
assign w11890 = b[18] & w6476;
assign w11891 = ~w1108 & w6469;
assign w11892 = ~w11889 & ~w11890;
assign w11893 = ~w11888 & w11892;
assign w11894 = ~w11891 & w11893;
assign w11895 = a[47] & ~w11894;
assign w11896 = ~a[47] & w11894;
assign w11897 = ~w11895 & ~w11896;
assign w11898 = ~w11602 & ~w11604;
assign w11899 = b[10] & w8515;
assign w11900 = b[12] & w8202;
assign w11901 = b[11] & w8200;
assign w11902 = w536 & w8195;
assign w11903 = ~w11900 & ~w11901;
assign w11904 = ~w11899 & w11903;
assign w11905 = ~w11902 & w11904;
assign w11906 = a[53] & ~w11905;
assign w11907 = ~a[53] & w11905;
assign w11908 = ~w11906 & ~w11907;
assign w11909 = ~w11585 & ~w11588;
assign w11910 = b[1] & w11561;
assign w11911 = b[2] & w11194;
assign w11912 = b[3] & w11196;
assign w11913 = w46 & w11189;
assign w11914 = ~w11911 & ~w11912;
assign w11915 = ~w11910 & w11914;
assign w11916 = ~w11913 & w11915;
assign w11917 = a[62] & ~w11916;
assign w11918 = ~a[62] & w11916;
assign w11919 = ~w11917 & ~w11918;
assign w11920 = w11555 & w11565;
assign w11921 = a[62] & a[63];
assign w11922 = ~a[62] & ~a[63];
assign w11923 = ~w11921 & ~w11922;
assign w11924 = b[0] & w11923;
assign w11925 = w11920 & w11924;
assign w11926 = ~w11920 & ~w11924;
assign w11927 = ~w11925 & ~w11926;
assign w11928 = w11919 & w11927;
assign w11929 = ~w11919 & ~w11927;
assign w11930 = ~w11928 & ~w11929;
assign w11931 = b[4] & w10496;
assign w11932 = b[6] & w10148;
assign w11933 = b[5] & w10146;
assign w11934 = w157 & w10141;
assign w11935 = ~w11932 & ~w11933;
assign w11936 = ~w11931 & w11935;
assign w11937 = ~w11934 & w11936;
assign w11938 = a[59] & ~w11937;
assign w11939 = ~a[59] & w11937;
assign w11940 = ~w11938 & ~w11939;
assign w11941 = w11930 & w11940;
assign w11942 = ~w11930 & ~w11940;
assign w11943 = ~w11941 & ~w11942;
assign w11944 = ~w11569 & ~w11572;
assign w11945 = w11943 & w11944;
assign w11946 = ~w11943 & ~w11944;
assign w11947 = ~w11945 & ~w11946;
assign w11948 = b[7] & w9482;
assign w11949 = b[8] & w9165;
assign w11950 = b[9] & w9160;
assign w11951 = w322 & w9158;
assign w11952 = ~w11949 & ~w11950;
assign w11953 = ~w11948 & w11952;
assign w11954 = ~w11951 & w11953;
assign w11955 = a[56] & ~w11954;
assign w11956 = ~a[56] & w11954;
assign w11957 = ~w11955 & ~w11956;
assign w11958 = w11947 & w11957;
assign w11959 = ~w11947 & ~w11957;
assign w11960 = ~w11958 & ~w11959;
assign w11961 = ~w11909 & w11960;
assign w11962 = w11909 & ~w11960;
assign w11963 = ~w11961 & ~w11962;
assign w11964 = w11908 & w11963;
assign w11965 = ~w11908 & ~w11963;
assign w11966 = ~w11964 & ~w11965;
assign w11967 = w11898 & ~w11966;
assign w11968 = ~w11898 & w11966;
assign w11969 = ~w11967 & ~w11968;
assign w11970 = b[13] & w7586;
assign w11971 = b[15] & w7314;
assign w11972 = b[14] & w7307;
assign w11973 = ~w799 & w7312;
assign w11974 = ~w11971 & ~w11972;
assign w11975 = ~w11970 & w11974;
assign w11976 = ~w11973 & w11975;
assign w11977 = a[50] & ~w11976;
assign w11978 = ~a[50] & w11976;
assign w11979 = ~w11977 & ~w11978;
assign w11980 = w11969 & w11979;
assign w11981 = ~w11969 & ~w11979;
assign w11982 = ~w11980 & ~w11981;
assign w11983 = (~w11617 & ~w11620) | (~w11617 & w24850) | (~w11620 & w24850);
assign w11984 = w11982 & ~w11983;
assign w11985 = ~w11982 & w11983;
assign w11986 = ~w11984 & ~w11985;
assign w11987 = w11897 & w11986;
assign w11988 = ~w11897 & ~w11986;
assign w11989 = ~w11987 & ~w11988;
assign w11990 = w11887 & ~w11989;
assign w11991 = ~w11887 & w11989;
assign w11992 = ~w11990 & ~w11991;
assign w11993 = ~w11886 & ~w11992;
assign w11994 = w11886 & w11992;
assign w11995 = ~w11993 & ~w11994;
assign w11996 = w11876 & ~w11995;
assign w11997 = ~w11876 & w11995;
assign w11998 = ~w11996 & ~w11997;
assign w11999 = b[22] & w5167;
assign w12000 = b[23] & w4918;
assign w12001 = b[24] & w4925;
assign w12002 = w1895 & w4923;
assign w12003 = ~w12000 & ~w12001;
assign w12004 = ~w11999 & w12003;
assign w12005 = ~w12002 & w12004;
assign w12006 = a[41] & ~w12005;
assign w12007 = ~a[41] & w12005;
assign w12008 = ~w12006 & ~w12007;
assign w12009 = w11998 & w12008;
assign w12010 = ~w11998 & ~w12008;
assign w12011 = ~w12009 & ~w12010;
assign w12012 = (~w11657 & w11529) | (~w11657 & w24699) | (w11529 & w24699);
assign w12013 = w12011 & ~w12012;
assign w12014 = ~w12011 & w12012;
assign w12015 = ~w12013 & ~w12014;
assign w12016 = w11875 & w12015;
assign w12017 = ~w11875 & ~w12015;
assign w12018 = ~w12016 & ~w12017;
assign w12019 = (~w11674 & ~w11676) | (~w11674 & w25191) | (~w11676 & w25191);
assign w12020 = w12018 & w12019;
assign w12021 = ~w12018 & ~w12019;
assign w12022 = ~w12020 & ~w12021;
assign w12023 = ~w11865 & ~w12022;
assign w12024 = w11865 & w12022;
assign w12025 = ~w12023 & ~w12024;
assign w12026 = ~w11680 & ~w11683;
assign w12027 = w12025 & ~w12026;
assign w12028 = ~w12025 & w12026;
assign w12029 = ~w12027 & ~w12028;
assign w12030 = b[31] & w3177;
assign w12031 = b[32] & w2973;
assign w12032 = b[33] & w2978;
assign w12033 = w2980 & w3499;
assign w12034 = ~w12031 & ~w12032;
assign w12035 = ~w12030 & w12034;
assign w12036 = ~w12033 & w12035;
assign w12037 = a[32] & ~w12036;
assign w12038 = ~a[32] & w12036;
assign w12039 = ~w12037 & ~w12038;
assign w12040 = w12029 & w12039;
assign w12041 = ~w12029 & ~w12039;
assign w12042 = ~w12040 & ~w12041;
assign w12043 = ~w11686 & ~w11691;
assign w12044 = w12042 & ~w12043;
assign w12045 = ~w12042 & w12043;
assign w12046 = ~w12044 & ~w12045;
assign w12047 = w11855 & w12046;
assign w12048 = ~w11855 & ~w12046;
assign w12049 = ~w12047 & ~w12048;
assign w12050 = (~w11694 & ~w11696) | (~w11694 & w24700) | (~w11696 & w24700);
assign w12051 = ~w12049 & ~w12050;
assign w12052 = w12049 & w12050;
assign w12053 = ~w12051 & ~w12052;
assign w12054 = b[38] & w1955;
assign w12055 = b[39] & w1957;
assign w12056 = b[37] & ~w2114;
assign w12057 = w1951 & ~w4812;
assign w12058 = ~w12054 & ~w12055;
assign w12059 = ~w12056 & w12058;
assign w12060 = ~w12057 & w12059;
assign w12061 = a[26] & ~w12060;
assign w12062 = ~a[26] & w12060;
assign w12063 = ~w12061 & ~w12062;
assign w12064 = ~w12053 & ~w12063;
assign w12065 = w12053 & w12063;
assign w12066 = ~w12064 & ~w12065;
assign w12067 = ~w11845 & w12066;
assign w12068 = w11845 & ~w12066;
assign w12069 = ~w12067 & ~w12068;
assign w12070 = ~w11844 & ~w12069;
assign w12071 = w11844 & w12069;
assign w12072 = ~w12070 & ~w12071;
assign w12073 = (~w11706 & ~w11476) | (~w11706 & w25555) | (~w11476 & w25555);
assign w12074 = w12072 & w12073;
assign w12075 = ~w12072 & ~w12073;
assign w12076 = ~w12074 & ~w12075;
assign w12077 = ~w11834 & ~w12076;
assign w12078 = w11834 & w12076;
assign w12079 = ~w12077 & ~w12078;
assign w12080 = ~w11824 & w12079;
assign w12081 = w11824 & ~w12079;
assign w12082 = ~w12080 & ~w12081;
assign w12083 = ~w11823 & ~w12082;
assign w12084 = w11823 & w12082;
assign w12085 = ~w12083 & ~w12084;
assign w12086 = (~w11730 & ~w11465) | (~w11730 & w24399) | (~w11465 & w24399);
assign w12087 = w12085 & w12086;
assign w12088 = ~w12085 & ~w12086;
assign w12089 = ~w12087 & ~w12088;
assign w12090 = b[50] & w573;
assign w12091 = b[51] & w575;
assign w12092 = b[49] & ~w649;
assign w12093 = w569 & ~w8058;
assign w12094 = ~w12090 & ~w12091;
assign w12095 = ~w12092 & w12094;
assign w12096 = ~w12093 & w12095;
assign w12097 = a[14] & ~w12096;
assign w12098 = ~a[14] & w12096;
assign w12099 = ~w12097 & ~w12098;
assign w12100 = w12089 & w12099;
assign w12101 = ~w12089 & ~w12099;
assign w12102 = ~w12100 & ~w12101;
assign w12103 = ~w11735 & ~w11739;
assign w12104 = w12102 & ~w12103;
assign w12105 = ~w12102 & w12103;
assign w12106 = ~w12104 & ~w12105;
assign w12107 = w11813 & w12106;
assign w12108 = ~w11813 & ~w12106;
assign w12109 = ~w12107 & ~w12108;
assign w12110 = ~w11742 & ~w11745;
assign w12111 = ~w12109 & ~w12110;
assign w12112 = w12109 & w12110;
assign w12113 = ~w12111 & ~w12112;
assign w12114 = ~w11803 & w12113;
assign w12115 = w11803 & ~w12113;
assign w12116 = ~w12114 & ~w12115;
assign w12117 = w11793 & w12116;
assign w12118 = ~w11793 & ~w12116;
assign w12119 = ~w12117 & ~w12118;
assign w12120 = ~w11441 & ~w11749;
assign w12121 = w12119 & ~w12120;
assign w12122 = ~w12119 & w12120;
assign w12123 = ~w12121 & ~w12122;
assign w12124 = b[63] & w11;
assign w12125 = b[62] & w9;
assign w12126 = (~w11759 & w11757) | (~w11759 & w24851) | (w11757 & w24851);
assign w12127 = ~b[62] & ~b[63];
assign w12128 = b[62] & b[63];
assign w12129 = ~w12127 & ~w12128;
assign w12130 = w12126 & ~w12129;
assign w12131 = ~w12126 & w12129;
assign w12132 = ~w12130 & ~w12131;
assign w12133 = w5 & w12132;
assign w12134 = ~w12124 & ~w12125;
assign w12135 = ~w12133 & w12134;
assign w12136 = b[61] & w24;
assign w12137 = a[2] & ~w12136;
assign w12138 = w12135 & ~w12137;
assign w12139 = a[2] & ~w12135;
assign w12140 = ~w12138 & ~w12139;
assign w12141 = w12123 & w12140;
assign w12142 = ~w12123 & ~w12140;
assign w12143 = ~w12141 & ~w12142;
assign w12144 = ~w11752 & ~w11773;
assign w12145 = w12143 & ~w12144;
assign w12146 = ~w12143 & w12144;
assign w12147 = ~w12145 & ~w12146;
assign w12148 = w11783 & w12147;
assign w12149 = ~w11783 & ~w12147;
assign w12150 = ~w12148 & ~w12149;
assign w12151 = (~w12121 & ~w12123) | (~w12121 & w24701) | (~w12123 & w24701);
assign w12152 = (~w12115 & ~w12116) | (~w12115 & w24702) | (~w12116 & w24702);
assign w12153 = ~b[63] & ~w12131;
assign w12154 = (~b[62] & w11757) | (~b[62] & w24852) | (w11757 & w24852);
assign w12155 = b[63] & ~w12154;
assign w12156 = ~w12153 & ~w12155;
assign w12157 = w5 & w12156;
assign w12158 = b[63] & w9;
assign w12159 = ~w12157 & ~w12158;
assign w12160 = b[62] & w24;
assign w12161 = a[2] & ~w12160;
assign w12162 = w12159 & ~w12161;
assign w12163 = a[2] & ~w12159;
assign w12164 = ~w12162 & ~w12163;
assign w12165 = ~w12152 & w12164;
assign w12166 = w12152 & ~w12164;
assign w12167 = ~w12165 & ~w12166;
assign w12168 = b[59] & w103;
assign w12169 = b[61] & w68;
assign w12170 = b[60] & w61;
assign w12171 = w66 & w11400;
assign w12172 = ~w12169 & ~w12170;
assign w12173 = ~w12168 & w12172;
assign w12174 = ~w12171 & w12173;
assign w12175 = a[5] & ~w12174;
assign w12176 = ~a[5] & w12174;
assign w12177 = ~w12175 & ~w12176;
assign w12178 = b[57] & w183;
assign w12179 = b[56] & ~w237;
assign w12180 = b[58] & w185;
assign w12181 = w179 & ~w10339;
assign w12182 = ~w12178 & ~w12179;
assign w12183 = ~w12180 & w12182;
assign w12184 = ~w12181 & w12183;
assign w12185 = a[8] & ~w12184;
assign w12186 = ~a[8] & w12184;
assign w12187 = ~w12185 & ~w12186;
assign w12188 = b[54] & w358;
assign w12189 = b[55] & w360;
assign w12190 = b[53] & ~w419;
assign w12191 = w354 & ~w9330;
assign w12192 = ~w12188 & ~w12189;
assign w12193 = ~w12190 & w12192;
assign w12194 = ~w12191 & w12193;
assign w12195 = a[11] & ~w12194;
assign w12196 = ~a[11] & w12194;
assign w12197 = ~w12195 & ~w12196;
assign w12198 = b[51] & w573;
assign w12199 = b[52] & w575;
assign w12200 = b[50] & ~w649;
assign w12201 = w569 & ~w8371;
assign w12202 = ~w12198 & ~w12199;
assign w12203 = ~w12200 & w12202;
assign w12204 = ~w12201 & w12203;
assign w12205 = a[14] & ~w12204;
assign w12206 = ~a[14] & w12204;
assign w12207 = ~w12205 & ~w12206;
assign w12208 = ~w12084 & ~w12087;
assign w12209 = b[47] & ~w934;
assign w12210 = b[48] & w838;
assign w12211 = b[49] & w834;
assign w12212 = w832 & ~w7468;
assign w12213 = ~w12209 & ~w12210;
assign w12214 = ~w12211 & w12213;
assign w12215 = ~w12212 & w12214;
assign w12216 = a[17] & ~w12215;
assign w12217 = ~a[17] & w12215;
assign w12218 = ~w12216 & ~w12217;
assign w12219 = (~w12078 & w11824) | (~w12078 & w25556) | (w11824 & w25556);
assign w12220 = b[45] & w1154;
assign w12221 = b[44] & ~w1272;
assign w12222 = b[46] & w1156;
assign w12223 = w1150 & ~w6613;
assign w12224 = ~w12220 & ~w12221;
assign w12225 = ~w12222 & w12224;
assign w12226 = ~w12223 & w12225;
assign w12227 = a[20] & ~w12226;
assign w12228 = ~a[20] & w12226;
assign w12229 = ~w12227 & ~w12228;
assign w12230 = (~w12071 & ~w12073) | (~w12071 & w25192) | (~w12073 & w25192);
assign w12231 = b[43] & w1519;
assign w12232 = b[41] & ~w1676;
assign w12233 = b[42] & w1517;
assign w12234 = w1513 & w5811;
assign w12235 = ~w12231 & ~w12232;
assign w12236 = ~w12233 & w12235;
assign w12237 = ~w12234 & w12236;
assign w12238 = a[23] & ~w12237;
assign w12239 = ~a[23] & w12237;
assign w12240 = ~w12238 & ~w12239;
assign w12241 = b[39] & w1955;
assign w12242 = b[40] & w1957;
assign w12243 = b[38] & ~w2114;
assign w12244 = w1951 & ~w5058;
assign w12245 = ~w12241 & ~w12242;
assign w12246 = ~w12243 & w12245;
assign w12247 = ~w12244 & w12246;
assign w12248 = a[26] & ~w12247;
assign w12249 = ~a[26] & w12247;
assign w12250 = ~w12248 & ~w12249;
assign w12251 = b[35] & ~w2622;
assign w12252 = b[36] & w2436;
assign w12253 = b[37] & w2438;
assign w12254 = w2432 & ~w4357;
assign w12255 = ~w12251 & ~w12252;
assign w12256 = ~w12253 & w12255;
assign w12257 = ~w12254 & w12256;
assign w12258 = a[29] & ~w12257;
assign w12259 = ~a[29] & w12257;
assign w12260 = ~w12258 & ~w12259;
assign w12261 = b[29] & w3785;
assign w12262 = b[31] & w3580;
assign w12263 = b[30] & w3578;
assign w12264 = ~w3112 & w3573;
assign w12265 = ~w12262 & ~w12263;
assign w12266 = ~w12261 & w12265;
assign w12267 = ~w12264 & w12266;
assign w12268 = a[35] & ~w12267;
assign w12269 = ~a[35] & w12267;
assign w12270 = ~w12268 & ~w12269;
assign w12271 = b[26] & w4453;
assign w12272 = b[27] & w4241;
assign w12273 = b[28] & w4243;
assign w12274 = w2559 & w4236;
assign w12275 = ~w12272 & ~w12273;
assign w12276 = ~w12271 & w12275;
assign w12277 = ~w12274 & w12276;
assign w12278 = a[38] & ~w12277;
assign w12279 = ~a[38] & w12277;
assign w12280 = ~w12278 & ~w12279;
assign w12281 = b[23] & w5167;
assign w12282 = b[24] & w4918;
assign w12283 = b[25] & w4925;
assign w12284 = w2061 & w4923;
assign w12285 = ~w12282 & ~w12283;
assign w12286 = ~w12281 & w12285;
assign w12287 = ~w12284 & w12286;
assign w12288 = a[41] & ~w12287;
assign w12289 = ~a[41] & w12287;
assign w12290 = ~w12288 & ~w12289;
assign w12291 = b[17] & w6732;
assign w12292 = b[19] & w6476;
assign w12293 = b[18] & w6474;
assign w12294 = ~w1231 & w6469;
assign w12295 = ~w12292 & ~w12293;
assign w12296 = ~w12291 & w12295;
assign w12297 = ~w12294 & w12296;
assign w12298 = a[47] & ~w12297;
assign w12299 = ~a[47] & w12297;
assign w12300 = ~w12298 & ~w12299;
assign w12301 = b[11] & w8515;
assign w12302 = b[13] & w8202;
assign w12303 = b[12] & w8200;
assign w12304 = w628 & w8195;
assign w12305 = ~w12302 & ~w12303;
assign w12306 = ~w12301 & w12305;
assign w12307 = ~w12304 & w12306;
assign w12308 = a[53] & ~w12307;
assign w12309 = ~a[53] & w12307;
assign w12310 = ~w12308 & ~w12309;
assign w12311 = ~w11941 & ~w11945;
assign w12312 = ~w11925 & ~w11928;
assign w12313 = b[0] & w11921;
assign w12314 = b[1] & w11923;
assign w12315 = ~w12313 & ~w12314;
assign w12316 = b[2] & w11561;
assign w12317 = b[3] & w11194;
assign w12318 = b[4] & w11196;
assign w12319 = w84 & w11189;
assign w12320 = ~w12317 & ~w12318;
assign w12321 = ~w12316 & w12320;
assign w12322 = ~w12319 & w12321;
assign w12323 = a[62] & ~w12322;
assign w12324 = ~a[62] & w12322;
assign w12325 = ~w12323 & ~w12324;
assign w12326 = ~w12315 & w12325;
assign w12327 = w12315 & ~w12325;
assign w12328 = ~w12326 & ~w12327;
assign w12329 = w12312 & ~w12328;
assign w12330 = ~w12312 & w12328;
assign w12331 = ~w12329 & ~w12330;
assign w12332 = b[5] & w10496;
assign w12333 = b[7] & w10148;
assign w12334 = b[6] & w10146;
assign w12335 = w216 & w10141;
assign w12336 = ~w12333 & ~w12334;
assign w12337 = ~w12332 & w12336;
assign w12338 = ~w12335 & w12337;
assign w12339 = a[59] & ~w12338;
assign w12340 = ~a[59] & w12338;
assign w12341 = ~w12339 & ~w12340;
assign w12342 = w12331 & w12341;
assign w12343 = ~w12331 & ~w12341;
assign w12344 = ~w12342 & ~w12343;
assign w12345 = ~w12311 & w12344;
assign w12346 = w12311 & ~w12344;
assign w12347 = ~w12345 & ~w12346;
assign w12348 = b[8] & w9482;
assign w12349 = b[9] & w9165;
assign w12350 = b[10] & w9160;
assign w12351 = w397 & w9158;
assign w12352 = ~w12349 & ~w12350;
assign w12353 = ~w12348 & w12352;
assign w12354 = ~w12351 & w12353;
assign w12355 = a[56] & ~w12354;
assign w12356 = ~a[56] & w12354;
assign w12357 = ~w12355 & ~w12356;
assign w12358 = w12347 & w12357;
assign w12359 = ~w12347 & ~w12357;
assign w12360 = ~w12358 & ~w12359;
assign w12361 = ~w11958 & ~w11961;
assign w12362 = w12360 & ~w12361;
assign w12363 = ~w12360 & w12361;
assign w12364 = ~w12362 & ~w12363;
assign w12365 = w12310 & w12364;
assign w12366 = ~w12310 & ~w12364;
assign w12367 = ~w12365 & ~w12366;
assign w12368 = ~w11964 & ~w11968;
assign w12369 = w12367 & ~w12368;
assign w12370 = ~w12367 & w12368;
assign w12371 = ~w12369 & ~w12370;
assign w12372 = b[14] & w7586;
assign w12373 = b[15] & w7307;
assign w12374 = b[16] & w7314;
assign w12375 = w905 & w7312;
assign w12376 = ~w12373 & ~w12374;
assign w12377 = ~w12372 & w12376;
assign w12378 = ~w12375 & w12377;
assign w12379 = a[50] & ~w12378;
assign w12380 = ~a[50] & w12378;
assign w12381 = ~w12379 & ~w12380;
assign w12382 = w12371 & w12381;
assign w12383 = ~w12371 & ~w12381;
assign w12384 = ~w12382 & ~w12383;
assign w12385 = ~w11980 & ~w11984;
assign w12386 = w12384 & ~w12385;
assign w12387 = ~w12384 & w12385;
assign w12388 = ~w12386 & ~w12387;
assign w12389 = w12300 & w12388;
assign w12390 = ~w12300 & ~w12388;
assign w12391 = ~w12389 & ~w12390;
assign w12392 = (~w11987 & w11887) | (~w11987 & w24853) | (w11887 & w24853);
assign w12393 = w12391 & ~w12392;
assign w12394 = ~w12391 & w12392;
assign w12395 = ~w12393 & ~w12394;
assign w12396 = b[20] & w5939;
assign w12397 = b[21] & w5670;
assign w12398 = b[22] & w5665;
assign w12399 = w1615 & w5663;
assign w12400 = ~w12397 & ~w12398;
assign w12401 = ~w12396 & w12400;
assign w12402 = ~w12399 & w12401;
assign w12403 = a[44] & ~w12402;
assign w12404 = ~a[44] & w12402;
assign w12405 = ~w12403 & ~w12404;
assign w12406 = w12395 & w12405;
assign w12407 = ~w12395 & ~w12405;
assign w12408 = ~w12406 & ~w12407;
assign w12409 = (~w11994 & w11876) | (~w11994 & w25305) | (w11876 & w25305);
assign w12410 = w12408 & ~w12409;
assign w12411 = ~w12408 & w12409;
assign w12412 = ~w12410 & ~w12411;
assign w12413 = w12290 & w12412;
assign w12414 = ~w12290 & ~w12412;
assign w12415 = ~w12413 & ~w12414;
assign w12416 = (~w12009 & w12012) | (~w12009 & w25193) | (w12012 & w25193);
assign w12417 = w12415 & ~w12416;
assign w12418 = ~w12415 & w12416;
assign w12419 = ~w12417 & ~w12418;
assign w12420 = w12280 & w12419;
assign w12421 = ~w12280 & ~w12419;
assign w12422 = ~w12420 & ~w12421;
assign w12423 = (~w12016 & ~w12019) | (~w12016 & w24703) | (~w12019 & w24703);
assign w12424 = w12422 & ~w12423;
assign w12425 = ~w12422 & w12423;
assign w12426 = ~w12424 & ~w12425;
assign w12427 = ~w12270 & ~w12426;
assign w12428 = w12270 & w12426;
assign w12429 = ~w12427 & ~w12428;
assign w12430 = (~w12024 & w12026) | (~w12024 & w25194) | (w12026 & w25194);
assign w12431 = w12429 & ~w12430;
assign w12432 = ~w12429 & w12430;
assign w12433 = ~w12431 & ~w12432;
assign w12434 = b[32] & w3177;
assign w12435 = b[34] & w2978;
assign w12436 = b[33] & w2973;
assign w12437 = w2980 & ~w3710;
assign w12438 = ~w12435 & ~w12436;
assign w12439 = ~w12434 & w12438;
assign w12440 = ~w12437 & w12439;
assign w12441 = a[32] & ~w12440;
assign w12442 = ~a[32] & w12440;
assign w12443 = ~w12441 & ~w12442;
assign w12444 = w12433 & w12443;
assign w12445 = ~w12433 & ~w12443;
assign w12446 = ~w12444 & ~w12445;
assign w12447 = ~w12040 & ~w12044;
assign w12448 = w12446 & ~w12447;
assign w12449 = ~w12446 & w12447;
assign w12450 = ~w12448 & ~w12449;
assign w12451 = w12260 & w12450;
assign w12452 = ~w12260 & ~w12450;
assign w12453 = ~w12451 & ~w12452;
assign w12454 = ~w12047 & ~w12052;
assign w12455 = w12453 & ~w12454;
assign w12456 = ~w12453 & w12454;
assign w12457 = ~w12455 & ~w12456;
assign w12458 = w12250 & w12457;
assign w12459 = ~w12250 & ~w12457;
assign w12460 = ~w12458 & ~w12459;
assign w12461 = (~w12065 & w11845) | (~w12065 & w24854) | (w11845 & w24854);
assign w12462 = w12460 & ~w12461;
assign w12463 = ~w12460 & w12461;
assign w12464 = ~w12462 & ~w12463;
assign w12465 = w12240 & w12464;
assign w12466 = ~w12240 & ~w12464;
assign w12467 = ~w12465 & ~w12466;
assign w12468 = w12230 & w12467;
assign w12469 = ~w12230 & ~w12467;
assign w12470 = ~w12468 & ~w12469;
assign w12471 = w12229 & ~w12470;
assign w12472 = ~w12229 & w12470;
assign w12473 = ~w12471 & ~w12472;
assign w12474 = ~w12219 & w12473;
assign w12475 = w12219 & ~w12473;
assign w12476 = ~w12474 & ~w12475;
assign w12477 = w12218 & w12476;
assign w12478 = ~w12218 & ~w12476;
assign w12479 = ~w12477 & ~w12478;
assign w12480 = w12208 & w12479;
assign w12481 = ~w12208 & ~w12479;
assign w12482 = ~w12480 & ~w12481;
assign w12483 = w12207 & ~w12482;
assign w12484 = ~w12207 & w12482;
assign w12485 = ~w12483 & ~w12484;
assign w12486 = (~w12100 & w12103) | (~w12100 & w24704) | (w12103 & w24704);
assign w12487 = ~w12485 & w12486;
assign w12488 = w12485 & ~w12486;
assign w12489 = ~w12487 & ~w12488;
assign w12490 = w12197 & w12489;
assign w12491 = ~w12197 & ~w12489;
assign w12492 = ~w12490 & ~w12491;
assign w12493 = ~w12108 & ~w12112;
assign w12494 = w12492 & w12493;
assign w12495 = ~w12492 & ~w12493;
assign w12496 = ~w12494 & ~w12495;
assign w12497 = w12187 & w12496;
assign w12498 = ~w12187 & ~w12496;
assign w12499 = ~w12497 & ~w12498;
assign w12500 = ~w12177 & w12499;
assign w12501 = w12177 & ~w12499;
assign w12502 = ~w12500 & ~w12501;
assign w12503 = ~w12167 & ~w12502;
assign w12504 = w12167 & w12502;
assign w12505 = ~w12503 & ~w12504;
assign w12506 = ~w12151 & ~w12505;
assign w12507 = w12151 & w12505;
assign w12508 = ~w12506 & ~w12507;
assign w12509 = (~w12146 & ~w12147) | (~w12146 & w24400) | (~w12147 & w24400);
assign w12510 = ~w12508 & w12509;
assign w12511 = w12508 & ~w12509;
assign w12512 = ~w12510 & ~w12511;
assign w12513 = b[60] & w103;
assign w12514 = b[62] & w68;
assign w12515 = b[61] & w61;
assign w12516 = w66 & w11763;
assign w12517 = ~w12514 & ~w12515;
assign w12518 = ~w12513 & w12517;
assign w12519 = ~w12516 & w12518;
assign w12520 = a[5] & ~w12519;
assign w12521 = ~a[5] & w12519;
assign w12522 = ~w12520 & ~w12521;
assign w12523 = (~w12490 & ~w12493) | (~w12490 & w24705) | (~w12493 & w24705);
assign w12524 = b[48] & ~w934;
assign w12525 = b[49] & w838;
assign w12526 = b[50] & w834;
assign w12527 = w832 & w7759;
assign w12528 = ~w12524 & ~w12525;
assign w12529 = ~w12526 & w12528;
assign w12530 = ~w12527 & w12529;
assign w12531 = a[17] & ~w12530;
assign w12532 = ~a[17] & w12530;
assign w12533 = ~w12531 & ~w12532;
assign w12534 = (~w12471 & w12219) | (~w12471 & w25195) | (w12219 & w25195);
assign w12535 = b[46] & w1154;
assign w12536 = b[45] & ~w1272;
assign w12537 = b[47] & w1156;
assign w12538 = w1150 & w6889;
assign w12539 = ~w12535 & ~w12536;
assign w12540 = ~w12537 & w12539;
assign w12541 = ~w12538 & w12540;
assign w12542 = a[20] & ~w12541;
assign w12543 = ~a[20] & w12541;
assign w12544 = ~w12542 & ~w12543;
assign w12545 = b[44] & w1519;
assign w12546 = b[42] & ~w1676;
assign w12547 = b[43] & w1517;
assign w12548 = w1513 & w6069;
assign w12549 = ~w12545 & ~w12546;
assign w12550 = ~w12547 & w12549;
assign w12551 = ~w12548 & w12550;
assign w12552 = a[23] & ~w12551;
assign w12553 = ~a[23] & w12551;
assign w12554 = ~w12552 & ~w12553;
assign w12555 = ~w12458 & ~w12462;
assign w12556 = (~w12444 & w12447) | (~w12444 & w25306) | (w12447 & w25306);
assign w12557 = b[33] & w3177;
assign w12558 = b[34] & w2973;
assign w12559 = b[35] & w2978;
assign w12560 = w2980 & w3918;
assign w12561 = ~w12558 & ~w12559;
assign w12562 = ~w12557 & w12561;
assign w12563 = ~w12560 & w12562;
assign w12564 = a[32] & ~w12563;
assign w12565 = ~a[32] & w12563;
assign w12566 = ~w12564 & ~w12565;
assign w12567 = (~w12428 & w12430) | (~w12428 & w24855) | (w12430 & w24855);
assign w12568 = (~w12406 & w12409) | (~w12406 & w24856) | (w12409 & w24856);
assign w12569 = b[21] & w5939;
assign w12570 = b[23] & w5665;
assign w12571 = b[22] & w5670;
assign w12572 = w1755 & w5663;
assign w12573 = ~w12570 & ~w12571;
assign w12574 = ~w12569 & w12573;
assign w12575 = ~w12572 & w12574;
assign w12576 = a[44] & ~w12575;
assign w12577 = ~a[44] & w12575;
assign w12578 = ~w12576 & ~w12577;
assign w12579 = ~w12389 & ~w12393;
assign w12580 = ~w12382 & ~w12386;
assign w12581 = b[15] & w7586;
assign w12582 = b[16] & w7307;
assign w12583 = b[17] & w7314;
assign w12584 = w1008 & w7312;
assign w12585 = ~w12582 & ~w12583;
assign w12586 = ~w12581 & w12585;
assign w12587 = ~w12584 & w12586;
assign w12588 = a[50] & ~w12587;
assign w12589 = ~a[50] & w12587;
assign w12590 = ~w12588 & ~w12589;
assign w12591 = ~w12365 & ~w12369;
assign w12592 = ~w12358 & ~w12362;
assign w12593 = ~w12342 & ~w12345;
assign w12594 = ~w12326 & ~w12330;
assign w12595 = b[1] & w11921;
assign w12596 = b[2] & w11923;
assign w12597 = ~w12595 & ~w12596;
assign w12598 = b[3] & w11561;
assign w12599 = b[5] & w11196;
assign w12600 = b[4] & w11194;
assign w12601 = w116 & w11189;
assign w12602 = ~w12599 & ~w12600;
assign w12603 = ~w12598 & w12602;
assign w12604 = ~w12601 & w12603;
assign w12605 = a[62] & ~w12604;
assign w12606 = ~a[62] & w12604;
assign w12607 = ~w12605 & ~w12606;
assign w12608 = ~w12597 & w12607;
assign w12609 = w12597 & ~w12607;
assign w12610 = ~w12608 & ~w12609;
assign w12611 = w12594 & ~w12610;
assign w12612 = ~w12594 & w12610;
assign w12613 = ~w12611 & ~w12612;
assign w12614 = b[6] & w10496;
assign w12615 = b[8] & w10148;
assign w12616 = b[7] & w10146;
assign w12617 = w270 & w10141;
assign w12618 = ~w12615 & ~w12616;
assign w12619 = ~w12614 & w12618;
assign w12620 = ~w12617 & w12619;
assign w12621 = a[59] & ~w12620;
assign w12622 = ~a[59] & w12620;
assign w12623 = ~w12621 & ~w12622;
assign w12624 = ~w12613 & ~w12623;
assign w12625 = w12613 & w12623;
assign w12626 = ~w12624 & ~w12625;
assign w12627 = w12593 & w12626;
assign w12628 = ~w12593 & ~w12626;
assign w12629 = ~w12627 & ~w12628;
assign w12630 = b[9] & w9482;
assign w12631 = b[11] & w9160;
assign w12632 = b[10] & w9165;
assign w12633 = w469 & w9158;
assign w12634 = ~w12631 & ~w12632;
assign w12635 = ~w12630 & w12634;
assign w12636 = ~w12633 & w12635;
assign w12637 = a[56] & ~w12636;
assign w12638 = ~a[56] & w12636;
assign w12639 = ~w12637 & ~w12638;
assign w12640 = ~w12629 & w12639;
assign w12641 = w12629 & ~w12639;
assign w12642 = ~w12640 & ~w12641;
assign w12643 = ~w12592 & w12642;
assign w12644 = w12592 & ~w12642;
assign w12645 = ~w12643 & ~w12644;
assign w12646 = b[12] & w8515;
assign w12647 = b[14] & w8202;
assign w12648 = b[13] & w8200;
assign w12649 = w714 & w8195;
assign w12650 = ~w12647 & ~w12648;
assign w12651 = ~w12646 & w12650;
assign w12652 = ~w12649 & w12651;
assign w12653 = a[53] & ~w12652;
assign w12654 = ~a[53] & w12652;
assign w12655 = ~w12653 & ~w12654;
assign w12656 = w12645 & w12655;
assign w12657 = ~w12645 & ~w12655;
assign w12658 = ~w12656 & ~w12657;
assign w12659 = ~w12591 & w12658;
assign w12660 = w12591 & ~w12658;
assign w12661 = ~w12659 & ~w12660;
assign w12662 = w12590 & w12661;
assign w12663 = ~w12590 & ~w12661;
assign w12664 = ~w12662 & ~w12663;
assign w12665 = w12580 & ~w12664;
assign w12666 = ~w12580 & w12664;
assign w12667 = ~w12665 & ~w12666;
assign w12668 = b[18] & w6732;
assign w12669 = b[20] & w6476;
assign w12670 = b[19] & w6474;
assign w12671 = w1347 & w6469;
assign w12672 = ~w12669 & ~w12670;
assign w12673 = ~w12668 & w12672;
assign w12674 = ~w12671 & w12673;
assign w12675 = a[47] & ~w12674;
assign w12676 = ~a[47] & w12674;
assign w12677 = ~w12675 & ~w12676;
assign w12678 = w12667 & w12677;
assign w12679 = ~w12667 & ~w12677;
assign w12680 = ~w12678 & ~w12679;
assign w12681 = ~w12579 & w12680;
assign w12682 = w12579 & ~w12680;
assign w12683 = ~w12681 & ~w12682;
assign w12684 = w12578 & w12683;
assign w12685 = ~w12578 & ~w12683;
assign w12686 = ~w12684 & ~w12685;
assign w12687 = w12568 & ~w12686;
assign w12688 = ~w12568 & w12686;
assign w12689 = ~w12687 & ~w12688;
assign w12690 = b[24] & w5167;
assign w12691 = b[25] & w4918;
assign w12692 = b[26] & w4925;
assign w12693 = w2219 & w4923;
assign w12694 = ~w12691 & ~w12692;
assign w12695 = ~w12690 & w12694;
assign w12696 = ~w12693 & w12695;
assign w12697 = a[41] & ~w12696;
assign w12698 = ~a[41] & w12696;
assign w12699 = ~w12697 & ~w12698;
assign w12700 = w12689 & w12699;
assign w12701 = ~w12689 & ~w12699;
assign w12702 = ~w12700 & ~w12701;
assign w12703 = (~w12413 & w12416) | (~w12413 & w25307) | (w12416 & w25307);
assign w12704 = ~w12702 & w12703;
assign w12705 = w12702 & ~w12703;
assign w12706 = ~w12704 & ~w12705;
assign w12707 = b[27] & w4453;
assign w12708 = b[29] & w4243;
assign w12709 = b[28] & w4241;
assign w12710 = w2734 & w4236;
assign w12711 = ~w12708 & ~w12709;
assign w12712 = ~w12707 & w12711;
assign w12713 = ~w12710 & w12712;
assign w12714 = a[38] & ~w12713;
assign w12715 = ~a[38] & w12713;
assign w12716 = ~w12714 & ~w12715;
assign w12717 = w12706 & w12716;
assign w12718 = ~w12706 & ~w12716;
assign w12719 = ~w12717 & ~w12718;
assign w12720 = (~w12420 & w12423) | (~w12420 & w25196) | (w12423 & w25196);
assign w12721 = ~w12719 & w12720;
assign w12722 = w12719 & ~w12720;
assign w12723 = ~w12721 & ~w12722;
assign w12724 = b[30] & w3785;
assign w12725 = b[32] & w3580;
assign w12726 = b[31] & w3578;
assign w12727 = w3304 & w3573;
assign w12728 = ~w12725 & ~w12726;
assign w12729 = ~w12724 & w12728;
assign w12730 = ~w12727 & w12729;
assign w12731 = a[35] & ~w12730;
assign w12732 = ~a[35] & w12730;
assign w12733 = ~w12731 & ~w12732;
assign w12734 = w12723 & w12733;
assign w12735 = ~w12723 & ~w12733;
assign w12736 = ~w12734 & ~w12735;
assign w12737 = w12567 & w12736;
assign w12738 = ~w12567 & ~w12736;
assign w12739 = ~w12737 & ~w12738;
assign w12740 = w12566 & ~w12739;
assign w12741 = ~w12566 & w12739;
assign w12742 = ~w12740 & ~w12741;
assign w12743 = w12556 & ~w12742;
assign w12744 = ~w12556 & w12742;
assign w12745 = ~w12743 & ~w12744;
assign w12746 = b[37] & w2436;
assign w12747 = b[36] & ~w2622;
assign w12748 = b[38] & w2438;
assign w12749 = w2432 & w4582;
assign w12750 = ~w12746 & ~w12747;
assign w12751 = ~w12748 & w12750;
assign w12752 = ~w12749 & w12751;
assign w12753 = a[29] & ~w12752;
assign w12754 = ~a[29] & w12752;
assign w12755 = ~w12753 & ~w12754;
assign w12756 = w12745 & w12755;
assign w12757 = ~w12745 & ~w12755;
assign w12758 = ~w12756 & ~w12757;
assign w12759 = ~w12451 & ~w12455;
assign w12760 = ~w12758 & w12759;
assign w12761 = w12758 & ~w12759;
assign w12762 = ~w12760 & ~w12761;
assign w12763 = b[40] & w1955;
assign w12764 = b[41] & w1957;
assign w12765 = b[39] & ~w2114;
assign w12766 = w1951 & w5302;
assign w12767 = ~w12763 & ~w12764;
assign w12768 = ~w12765 & w12767;
assign w12769 = ~w12766 & w12768;
assign w12770 = a[26] & ~w12769;
assign w12771 = ~a[26] & w12769;
assign w12772 = ~w12770 & ~w12771;
assign w12773 = w12762 & w12772;
assign w12774 = ~w12762 & ~w12772;
assign w12775 = ~w12773 & ~w12774;
assign w12776 = w12555 & w12775;
assign w12777 = ~w12555 & ~w12775;
assign w12778 = ~w12776 & ~w12777;
assign w12779 = w12554 & ~w12778;
assign w12780 = ~w12554 & w12778;
assign w12781 = ~w12779 & ~w12780;
assign w12782 = (~w12466 & ~w12230) | (~w12466 & w24857) | (~w12230 & w24857);
assign w12783 = w12781 & w12782;
assign w12784 = ~w12781 & ~w12782;
assign w12785 = ~w12783 & ~w12784;
assign w12786 = ~w12544 & ~w12785;
assign w12787 = w12544 & w12785;
assign w12788 = ~w12786 & ~w12787;
assign w12789 = ~w12534 & w12788;
assign w12790 = w12534 & ~w12788;
assign w12791 = ~w12789 & ~w12790;
assign w12792 = w12533 & w12791;
assign w12793 = ~w12533 & ~w12791;
assign w12794 = ~w12792 & ~w12793;
assign w12795 = (~w12478 & ~w12208) | (~w12478 & w25557) | (~w12208 & w25557);
assign w12796 = ~w12794 & ~w12795;
assign w12797 = w12794 & w12795;
assign w12798 = ~w12796 & ~w12797;
assign w12799 = b[51] & ~w649;
assign w12800 = b[52] & w573;
assign w12801 = b[53] & w575;
assign w12802 = w569 & w8683;
assign w12803 = ~w12799 & ~w12800;
assign w12804 = ~w12801 & w12803;
assign w12805 = ~w12802 & w12804;
assign w12806 = a[14] & ~w12805;
assign w12807 = ~a[14] & w12805;
assign w12808 = ~w12806 & ~w12807;
assign w12809 = w12798 & w12808;
assign w12810 = ~w12798 & ~w12808;
assign w12811 = ~w12809 & ~w12810;
assign w12812 = ~w12483 & ~w12488;
assign w12813 = ~w12811 & w12812;
assign w12814 = w12811 & ~w12812;
assign w12815 = ~w12813 & ~w12814;
assign w12816 = b[56] & w360;
assign w12817 = b[55] & w358;
assign w12818 = b[54] & ~w419;
assign w12819 = w354 & w9657;
assign w12820 = ~w12816 & ~w12817;
assign w12821 = ~w12818 & w12820;
assign w12822 = ~w12819 & w12821;
assign w12823 = a[11] & ~w12822;
assign w12824 = ~a[11] & w12822;
assign w12825 = ~w12823 & ~w12824;
assign w12826 = b[57] & ~w237;
assign w12827 = b[59] & w185;
assign w12828 = b[58] & w183;
assign w12829 = w179 & w10371;
assign w12830 = ~w12826 & ~w12827;
assign w12831 = ~w12828 & w12830;
assign w12832 = ~w12829 & w12831;
assign w12833 = a[8] & ~w12832;
assign w12834 = ~a[8] & w12832;
assign w12835 = ~w12833 & ~w12834;
assign w12836 = w12825 & w12835;
assign w12837 = ~w12825 & ~w12835;
assign w12838 = ~w12836 & ~w12837;
assign w12839 = w12815 & ~w12838;
assign w12840 = ~w12815 & w12838;
assign w12841 = ~w12839 & ~w12840;
assign w12842 = ~w12523 & ~w12841;
assign w12843 = w12523 & w12841;
assign w12844 = ~w12842 & ~w12843;
assign w12845 = w12522 & w12844;
assign w12846 = ~w12522 & ~w12844;
assign w12847 = ~w12845 & ~w12846;
assign w12848 = ~a[2] & ~w12155;
assign w12849 = ~w117 & ~w10378;
assign w12850 = ~w12154 & ~w12849;
assign w12851 = ~w25 & ~w12850;
assign w12852 = b[63] & ~w12851;
assign w12853 = ~w12848 & ~w12852;
assign w12854 = (w12499 & w24858) | (w12499 & w24859) | (w24858 & w24859);
assign w12855 = (~w12499 & w24860) | (~w12499 & w24861) | (w24860 & w24861);
assign w12856 = ~w12854 & ~w12855;
assign w12857 = ~w12847 & ~w12856;
assign w12858 = w12847 & w12856;
assign w12859 = ~w12857 & ~w12858;
assign w12860 = ~w12166 & ~w12504;
assign w12861 = ~w12859 & ~w12860;
assign w12862 = w12859 & w12860;
assign w12863 = ~w12861 & ~w12862;
assign w12864 = (~w12507 & w12509) | (~w12507 & w24401) | (w12509 & w24401);
assign w12865 = (w12509 & w25010) | (w12509 & w25011) | (w25010 & w25011);
assign w12866 = ~w12863 & ~w12864;
assign w12867 = ~w12865 & ~w12866;
assign w12868 = (~w12855 & ~w12856) | (~w12855 & w25558) | (~w12856 & w25558);
assign w12869 = (~w12842 & ~w12844) | (~w12842 & w24862) | (~w12844 & w24862);
assign w12870 = b[61] & w103;
assign w12871 = b[62] & w61;
assign w12872 = b[63] & w68;
assign w12873 = w66 & w12132;
assign w12874 = ~w12871 & ~w12872;
assign w12875 = ~w12870 & w12874;
assign w12876 = ~w12873 & w12875;
assign w12877 = a[5] & ~w12876;
assign w12878 = ~a[5] & w12876;
assign w12879 = ~w12877 & ~w12878;
assign w12880 = ~w12869 & w12879;
assign w12881 = w12869 & ~w12879;
assign w12882 = ~w12880 & ~w12881;
assign w12883 = b[57] & w360;
assign w12884 = b[55] & ~w419;
assign w12885 = b[56] & w358;
assign w12886 = w354 & ~w9992;
assign w12887 = ~w12883 & ~w12884;
assign w12888 = ~w12885 & w12887;
assign w12889 = ~w12886 & w12888;
assign w12890 = a[11] & ~w12889;
assign w12891 = ~a[11] & w12889;
assign w12892 = ~w12890 & ~w12891;
assign w12893 = (w12892 & w24863) | (w12892 & w12814) | (w24863 & w12814);
assign w12894 = (w24864 & w12812) | (w24864 & w25559) | (w12812 & w25559);
assign w12895 = ~w12893 & ~w12894;
assign w12896 = b[25] & w5167;
assign w12897 = b[27] & w4925;
assign w12898 = b[26] & w4918;
assign w12899 = w2378 & w4923;
assign w12900 = ~w12897 & ~w12898;
assign w12901 = ~w12896 & w12900;
assign w12902 = ~w12899 & w12901;
assign w12903 = a[41] & ~w12902;
assign w12904 = ~a[41] & w12902;
assign w12905 = ~w12903 & ~w12904;
assign w12906 = b[19] & w6732;
assign w12907 = b[20] & w6474;
assign w12908 = b[21] & w6476;
assign w12909 = w1467 & w6469;
assign w12910 = ~w12907 & ~w12908;
assign w12911 = ~w12906 & w12910;
assign w12912 = ~w12909 & w12911;
assign w12913 = a[47] & ~w12912;
assign w12914 = ~a[47] & w12912;
assign w12915 = ~w12913 & ~w12914;
assign w12916 = b[16] & w7586;
assign w12917 = b[17] & w7307;
assign w12918 = b[18] & w7314;
assign w12919 = ~w1108 & w7312;
assign w12920 = ~w12917 & ~w12918;
assign w12921 = ~w12916 & w12920;
assign w12922 = ~w12919 & w12921;
assign w12923 = a[50] & ~w12922;
assign w12924 = ~a[50] & w12922;
assign w12925 = ~w12923 & ~w12924;
assign w12926 = ~w12640 & ~w12643;
assign w12927 = ~w12608 & ~w12612;
assign w12928 = b[2] & w11921;
assign w12929 = b[3] & w11923;
assign w12930 = ~w12928 & ~w12929;
assign w12931 = a[2] & ~w12930;
assign w12932 = ~a[2] & w12930;
assign w12933 = ~w12931 & ~w12932;
assign w12934 = b[4] & w11561;
assign w12935 = b[6] & w11196;
assign w12936 = b[5] & w11194;
assign w12937 = w157 & w11189;
assign w12938 = ~w12935 & ~w12936;
assign w12939 = ~w12934 & w12938;
assign w12940 = ~w12937 & w12939;
assign w12941 = a[62] & ~w12940;
assign w12942 = ~a[62] & w12940;
assign w12943 = ~w12941 & ~w12942;
assign w12944 = w12933 & w12943;
assign w12945 = ~w12933 & ~w12943;
assign w12946 = ~w12944 & ~w12945;
assign w12947 = w12927 & ~w12946;
assign w12948 = ~w12927 & w12946;
assign w12949 = ~w12947 & ~w12948;
assign w12950 = b[7] & w10496;
assign w12951 = b[8] & w10146;
assign w12952 = b[9] & w10148;
assign w12953 = w322 & w10141;
assign w12954 = ~w12951 & ~w12952;
assign w12955 = ~w12950 & w12954;
assign w12956 = ~w12953 & w12955;
assign w12957 = a[59] & ~w12956;
assign w12958 = ~a[59] & w12956;
assign w12959 = ~w12957 & ~w12958;
assign w12960 = w12949 & w12959;
assign w12961 = ~w12949 & ~w12959;
assign w12962 = ~w12960 & ~w12961;
assign w12963 = ~w12624 & ~w12627;
assign w12964 = w12962 & w12963;
assign w12965 = ~w12962 & ~w12963;
assign w12966 = ~w12964 & ~w12965;
assign w12967 = b[10] & w9482;
assign w12968 = b[11] & w9165;
assign w12969 = b[12] & w9160;
assign w12970 = w536 & w9158;
assign w12971 = ~w12968 & ~w12969;
assign w12972 = ~w12967 & w12971;
assign w12973 = ~w12970 & w12972;
assign w12974 = a[56] & ~w12973;
assign w12975 = ~a[56] & w12973;
assign w12976 = ~w12974 & ~w12975;
assign w12977 = w12966 & w12976;
assign w12978 = ~w12966 & ~w12976;
assign w12979 = ~w12977 & ~w12978;
assign w12980 = w12926 & ~w12979;
assign w12981 = ~w12926 & w12979;
assign w12982 = ~w12980 & ~w12981;
assign w12983 = b[13] & w8515;
assign w12984 = b[14] & w8200;
assign w12985 = b[15] & w8202;
assign w12986 = ~w799 & w8195;
assign w12987 = ~w12984 & ~w12985;
assign w12988 = ~w12983 & w12987;
assign w12989 = ~w12986 & w12988;
assign w12990 = a[53] & ~w12989;
assign w12991 = ~a[53] & w12989;
assign w12992 = ~w12990 & ~w12991;
assign w12993 = w12982 & w12992;
assign w12994 = ~w12982 & ~w12992;
assign w12995 = ~w12993 & ~w12994;
assign w12996 = (~w12656 & w12591) | (~w12656 & w25012) | (w12591 & w25012);
assign w12997 = w12995 & ~w12996;
assign w12998 = ~w12995 & w12996;
assign w12999 = ~w12997 & ~w12998;
assign w13000 = w12925 & w12999;
assign w13001 = ~w12925 & ~w12999;
assign w13002 = ~w13000 & ~w13001;
assign w13003 = ~w12662 & ~w12666;
assign w13004 = w13002 & ~w13003;
assign w13005 = ~w13002 & w13003;
assign w13006 = ~w13004 & ~w13005;
assign w13007 = ~w12915 & ~w13006;
assign w13008 = w12915 & w13006;
assign w13009 = ~w13007 & ~w13008;
assign w13010 = ~w12678 & ~w12681;
assign w13011 = w13009 & ~w13010;
assign w13012 = ~w13009 & w13010;
assign w13013 = ~w13011 & ~w13012;
assign w13014 = b[22] & w5939;
assign w13015 = b[23] & w5670;
assign w13016 = b[24] & w5665;
assign w13017 = w1895 & w5663;
assign w13018 = ~w13015 & ~w13016;
assign w13019 = ~w13014 & w13018;
assign w13020 = ~w13017 & w13019;
assign w13021 = a[44] & ~w13020;
assign w13022 = ~a[44] & w13020;
assign w13023 = ~w13021 & ~w13022;
assign w13024 = w13013 & w13023;
assign w13025 = ~w13013 & ~w13023;
assign w13026 = ~w13024 & ~w13025;
assign w13027 = ~w12684 & ~w12688;
assign w13028 = w13026 & ~w13027;
assign w13029 = ~w13026 & w13027;
assign w13030 = ~w13028 & ~w13029;
assign w13031 = w12905 & w13030;
assign w13032 = ~w12905 & ~w13030;
assign w13033 = ~w13031 & ~w13032;
assign w13034 = (~w12700 & w12703) | (~w12700 & w24865) | (w12703 & w24865);
assign w13035 = w13033 & ~w13034;
assign w13036 = ~w13033 & w13034;
assign w13037 = ~w13035 & ~w13036;
assign w13038 = b[28] & w4453;
assign w13039 = b[30] & w4243;
assign w13040 = b[29] & w4241;
assign w13041 = ~w2908 & w4236;
assign w13042 = ~w13039 & ~w13040;
assign w13043 = ~w13038 & w13042;
assign w13044 = ~w13041 & w13043;
assign w13045 = a[38] & ~w13044;
assign w13046 = ~a[38] & w13044;
assign w13047 = ~w13045 & ~w13046;
assign w13048 = ~w13037 & ~w13047;
assign w13049 = w13037 & w13047;
assign w13050 = ~w13048 & ~w13049;
assign w13051 = (~w12717 & w12720) | (~w12717 & w25308) | (w12720 & w25308);
assign w13052 = w13050 & ~w13051;
assign w13053 = ~w13050 & w13051;
assign w13054 = ~w13052 & ~w13053;
assign w13055 = b[31] & w3785;
assign w13056 = b[32] & w3578;
assign w13057 = b[33] & w3580;
assign w13058 = w3499 & w3573;
assign w13059 = ~w13056 & ~w13057;
assign w13060 = ~w13055 & w13059;
assign w13061 = ~w13058 & w13060;
assign w13062 = a[35] & ~w13061;
assign w13063 = ~a[35] & w13061;
assign w13064 = ~w13062 & ~w13063;
assign w13065 = w13054 & w13064;
assign w13066 = ~w13054 & ~w13064;
assign w13067 = ~w13065 & ~w13066;
assign w13068 = b[34] & w3177;
assign w13069 = b[35] & w2973;
assign w13070 = b[36] & w2978;
assign w13071 = w2980 & w4129;
assign w13072 = ~w13069 & ~w13070;
assign w13073 = ~w13068 & w13072;
assign w13074 = ~w13071 & w13073;
assign w13075 = a[32] & ~w13074;
assign w13076 = ~a[32] & w13074;
assign w13077 = ~w13075 & ~w13076;
assign w13078 = (w25013 & ~w12567) | (w25013 & w25197) | (~w12567 & w25197);
assign w13079 = (w12567 & w25198) | (w12567 & w25199) | (w25198 & w25199);
assign w13080 = ~w13078 & ~w13079;
assign w13081 = w13067 & w13080;
assign w13082 = ~w13067 & ~w13080;
assign w13083 = ~w13081 & ~w13082;
assign w13084 = ~w12740 & ~w12744;
assign w13085 = b[37] & ~w2622;
assign w13086 = b[38] & w2436;
assign w13087 = b[39] & w2438;
assign w13088 = w2432 & ~w4812;
assign w13089 = ~w13085 & ~w13086;
assign w13090 = ~w13087 & w13089;
assign w13091 = ~w13088 & w13090;
assign w13092 = a[29] & ~w13091;
assign w13093 = ~a[29] & w13091;
assign w13094 = ~w13092 & ~w13093;
assign w13095 = ~w13084 & w13094;
assign w13096 = w13084 & ~w13094;
assign w13097 = ~w13095 & ~w13096;
assign w13098 = w13083 & w13097;
assign w13099 = ~w13083 & ~w13097;
assign w13100 = ~w13098 & ~w13099;
assign w13101 = b[40] & ~w2114;
assign w13102 = b[42] & w1957;
assign w13103 = b[41] & w1955;
assign w13104 = w1951 & w5548;
assign w13105 = ~w13101 & ~w13102;
assign w13106 = ~w13103 & w13105;
assign w13107 = ~w13104 & w13106;
assign w13108 = a[26] & ~w13107;
assign w13109 = ~a[26] & w13107;
assign w13110 = ~w13108 & ~w13109;
assign w13111 = (~w12756 & w12759) | (~w12756 & w25309) | (w12759 & w25309);
assign w13112 = w13110 & ~w13111;
assign w13113 = ~w13110 & w13111;
assign w13114 = ~w13112 & ~w13113;
assign w13115 = w13100 & w13114;
assign w13116 = ~w13100 & ~w13114;
assign w13117 = ~w13115 & ~w13116;
assign w13118 = b[45] & w1519;
assign w13119 = b[43] & ~w1676;
assign w13120 = b[44] & w1517;
assign w13121 = w1513 & w6334;
assign w13122 = ~w13118 & ~w13119;
assign w13123 = ~w13120 & w13122;
assign w13124 = ~w13121 & w13123;
assign w13125 = a[23] & ~w13124;
assign w13126 = ~a[23] & w13124;
assign w13127 = ~w13125 & ~w13126;
assign w13128 = ~w12774 & ~w12776;
assign w13129 = w13127 & w13128;
assign w13130 = ~w13127 & ~w13128;
assign w13131 = ~w13129 & ~w13130;
assign w13132 = ~w13117 & ~w13131;
assign w13133 = w13117 & w13131;
assign w13134 = ~w13132 & ~w13133;
assign w13135 = b[46] & ~w1272;
assign w13136 = b[47] & w1154;
assign w13137 = b[48] & w1156;
assign w13138 = w1150 & ~w7170;
assign w13139 = ~w13135 & ~w13136;
assign w13140 = ~w13137 & w13139;
assign w13141 = ~w13138 & w13140;
assign w13142 = a[20] & ~w13141;
assign w13143 = ~a[20] & w13141;
assign w13144 = ~w13142 & ~w13143;
assign w13145 = ~w12779 & ~w12783;
assign w13146 = w13144 & ~w13145;
assign w13147 = ~w13144 & w13145;
assign w13148 = ~w13146 & ~w13147;
assign w13149 = w13134 & w13148;
assign w13150 = ~w13134 & ~w13148;
assign w13151 = ~w13149 & ~w13150;
assign w13152 = b[49] & ~w934;
assign w13153 = b[51] & w834;
assign w13154 = b[50] & w838;
assign w13155 = w832 & ~w8058;
assign w13156 = ~w13152 & ~w13153;
assign w13157 = ~w13154 & w13156;
assign w13158 = ~w13155 & w13157;
assign w13159 = a[17] & ~w13158;
assign w13160 = ~a[17] & w13158;
assign w13161 = ~w13159 & ~w13160;
assign w13162 = (~w12787 & w12534) | (~w12787 & w25310) | (w12534 & w25310);
assign w13163 = w13161 & ~w13162;
assign w13164 = ~w13161 & w13162;
assign w13165 = ~w13163 & ~w13164;
assign w13166 = w13151 & w13165;
assign w13167 = ~w13151 & ~w13165;
assign w13168 = ~w13166 & ~w13167;
assign w13169 = b[54] & w575;
assign w13170 = b[52] & ~w649;
assign w13171 = b[53] & w573;
assign w13172 = w569 & ~w8998;
assign w13173 = ~w13169 & ~w13170;
assign w13174 = ~w13171 & w13173;
assign w13175 = ~w13172 & w13174;
assign w13176 = a[14] & ~w13175;
assign w13177 = ~a[14] & w13175;
assign w13178 = ~w13176 & ~w13177;
assign w13179 = w13178 & w25726;
assign w13180 = ~w12792 & w25727;
assign w13181 = ~w13179 & ~w13180;
assign w13182 = w13168 & w13181;
assign w13183 = ~w13168 & ~w13181;
assign w13184 = ~w13182 & ~w13183;
assign w13185 = w12895 & w13184;
assign w13186 = ~w12895 & ~w13184;
assign w13187 = ~w13185 & ~w13186;
assign w13188 = b[60] & w185;
assign w13189 = b[58] & ~w237;
assign w13190 = b[59] & w183;
assign w13191 = w179 & w11035;
assign w13192 = ~w13188 & ~w13189;
assign w13193 = ~w13190 & w13192;
assign w13194 = ~w13191 & w13193;
assign w13195 = a[8] & ~w13194;
assign w13196 = ~a[8] & w13194;
assign w13197 = ~w13195 & ~w13196;
assign w13198 = (w12815 & w25201) | (w12815 & w25202) | (w25201 & w25202);
assign w13199 = (~w12815 & w25203) | (~w12815 & w25204) | (w25203 & w25204);
assign w13200 = ~w13198 & ~w13199;
assign w13201 = w13187 & w13200;
assign w13202 = ~w13187 & ~w13200;
assign w13203 = ~w13201 & ~w13202;
assign w13204 = w12882 & w13203;
assign w13205 = ~w12882 & ~w13203;
assign w13206 = ~w13204 & ~w13205;
assign w13207 = w12868 & ~w13206;
assign w13208 = ~w12868 & w13206;
assign w13209 = ~w13207 & ~w13208;
assign w13210 = ~w12862 & ~w12865;
assign w13211 = ~w13209 & ~w13210;
assign w13212 = ~w12865 & w24402;
assign w13213 = ~w13211 & ~w13212;
assign w13214 = (~w12880 & ~w12882) | (~w12880 & w25205) | (~w12882 & w25205);
assign w13215 = b[54] & w573;
assign w13216 = b[55] & w575;
assign w13217 = b[53] & ~w649;
assign w13218 = w569 & ~w9330;
assign w13219 = ~w13215 & ~w13216;
assign w13220 = ~w13217 & w13219;
assign w13221 = ~w13218 & w13220;
assign w13222 = a[14] & ~w13221;
assign w13223 = ~a[14] & w13221;
assign w13224 = ~w13222 & ~w13223;
assign w13225 = ~w13163 & ~w13166;
assign w13226 = w13224 & ~w13225;
assign w13227 = ~w13224 & w13225;
assign w13228 = ~w13226 & ~w13227;
assign w13229 = b[49] & w1156;
assign w13230 = b[47] & ~w1272;
assign w13231 = b[48] & w1154;
assign w13232 = w1150 & ~w7468;
assign w13233 = ~w13229 & ~w13230;
assign w13234 = ~w13231 & w13233;
assign w13235 = ~w13232 & w13234;
assign w13236 = a[20] & ~w13235;
assign w13237 = ~a[20] & w13235;
assign w13238 = ~w13236 & ~w13237;
assign w13239 = ~w13129 & ~w13133;
assign w13240 = w13238 & ~w13239;
assign w13241 = ~w13238 & w13239;
assign w13242 = ~w13240 & ~w13241;
assign w13243 = b[32] & w3785;
assign w13244 = b[33] & w3578;
assign w13245 = b[34] & w3580;
assign w13246 = w3573 & ~w3710;
assign w13247 = ~w13244 & ~w13245;
assign w13248 = ~w13243 & w13247;
assign w13249 = ~w13246 & w13248;
assign w13250 = a[35] & ~w13249;
assign w13251 = ~a[35] & w13249;
assign w13252 = ~w13250 & ~w13251;
assign w13253 = (~w13035 & ~w13037) | (~w13035 & w25015) | (~w13037 & w25015);
assign w13254 = b[29] & w4453;
assign w13255 = b[30] & w4241;
assign w13256 = b[31] & w4243;
assign w13257 = ~w3112 & w4236;
assign w13258 = ~w13255 & ~w13256;
assign w13259 = ~w13254 & w13258;
assign w13260 = ~w13257 & w13259;
assign w13261 = a[38] & ~w13260;
assign w13262 = ~a[38] & w13260;
assign w13263 = ~w13261 & ~w13262;
assign w13264 = b[26] & w5167;
assign w13265 = b[28] & w4925;
assign w13266 = b[27] & w4918;
assign w13267 = w2559 & w4923;
assign w13268 = ~w13265 & ~w13266;
assign w13269 = ~w13264 & w13268;
assign w13270 = ~w13267 & w13269;
assign w13271 = a[41] & ~w13270;
assign w13272 = ~a[41] & w13270;
assign w13273 = ~w13271 & ~w13272;
assign w13274 = (~w13011 & ~w13013) | (~w13011 & w25016) | (~w13013 & w25016);
assign w13275 = b[23] & w5939;
assign w13276 = b[25] & w5665;
assign w13277 = b[24] & w5670;
assign w13278 = w2061 & w5663;
assign w13279 = ~w13276 & ~w13277;
assign w13280 = ~w13275 & w13279;
assign w13281 = ~w13278 & w13280;
assign w13282 = a[44] & ~w13281;
assign w13283 = ~a[44] & w13281;
assign w13284 = ~w13282 & ~w13283;
assign w13285 = b[20] & w6732;
assign w13286 = b[21] & w6474;
assign w13287 = b[22] & w6476;
assign w13288 = w1615 & w6469;
assign w13289 = ~w13286 & ~w13287;
assign w13290 = ~w13285 & w13289;
assign w13291 = ~w13288 & w13290;
assign w13292 = a[47] & ~w13291;
assign w13293 = ~a[47] & w13291;
assign w13294 = ~w13292 & ~w13293;
assign w13295 = b[17] & w7586;
assign w13296 = b[19] & w7314;
assign w13297 = b[18] & w7307;
assign w13298 = ~w1231 & w7312;
assign w13299 = ~w13296 & ~w13297;
assign w13300 = ~w13295 & w13299;
assign w13301 = ~w13298 & w13300;
assign w13302 = a[50] & ~w13301;
assign w13303 = ~a[50] & w13301;
assign w13304 = ~w13302 & ~w13303;
assign w13305 = b[11] & w9482;
assign w13306 = b[13] & w9160;
assign w13307 = b[12] & w9165;
assign w13308 = w628 & w9158;
assign w13309 = ~w13306 & ~w13307;
assign w13310 = ~w13305 & w13309;
assign w13311 = ~w13308 & w13310;
assign w13312 = a[56] & ~w13311;
assign w13313 = ~a[56] & w13311;
assign w13314 = ~w13312 & ~w13313;
assign w13315 = b[8] & w10496;
assign w13316 = b[10] & w10148;
assign w13317 = b[9] & w10146;
assign w13318 = w397 & w10141;
assign w13319 = ~w13316 & ~w13317;
assign w13320 = ~w13315 & w13319;
assign w13321 = ~w13318 & w13320;
assign w13322 = a[59] & ~w13321;
assign w13323 = ~a[59] & w13321;
assign w13324 = ~w13322 & ~w13323;
assign w13325 = ~w12931 & ~w12944;
assign w13326 = b[3] & w11921;
assign w13327 = b[4] & w11923;
assign w13328 = ~w13326 & ~w13327;
assign w13329 = a[2] & ~w13328;
assign w13330 = ~a[2] & w13328;
assign w13331 = ~w13329 & ~w13330;
assign w13332 = b[5] & w11561;
assign w13333 = b[6] & w11194;
assign w13334 = b[7] & w11196;
assign w13335 = w216 & w11189;
assign w13336 = ~w13333 & ~w13334;
assign w13337 = ~w13332 & w13336;
assign w13338 = ~w13335 & w13337;
assign w13339 = a[62] & ~w13338;
assign w13340 = ~a[62] & w13338;
assign w13341 = ~w13339 & ~w13340;
assign w13342 = w13331 & w13341;
assign w13343 = ~w13331 & ~w13341;
assign w13344 = ~w13342 & ~w13343;
assign w13345 = ~w13325 & w13344;
assign w13346 = w13325 & ~w13344;
assign w13347 = ~w13345 & ~w13346;
assign w13348 = w13324 & w13347;
assign w13349 = ~w13324 & ~w13347;
assign w13350 = ~w13348 & ~w13349;
assign w13351 = ~w12948 & ~w12960;
assign w13352 = w13350 & ~w13351;
assign w13353 = ~w13350 & w13351;
assign w13354 = ~w13352 & ~w13353;
assign w13355 = ~w13314 & ~w13354;
assign w13356 = w13314 & w13354;
assign w13357 = ~w13355 & ~w13356;
assign w13358 = ~w12964 & ~w12977;
assign w13359 = w13357 & ~w13358;
assign w13360 = ~w13357 & w13358;
assign w13361 = ~w13359 & ~w13360;
assign w13362 = b[14] & w8515;
assign w13363 = b[16] & w8202;
assign w13364 = b[15] & w8200;
assign w13365 = w905 & w8195;
assign w13366 = ~w13363 & ~w13364;
assign w13367 = ~w13362 & w13366;
assign w13368 = ~w13365 & w13367;
assign w13369 = a[53] & ~w13368;
assign w13370 = ~a[53] & w13368;
assign w13371 = ~w13369 & ~w13370;
assign w13372 = w13361 & w13371;
assign w13373 = ~w13361 & ~w13371;
assign w13374 = ~w13372 & ~w13373;
assign w13375 = ~w12981 & ~w12993;
assign w13376 = w13374 & ~w13375;
assign w13377 = ~w13374 & w13375;
assign w13378 = ~w13376 & ~w13377;
assign w13379 = w13304 & w13378;
assign w13380 = ~w13304 & ~w13378;
assign w13381 = ~w13379 & ~w13380;
assign w13382 = ~w12997 & ~w13000;
assign w13383 = w13381 & ~w13382;
assign w13384 = ~w13381 & w13382;
assign w13385 = ~w13383 & ~w13384;
assign w13386 = w13294 & w13385;
assign w13387 = ~w13294 & ~w13385;
assign w13388 = ~w13386 & ~w13387;
assign w13389 = (~w13004 & ~w13006) | (~w13004 & w25017) | (~w13006 & w25017);
assign w13390 = w13388 & ~w13389;
assign w13391 = ~w13388 & w13389;
assign w13392 = ~w13390 & ~w13391;
assign w13393 = w13284 & w13392;
assign w13394 = ~w13284 & ~w13392;
assign w13395 = ~w13393 & ~w13394;
assign w13396 = ~w13274 & w13395;
assign w13397 = w13274 & ~w13395;
assign w13398 = ~w13396 & ~w13397;
assign w13399 = w13273 & w13398;
assign w13400 = ~w13273 & ~w13398;
assign w13401 = ~w13399 & ~w13400;
assign w13402 = (~w13028 & ~w13030) | (~w13028 & w25018) | (~w13030 & w25018);
assign w13403 = w13401 & ~w13402;
assign w13404 = ~w13401 & w13402;
assign w13405 = ~w13403 & ~w13404;
assign w13406 = ~w13263 & ~w13405;
assign w13407 = w13263 & w13405;
assign w13408 = ~w13406 & ~w13407;
assign w13409 = w13253 & ~w13408;
assign w13410 = ~w13253 & w13408;
assign w13411 = ~w13409 & ~w13410;
assign w13412 = w13252 & w13411;
assign w13413 = ~w13252 & ~w13411;
assign w13414 = ~w13412 & ~w13413;
assign w13415 = (~w13052 & ~w13054) | (~w13052 & w24867) | (~w13054 & w24867);
assign w13416 = b[35] & w3177;
assign w13417 = b[36] & w2973;
assign w13418 = b[37] & w2978;
assign w13419 = w2980 & ~w4357;
assign w13420 = ~w13417 & ~w13418;
assign w13421 = ~w13416 & w13420;
assign w13422 = ~w13419 & w13421;
assign w13423 = a[32] & ~w13422;
assign w13424 = ~a[32] & w13422;
assign w13425 = ~w13423 & ~w13424;
assign w13426 = ~w13415 & w13425;
assign w13427 = w13415 & ~w13425;
assign w13428 = ~w13426 & ~w13427;
assign w13429 = ~w13414 & ~w13428;
assign w13430 = w13414 & w13428;
assign w13431 = ~w13429 & ~w13430;
assign w13432 = (~w13078 & ~w13080) | (~w13078 & w25312) | (~w13080 & w25312);
assign w13433 = b[40] & w2438;
assign w13434 = b[39] & w2436;
assign w13435 = b[38] & ~w2622;
assign w13436 = w2432 & ~w5058;
assign w13437 = ~w13433 & ~w13434;
assign w13438 = ~w13435 & w13437;
assign w13439 = ~w13436 & w13438;
assign w13440 = a[29] & ~w13439;
assign w13441 = ~a[29] & w13439;
assign w13442 = ~w13440 & ~w13441;
assign w13443 = ~w13432 & w13442;
assign w13444 = w13432 & ~w13442;
assign w13445 = ~w13443 & ~w13444;
assign w13446 = w13431 & w13445;
assign w13447 = ~w13431 & ~w13445;
assign w13448 = ~w13446 & ~w13447;
assign w13449 = b[43] & w1957;
assign w13450 = b[42] & w1955;
assign w13451 = b[41] & ~w2114;
assign w13452 = w1951 & w5811;
assign w13453 = ~w13449 & ~w13450;
assign w13454 = ~w13451 & w13453;
assign w13455 = ~w13452 & w13454;
assign w13456 = a[26] & ~w13455;
assign w13457 = ~a[26] & w13455;
assign w13458 = ~w13456 & ~w13457;
assign w13459 = ~w13095 & ~w13098;
assign w13460 = w13458 & ~w13459;
assign w13461 = ~w13458 & w13459;
assign w13462 = ~w13460 & ~w13461;
assign w13463 = w13448 & w13462;
assign w13464 = ~w13448 & ~w13462;
assign w13465 = ~w13463 & ~w13464;
assign w13466 = b[46] & w1519;
assign w13467 = b[44] & ~w1676;
assign w13468 = b[45] & w1517;
assign w13469 = w1513 & ~w6613;
assign w13470 = ~w13466 & ~w13467;
assign w13471 = ~w13468 & w13470;
assign w13472 = ~w13469 & w13471;
assign w13473 = a[23] & ~w13472;
assign w13474 = ~a[23] & w13472;
assign w13475 = ~w13473 & ~w13474;
assign w13476 = ~w13112 & ~w13115;
assign w13477 = w13475 & ~w13476;
assign w13478 = ~w13475 & w13476;
assign w13479 = ~w13477 & ~w13478;
assign w13480 = w13465 & w13479;
assign w13481 = ~w13465 & ~w13479;
assign w13482 = ~w13480 & ~w13481;
assign w13483 = w13242 & w13482;
assign w13484 = ~w13242 & ~w13482;
assign w13485 = ~w13483 & ~w13484;
assign w13486 = b[52] & w834;
assign w13487 = b[51] & w838;
assign w13488 = b[50] & ~w934;
assign w13489 = w832 & ~w8371;
assign w13490 = ~w13486 & ~w13487;
assign w13491 = ~w13488 & w13490;
assign w13492 = ~w13489 & w13491;
assign w13493 = a[17] & ~w13492;
assign w13494 = ~a[17] & w13492;
assign w13495 = ~w13493 & ~w13494;
assign w13496 = ~w13146 & ~w13149;
assign w13497 = w13495 & ~w13496;
assign w13498 = ~w13495 & w13496;
assign w13499 = ~w13497 & ~w13498;
assign w13500 = w13485 & w13499;
assign w13501 = ~w13485 & ~w13499;
assign w13502 = ~w13500 & ~w13501;
assign w13503 = w13228 & w13502;
assign w13504 = ~w13228 & ~w13502;
assign w13505 = ~w13503 & ~w13504;
assign w13506 = ~w13179 & ~w13182;
assign w13507 = b[58] & w360;
assign w13508 = b[56] & ~w419;
assign w13509 = b[57] & w358;
assign w13510 = w354 & ~w10339;
assign w13511 = ~w13507 & ~w13508;
assign w13512 = ~w13509 & w13511;
assign w13513 = ~w13510 & w13512;
assign w13514 = a[11] & ~w13513;
assign w13515 = ~a[11] & w13513;
assign w13516 = ~w13514 & ~w13515;
assign w13517 = ~w13506 & w13516;
assign w13518 = w13506 & ~w13516;
assign w13519 = ~w13517 & ~w13518;
assign w13520 = w13505 & w13519;
assign w13521 = ~w13505 & ~w13519;
assign w13522 = ~w13520 & ~w13521;
assign w13523 = (~w12893 & ~w12895) | (~w12893 & w25206) | (~w12895 & w25206);
assign w13524 = b[59] & ~w237;
assign w13525 = b[60] & w183;
assign w13526 = b[61] & w185;
assign w13527 = w179 & w11400;
assign w13528 = ~w13524 & ~w13525;
assign w13529 = ~w13526 & w13528;
assign w13530 = ~w13527 & w13529;
assign w13531 = a[8] & ~w13530;
assign w13532 = ~a[8] & w13530;
assign w13533 = ~w13531 & ~w13532;
assign w13534 = ~w13523 & w13533;
assign w13535 = w13523 & ~w13533;
assign w13536 = ~w13534 & ~w13535;
assign w13537 = w13522 & w13536;
assign w13538 = ~w13522 & ~w13536;
assign w13539 = ~w13537 & ~w13538;
assign w13540 = (~w13198 & ~w13187) | (~w13198 & w25207) | (~w13187 & w25207);
assign w13541 = b[62] & w103;
assign w13542 = b[63] & w61;
assign w13543 = w66 & w12156;
assign w13544 = ~w13541 & ~w13542;
assign w13545 = ~w13543 & w13544;
assign w13546 = a[5] & w13545;
assign w13547 = ~a[5] & ~w13545;
assign w13548 = ~w13546 & ~w13547;
assign w13549 = ~w13540 & ~w13548;
assign w13550 = w13540 & w13548;
assign w13551 = ~w13549 & ~w13550;
assign w13552 = w13539 & w13551;
assign w13553 = ~w13539 & ~w13551;
assign w13554 = ~w13552 & ~w13553;
assign w13555 = w13214 & ~w13554;
assign w13556 = ~w13214 & w13554;
assign w13557 = ~w13555 & ~w13556;
assign w13558 = ~w13207 & ~w13212;
assign w13559 = ~w13212 & w24403;
assign w13560 = ~w13557 & ~w13558;
assign w13561 = ~w13559 & ~w13560;
assign w13562 = ~w13549 & ~w13552;
assign w13563 = b[57] & ~w419;
assign w13564 = b[59] & w360;
assign w13565 = b[58] & w358;
assign w13566 = w354 & w10371;
assign w13567 = ~w13563 & ~w13564;
assign w13568 = ~w13565 & w13567;
assign w13569 = ~w13566 & w13568;
assign w13570 = a[11] & ~w13569;
assign w13571 = ~a[11] & w13569;
assign w13572 = ~w13570 & ~w13571;
assign w13573 = ~w13226 & ~w13503;
assign w13574 = w13572 & ~w13573;
assign w13575 = ~w13572 & w13573;
assign w13576 = ~w13574 & ~w13575;
assign w13577 = b[46] & w1517;
assign w13578 = b[47] & w1519;
assign w13579 = b[45] & ~w1676;
assign w13580 = w1513 & w6889;
assign w13581 = ~w13577 & ~w13578;
assign w13582 = ~w13579 & w13581;
assign w13583 = ~w13580 & w13582;
assign w13584 = a[23] & ~w13583;
assign w13585 = ~a[23] & w13583;
assign w13586 = ~w13584 & ~w13585;
assign w13587 = ~w13460 & ~w13463;
assign w13588 = w13586 & ~w13587;
assign w13589 = ~w13586 & w13587;
assign w13590 = ~w13588 & ~w13589;
assign w13591 = b[30] & w4453;
assign w13592 = b[32] & w4243;
assign w13593 = b[31] & w4241;
assign w13594 = w3304 & w4236;
assign w13595 = ~w13592 & ~w13593;
assign w13596 = ~w13591 & w13595;
assign w13597 = ~w13594 & w13596;
assign w13598 = a[38] & ~w13597;
assign w13599 = ~a[38] & w13597;
assign w13600 = ~w13598 & ~w13599;
assign w13601 = b[24] & w5939;
assign w13602 = b[26] & w5665;
assign w13603 = b[25] & w5670;
assign w13604 = w2219 & w5663;
assign w13605 = ~w13602 & ~w13603;
assign w13606 = ~w13601 & w13605;
assign w13607 = ~w13604 & w13606;
assign w13608 = a[44] & ~w13607;
assign w13609 = ~a[44] & w13607;
assign w13610 = ~w13608 & ~w13609;
assign w13611 = ~w13359 & ~w13372;
assign w13612 = b[15] & w8515;
assign w13613 = b[16] & w8200;
assign w13614 = b[17] & w8202;
assign w13615 = w1008 & w8195;
assign w13616 = ~w13613 & ~w13614;
assign w13617 = ~w13612 & w13616;
assign w13618 = ~w13615 & w13617;
assign w13619 = a[53] & ~w13618;
assign w13620 = ~a[53] & w13618;
assign w13621 = ~w13619 & ~w13620;
assign w13622 = ~w13329 & ~w13342;
assign w13623 = b[4] & w11921;
assign w13624 = b[5] & w11923;
assign w13625 = ~w13623 & ~w13624;
assign w13626 = a[2] & ~w13625;
assign w13627 = ~a[2] & w13625;
assign w13628 = ~w13626 & ~w13627;
assign w13629 = b[6] & w11561;
assign w13630 = b[7] & w11194;
assign w13631 = b[8] & w11196;
assign w13632 = w270 & w11189;
assign w13633 = ~w13630 & ~w13631;
assign w13634 = ~w13629 & w13633;
assign w13635 = ~w13632 & w13634;
assign w13636 = a[62] & ~w13635;
assign w13637 = ~a[62] & w13635;
assign w13638 = ~w13636 & ~w13637;
assign w13639 = w13628 & w13638;
assign w13640 = ~w13628 & ~w13638;
assign w13641 = ~w13639 & ~w13640;
assign w13642 = ~w13622 & w13641;
assign w13643 = w13622 & ~w13641;
assign w13644 = ~w13642 & ~w13643;
assign w13645 = b[9] & w10496;
assign w13646 = b[10] & w10146;
assign w13647 = b[11] & w10148;
assign w13648 = w469 & w10141;
assign w13649 = ~w13646 & ~w13647;
assign w13650 = ~w13645 & w13649;
assign w13651 = ~w13648 & w13650;
assign w13652 = a[59] & ~w13651;
assign w13653 = ~a[59] & w13651;
assign w13654 = ~w13652 & ~w13653;
assign w13655 = ~w13644 & ~w13654;
assign w13656 = w13644 & w13654;
assign w13657 = ~w13655 & ~w13656;
assign w13658 = ~w13345 & ~w13348;
assign w13659 = w13657 & ~w13658;
assign w13660 = ~w13657 & w13658;
assign w13661 = ~w13659 & ~w13660;
assign w13662 = b[12] & w9482;
assign w13663 = b[14] & w9160;
assign w13664 = b[13] & w9165;
assign w13665 = w714 & w9158;
assign w13666 = ~w13663 & ~w13664;
assign w13667 = ~w13662 & w13666;
assign w13668 = ~w13665 & w13667;
assign w13669 = a[56] & ~w13668;
assign w13670 = ~a[56] & w13668;
assign w13671 = ~w13669 & ~w13670;
assign w13672 = w13661 & w13671;
assign w13673 = ~w13661 & ~w13671;
assign w13674 = ~w13672 & ~w13673;
assign w13675 = ~w13352 & ~w13356;
assign w13676 = w13674 & ~w13675;
assign w13677 = ~w13674 & w13675;
assign w13678 = ~w13676 & ~w13677;
assign w13679 = w13621 & w13678;
assign w13680 = ~w13621 & ~w13678;
assign w13681 = ~w13679 & ~w13680;
assign w13682 = ~w13611 & w13681;
assign w13683 = w13611 & ~w13681;
assign w13684 = ~w13682 & ~w13683;
assign w13685 = b[18] & w7586;
assign w13686 = b[19] & w7307;
assign w13687 = b[20] & w7314;
assign w13688 = w1347 & w7312;
assign w13689 = ~w13686 & ~w13687;
assign w13690 = ~w13685 & w13689;
assign w13691 = ~w13688 & w13690;
assign w13692 = a[50] & ~w13691;
assign w13693 = ~a[50] & w13691;
assign w13694 = ~w13692 & ~w13693;
assign w13695 = ~w13684 & ~w13694;
assign w13696 = w13684 & w13694;
assign w13697 = ~w13695 & ~w13696;
assign w13698 = ~w13376 & ~w13379;
assign w13699 = w13697 & ~w13698;
assign w13700 = ~w13697 & w13698;
assign w13701 = ~w13699 & ~w13700;
assign w13702 = b[21] & w6732;
assign w13703 = b[22] & w6474;
assign w13704 = b[23] & w6476;
assign w13705 = w1755 & w6469;
assign w13706 = ~w13703 & ~w13704;
assign w13707 = ~w13702 & w13706;
assign w13708 = ~w13705 & w13707;
assign w13709 = a[47] & ~w13708;
assign w13710 = ~a[47] & w13708;
assign w13711 = ~w13709 & ~w13710;
assign w13712 = w13701 & w13711;
assign w13713 = ~w13701 & ~w13711;
assign w13714 = ~w13712 & ~w13713;
assign w13715 = ~w13383 & ~w13386;
assign w13716 = w13714 & ~w13715;
assign w13717 = ~w13714 & w13715;
assign w13718 = ~w13716 & ~w13717;
assign w13719 = w13610 & w13718;
assign w13720 = ~w13610 & ~w13718;
assign w13721 = ~w13719 & ~w13720;
assign w13722 = ~w13390 & ~w13393;
assign w13723 = w13721 & ~w13722;
assign w13724 = ~w13721 & w13722;
assign w13725 = ~w13723 & ~w13724;
assign w13726 = b[27] & w5167;
assign w13727 = b[29] & w4925;
assign w13728 = b[28] & w4918;
assign w13729 = w2734 & w4923;
assign w13730 = ~w13727 & ~w13728;
assign w13731 = ~w13726 & w13730;
assign w13732 = ~w13729 & w13731;
assign w13733 = a[41] & ~w13732;
assign w13734 = ~a[41] & w13732;
assign w13735 = ~w13733 & ~w13734;
assign w13736 = w13725 & w13735;
assign w13737 = ~w13725 & ~w13735;
assign w13738 = ~w13736 & ~w13737;
assign w13739 = ~w13396 & ~w13399;
assign w13740 = w13738 & ~w13739;
assign w13741 = ~w13738 & w13739;
assign w13742 = ~w13740 & ~w13741;
assign w13743 = ~w13600 & ~w13742;
assign w13744 = w13600 & w13742;
assign w13745 = ~w13743 & ~w13744;
assign w13746 = ~w13403 & ~w13407;
assign w13747 = w13745 & ~w13746;
assign w13748 = ~w13745 & w13746;
assign w13749 = ~w13747 & ~w13748;
assign w13750 = b[33] & w3785;
assign w13751 = b[35] & w3580;
assign w13752 = b[34] & w3578;
assign w13753 = w3573 & w3918;
assign w13754 = ~w13751 & ~w13752;
assign w13755 = ~w13750 & w13754;
assign w13756 = ~w13753 & w13755;
assign w13757 = a[35] & ~w13756;
assign w13758 = ~a[35] & w13756;
assign w13759 = ~w13757 & ~w13758;
assign w13760 = w13749 & w13759;
assign w13761 = ~w13749 & ~w13759;
assign w13762 = ~w13760 & ~w13761;
assign w13763 = ~w13410 & ~w13412;
assign w13764 = b[36] & w3177;
assign w13765 = b[37] & w2973;
assign w13766 = b[38] & w2978;
assign w13767 = w2980 & w4582;
assign w13768 = ~w13765 & ~w13766;
assign w13769 = ~w13764 & w13768;
assign w13770 = ~w13767 & w13769;
assign w13771 = a[32] & ~w13770;
assign w13772 = ~a[32] & w13770;
assign w13773 = ~w13771 & ~w13772;
assign w13774 = ~w13763 & w13773;
assign w13775 = w13763 & ~w13773;
assign w13776 = ~w13774 & ~w13775;
assign w13777 = ~w13762 & ~w13776;
assign w13778 = w13762 & w13776;
assign w13779 = ~w13777 & ~w13778;
assign w13780 = b[40] & w2436;
assign w13781 = b[39] & ~w2622;
assign w13782 = b[41] & w2438;
assign w13783 = w2432 & w5302;
assign w13784 = ~w13780 & ~w13781;
assign w13785 = ~w13782 & w13784;
assign w13786 = ~w13783 & w13785;
assign w13787 = a[29] & ~w13786;
assign w13788 = ~a[29] & w13786;
assign w13789 = ~w13787 & ~w13788;
assign w13790 = (~w13426 & ~w13428) | (~w13426 & w25019) | (~w13428 & w25019);
assign w13791 = w13789 & ~w13790;
assign w13792 = ~w13789 & w13790;
assign w13793 = ~w13791 & ~w13792;
assign w13794 = w13779 & w13793;
assign w13795 = ~w13779 & ~w13793;
assign w13796 = ~w13794 & ~w13795;
assign w13797 = ~w13443 & ~w13446;
assign w13798 = b[44] & w1957;
assign w13799 = b[42] & ~w2114;
assign w13800 = b[43] & w1955;
assign w13801 = w1951 & w6069;
assign w13802 = ~w13798 & ~w13799;
assign w13803 = ~w13800 & w13802;
assign w13804 = ~w13801 & w13803;
assign w13805 = a[26] & ~w13804;
assign w13806 = ~a[26] & w13804;
assign w13807 = ~w13805 & ~w13806;
assign w13808 = ~w13797 & w13807;
assign w13809 = w13797 & ~w13807;
assign w13810 = ~w13808 & ~w13809;
assign w13811 = w13796 & w13810;
assign w13812 = ~w13796 & ~w13810;
assign w13813 = ~w13811 & ~w13812;
assign w13814 = w13590 & w13813;
assign w13815 = ~w13590 & ~w13813;
assign w13816 = ~w13814 & ~w13815;
assign w13817 = b[48] & ~w1272;
assign w13818 = b[49] & w1154;
assign w13819 = b[50] & w1156;
assign w13820 = w1150 & w7759;
assign w13821 = ~w13817 & ~w13818;
assign w13822 = ~w13819 & w13821;
assign w13823 = ~w13820 & w13822;
assign w13824 = a[20] & ~w13823;
assign w13825 = ~a[20] & w13823;
assign w13826 = ~w13824 & ~w13825;
assign w13827 = ~w13477 & ~w13480;
assign w13828 = w13826 & ~w13827;
assign w13829 = ~w13826 & w13827;
assign w13830 = ~w13828 & ~w13829;
assign w13831 = w13816 & w13830;
assign w13832 = ~w13816 & ~w13830;
assign w13833 = ~w13831 & ~w13832;
assign w13834 = ~w13240 & ~w13483;
assign w13835 = b[53] & w834;
assign w13836 = b[51] & ~w934;
assign w13837 = b[52] & w838;
assign w13838 = w832 & w8683;
assign w13839 = ~w13835 & ~w13836;
assign w13840 = ~w13837 & w13839;
assign w13841 = ~w13838 & w13840;
assign w13842 = a[17] & ~w13841;
assign w13843 = ~a[17] & w13841;
assign w13844 = ~w13842 & ~w13843;
assign w13845 = ~w13834 & w13844;
assign w13846 = w13834 & ~w13844;
assign w13847 = ~w13845 & ~w13846;
assign w13848 = w13833 & w13847;
assign w13849 = ~w13833 & ~w13847;
assign w13850 = ~w13848 & ~w13849;
assign w13851 = b[55] & w573;
assign w13852 = b[54] & ~w649;
assign w13853 = b[56] & w575;
assign w13854 = w569 & w9657;
assign w13855 = ~w13851 & ~w13852;
assign w13856 = ~w13853 & w13855;
assign w13857 = ~w13854 & w13856;
assign w13858 = a[14] & ~w13857;
assign w13859 = ~a[14] & w13857;
assign w13860 = ~w13858 & ~w13859;
assign w13861 = ~w13497 & ~w13500;
assign w13862 = w13860 & ~w13861;
assign w13863 = ~w13860 & w13861;
assign w13864 = ~w13862 & ~w13863;
assign w13865 = w13850 & w13864;
assign w13866 = ~w13850 & ~w13864;
assign w13867 = ~w13865 & ~w13866;
assign w13868 = w13576 & w13867;
assign w13869 = ~w13576 & ~w13867;
assign w13870 = ~w13868 & ~w13869;
assign w13871 = ~w13517 & ~w13520;
assign w13872 = b[62] & w185;
assign w13873 = b[60] & ~w237;
assign w13874 = b[61] & w183;
assign w13875 = w179 & w11763;
assign w13876 = ~w13872 & ~w13873;
assign w13877 = ~w13874 & w13876;
assign w13878 = ~w13875 & w13877;
assign w13879 = a[8] & ~w13878;
assign w13880 = ~a[8] & w13878;
assign w13881 = ~w13879 & ~w13880;
assign w13882 = ~w13871 & w13881;
assign w13883 = w13871 & ~w13881;
assign w13884 = ~w13882 & ~w13883;
assign w13885 = w13870 & w13884;
assign w13886 = ~w13870 & ~w13884;
assign w13887 = ~w13885 & ~w13886;
assign w13888 = ~w13534 & ~w13537;
assign w13889 = w66 & ~w12154;
assign w13890 = ~w103 & ~w13889;
assign w13891 = b[63] & ~w13890;
assign w13892 = ~a[5] & ~w13891;
assign w13893 = a[5] & w13891;
assign w13894 = ~w13892 & ~w13893;
assign w13895 = ~w13888 & w13894;
assign w13896 = w13888 & ~w13894;
assign w13897 = ~w13895 & ~w13896;
assign w13898 = w13887 & w13897;
assign w13899 = ~w13887 & ~w13897;
assign w13900 = ~w13898 & ~w13899;
assign w13901 = w13562 & ~w13900;
assign w13902 = ~w13562 & w13900;
assign w13903 = ~w13901 & ~w13902;
assign w13904 = (~w12865 & w24706) | (~w12865 & w24707) | (w24706 & w24707);
assign w13905 = w13903 & ~w13904;
assign w13906 = ~w13903 & w13904;
assign w13907 = ~w13905 & ~w13906;
assign w13908 = (~w12865 & w25437) | (~w12865 & w25438) | (w25437 & w25438);
assign w13909 = ~w13895 & ~w13898;
assign w13910 = ~w13747 & ~w13760;
assign w13911 = b[34] & w3785;
assign w13912 = b[35] & w3578;
assign w13913 = b[36] & w3580;
assign w13914 = w3573 & w4129;
assign w13915 = ~w13912 & ~w13913;
assign w13916 = ~w13911 & w13915;
assign w13917 = ~w13914 & w13916;
assign w13918 = a[35] & ~w13917;
assign w13919 = ~a[35] & w13917;
assign w13920 = ~w13918 & ~w13919;
assign w13921 = ~w13740 & ~w13744;
assign w13922 = b[31] & w4453;
assign w13923 = b[32] & w4241;
assign w13924 = b[33] & w4243;
assign w13925 = w3499 & w4236;
assign w13926 = ~w13923 & ~w13924;
assign w13927 = ~w13922 & w13926;
assign w13928 = ~w13925 & w13927;
assign w13929 = a[38] & ~w13928;
assign w13930 = ~a[38] & w13928;
assign w13931 = ~w13929 & ~w13930;
assign w13932 = ~w13723 & ~w13736;
assign w13933 = ~w13699 & ~w13712;
assign w13934 = b[22] & w6732;
assign w13935 = b[23] & w6474;
assign w13936 = b[24] & w6476;
assign w13937 = w1895 & w6469;
assign w13938 = ~w13935 & ~w13936;
assign w13939 = ~w13934 & w13938;
assign w13940 = ~w13937 & w13939;
assign w13941 = a[47] & ~w13940;
assign w13942 = ~a[47] & w13940;
assign w13943 = ~w13941 & ~w13942;
assign w13944 = ~w13682 & ~w13696;
assign w13945 = ~w13659 & ~w13672;
assign w13946 = b[13] & w9482;
assign w13947 = b[14] & w9165;
assign w13948 = b[15] & w9160;
assign w13949 = ~w799 & w9158;
assign w13950 = ~w13947 & ~w13948;
assign w13951 = ~w13946 & w13950;
assign w13952 = ~w13949 & w13951;
assign w13953 = a[56] & ~w13952;
assign w13954 = ~a[56] & w13952;
assign w13955 = ~w13953 & ~w13954;
assign w13956 = ~w13642 & ~w13656;
assign w13957 = ~w13626 & ~w13639;
assign w13958 = b[5] & w11921;
assign w13959 = b[6] & w11923;
assign w13960 = ~w13958 & ~w13959;
assign w13961 = ~a[2] & ~a[5];
assign w13962 = a[2] & a[5];
assign w13963 = ~w13961 & ~w13962;
assign w13964 = ~w13960 & w13963;
assign w13965 = w13960 & ~w13963;
assign w13966 = ~w13964 & ~w13965;
assign w13967 = w13957 & ~w13966;
assign w13968 = ~w13957 & w13966;
assign w13969 = ~w13967 & ~w13968;
assign w13970 = b[7] & w11561;
assign w13971 = b[9] & w11196;
assign w13972 = b[8] & w11194;
assign w13973 = w322 & w11189;
assign w13974 = ~w13971 & ~w13972;
assign w13975 = ~w13970 & w13974;
assign w13976 = ~w13973 & w13975;
assign w13977 = a[62] & ~w13976;
assign w13978 = ~a[62] & w13976;
assign w13979 = ~w13977 & ~w13978;
assign w13980 = ~w13969 & ~w13979;
assign w13981 = w13969 & w13979;
assign w13982 = ~w13980 & ~w13981;
assign w13983 = b[10] & w10496;
assign w13984 = b[11] & w10146;
assign w13985 = b[12] & w10148;
assign w13986 = w536 & w10141;
assign w13987 = ~w13984 & ~w13985;
assign w13988 = ~w13983 & w13987;
assign w13989 = ~w13986 & w13988;
assign w13990 = a[59] & ~w13989;
assign w13991 = ~a[59] & w13989;
assign w13992 = ~w13990 & ~w13991;
assign w13993 = ~w13982 & ~w13992;
assign w13994 = w13982 & w13992;
assign w13995 = ~w13993 & ~w13994;
assign w13996 = ~w13956 & w13995;
assign w13997 = w13956 & ~w13995;
assign w13998 = ~w13996 & ~w13997;
assign w13999 = w13955 & w13998;
assign w14000 = ~w13955 & ~w13998;
assign w14001 = ~w13999 & ~w14000;
assign w14002 = w13945 & ~w14001;
assign w14003 = ~w13945 & w14001;
assign w14004 = ~w14002 & ~w14003;
assign w14005 = b[16] & w8515;
assign w14006 = b[17] & w8200;
assign w14007 = b[18] & w8202;
assign w14008 = ~w1108 & w8195;
assign w14009 = ~w14006 & ~w14007;
assign w14010 = ~w14005 & w14009;
assign w14011 = ~w14008 & w14010;
assign w14012 = a[53] & ~w14011;
assign w14013 = ~a[53] & w14011;
assign w14014 = ~w14012 & ~w14013;
assign w14015 = w14004 & w14014;
assign w14016 = ~w14004 & ~w14014;
assign w14017 = ~w14015 & ~w14016;
assign w14018 = ~w13676 & ~w13679;
assign w14019 = ~w14017 & w14018;
assign w14020 = w14017 & ~w14018;
assign w14021 = ~w14019 & ~w14020;
assign w14022 = b[19] & w7586;
assign w14023 = b[20] & w7307;
assign w14024 = b[21] & w7314;
assign w14025 = w1467 & w7312;
assign w14026 = ~w14023 & ~w14024;
assign w14027 = ~w14022 & w14026;
assign w14028 = ~w14025 & w14027;
assign w14029 = a[50] & ~w14028;
assign w14030 = ~a[50] & w14028;
assign w14031 = ~w14029 & ~w14030;
assign w14032 = w14021 & w14031;
assign w14033 = ~w14021 & ~w14031;
assign w14034 = ~w14032 & ~w14033;
assign w14035 = ~w13944 & w14034;
assign w14036 = w13944 & ~w14034;
assign w14037 = ~w14035 & ~w14036;
assign w14038 = w13943 & w14037;
assign w14039 = ~w13943 & ~w14037;
assign w14040 = ~w14038 & ~w14039;
assign w14041 = w13933 & ~w14040;
assign w14042 = ~w13933 & w14040;
assign w14043 = ~w14041 & ~w14042;
assign w14044 = b[25] & w5939;
assign w14045 = b[26] & w5670;
assign w14046 = b[27] & w5665;
assign w14047 = w2378 & w5663;
assign w14048 = ~w14045 & ~w14046;
assign w14049 = ~w14044 & w14048;
assign w14050 = ~w14047 & w14049;
assign w14051 = a[44] & ~w14050;
assign w14052 = ~a[44] & w14050;
assign w14053 = ~w14051 & ~w14052;
assign w14054 = w14043 & w14053;
assign w14055 = ~w14043 & ~w14053;
assign w14056 = ~w14054 & ~w14055;
assign w14057 = ~w13716 & ~w13719;
assign w14058 = ~w14056 & w14057;
assign w14059 = w14056 & ~w14057;
assign w14060 = ~w14058 & ~w14059;
assign w14061 = b[28] & w5167;
assign w14062 = b[29] & w4918;
assign w14063 = b[30] & w4925;
assign w14064 = ~w2908 & w4923;
assign w14065 = ~w14062 & ~w14063;
assign w14066 = ~w14061 & w14065;
assign w14067 = ~w14064 & w14066;
assign w14068 = a[41] & ~w14067;
assign w14069 = ~a[41] & w14067;
assign w14070 = ~w14068 & ~w14069;
assign w14071 = ~w14060 & ~w14070;
assign w14072 = w14060 & w14070;
assign w14073 = ~w14071 & ~w14072;
assign w14074 = w13932 & w14073;
assign w14075 = ~w13932 & ~w14073;
assign w14076 = ~w14074 & ~w14075;
assign w14077 = w13931 & ~w14076;
assign w14078 = ~w13931 & w14076;
assign w14079 = ~w14077 & ~w14078;
assign w14080 = ~w13921 & w14079;
assign w14081 = w13921 & ~w14079;
assign w14082 = ~w14080 & ~w14081;
assign w14083 = w13920 & w14082;
assign w14084 = ~w13920 & ~w14082;
assign w14085 = ~w14083 & ~w14084;
assign w14086 = w13910 & ~w14085;
assign w14087 = ~w13910 & w14085;
assign w14088 = ~w14086 & ~w14087;
assign w14089 = b[37] & w3177;
assign w14090 = b[38] & w2973;
assign w14091 = b[39] & w2978;
assign w14092 = w2980 & ~w4812;
assign w14093 = ~w14090 & ~w14091;
assign w14094 = ~w14089 & w14093;
assign w14095 = ~w14092 & w14094;
assign w14096 = a[32] & ~w14095;
assign w14097 = ~a[32] & w14095;
assign w14098 = ~w14096 & ~w14097;
assign w14099 = (~w13774 & ~w13776) | (~w13774 & w24708) | (~w13776 & w24708);
assign w14100 = w14098 & ~w14099;
assign w14101 = ~w14098 & w14099;
assign w14102 = ~w14100 & ~w14101;
assign w14103 = w14088 & w14102;
assign w14104 = ~w14088 & ~w14102;
assign w14105 = ~w14103 & ~w14104;
assign w14106 = b[41] & w2436;
assign w14107 = b[42] & w2438;
assign w14108 = b[40] & ~w2622;
assign w14109 = w2432 & w5548;
assign w14110 = ~w14106 & ~w14107;
assign w14111 = ~w14108 & w14110;
assign w14112 = ~w14109 & w14111;
assign w14113 = a[29] & ~w14112;
assign w14114 = ~a[29] & w14112;
assign w14115 = ~w14113 & ~w14114;
assign w14116 = (~w13791 & ~w13793) | (~w13791 & w24709) | (~w13793 & w24709);
assign w14117 = w14115 & ~w14116;
assign w14118 = ~w14115 & w14116;
assign w14119 = ~w14117 & ~w14118;
assign w14120 = w14105 & w14119;
assign w14121 = ~w14105 & ~w14119;
assign w14122 = ~w14120 & ~w14121;
assign w14123 = (~w13808 & ~w13810) | (~w13808 & w24710) | (~w13810 & w24710);
assign w14124 = b[44] & w1955;
assign w14125 = b[43] & ~w2114;
assign w14126 = b[45] & w1957;
assign w14127 = w1951 & w6334;
assign w14128 = ~w14124 & ~w14125;
assign w14129 = ~w14126 & w14128;
assign w14130 = ~w14127 & w14129;
assign w14131 = a[26] & ~w14130;
assign w14132 = ~a[26] & w14130;
assign w14133 = ~w14131 & ~w14132;
assign w14134 = ~w14123 & w14133;
assign w14135 = w14123 & ~w14133;
assign w14136 = ~w14134 & ~w14135;
assign w14137 = ~w14122 & ~w14136;
assign w14138 = w14122 & w14136;
assign w14139 = ~w14137 & ~w14138;
assign w14140 = b[46] & ~w1676;
assign w14141 = b[48] & w1519;
assign w14142 = b[47] & w1517;
assign w14143 = w1513 & ~w7170;
assign w14144 = ~w14140 & ~w14141;
assign w14145 = ~w14142 & w14144;
assign w14146 = ~w14143 & w14145;
assign w14147 = a[23] & ~w14146;
assign w14148 = ~a[23] & w14146;
assign w14149 = ~w14147 & ~w14148;
assign w14150 = (~w13588 & ~w13590) | (~w13588 & w24711) | (~w13590 & w24711);
assign w14151 = w14149 & ~w14150;
assign w14152 = ~w14149 & w14150;
assign w14153 = ~w14151 & ~w14152;
assign w14154 = w14139 & w14153;
assign w14155 = ~w14139 & ~w14153;
assign w14156 = ~w14154 & ~w14155;
assign w14157 = b[49] & ~w1272;
assign w14158 = b[50] & w1154;
assign w14159 = b[51] & w1156;
assign w14160 = w1150 & ~w8058;
assign w14161 = ~w14157 & ~w14158;
assign w14162 = ~w14159 & w14161;
assign w14163 = ~w14160 & w14162;
assign w14164 = a[20] & ~w14163;
assign w14165 = ~a[20] & w14163;
assign w14166 = ~w14164 & ~w14165;
assign w14167 = (~w13828 & ~w13830) | (~w13828 & w24712) | (~w13830 & w24712);
assign w14168 = w14166 & ~w14167;
assign w14169 = ~w14166 & w14167;
assign w14170 = ~w14168 & ~w14169;
assign w14171 = ~w14156 & ~w14170;
assign w14172 = w14156 & w14170;
assign w14173 = ~w14171 & ~w14172;
assign w14174 = (~w13845 & ~w13847) | (~w13845 & w24713) | (~w13847 & w24713);
assign w14175 = b[52] & ~w934;
assign w14176 = b[54] & w834;
assign w14177 = b[53] & w838;
assign w14178 = w832 & ~w8998;
assign w14179 = ~w14175 & ~w14176;
assign w14180 = ~w14177 & w14179;
assign w14181 = ~w14178 & w14180;
assign w14182 = a[17] & ~w14181;
assign w14183 = ~a[17] & w14181;
assign w14184 = ~w14182 & ~w14183;
assign w14185 = ~w14174 & w14184;
assign w14186 = w14174 & ~w14184;
assign w14187 = ~w14185 & ~w14186;
assign w14188 = w14173 & w14187;
assign w14189 = ~w14173 & ~w14187;
assign w14190 = ~w14188 & ~w14189;
assign w14191 = b[57] & w575;
assign w14192 = b[56] & w573;
assign w14193 = b[55] & ~w649;
assign w14194 = w569 & ~w9992;
assign w14195 = ~w14191 & ~w14192;
assign w14196 = ~w14193 & w14195;
assign w14197 = ~w14194 & w14196;
assign w14198 = a[14] & ~w14197;
assign w14199 = ~a[14] & w14197;
assign w14200 = ~w14198 & ~w14199;
assign w14201 = (~w13862 & ~w13864) | (~w13862 & w24714) | (~w13864 & w24714);
assign w14202 = w14200 & ~w14201;
assign w14203 = ~w14200 & w14201;
assign w14204 = ~w14202 & ~w14203;
assign w14205 = ~w14190 & ~w14204;
assign w14206 = w14190 & w14204;
assign w14207 = ~w14205 & ~w14206;
assign w14208 = b[59] & w358;
assign w14209 = b[60] & w360;
assign w14210 = b[58] & ~w419;
assign w14211 = w354 & w11035;
assign w14212 = ~w14208 & ~w14209;
assign w14213 = ~w14210 & w14212;
assign w14214 = ~w14211 & w14213;
assign w14215 = a[11] & ~w14214;
assign w14216 = ~a[11] & w14214;
assign w14217 = ~w14215 & ~w14216;
assign w14218 = (~w13574 & ~w13576) | (~w13574 & w24715) | (~w13576 & w24715);
assign w14219 = w14217 & ~w14218;
assign w14220 = ~w14217 & w14218;
assign w14221 = ~w14219 & ~w14220;
assign w14222 = w14207 & w14221;
assign w14223 = ~w14207 & ~w14221;
assign w14224 = ~w14222 & ~w14223;
assign w14225 = (~w13882 & ~w13884) | (~w13882 & w24716) | (~w13884 & w24716);
assign w14226 = b[61] & ~w237;
assign w14227 = b[62] & w183;
assign w14228 = b[63] & w185;
assign w14229 = w179 & w12132;
assign w14230 = ~w14226 & ~w14227;
assign w14231 = ~w14228 & w14230;
assign w14232 = ~w14229 & w14231;
assign w14233 = a[8] & ~w14232;
assign w14234 = ~a[8] & w14232;
assign w14235 = ~w14233 & ~w14234;
assign w14236 = ~w14225 & w14235;
assign w14237 = w14225 & ~w14235;
assign w14238 = ~w14236 & ~w14237;
assign w14239 = w14224 & w14238;
assign w14240 = ~w14224 & ~w14238;
assign w14241 = ~w14239 & ~w14240;
assign w14242 = ~w13909 & w14241;
assign w14243 = w13909 & ~w14241;
assign w14244 = ~w14242 & ~w14243;
assign w14245 = ~w13908 & ~w14244;
assign w14246 = w13908 & w14244;
assign w14247 = ~w14245 & ~w14246;
assign w14248 = ~w14236 & ~w14239;
assign w14249 = b[59] & ~w419;
assign w14250 = b[61] & w360;
assign w14251 = b[60] & w358;
assign w14252 = w354 & w11400;
assign w14253 = ~w14249 & ~w14250;
assign w14254 = ~w14251 & w14253;
assign w14255 = ~w14252 & w14254;
assign w14256 = a[11] & ~w14255;
assign w14257 = ~a[11] & w14255;
assign w14258 = ~w14256 & ~w14257;
assign w14259 = (~w14202 & ~w14204) | (~w14202 & w25439) | (~w14204 & w25439);
assign w14260 = w14258 & ~w14259;
assign w14261 = ~w14258 & w14259;
assign w14262 = ~w14260 & ~w14261;
assign w14263 = b[50] & ~w1272;
assign w14264 = b[52] & w1156;
assign w14265 = b[51] & w1154;
assign w14266 = w1150 & ~w8371;
assign w14267 = ~w14263 & ~w14264;
assign w14268 = ~w14265 & w14267;
assign w14269 = ~w14266 & w14268;
assign w14270 = a[20] & ~w14269;
assign w14271 = ~a[20] & w14269;
assign w14272 = ~w14270 & ~w14271;
assign w14273 = (~w14151 & ~w14153) | (~w14151 & w25440) | (~w14153 & w25440);
assign w14274 = w14272 & ~w14273;
assign w14275 = ~w14272 & w14273;
assign w14276 = ~w14274 & ~w14275;
assign w14277 = b[35] & w3785;
assign w14278 = b[36] & w3578;
assign w14279 = b[37] & w3580;
assign w14280 = w3573 & ~w4357;
assign w14281 = ~w14278 & ~w14279;
assign w14282 = ~w14277 & w14281;
assign w14283 = ~w14280 & w14282;
assign w14284 = a[35] & ~w14283;
assign w14285 = ~a[35] & w14283;
assign w14286 = ~w14284 & ~w14285;
assign w14287 = ~w14077 & ~w14080;
assign w14288 = b[32] & w4453;
assign w14289 = b[34] & w4243;
assign w14290 = b[33] & w4241;
assign w14291 = ~w3710 & w4236;
assign w14292 = ~w14289 & ~w14290;
assign w14293 = ~w14288 & w14292;
assign w14294 = ~w14291 & w14293;
assign w14295 = a[38] & ~w14294;
assign w14296 = ~a[38] & w14294;
assign w14297 = ~w14295 & ~w14296;
assign w14298 = b[29] & w5167;
assign w14299 = b[31] & w4925;
assign w14300 = b[30] & w4918;
assign w14301 = ~w3112 & w4923;
assign w14302 = ~w14299 & ~w14300;
assign w14303 = ~w14298 & w14302;
assign w14304 = ~w14301 & w14303;
assign w14305 = a[41] & ~w14304;
assign w14306 = ~a[41] & w14304;
assign w14307 = ~w14305 & ~w14306;
assign w14308 = b[26] & w5939;
assign w14309 = b[27] & w5670;
assign w14310 = b[28] & w5665;
assign w14311 = w2559 & w5663;
assign w14312 = ~w14309 & ~w14310;
assign w14313 = ~w14308 & w14312;
assign w14314 = ~w14311 & w14313;
assign w14315 = a[44] & ~w14314;
assign w14316 = ~a[44] & w14314;
assign w14317 = ~w14315 & ~w14316;
assign w14318 = b[23] & w6732;
assign w14319 = b[24] & w6474;
assign w14320 = b[25] & w6476;
assign w14321 = w2061 & w6469;
assign w14322 = ~w14319 & ~w14320;
assign w14323 = ~w14318 & w14322;
assign w14324 = ~w14321 & w14323;
assign w14325 = a[47] & ~w14324;
assign w14326 = ~a[47] & w14324;
assign w14327 = ~w14325 & ~w14326;
assign w14328 = b[20] & w7586;
assign w14329 = b[22] & w7314;
assign w14330 = b[21] & w7307;
assign w14331 = w1615 & w7312;
assign w14332 = ~w14329 & ~w14330;
assign w14333 = ~w14328 & w14332;
assign w14334 = ~w14331 & w14333;
assign w14335 = a[50] & ~w14334;
assign w14336 = ~a[50] & w14334;
assign w14337 = ~w14335 & ~w14336;
assign w14338 = b[17] & w8515;
assign w14339 = b[18] & w8200;
assign w14340 = b[19] & w8202;
assign w14341 = ~w1231 & w8195;
assign w14342 = ~w14339 & ~w14340;
assign w14343 = ~w14338 & w14342;
assign w14344 = ~w14341 & w14343;
assign w14345 = a[53] & ~w14344;
assign w14346 = ~a[53] & w14344;
assign w14347 = ~w14345 & ~w14346;
assign w14348 = b[14] & w9482;
assign w14349 = b[16] & w9160;
assign w14350 = b[15] & w9165;
assign w14351 = w905 & w9158;
assign w14352 = ~w14349 & ~w14350;
assign w14353 = ~w14348 & w14352;
assign w14354 = ~w14351 & w14353;
assign w14355 = a[56] & ~w14354;
assign w14356 = ~a[56] & w14354;
assign w14357 = ~w14355 & ~w14356;
assign w14358 = ~w13968 & ~w13981;
assign w14359 = ~w13961 & ~w13964;
assign w14360 = b[6] & w11921;
assign w14361 = b[7] & w11923;
assign w14362 = ~w14360 & ~w14361;
assign w14363 = w14359 & ~w14362;
assign w14364 = ~w14359 & w14362;
assign w14365 = ~w14363 & ~w14364;
assign w14366 = b[8] & w11561;
assign w14367 = b[9] & w11194;
assign w14368 = b[10] & w11196;
assign w14369 = w397 & w11189;
assign w14370 = ~w14367 & ~w14368;
assign w14371 = ~w14366 & w14370;
assign w14372 = ~w14369 & w14371;
assign w14373 = a[62] & ~w14372;
assign w14374 = ~a[62] & w14372;
assign w14375 = ~w14373 & ~w14374;
assign w14376 = w14365 & w14375;
assign w14377 = ~w14365 & ~w14375;
assign w14378 = ~w14376 & ~w14377;
assign w14379 = w14358 & ~w14378;
assign w14380 = ~w14358 & w14378;
assign w14381 = ~w14379 & ~w14380;
assign w14382 = b[11] & w10496;
assign w14383 = b[12] & w10146;
assign w14384 = b[13] & w10148;
assign w14385 = w628 & w10141;
assign w14386 = ~w14383 & ~w14384;
assign w14387 = ~w14382 & w14386;
assign w14388 = ~w14385 & w14387;
assign w14389 = a[59] & ~w14388;
assign w14390 = ~a[59] & w14388;
assign w14391 = ~w14389 & ~w14390;
assign w14392 = w14381 & w14391;
assign w14393 = ~w14381 & ~w14391;
assign w14394 = ~w14392 & ~w14393;
assign w14395 = ~w13994 & ~w13996;
assign w14396 = w14394 & ~w14395;
assign w14397 = ~w14394 & w14395;
assign w14398 = ~w14396 & ~w14397;
assign w14399 = w14357 & w14398;
assign w14400 = ~w14357 & ~w14398;
assign w14401 = ~w14399 & ~w14400;
assign w14402 = ~w13999 & ~w14003;
assign w14403 = w14401 & ~w14402;
assign w14404 = ~w14401 & w14402;
assign w14405 = ~w14403 & ~w14404;
assign w14406 = w14347 & w14405;
assign w14407 = ~w14347 & ~w14405;
assign w14408 = ~w14406 & ~w14407;
assign w14409 = ~w14015 & ~w14020;
assign w14410 = w14408 & ~w14409;
assign w14411 = ~w14408 & w14409;
assign w14412 = ~w14410 & ~w14411;
assign w14413 = w14337 & w14412;
assign w14414 = ~w14337 & ~w14412;
assign w14415 = ~w14413 & ~w14414;
assign w14416 = ~w14032 & ~w14035;
assign w14417 = w14415 & ~w14416;
assign w14418 = ~w14415 & w14416;
assign w14419 = ~w14417 & ~w14418;
assign w14420 = w14327 & w14419;
assign w14421 = ~w14327 & ~w14419;
assign w14422 = ~w14420 & ~w14421;
assign w14423 = ~w14038 & ~w14042;
assign w14424 = w14422 & ~w14423;
assign w14425 = ~w14422 & w14423;
assign w14426 = ~w14424 & ~w14425;
assign w14427 = w14317 & w14426;
assign w14428 = ~w14317 & ~w14426;
assign w14429 = ~w14427 & ~w14428;
assign w14430 = ~w14054 & ~w14059;
assign w14431 = w14429 & ~w14430;
assign w14432 = ~w14429 & w14430;
assign w14433 = ~w14431 & ~w14432;
assign w14434 = ~w14307 & ~w14433;
assign w14435 = w14307 & w14433;
assign w14436 = ~w14434 & ~w14435;
assign w14437 = ~w14071 & ~w14074;
assign w14438 = ~w14436 & ~w14437;
assign w14439 = w14436 & w14437;
assign w14440 = ~w14438 & ~w14439;
assign w14441 = w14297 & w14440;
assign w14442 = ~w14297 & ~w14440;
assign w14443 = ~w14441 & ~w14442;
assign w14444 = w14287 & ~w14443;
assign w14445 = ~w14287 & w14443;
assign w14446 = ~w14444 & ~w14445;
assign w14447 = ~w14286 & ~w14446;
assign w14448 = w14286 & w14446;
assign w14449 = ~w14447 & ~w14448;
assign w14450 = b[38] & w3177;
assign w14451 = b[40] & w2978;
assign w14452 = b[39] & w2973;
assign w14453 = w2980 & ~w5058;
assign w14454 = ~w14451 & ~w14452;
assign w14455 = ~w14450 & w14454;
assign w14456 = ~w14453 & w14455;
assign w14457 = a[32] & ~w14456;
assign w14458 = ~a[32] & w14456;
assign w14459 = ~w14457 & ~w14458;
assign w14460 = ~w14083 & ~w14087;
assign w14461 = w14459 & ~w14460;
assign w14462 = ~w14459 & w14460;
assign w14463 = ~w14461 & ~w14462;
assign w14464 = w14449 & w14463;
assign w14465 = ~w14449 & ~w14463;
assign w14466 = ~w14464 & ~w14465;
assign w14467 = b[43] & w2438;
assign w14468 = b[41] & ~w2622;
assign w14469 = b[42] & w2436;
assign w14470 = w2432 & w5811;
assign w14471 = ~w14467 & ~w14468;
assign w14472 = ~w14469 & w14471;
assign w14473 = ~w14470 & w14472;
assign w14474 = a[29] & ~w14473;
assign w14475 = ~a[29] & w14473;
assign w14476 = ~w14474 & ~w14475;
assign w14477 = (~w14100 & ~w14102) | (~w14100 & w25441) | (~w14102 & w25441);
assign w14478 = w14476 & ~w14477;
assign w14479 = ~w14476 & w14477;
assign w14480 = ~w14478 & ~w14479;
assign w14481 = w14466 & w14480;
assign w14482 = ~w14466 & ~w14480;
assign w14483 = ~w14481 & ~w14482;
assign w14484 = (~w14117 & ~w14119) | (~w14117 & w25442) | (~w14119 & w25442);
assign w14485 = b[46] & w1957;
assign w14486 = b[45] & w1955;
assign w14487 = b[44] & ~w2114;
assign w14488 = w1951 & ~w6613;
assign w14489 = ~w14485 & ~w14486;
assign w14490 = ~w14487 & w14489;
assign w14491 = ~w14488 & w14490;
assign w14492 = a[26] & ~w14491;
assign w14493 = ~a[26] & w14491;
assign w14494 = ~w14492 & ~w14493;
assign w14495 = ~w14484 & w14494;
assign w14496 = w14484 & ~w14494;
assign w14497 = ~w14495 & ~w14496;
assign w14498 = w14483 & w14497;
assign w14499 = ~w14483 & ~w14497;
assign w14500 = ~w14498 & ~w14499;
assign w14501 = b[49] & w1519;
assign w14502 = b[48] & w1517;
assign w14503 = b[47] & ~w1676;
assign w14504 = w1513 & ~w7468;
assign w14505 = ~w14501 & ~w14502;
assign w14506 = ~w14503 & w14505;
assign w14507 = ~w14504 & w14506;
assign w14508 = a[23] & ~w14507;
assign w14509 = ~a[23] & w14507;
assign w14510 = ~w14508 & ~w14509;
assign w14511 = (~w14134 & ~w14136) | (~w14134 & w25443) | (~w14136 & w25443);
assign w14512 = w14510 & ~w14511;
assign w14513 = ~w14510 & w14511;
assign w14514 = ~w14512 & ~w14513;
assign w14515 = w14500 & w14514;
assign w14516 = ~w14500 & ~w14514;
assign w14517 = ~w14515 & ~w14516;
assign w14518 = w14276 & w14517;
assign w14519 = ~w14276 & ~w14517;
assign w14520 = ~w14518 & ~w14519;
assign w14521 = b[53] & ~w934;
assign w14522 = b[54] & w838;
assign w14523 = b[55] & w834;
assign w14524 = w832 & ~w9330;
assign w14525 = ~w14521 & ~w14522;
assign w14526 = ~w14523 & w14525;
assign w14527 = ~w14524 & w14526;
assign w14528 = a[17] & ~w14527;
assign w14529 = ~a[17] & w14527;
assign w14530 = ~w14528 & ~w14529;
assign w14531 = (~w14168 & ~w14170) | (~w14168 & w25444) | (~w14170 & w25444);
assign w14532 = w14530 & ~w14531;
assign w14533 = ~w14530 & w14531;
assign w14534 = ~w14532 & ~w14533;
assign w14535 = w14520 & w14534;
assign w14536 = ~w14520 & ~w14534;
assign w14537 = ~w14535 & ~w14536;
assign w14538 = (~w14185 & ~w14187) | (~w14185 & w25445) | (~w14187 & w25445);
assign w14539 = b[57] & w573;
assign w14540 = b[58] & w575;
assign w14541 = b[56] & ~w649;
assign w14542 = w569 & ~w10339;
assign w14543 = ~w14539 & ~w14540;
assign w14544 = ~w14541 & w14543;
assign w14545 = ~w14542 & w14544;
assign w14546 = a[14] & ~w14545;
assign w14547 = ~a[14] & w14545;
assign w14548 = ~w14546 & ~w14547;
assign w14549 = ~w14538 & w14548;
assign w14550 = w14538 & ~w14548;
assign w14551 = ~w14549 & ~w14550;
assign w14552 = w14537 & w14551;
assign w14553 = ~w14537 & ~w14551;
assign w14554 = ~w14552 & ~w14553;
assign w14555 = w14262 & w14554;
assign w14556 = ~w14262 & ~w14554;
assign w14557 = ~w14555 & ~w14556;
assign w14558 = (~w14219 & ~w14221) | (~w14219 & w25446) | (~w14221 & w25446);
assign w14559 = b[62] & ~w237;
assign w14560 = b[63] & w183;
assign w14561 = w179 & w12156;
assign w14562 = ~w14559 & ~w14560;
assign w14563 = ~w14561 & w14562;
assign w14564 = ~a[8] & w14563;
assign w14565 = a[8] & ~w14563;
assign w14566 = ~w14564 & ~w14565;
assign w14567 = ~w14558 & w14566;
assign w14568 = w14558 & ~w14566;
assign w14569 = ~w14567 & ~w14568;
assign w14570 = w14557 & w14569;
assign w14571 = ~w14557 & ~w14569;
assign w14572 = ~w14570 & ~w14571;
assign w14573 = ~w14248 & w14572;
assign w14574 = w14248 & ~w14572;
assign w14575 = ~w14573 & ~w14574;
assign w14576 = (~w14243 & ~w13908) | (~w14243 & w24406) | (~w13908 & w24406);
assign w14577 = (~w13908 & w24407) | (~w13908 & w24408) | (w24407 & w24408);
assign w14578 = ~w14575 & ~w14576;
assign w14579 = ~w14577 & ~w14578;
assign w14580 = ~w14567 & ~w14570;
assign w14581 = b[50] & w1519;
assign w14582 = b[49] & w1517;
assign w14583 = b[48] & ~w1676;
assign w14584 = w1513 & w7759;
assign w14585 = ~w14581 & ~w14582;
assign w14586 = ~w14583 & w14585;
assign w14587 = ~w14584 & w14586;
assign w14588 = a[23] & ~w14587;
assign w14589 = ~a[23] & w14587;
assign w14590 = ~w14588 & ~w14589;
assign w14591 = ~w14495 & ~w14498;
assign w14592 = w14590 & ~w14591;
assign w14593 = ~w14590 & w14591;
assign w14594 = ~w14592 & ~w14593;
assign w14595 = b[46] & w1955;
assign w14596 = b[45] & ~w2114;
assign w14597 = b[47] & w1957;
assign w14598 = w1951 & w6889;
assign w14599 = ~w14595 & ~w14596;
assign w14600 = ~w14597 & w14599;
assign w14601 = ~w14598 & w14600;
assign w14602 = a[26] & ~w14601;
assign w14603 = ~a[26] & w14601;
assign w14604 = ~w14602 & ~w14603;
assign w14605 = ~w14478 & ~w14481;
assign w14606 = w14604 & ~w14605;
assign w14607 = ~w14604 & w14605;
assign w14608 = ~w14606 & ~w14607;
assign w14609 = b[36] & w3785;
assign w14610 = b[38] & w3580;
assign w14611 = b[37] & w3578;
assign w14612 = w3573 & w4582;
assign w14613 = ~w14610 & ~w14611;
assign w14614 = ~w14609 & w14613;
assign w14615 = ~w14612 & w14614;
assign w14616 = a[35] & ~w14615;
assign w14617 = ~a[35] & w14615;
assign w14618 = ~w14616 & ~w14617;
assign w14619 = b[30] & w5167;
assign w14620 = b[32] & w4925;
assign w14621 = b[31] & w4918;
assign w14622 = w3304 & w4923;
assign w14623 = ~w14620 & ~w14621;
assign w14624 = ~w14619 & w14623;
assign w14625 = ~w14622 & w14624;
assign w14626 = a[41] & ~w14625;
assign w14627 = ~a[41] & w14625;
assign w14628 = ~w14626 & ~w14627;
assign w14629 = ~w14410 & ~w14413;
assign w14630 = b[21] & w7586;
assign w14631 = b[23] & w7314;
assign w14632 = b[22] & w7307;
assign w14633 = w1755 & w7312;
assign w14634 = ~w14631 & ~w14632;
assign w14635 = ~w14630 & w14634;
assign w14636 = ~w14633 & w14635;
assign w14637 = a[50] & ~w14636;
assign w14638 = ~a[50] & w14636;
assign w14639 = ~w14637 & ~w14638;
assign w14640 = ~w14403 & ~w14406;
assign w14641 = b[18] & w8515;
assign w14642 = b[20] & w8202;
assign w14643 = b[19] & w8200;
assign w14644 = w1347 & w8195;
assign w14645 = ~w14642 & ~w14643;
assign w14646 = ~w14641 & w14645;
assign w14647 = ~w14644 & w14646;
assign w14648 = a[53] & ~w14647;
assign w14649 = ~a[53] & w14647;
assign w14650 = ~w14648 & ~w14649;
assign w14651 = ~w14380 & ~w14392;
assign w14652 = b[9] & w11561;
assign w14653 = b[10] & w11194;
assign w14654 = b[11] & w11196;
assign w14655 = w469 & w11189;
assign w14656 = ~w14653 & ~w14654;
assign w14657 = ~w14652 & w14656;
assign w14658 = ~w14655 & w14657;
assign w14659 = a[62] & ~w14658;
assign w14660 = ~a[62] & w14658;
assign w14661 = ~w14659 & ~w14660;
assign w14662 = ~w14364 & ~w14376;
assign w14663 = b[7] & w11921;
assign w14664 = b[8] & w11923;
assign w14665 = ~w14663 & ~w14664;
assign w14666 = w14362 & ~w14665;
assign w14667 = ~w14362 & w14665;
assign w14668 = ~w14666 & ~w14667;
assign w14669 = w14662 & w14668;
assign w14670 = ~w14662 & ~w14668;
assign w14671 = ~w14669 & ~w14670;
assign w14672 = w14661 & ~w14671;
assign w14673 = ~w14661 & w14671;
assign w14674 = ~w14672 & ~w14673;
assign w14675 = b[12] & w10496;
assign w14676 = b[13] & w10146;
assign w14677 = b[14] & w10148;
assign w14678 = w714 & w10141;
assign w14679 = ~w14676 & ~w14677;
assign w14680 = ~w14675 & w14679;
assign w14681 = ~w14678 & w14680;
assign w14682 = a[59] & ~w14681;
assign w14683 = ~a[59] & w14681;
assign w14684 = ~w14682 & ~w14683;
assign w14685 = w14674 & w14684;
assign w14686 = ~w14674 & ~w14684;
assign w14687 = ~w14685 & ~w14686;
assign w14688 = w14651 & ~w14687;
assign w14689 = ~w14651 & w14687;
assign w14690 = ~w14688 & ~w14689;
assign w14691 = b[15] & w9482;
assign w14692 = b[16] & w9165;
assign w14693 = b[17] & w9160;
assign w14694 = w1008 & w9158;
assign w14695 = ~w14692 & ~w14693;
assign w14696 = ~w14691 & w14695;
assign w14697 = ~w14694 & w14696;
assign w14698 = a[56] & ~w14697;
assign w14699 = ~a[56] & w14697;
assign w14700 = ~w14698 & ~w14699;
assign w14701 = w14690 & w14700;
assign w14702 = ~w14690 & ~w14700;
assign w14703 = ~w14701 & ~w14702;
assign w14704 = ~w14396 & ~w14399;
assign w14705 = w14703 & ~w14704;
assign w14706 = ~w14703 & w14704;
assign w14707 = ~w14705 & ~w14706;
assign w14708 = ~w14650 & ~w14707;
assign w14709 = w14650 & w14707;
assign w14710 = ~w14708 & ~w14709;
assign w14711 = w14640 & ~w14710;
assign w14712 = ~w14640 & w14710;
assign w14713 = ~w14711 & ~w14712;
assign w14714 = w14639 & w14713;
assign w14715 = ~w14639 & ~w14713;
assign w14716 = ~w14714 & ~w14715;
assign w14717 = w14629 & ~w14716;
assign w14718 = ~w14629 & w14716;
assign w14719 = ~w14717 & ~w14718;
assign w14720 = b[24] & w6732;
assign w14721 = b[26] & w6476;
assign w14722 = b[25] & w6474;
assign w14723 = w2219 & w6469;
assign w14724 = ~w14721 & ~w14722;
assign w14725 = ~w14720 & w14724;
assign w14726 = ~w14723 & w14725;
assign w14727 = a[47] & ~w14726;
assign w14728 = ~a[47] & w14726;
assign w14729 = ~w14727 & ~w14728;
assign w14730 = w14719 & w14729;
assign w14731 = ~w14719 & ~w14729;
assign w14732 = ~w14730 & ~w14731;
assign w14733 = ~w14417 & ~w14420;
assign w14734 = w14732 & ~w14733;
assign w14735 = ~w14732 & w14733;
assign w14736 = ~w14734 & ~w14735;
assign w14737 = b[27] & w5939;
assign w14738 = b[29] & w5665;
assign w14739 = b[28] & w5670;
assign w14740 = w2734 & w5663;
assign w14741 = ~w14738 & ~w14739;
assign w14742 = ~w14737 & w14741;
assign w14743 = ~w14740 & w14742;
assign w14744 = a[44] & ~w14743;
assign w14745 = ~a[44] & w14743;
assign w14746 = ~w14744 & ~w14745;
assign w14747 = w14736 & w14746;
assign w14748 = ~w14736 & ~w14746;
assign w14749 = ~w14747 & ~w14748;
assign w14750 = ~w14424 & ~w14427;
assign w14751 = w14749 & ~w14750;
assign w14752 = ~w14749 & w14750;
assign w14753 = ~w14751 & ~w14752;
assign w14754 = ~w14628 & ~w14753;
assign w14755 = w14628 & w14753;
assign w14756 = ~w14754 & ~w14755;
assign w14757 = ~w14431 & ~w14435;
assign w14758 = w14756 & ~w14757;
assign w14759 = ~w14756 & w14757;
assign w14760 = ~w14758 & ~w14759;
assign w14761 = b[33] & w4453;
assign w14762 = b[35] & w4243;
assign w14763 = b[34] & w4241;
assign w14764 = w3918 & w4236;
assign w14765 = ~w14762 & ~w14763;
assign w14766 = ~w14761 & w14765;
assign w14767 = ~w14764 & w14766;
assign w14768 = a[38] & ~w14767;
assign w14769 = ~a[38] & w14767;
assign w14770 = ~w14768 & ~w14769;
assign w14771 = w14760 & w14770;
assign w14772 = ~w14760 & ~w14770;
assign w14773 = ~w14771 & ~w14772;
assign w14774 = ~w14439 & ~w14441;
assign w14775 = w14773 & ~w14774;
assign w14776 = ~w14773 & w14774;
assign w14777 = ~w14775 & ~w14776;
assign w14778 = w14618 & w14777;
assign w14779 = ~w14618 & ~w14777;
assign w14780 = ~w14778 & ~w14779;
assign w14781 = b[39] & w3177;
assign w14782 = b[41] & w2978;
assign w14783 = b[40] & w2973;
assign w14784 = w2980 & w5302;
assign w14785 = ~w14782 & ~w14783;
assign w14786 = ~w14781 & w14785;
assign w14787 = ~w14784 & w14786;
assign w14788 = a[32] & ~w14787;
assign w14789 = ~a[32] & w14787;
assign w14790 = ~w14788 & ~w14789;
assign w14791 = ~w14445 & ~w14448;
assign w14792 = w14790 & ~w14791;
assign w14793 = ~w14790 & w14791;
assign w14794 = ~w14792 & ~w14793;
assign w14795 = w14780 & w14794;
assign w14796 = ~w14780 & ~w14794;
assign w14797 = ~w14795 & ~w14796;
assign w14798 = ~w14461 & ~w14464;
assign w14799 = b[44] & w2438;
assign w14800 = b[43] & w2436;
assign w14801 = b[42] & ~w2622;
assign w14802 = w2432 & w6069;
assign w14803 = ~w14799 & ~w14800;
assign w14804 = ~w14801 & w14803;
assign w14805 = ~w14802 & w14804;
assign w14806 = a[29] & ~w14805;
assign w14807 = ~a[29] & w14805;
assign w14808 = ~w14806 & ~w14807;
assign w14809 = ~w14798 & w14808;
assign w14810 = w14798 & ~w14808;
assign w14811 = ~w14809 & ~w14810;
assign w14812 = w14797 & w14811;
assign w14813 = ~w14797 & ~w14811;
assign w14814 = ~w14812 & ~w14813;
assign w14815 = w14608 & w14814;
assign w14816 = ~w14608 & ~w14814;
assign w14817 = ~w14815 & ~w14816;
assign w14818 = ~w14594 & ~w14817;
assign w14819 = w14594 & w14817;
assign w14820 = ~w14818 & ~w14819;
assign w14821 = ~w14512 & ~w14515;
assign w14822 = b[52] & w1154;
assign w14823 = b[51] & ~w1272;
assign w14824 = b[53] & w1156;
assign w14825 = w1150 & w8683;
assign w14826 = ~w14822 & ~w14823;
assign w14827 = ~w14824 & w14826;
assign w14828 = ~w14825 & w14827;
assign w14829 = a[20] & ~w14828;
assign w14830 = ~a[20] & w14828;
assign w14831 = ~w14829 & ~w14830;
assign w14832 = ~w14821 & w14831;
assign w14833 = w14821 & ~w14831;
assign w14834 = ~w14832 & ~w14833;
assign w14835 = w14820 & w14834;
assign w14836 = ~w14820 & ~w14834;
assign w14837 = ~w14835 & ~w14836;
assign w14838 = b[54] & ~w934;
assign w14839 = b[55] & w838;
assign w14840 = b[56] & w834;
assign w14841 = w832 & w9657;
assign w14842 = ~w14838 & ~w14839;
assign w14843 = ~w14840 & w14842;
assign w14844 = ~w14841 & w14843;
assign w14845 = a[17] & ~w14844;
assign w14846 = ~a[17] & w14844;
assign w14847 = ~w14845 & ~w14846;
assign w14848 = ~w14274 & ~w14518;
assign w14849 = w14847 & ~w14848;
assign w14850 = ~w14847 & w14848;
assign w14851 = ~w14849 & ~w14850;
assign w14852 = w14837 & w14851;
assign w14853 = ~w14837 & ~w14851;
assign w14854 = ~w14852 & ~w14853;
assign w14855 = b[58] & w573;
assign w14856 = b[59] & w575;
assign w14857 = b[57] & ~w649;
assign w14858 = w569 & w10371;
assign w14859 = ~w14855 & ~w14856;
assign w14860 = ~w14857 & w14859;
assign w14861 = ~w14858 & w14860;
assign w14862 = a[14] & ~w14861;
assign w14863 = ~a[14] & w14861;
assign w14864 = ~w14862 & ~w14863;
assign w14865 = ~w14532 & ~w14535;
assign w14866 = w14864 & ~w14865;
assign w14867 = ~w14864 & w14865;
assign w14868 = ~w14866 & ~w14867;
assign w14869 = w14854 & w14868;
assign w14870 = ~w14854 & ~w14868;
assign w14871 = ~w14869 & ~w14870;
assign w14872 = ~w14549 & ~w14552;
assign w14873 = b[62] & w360;
assign w14874 = b[60] & ~w419;
assign w14875 = b[61] & w358;
assign w14876 = w354 & w11763;
assign w14877 = ~w14873 & ~w14874;
assign w14878 = ~w14875 & w14877;
assign w14879 = ~w14876 & w14878;
assign w14880 = a[11] & ~w14879;
assign w14881 = ~a[11] & w14879;
assign w14882 = ~w14880 & ~w14881;
assign w14883 = ~w14872 & w14882;
assign w14884 = w14872 & ~w14882;
assign w14885 = ~w14883 & ~w14884;
assign w14886 = w14871 & w14885;
assign w14887 = ~w14871 & ~w14885;
assign w14888 = ~w14886 & ~w14887;
assign w14889 = ~w14260 & ~w14555;
assign w14890 = w179 & ~w12154;
assign w14891 = w237 & ~w14890;
assign w14892 = b[63] & ~w14891;
assign w14893 = ~a[8] & ~w14892;
assign w14894 = a[8] & w14892;
assign w14895 = ~w14893 & ~w14894;
assign w14896 = ~w14889 & w14895;
assign w14897 = w14889 & ~w14895;
assign w14898 = ~w14896 & ~w14897;
assign w14899 = w14888 & w14898;
assign w14900 = ~w14888 & ~w14898;
assign w14901 = ~w14899 & ~w14900;
assign w14902 = w14580 & ~w14901;
assign w14903 = ~w14580 & w14901;
assign w14904 = ~w14902 & ~w14903;
assign w14905 = ~w14573 & ~w14577;
assign w14906 = (w14904 & w14577) | (w14904 & w24409) | (w14577 & w24409);
assign w14907 = ~w14904 & w14905;
assign w14908 = ~w14906 & ~w14907;
assign w14909 = ~w14896 & ~w14899;
assign w14910 = b[57] & w834;
assign w14911 = b[56] & w838;
assign w14912 = b[55] & ~w934;
assign w14913 = w832 & ~w9992;
assign w14914 = ~w14910 & ~w14911;
assign w14915 = ~w14912 & w14914;
assign w14916 = ~w14913 & w14915;
assign w14917 = a[17] & ~w14916;
assign w14918 = ~a[17] & w14916;
assign w14919 = ~w14917 & ~w14918;
assign w14920 = ~w14849 & ~w14852;
assign w14921 = w14919 & ~w14920;
assign w14922 = ~w14919 & w14920;
assign w14923 = ~w14921 & ~w14922;
assign w14924 = b[46] & ~w2114;
assign w14925 = b[48] & w1957;
assign w14926 = b[47] & w1955;
assign w14927 = w1951 & ~w7170;
assign w14928 = ~w14924 & ~w14925;
assign w14929 = ~w14926 & w14928;
assign w14930 = ~w14927 & w14929;
assign w14931 = a[26] & ~w14930;
assign w14932 = ~a[26] & w14930;
assign w14933 = ~w14931 & ~w14932;
assign w14934 = ~w14606 & ~w14815;
assign w14935 = w14933 & ~w14934;
assign w14936 = ~w14933 & w14934;
assign w14937 = ~w14935 & ~w14936;
assign w14938 = ~w14809 & ~w14812;
assign w14939 = b[43] & ~w2622;
assign w14940 = b[44] & w2436;
assign w14941 = b[45] & w2438;
assign w14942 = w2432 & w6334;
assign w14943 = ~w14939 & ~w14940;
assign w14944 = ~w14941 & w14943;
assign w14945 = ~w14942 & w14944;
assign w14946 = a[29] & ~w14945;
assign w14947 = ~a[29] & w14945;
assign w14948 = ~w14946 & ~w14947;
assign w14949 = ~w14938 & w14948;
assign w14950 = w14938 & ~w14948;
assign w14951 = ~w14949 & ~w14950;
assign w14952 = ~w14792 & ~w14795;
assign w14953 = b[40] & w3177;
assign w14954 = b[42] & w2978;
assign w14955 = b[41] & w2973;
assign w14956 = w2980 & w5548;
assign w14957 = ~w14954 & ~w14955;
assign w14958 = ~w14953 & w14957;
assign w14959 = ~w14956 & w14958;
assign w14960 = a[32] & ~w14959;
assign w14961 = ~a[32] & w14959;
assign w14962 = ~w14960 & ~w14961;
assign w14963 = ~w14952 & w14962;
assign w14964 = w14952 & ~w14962;
assign w14965 = ~w14963 & ~w14964;
assign w14966 = ~w14758 & ~w14771;
assign w14967 = b[34] & w4453;
assign w14968 = b[35] & w4241;
assign w14969 = b[36] & w4243;
assign w14970 = w4129 & w4236;
assign w14971 = ~w14968 & ~w14969;
assign w14972 = ~w14967 & w14971;
assign w14973 = ~w14970 & w14972;
assign w14974 = a[38] & ~w14973;
assign w14975 = ~a[38] & w14973;
assign w14976 = ~w14974 & ~w14975;
assign w14977 = ~w14751 & ~w14755;
assign w14978 = b[31] & w5167;
assign w14979 = b[32] & w4918;
assign w14980 = b[33] & w4925;
assign w14981 = w3499 & w4923;
assign w14982 = ~w14979 & ~w14980;
assign w14983 = ~w14978 & w14982;
assign w14984 = ~w14981 & w14983;
assign w14985 = a[41] & ~w14984;
assign w14986 = ~a[41] & w14984;
assign w14987 = ~w14985 & ~w14986;
assign w14988 = ~w14734 & ~w14747;
assign w14989 = ~w14718 & ~w14730;
assign w14990 = b[25] & w6732;
assign w14991 = b[27] & w6476;
assign w14992 = b[26] & w6474;
assign w14993 = w2378 & w6469;
assign w14994 = ~w14991 & ~w14992;
assign w14995 = ~w14990 & w14994;
assign w14996 = ~w14993 & w14995;
assign w14997 = a[47] & ~w14996;
assign w14998 = ~a[47] & w14996;
assign w14999 = ~w14997 & ~w14998;
assign w15000 = ~w14712 & ~w14714;
assign w15001 = b[22] & w7586;
assign w15002 = b[24] & w7314;
assign w15003 = b[23] & w7307;
assign w15004 = w1895 & w7312;
assign w15005 = ~w15002 & ~w15003;
assign w15006 = ~w15001 & w15005;
assign w15007 = ~w15004 & w15006;
assign w15008 = a[50] & ~w15007;
assign w15009 = ~a[50] & w15007;
assign w15010 = ~w15008 & ~w15009;
assign w15011 = ~w14672 & ~w14685;
assign w15012 = b[8] & w11921;
assign w15013 = b[9] & w11923;
assign w15014 = ~w15012 & ~w15013;
assign w15015 = ~a[8] & ~w14665;
assign w15016 = a[8] & w14665;
assign w15017 = ~w15015 & ~w15016;
assign w15018 = ~w15014 & w15017;
assign w15019 = w15014 & ~w15017;
assign w15020 = ~w15018 & ~w15019;
assign w15021 = ~w14666 & ~w14669;
assign w15022 = ~w15020 & ~w15021;
assign w15023 = w15020 & w15021;
assign w15024 = ~w15022 & ~w15023;
assign w15025 = b[10] & w11561;
assign w15026 = b[12] & w11196;
assign w15027 = b[11] & w11194;
assign w15028 = w536 & w11189;
assign w15029 = ~w15026 & ~w15027;
assign w15030 = ~w15025 & w15029;
assign w15031 = ~w15028 & w15030;
assign w15032 = a[62] & ~w15031;
assign w15033 = ~a[62] & w15031;
assign w15034 = ~w15032 & ~w15033;
assign w15035 = ~w15024 & ~w15034;
assign w15036 = w15024 & w15034;
assign w15037 = ~w15035 & ~w15036;
assign w15038 = b[13] & w10496;
assign w15039 = b[14] & w10146;
assign w15040 = b[15] & w10148;
assign w15041 = ~w799 & w10141;
assign w15042 = ~w15039 & ~w15040;
assign w15043 = ~w15038 & w15042;
assign w15044 = ~w15041 & w15043;
assign w15045 = a[59] & ~w15044;
assign w15046 = ~a[59] & w15044;
assign w15047 = ~w15045 & ~w15046;
assign w15048 = w15037 & w15047;
assign w15049 = ~w15037 & ~w15047;
assign w15050 = ~w15048 & ~w15049;
assign w15051 = ~w15011 & w15050;
assign w15052 = w15011 & ~w15050;
assign w15053 = ~w15051 & ~w15052;
assign w15054 = b[16] & w9482;
assign w15055 = b[17] & w9165;
assign w15056 = b[18] & w9160;
assign w15057 = ~w1108 & w9158;
assign w15058 = ~w15055 & ~w15056;
assign w15059 = ~w15054 & w15058;
assign w15060 = ~w15057 & w15059;
assign w15061 = a[56] & ~w15060;
assign w15062 = ~a[56] & w15060;
assign w15063 = ~w15061 & ~w15062;
assign w15064 = w15053 & w15063;
assign w15065 = ~w15053 & ~w15063;
assign w15066 = ~w15064 & ~w15065;
assign w15067 = ~w14689 & ~w14701;
assign w15068 = ~w15066 & w15067;
assign w15069 = w15066 & ~w15067;
assign w15070 = ~w15068 & ~w15069;
assign w15071 = b[19] & w8515;
assign w15072 = b[21] & w8202;
assign w15073 = b[20] & w8200;
assign w15074 = w1467 & w8195;
assign w15075 = ~w15072 & ~w15073;
assign w15076 = ~w15071 & w15075;
assign w15077 = ~w15074 & w15076;
assign w15078 = a[53] & ~w15077;
assign w15079 = ~a[53] & w15077;
assign w15080 = ~w15078 & ~w15079;
assign w15081 = w15070 & w15080;
assign w15082 = ~w15070 & ~w15080;
assign w15083 = ~w15081 & ~w15082;
assign w15084 = ~w14705 & ~w14709;
assign w15085 = w15083 & ~w15084;
assign w15086 = ~w15083 & w15084;
assign w15087 = ~w15085 & ~w15086;
assign w15088 = ~w15010 & ~w15087;
assign w15089 = w15010 & w15087;
assign w15090 = ~w15088 & ~w15089;
assign w15091 = ~w15000 & w15090;
assign w15092 = w15000 & ~w15090;
assign w15093 = ~w15091 & ~w15092;
assign w15094 = w14999 & w15093;
assign w15095 = ~w14999 & ~w15093;
assign w15096 = ~w15094 & ~w15095;
assign w15097 = w14989 & ~w15096;
assign w15098 = ~w14989 & w15096;
assign w15099 = ~w15097 & ~w15098;
assign w15100 = b[28] & w5939;
assign w15101 = b[29] & w5670;
assign w15102 = b[30] & w5665;
assign w15103 = ~w2908 & w5663;
assign w15104 = ~w15101 & ~w15102;
assign w15105 = ~w15100 & w15104;
assign w15106 = ~w15103 & w15105;
assign w15107 = a[44] & ~w15106;
assign w15108 = ~a[44] & w15106;
assign w15109 = ~w15107 & ~w15108;
assign w15110 = ~w15099 & ~w15109;
assign w15111 = w15099 & w15109;
assign w15112 = ~w15110 & ~w15111;
assign w15113 = w14988 & w15112;
assign w15114 = ~w14988 & ~w15112;
assign w15115 = ~w15113 & ~w15114;
assign w15116 = w14987 & ~w15115;
assign w15117 = ~w14987 & w15115;
assign w15118 = ~w15116 & ~w15117;
assign w15119 = ~w14977 & w15118;
assign w15120 = w14977 & ~w15118;
assign w15121 = ~w15119 & ~w15120;
assign w15122 = w14976 & w15121;
assign w15123 = ~w14976 & ~w15121;
assign w15124 = ~w15122 & ~w15123;
assign w15125 = w14966 & ~w15124;
assign w15126 = ~w14966 & w15124;
assign w15127 = ~w15125 & ~w15126;
assign w15128 = b[37] & w3785;
assign w15129 = b[38] & w3578;
assign w15130 = b[39] & w3580;
assign w15131 = w3573 & ~w4812;
assign w15132 = ~w15129 & ~w15130;
assign w15133 = ~w15128 & w15132;
assign w15134 = ~w15131 & w15133;
assign w15135 = a[35] & ~w15134;
assign w15136 = ~a[35] & w15134;
assign w15137 = ~w15135 & ~w15136;
assign w15138 = w15127 & w15137;
assign w15139 = ~w15127 & ~w15137;
assign w15140 = ~w15138 & ~w15139;
assign w15141 = ~w14775 & ~w14778;
assign w15142 = w15140 & ~w15141;
assign w15143 = ~w15140 & w15141;
assign w15144 = ~w15142 & ~w15143;
assign w15145 = w14965 & w15144;
assign w15146 = ~w14965 & ~w15144;
assign w15147 = ~w15145 & ~w15146;
assign w15148 = w14951 & w15147;
assign w15149 = ~w14951 & ~w15147;
assign w15150 = ~w15148 & ~w15149;
assign w15151 = w14937 & w15150;
assign w15152 = ~w14937 & ~w15150;
assign w15153 = ~w15151 & ~w15152;
assign w15154 = b[49] & ~w1676;
assign w15155 = b[50] & w1517;
assign w15156 = b[51] & w1519;
assign w15157 = w1513 & ~w8058;
assign w15158 = ~w15154 & ~w15155;
assign w15159 = ~w15156 & w15158;
assign w15160 = ~w15157 & w15159;
assign w15161 = a[23] & ~w15160;
assign w15162 = ~a[23] & w15160;
assign w15163 = ~w15161 & ~w15162;
assign w15164 = ~w14592 & ~w14819;
assign w15165 = w15163 & ~w15164;
assign w15166 = ~w15163 & w15164;
assign w15167 = ~w15165 & ~w15166;
assign w15168 = ~w15153 & ~w15167;
assign w15169 = w15153 & w15167;
assign w15170 = ~w15168 & ~w15169;
assign w15171 = ~w14832 & ~w14835;
assign w15172 = b[54] & w1156;
assign w15173 = b[52] & ~w1272;
assign w15174 = b[53] & w1154;
assign w15175 = w1150 & ~w8998;
assign w15176 = ~w15172 & ~w15173;
assign w15177 = ~w15174 & w15176;
assign w15178 = ~w15175 & w15177;
assign w15179 = a[20] & ~w15178;
assign w15180 = ~a[20] & w15178;
assign w15181 = ~w15179 & ~w15180;
assign w15182 = ~w15171 & w15181;
assign w15183 = w15171 & ~w15181;
assign w15184 = ~w15182 & ~w15183;
assign w15185 = w15170 & w15184;
assign w15186 = ~w15170 & ~w15184;
assign w15187 = ~w15185 & ~w15186;
assign w15188 = w14923 & w15187;
assign w15189 = ~w14923 & ~w15187;
assign w15190 = ~w15188 & ~w15189;
assign w15191 = ~w14866 & ~w14869;
assign w15192 = b[58] & ~w649;
assign w15193 = b[60] & w575;
assign w15194 = b[59] & w573;
assign w15195 = w569 & w11035;
assign w15196 = ~w15192 & ~w15193;
assign w15197 = ~w15194 & w15196;
assign w15198 = ~w15195 & w15197;
assign w15199 = a[14] & ~w15198;
assign w15200 = ~a[14] & w15198;
assign w15201 = ~w15199 & ~w15200;
assign w15202 = ~w15191 & w15201;
assign w15203 = w15191 & ~w15201;
assign w15204 = ~w15202 & ~w15203;
assign w15205 = ~w15190 & ~w15204;
assign w15206 = w15190 & w15204;
assign w15207 = ~w15205 & ~w15206;
assign w15208 = ~w14883 & ~w14886;
assign w15209 = b[62] & w358;
assign w15210 = b[63] & w360;
assign w15211 = b[61] & ~w419;
assign w15212 = w354 & w12132;
assign w15213 = ~w15209 & ~w15210;
assign w15214 = ~w15211 & w15213;
assign w15215 = ~w15212 & w15214;
assign w15216 = a[11] & ~w15215;
assign w15217 = ~a[11] & w15215;
assign w15218 = ~w15216 & ~w15217;
assign w15219 = ~w15208 & w15218;
assign w15220 = w15208 & ~w15218;
assign w15221 = ~w15219 & ~w15220;
assign w15222 = w15207 & w15221;
assign w15223 = ~w15207 & ~w15221;
assign w15224 = ~w15222 & ~w15223;
assign w15225 = ~w14909 & w15224;
assign w15226 = w14909 & ~w15224;
assign w15227 = ~w15225 & ~w15226;
assign w15228 = w15227 & w25729;
assign w15229 = ~w25729 & ~w15227;
assign w15230 = ~w15228 & ~w15229;
assign w15231 = ~w15219 & ~w15222;
assign w15232 = b[60] & w573;
assign w15233 = b[59] & ~w649;
assign w15234 = b[61] & w575;
assign w15235 = w569 & w11400;
assign w15236 = ~w15232 & ~w15233;
assign w15237 = ~w15234 & w15236;
assign w15238 = ~w15235 & w15237;
assign w15239 = a[14] & ~w15238;
assign w15240 = ~a[14] & w15238;
assign w15241 = ~w15239 & ~w15240;
assign w15242 = ~w14921 & ~w15188;
assign w15243 = w15241 & ~w15242;
assign w15244 = ~w15241 & w15242;
assign w15245 = ~w15243 & ~w15244;
assign w15246 = b[51] & w1517;
assign w15247 = b[52] & w1519;
assign w15248 = b[50] & ~w1676;
assign w15249 = w1513 & ~w8371;
assign w15250 = ~w15246 & ~w15247;
assign w15251 = ~w15248 & w15250;
assign w15252 = ~w15249 & w15251;
assign w15253 = a[23] & ~w15252;
assign w15254 = ~a[23] & w15252;
assign w15255 = ~w15253 & ~w15254;
assign w15256 = ~w14935 & ~w15151;
assign w15257 = w15255 & ~w15256;
assign w15258 = ~w15255 & w15256;
assign w15259 = ~w15257 & ~w15258;
assign w15260 = b[49] & w1957;
assign w15261 = b[48] & w1955;
assign w15262 = b[47] & ~w2114;
assign w15263 = w1951 & ~w7468;
assign w15264 = ~w15260 & ~w15261;
assign w15265 = ~w15262 & w15264;
assign w15266 = ~w15263 & w15265;
assign w15267 = a[26] & ~w15266;
assign w15268 = ~a[26] & w15266;
assign w15269 = ~w15267 & ~w15268;
assign w15270 = ~w14949 & ~w15148;
assign w15271 = w15269 & ~w15270;
assign w15272 = ~w15269 & w15270;
assign w15273 = ~w15271 & ~w15272;
assign w15274 = b[41] & w3177;
assign w15275 = b[43] & w2978;
assign w15276 = b[42] & w2973;
assign w15277 = w2980 & w5811;
assign w15278 = ~w15275 & ~w15276;
assign w15279 = ~w15274 & w15278;
assign w15280 = ~w15277 & w15279;
assign w15281 = a[32] & ~w15280;
assign w15282 = ~a[32] & w15280;
assign w15283 = ~w15281 & ~w15282;
assign w15284 = ~w15138 & ~w15142;
assign w15285 = w15283 & ~w15284;
assign w15286 = ~w15283 & w15284;
assign w15287 = ~w15285 & ~w15286;
assign w15288 = b[38] & w3785;
assign w15289 = b[40] & w3580;
assign w15290 = b[39] & w3578;
assign w15291 = w3573 & ~w5058;
assign w15292 = ~w15289 & ~w15290;
assign w15293 = ~w15288 & w15292;
assign w15294 = ~w15291 & w15293;
assign w15295 = a[35] & ~w15294;
assign w15296 = ~a[35] & w15294;
assign w15297 = ~w15295 & ~w15296;
assign w15298 = ~w15122 & ~w15126;
assign w15299 = b[35] & w4453;
assign w15300 = b[36] & w4241;
assign w15301 = b[37] & w4243;
assign w15302 = w4236 & ~w4357;
assign w15303 = ~w15300 & ~w15301;
assign w15304 = ~w15299 & w15303;
assign w15305 = ~w15302 & w15304;
assign w15306 = a[38] & ~w15305;
assign w15307 = ~a[38] & w15305;
assign w15308 = ~w15306 & ~w15307;
assign w15309 = ~w15116 & ~w15119;
assign w15310 = b[32] & w5167;
assign w15311 = b[33] & w4918;
assign w15312 = b[34] & w4925;
assign w15313 = ~w3710 & w4923;
assign w15314 = ~w15311 & ~w15312;
assign w15315 = ~w15310 & w15314;
assign w15316 = ~w15313 & w15315;
assign w15317 = a[41] & ~w15316;
assign w15318 = ~a[41] & w15316;
assign w15319 = ~w15317 & ~w15318;
assign w15320 = b[29] & w5939;
assign w15321 = b[30] & w5670;
assign w15322 = b[31] & w5665;
assign w15323 = ~w3112 & w5663;
assign w15324 = ~w15321 & ~w15322;
assign w15325 = ~w15320 & w15324;
assign w15326 = ~w15323 & w15325;
assign w15327 = a[44] & ~w15326;
assign w15328 = ~a[44] & w15326;
assign w15329 = ~w15327 & ~w15328;
assign w15330 = b[26] & w6732;
assign w15331 = b[27] & w6474;
assign w15332 = b[28] & w6476;
assign w15333 = w2559 & w6469;
assign w15334 = ~w15331 & ~w15332;
assign w15335 = ~w15330 & w15334;
assign w15336 = ~w15333 & w15335;
assign w15337 = a[47] & ~w15336;
assign w15338 = ~a[47] & w15336;
assign w15339 = ~w15337 & ~w15338;
assign w15340 = b[23] & w7586;
assign w15341 = b[24] & w7307;
assign w15342 = b[25] & w7314;
assign w15343 = w2061 & w7312;
assign w15344 = ~w15341 & ~w15342;
assign w15345 = ~w15340 & w15344;
assign w15346 = ~w15343 & w15345;
assign w15347 = a[50] & ~w15346;
assign w15348 = ~a[50] & w15346;
assign w15349 = ~w15347 & ~w15348;
assign w15350 = b[20] & w8515;
assign w15351 = b[21] & w8200;
assign w15352 = b[22] & w8202;
assign w15353 = w1615 & w8195;
assign w15354 = ~w15351 & ~w15352;
assign w15355 = ~w15350 & w15354;
assign w15356 = ~w15353 & w15355;
assign w15357 = a[53] & ~w15356;
assign w15358 = ~a[53] & w15356;
assign w15359 = ~w15357 & ~w15358;
assign w15360 = b[17] & w9482;
assign w15361 = b[18] & w9165;
assign w15362 = b[19] & w9160;
assign w15363 = ~w1231 & w9158;
assign w15364 = ~w15361 & ~w15362;
assign w15365 = ~w15360 & w15364;
assign w15366 = ~w15363 & w15365;
assign w15367 = a[56] & ~w15366;
assign w15368 = ~a[56] & w15366;
assign w15369 = ~w15367 & ~w15368;
assign w15370 = ~w15048 & ~w15051;
assign w15371 = b[14] & w10496;
assign w15372 = b[16] & w10148;
assign w15373 = b[15] & w10146;
assign w15374 = w905 & w10141;
assign w15375 = ~w15372 & ~w15373;
assign w15376 = ~w15371 & w15375;
assign w15377 = ~w15374 & w15376;
assign w15378 = a[59] & ~w15377;
assign w15379 = ~a[59] & w15377;
assign w15380 = ~w15378 & ~w15379;
assign w15381 = ~w15023 & ~w15036;
assign w15382 = b[11] & w11561;
assign w15383 = b[13] & w11196;
assign w15384 = b[12] & w11194;
assign w15385 = w628 & w11189;
assign w15386 = ~w15383 & ~w15384;
assign w15387 = ~w15382 & w15386;
assign w15388 = ~w15385 & w15387;
assign w15389 = a[62] & ~w15388;
assign w15390 = ~a[62] & w15388;
assign w15391 = ~w15389 & ~w15390;
assign w15392 = b[9] & w11921;
assign w15393 = b[10] & w11923;
assign w15394 = ~w15392 & ~w15393;
assign w15395 = ~w15015 & ~w15018;
assign w15396 = w15394 & ~w15395;
assign w15397 = ~w15394 & w15395;
assign w15398 = ~w15396 & ~w15397;
assign w15399 = w15391 & w15398;
assign w15400 = ~w15391 & ~w15398;
assign w15401 = ~w15399 & ~w15400;
assign w15402 = ~w15381 & w15401;
assign w15403 = w15381 & ~w15401;
assign w15404 = ~w15402 & ~w15403;
assign w15405 = w15380 & w15404;
assign w15406 = ~w15380 & ~w15404;
assign w15407 = ~w15405 & ~w15406;
assign w15408 = ~w15370 & w15407;
assign w15409 = w15370 & ~w15407;
assign w15410 = ~w15408 & ~w15409;
assign w15411 = w15369 & w15410;
assign w15412 = ~w15369 & ~w15410;
assign w15413 = ~w15411 & ~w15412;
assign w15414 = ~w15064 & ~w15069;
assign w15415 = w15413 & ~w15414;
assign w15416 = ~w15413 & w15414;
assign w15417 = ~w15415 & ~w15416;
assign w15418 = w15359 & w15417;
assign w15419 = ~w15359 & ~w15417;
assign w15420 = ~w15418 & ~w15419;
assign w15421 = ~w15081 & ~w15085;
assign w15422 = w15420 & ~w15421;
assign w15423 = ~w15420 & w15421;
assign w15424 = ~w15422 & ~w15423;
assign w15425 = w15349 & w15424;
assign w15426 = ~w15349 & ~w15424;
assign w15427 = ~w15425 & ~w15426;
assign w15428 = ~w15089 & ~w15091;
assign w15429 = w15427 & ~w15428;
assign w15430 = ~w15427 & w15428;
assign w15431 = ~w15429 & ~w15430;
assign w15432 = w15339 & w15431;
assign w15433 = ~w15339 & ~w15431;
assign w15434 = ~w15432 & ~w15433;
assign w15435 = ~w15094 & ~w15098;
assign w15436 = w15434 & ~w15435;
assign w15437 = ~w15434 & w15435;
assign w15438 = ~w15436 & ~w15437;
assign w15439 = ~w15329 & ~w15438;
assign w15440 = w15329 & w15438;
assign w15441 = ~w15439 & ~w15440;
assign w15442 = ~w15110 & ~w15113;
assign w15443 = ~w15441 & ~w15442;
assign w15444 = w15441 & w15442;
assign w15445 = ~w15443 & ~w15444;
assign w15446 = w15319 & w15445;
assign w15447 = ~w15319 & ~w15445;
assign w15448 = ~w15446 & ~w15447;
assign w15449 = w15309 & ~w15448;
assign w15450 = ~w15309 & w15448;
assign w15451 = ~w15449 & ~w15450;
assign w15452 = w15308 & w15451;
assign w15453 = ~w15308 & ~w15451;
assign w15454 = ~w15452 & ~w15453;
assign w15455 = w15298 & ~w15454;
assign w15456 = ~w15298 & w15454;
assign w15457 = ~w15455 & ~w15456;
assign w15458 = w15297 & w15457;
assign w15459 = ~w15297 & ~w15457;
assign w15460 = ~w15458 & ~w15459;
assign w15461 = w15287 & w15460;
assign w15462 = ~w15287 & ~w15460;
assign w15463 = ~w15461 & ~w15462;
assign w15464 = ~w14963 & ~w15145;
assign w15465 = b[44] & ~w2622;
assign w15466 = b[45] & w2436;
assign w15467 = b[46] & w2438;
assign w15468 = w2432 & ~w6613;
assign w15469 = ~w15465 & ~w15466;
assign w15470 = ~w15467 & w15469;
assign w15471 = ~w15468 & w15470;
assign w15472 = a[29] & ~w15471;
assign w15473 = ~a[29] & w15471;
assign w15474 = ~w15472 & ~w15473;
assign w15475 = ~w15464 & w15474;
assign w15476 = w15464 & ~w15474;
assign w15477 = ~w15475 & ~w15476;
assign w15478 = w15463 & w15477;
assign w15479 = ~w15463 & ~w15477;
assign w15480 = ~w15478 & ~w15479;
assign w15481 = w15273 & w15480;
assign w15482 = ~w15273 & ~w15480;
assign w15483 = ~w15481 & ~w15482;
assign w15484 = w15259 & w15483;
assign w15485 = ~w15259 & ~w15483;
assign w15486 = ~w15484 & ~w15485;
assign w15487 = b[55] & w1156;
assign w15488 = b[53] & ~w1272;
assign w15489 = b[54] & w1154;
assign w15490 = w1150 & ~w9330;
assign w15491 = ~w15487 & ~w15488;
assign w15492 = ~w15489 & w15491;
assign w15493 = ~w15490 & w15492;
assign w15494 = a[20] & ~w15493;
assign w15495 = ~a[20] & w15493;
assign w15496 = ~w15494 & ~w15495;
assign w15497 = ~w15165 & ~w15169;
assign w15498 = w15496 & ~w15497;
assign w15499 = ~w15496 & w15497;
assign w15500 = ~w15498 & ~w15499;
assign w15501 = w15486 & w15500;
assign w15502 = ~w15486 & ~w15500;
assign w15503 = ~w15501 & ~w15502;
assign w15504 = ~w15182 & ~w15185;
assign w15505 = b[56] & ~w934;
assign w15506 = b[57] & w838;
assign w15507 = b[58] & w834;
assign w15508 = w832 & ~w10339;
assign w15509 = ~w15505 & ~w15506;
assign w15510 = ~w15507 & w15509;
assign w15511 = ~w15508 & w15510;
assign w15512 = a[17] & ~w15511;
assign w15513 = ~a[17] & w15511;
assign w15514 = ~w15512 & ~w15513;
assign w15515 = ~w15504 & w15514;
assign w15516 = w15504 & ~w15514;
assign w15517 = ~w15515 & ~w15516;
assign w15518 = w15503 & w15517;
assign w15519 = ~w15503 & ~w15517;
assign w15520 = ~w15518 & ~w15519;
assign w15521 = w15245 & w15520;
assign w15522 = ~w15245 & ~w15520;
assign w15523 = ~w15521 & ~w15522;
assign w15524 = ~w15202 & ~w15206;
assign w15525 = b[62] & ~w419;
assign w15526 = b[63] & w358;
assign w15527 = w354 & w12156;
assign w15528 = ~w15525 & ~w15526;
assign w15529 = ~w15527 & w15528;
assign w15530 = a[11] & ~w15529;
assign w15531 = ~a[11] & w15529;
assign w15532 = ~w15530 & ~w15531;
assign w15533 = ~w15524 & w15532;
assign w15534 = w15524 & ~w15532;
assign w15535 = ~w15533 & ~w15534;
assign w15536 = w15523 & w15535;
assign w15537 = ~w15523 & ~w15535;
assign w15538 = ~w15536 & ~w15537;
assign w15539 = w15231 & ~w15538;
assign w15540 = ~w15231 & w15538;
assign w15541 = ~w15539 & ~w15540;
assign w15542 = (~w13908 & w25560) | (~w13908 & w25561) | (w25560 & w25561);
assign w15543 = w15541 & w15542;
assign w15544 = ~w15541 & ~w15542;
assign w15545 = ~w15543 & ~w15544;
assign w15546 = (~w15533 & ~w15535) | (~w15533 & w25562) | (~w15535 & w25562);
assign w15547 = (~w15243 & ~w15245) | (~w15243 & w25563) | (~w15245 & w25563);
assign w15548 = w354 & ~w12154;
assign w15549 = w419 & ~w15548;
assign w15550 = b[63] & ~w15549;
assign w15551 = ~a[11] & ~w15550;
assign w15552 = a[11] & w15550;
assign w15553 = ~w15551 & ~w15552;
assign w15554 = ~w15547 & w15553;
assign w15555 = w15547 & ~w15553;
assign w15556 = ~w15554 & ~w15555;
assign w15557 = b[57] & ~w934;
assign w15558 = b[58] & w838;
assign w15559 = b[59] & w834;
assign w15560 = ~w15557 & ~w15558;
assign w15561 = ~w15559 & w15560;
assign w15562 = (w10371 & w25313) | (w10371 & w25314) | (w25313 & w25314);
assign w15563 = (~w10371 & w25315) | (~w10371 & w25316) | (w25315 & w25316);
assign w15564 = ~w15562 & ~w15563;
assign w15565 = ~w15498 & ~w15501;
assign w15566 = w15564 & ~w15565;
assign w15567 = ~w15564 & w15565;
assign w15568 = ~w15566 & ~w15567;
assign w15569 = b[56] & w1156;
assign w15570 = b[54] & ~w1272;
assign w15571 = b[55] & w1154;
assign w15572 = ~w15569 & ~w15570;
assign w15573 = ~w15571 & w15572;
assign w15574 = (w9657 & w25564) | (w9657 & w25565) | (w25564 & w25565);
assign w15575 = ~a[20] & w25730;
assign w15576 = ~w15574 & ~w15575;
assign w15577 = (~w15257 & ~w15259) | (~w15257 & w25566) | (~w15259 & w25566);
assign w15578 = w15576 & ~w15577;
assign w15579 = ~w15576 & w15577;
assign w15580 = ~w15578 & ~w15579;
assign w15581 = b[39] & w3785;
assign w15582 = b[40] & w3578;
assign w15583 = b[41] & w3580;
assign w15584 = w3573 & w5302;
assign w15585 = ~w15582 & ~w15583;
assign w15586 = ~w15581 & w15585;
assign w15587 = ~w15584 & w15586;
assign w15588 = a[35] & ~w15587;
assign w15589 = ~a[35] & w15587;
assign w15590 = ~w15588 & ~w15589;
assign w15591 = ~w15450 & ~w15452;
assign w15592 = b[36] & w4453;
assign w15593 = b[37] & w4241;
assign w15594 = b[38] & w4243;
assign w15595 = w4236 & w4582;
assign w15596 = ~w15593 & ~w15594;
assign w15597 = ~w15592 & w15596;
assign w15598 = ~w15595 & w15597;
assign w15599 = a[38] & ~w15598;
assign w15600 = ~a[38] & w15598;
assign w15601 = ~w15599 & ~w15600;
assign w15602 = b[30] & w5939;
assign w15603 = b[31] & w5670;
assign w15604 = b[32] & w5665;
assign w15605 = w3304 & w5663;
assign w15606 = ~w15603 & ~w15604;
assign w15607 = ~w15602 & w15606;
assign w15608 = ~w15605 & w15607;
assign w15609 = a[44] & ~w15608;
assign w15610 = ~a[44] & w15608;
assign w15611 = ~w15609 & ~w15610;
assign w15612 = ~w15422 & ~w15425;
assign w15613 = ~w15415 & ~w15418;
assign w15614 = b[21] & w8515;
assign w15615 = b[23] & w8202;
assign w15616 = b[22] & w8200;
assign w15617 = w1755 & w8195;
assign w15618 = ~w15615 & ~w15616;
assign w15619 = ~w15614 & w15618;
assign w15620 = ~w15617 & w15619;
assign w15621 = a[53] & ~w15620;
assign w15622 = ~a[53] & w15620;
assign w15623 = ~w15621 & ~w15622;
assign w15624 = ~w15408 & ~w15411;
assign w15625 = ~w15402 & ~w15405;
assign w15626 = b[15] & w10496;
assign w15627 = b[16] & w10146;
assign w15628 = b[17] & w10148;
assign w15629 = w1008 & w10141;
assign w15630 = ~w15627 & ~w15628;
assign w15631 = ~w15626 & w15630;
assign w15632 = ~w15629 & w15631;
assign w15633 = a[59] & ~w15632;
assign w15634 = ~a[59] & w15632;
assign w15635 = ~w15633 & ~w15634;
assign w15636 = b[12] & w11561;
assign w15637 = b[13] & w11194;
assign w15638 = b[14] & w11196;
assign w15639 = w714 & w11189;
assign w15640 = ~w15637 & ~w15638;
assign w15641 = ~w15636 & w15640;
assign w15642 = ~w15639 & w15641;
assign w15643 = a[62] & ~w15642;
assign w15644 = ~a[62] & w15642;
assign w15645 = ~w15643 & ~w15644;
assign w15646 = ~w15396 & ~w15399;
assign w15647 = b[10] & w11921;
assign w15648 = b[11] & w11923;
assign w15649 = ~w15647 & ~w15648;
assign w15650 = w15394 & ~w15649;
assign w15651 = ~w15394 & w15649;
assign w15652 = ~w15650 & ~w15651;
assign w15653 = ~w15646 & w15652;
assign w15654 = w15646 & ~w15652;
assign w15655 = ~w15653 & ~w15654;
assign w15656 = w15645 & w15655;
assign w15657 = ~w15645 & ~w15655;
assign w15658 = ~w15656 & ~w15657;
assign w15659 = w15635 & w15658;
assign w15660 = ~w15635 & ~w15658;
assign w15661 = ~w15659 & ~w15660;
assign w15662 = ~w15625 & w15661;
assign w15663 = w15625 & ~w15661;
assign w15664 = ~w15662 & ~w15663;
assign w15665 = b[18] & w9482;
assign w15666 = b[20] & w9160;
assign w15667 = b[19] & w9165;
assign w15668 = w1347 & w9158;
assign w15669 = ~w15666 & ~w15667;
assign w15670 = ~w15665 & w15669;
assign w15671 = ~w15668 & w15670;
assign w15672 = a[56] & ~w15671;
assign w15673 = ~a[56] & w15671;
assign w15674 = ~w15672 & ~w15673;
assign w15675 = ~w15664 & ~w15674;
assign w15676 = w15664 & w15674;
assign w15677 = ~w15675 & ~w15676;
assign w15678 = w15624 & ~w15677;
assign w15679 = ~w15624 & w15677;
assign w15680 = ~w15678 & ~w15679;
assign w15681 = w15623 & w15680;
assign w15682 = ~w15623 & ~w15680;
assign w15683 = ~w15681 & ~w15682;
assign w15684 = w15613 & ~w15683;
assign w15685 = ~w15613 & w15683;
assign w15686 = ~w15684 & ~w15685;
assign w15687 = b[24] & w7586;
assign w15688 = b[25] & w7307;
assign w15689 = b[26] & w7314;
assign w15690 = w2219 & w7312;
assign w15691 = ~w15688 & ~w15689;
assign w15692 = ~w15687 & w15691;
assign w15693 = ~w15690 & w15692;
assign w15694 = a[50] & ~w15693;
assign w15695 = ~a[50] & w15693;
assign w15696 = ~w15694 & ~w15695;
assign w15697 = w15686 & w15696;
assign w15698 = ~w15686 & ~w15696;
assign w15699 = ~w15697 & ~w15698;
assign w15700 = w15612 & ~w15699;
assign w15701 = ~w15612 & w15699;
assign w15702 = ~w15700 & ~w15701;
assign w15703 = b[27] & w6732;
assign w15704 = b[29] & w6476;
assign w15705 = b[28] & w6474;
assign w15706 = w2734 & w6469;
assign w15707 = ~w15704 & ~w15705;
assign w15708 = ~w15703 & w15707;
assign w15709 = ~w15706 & w15708;
assign w15710 = a[47] & ~w15709;
assign w15711 = ~a[47] & w15709;
assign w15712 = ~w15710 & ~w15711;
assign w15713 = w15702 & w15712;
assign w15714 = ~w15702 & ~w15712;
assign w15715 = ~w15713 & ~w15714;
assign w15716 = ~w15429 & ~w15432;
assign w15717 = w15715 & ~w15716;
assign w15718 = ~w15715 & w15716;
assign w15719 = ~w15717 & ~w15718;
assign w15720 = ~w15611 & ~w15719;
assign w15721 = w15611 & w15719;
assign w15722 = ~w15720 & ~w15721;
assign w15723 = ~w15436 & ~w15440;
assign w15724 = w15722 & ~w15723;
assign w15725 = ~w15722 & w15723;
assign w15726 = ~w15724 & ~w15725;
assign w15727 = b[33] & w5167;
assign w15728 = b[35] & w4925;
assign w15729 = b[34] & w4918;
assign w15730 = w3918 & w4923;
assign w15731 = ~w15728 & ~w15729;
assign w15732 = ~w15727 & w15731;
assign w15733 = ~w15730 & w15732;
assign w15734 = a[41] & ~w15733;
assign w15735 = ~a[41] & w15733;
assign w15736 = ~w15734 & ~w15735;
assign w15737 = w15726 & w15736;
assign w15738 = ~w15726 & ~w15736;
assign w15739 = ~w15737 & ~w15738;
assign w15740 = ~w15444 & ~w15446;
assign w15741 = w15739 & ~w15740;
assign w15742 = ~w15739 & w15740;
assign w15743 = ~w15741 & ~w15742;
assign w15744 = ~w15601 & ~w15743;
assign w15745 = w15601 & w15743;
assign w15746 = ~w15744 & ~w15745;
assign w15747 = w15591 & ~w15746;
assign w15748 = ~w15591 & w15746;
assign w15749 = ~w15747 & ~w15748;
assign w15750 = ~w15590 & ~w15749;
assign w15751 = w15590 & w15749;
assign w15752 = ~w15750 & ~w15751;
assign w15753 = ~w15456 & ~w15458;
assign w15754 = b[42] & w3177;
assign w15755 = b[44] & w2978;
assign w15756 = b[43] & w2973;
assign w15757 = w2980 & w6069;
assign w15758 = ~w15755 & ~w15756;
assign w15759 = ~w15754 & w15758;
assign w15760 = ~w15757 & w15759;
assign w15761 = a[32] & ~w15760;
assign w15762 = ~a[32] & w15760;
assign w15763 = ~w15761 & ~w15762;
assign w15764 = ~w15753 & w15763;
assign w15765 = w15753 & ~w15763;
assign w15766 = ~w15764 & ~w15765;
assign w15767 = w15752 & w15766;
assign w15768 = ~w15752 & ~w15766;
assign w15769 = ~w15767 & ~w15768;
assign w15770 = b[47] & w2438;
assign w15771 = b[45] & ~w2622;
assign w15772 = b[46] & w2436;
assign w15773 = w2432 & w6889;
assign w15774 = ~w15770 & ~w15771;
assign w15775 = ~w15772 & w15774;
assign w15776 = ~w15773 & w15775;
assign w15777 = a[29] & ~w15776;
assign w15778 = ~a[29] & w15776;
assign w15779 = ~w15777 & ~w15778;
assign w15780 = ~w15285 & ~w15461;
assign w15781 = w15779 & ~w15780;
assign w15782 = ~w15779 & w15780;
assign w15783 = ~w15781 & ~w15782;
assign w15784 = w15769 & w15783;
assign w15785 = ~w15769 & ~w15783;
assign w15786 = ~w15784 & ~w15785;
assign w15787 = ~w15475 & ~w15478;
assign w15788 = b[48] & ~w2114;
assign w15789 = b[50] & w1957;
assign w15790 = b[49] & w1955;
assign w15791 = w1951 & w7759;
assign w15792 = ~w15788 & ~w15789;
assign w15793 = ~w15790 & w15792;
assign w15794 = ~w15791 & w15793;
assign w15795 = a[26] & ~w15794;
assign w15796 = ~a[26] & w15794;
assign w15797 = ~w15795 & ~w15796;
assign w15798 = ~w15787 & w15797;
assign w15799 = w15787 & ~w15797;
assign w15800 = ~w15798 & ~w15799;
assign w15801 = w15786 & w15800;
assign w15802 = ~w15786 & ~w15800;
assign w15803 = ~w15801 & ~w15802;
assign w15804 = (~w15271 & ~w15273) | (~w15271 & w25567) | (~w15273 & w25567);
assign w15805 = b[51] & ~w1676;
assign w15806 = b[53] & w1519;
assign w15807 = b[52] & w1517;
assign w15808 = ~w15805 & ~w15806;
assign w15809 = ~w15807 & w15808;
assign w15810 = (w15809 & ~w8683) | (w15809 & w25568) | (~w8683 & w25568);
assign w15811 = a[23] & ~w15810;
assign w15812 = ~a[23] & w15810;
assign w15813 = ~w15811 & ~w15812;
assign w15814 = ~w15804 & w15813;
assign w15815 = w15804 & ~w15813;
assign w15816 = ~w15814 & ~w15815;
assign w15817 = w15803 & w15816;
assign w15818 = ~w15803 & ~w15816;
assign w15819 = ~w15817 & ~w15818;
assign w15820 = w15580 & w15819;
assign w15821 = ~w15580 & ~w15819;
assign w15822 = ~w15820 & ~w15821;
assign w15823 = w15568 & w15822;
assign w15824 = ~w15568 & ~w15822;
assign w15825 = ~w15823 & ~w15824;
assign w15826 = (~w15515 & ~w15517) | (~w15515 & w25569) | (~w15517 & w25569);
assign w15827 = b[60] & ~w649;
assign w15828 = b[62] & w575;
assign w15829 = b[61] & w573;
assign w15830 = ~w15827 & ~w15828;
assign w15831 = ~w15829 & w15830;
assign w15832 = (w11763 & w25570) | (w11763 & w25571) | (w25570 & w25571);
assign w15833 = (~w11763 & w25572) | (~w11763 & w25573) | (w25572 & w25573);
assign w15834 = ~w15832 & ~w15833;
assign w15835 = ~w15826 & w15834;
assign w15836 = w15826 & ~w15834;
assign w15837 = ~w15835 & ~w15836;
assign w15838 = w15825 & w15837;
assign w15839 = ~w15825 & ~w15837;
assign w15840 = ~w15838 & ~w15839;
assign w15841 = w15556 & w15840;
assign w15842 = ~w15556 & ~w15840;
assign w15843 = ~w15841 & ~w15842;
assign w15844 = ~w15546 & w15843;
assign w15845 = w15546 & ~w15843;
assign w15846 = ~w15844 & ~w15845;
assign w15847 = ~w15539 & w15846;
assign w15848 = (w15847 & w15542) | (w15847 & w24414) | (w15542 & w24414);
assign w15849 = ~w15540 & ~w15846;
assign w15850 = ~w15543 & w15849;
assign w15851 = ~w15848 & ~w15850;
assign w15852 = (~w15844 & ~w15847) | (~w15844 & w25731) | (~w15847 & w25731);
assign w15853 = ~w15554 & ~w15841;
assign w15854 = ~w15748 & ~w15751;
assign w15855 = b[40] & w3785;
assign w15856 = b[42] & w3580;
assign w15857 = b[41] & w3578;
assign w15858 = w3573 & w5548;
assign w15859 = ~w15856 & ~w15857;
assign w15860 = ~w15855 & w15859;
assign w15861 = ~w15858 & w15860;
assign w15862 = a[35] & ~w15861;
assign w15863 = ~a[35] & w15861;
assign w15864 = ~w15862 & ~w15863;
assign w15865 = ~w15741 & ~w15745;
assign w15866 = ~w15724 & ~w15737;
assign w15867 = b[34] & w5167;
assign w15868 = b[35] & w4918;
assign w15869 = b[36] & w4925;
assign w15870 = w4129 & w4923;
assign w15871 = ~w15868 & ~w15869;
assign w15872 = ~w15867 & w15871;
assign w15873 = ~w15870 & w15872;
assign w15874 = a[41] & ~w15873;
assign w15875 = ~a[41] & w15873;
assign w15876 = ~w15874 & ~w15875;
assign w15877 = ~w15717 & ~w15721;
assign w15878 = b[31] & w5939;
assign w15879 = b[33] & w5665;
assign w15880 = b[32] & w5670;
assign w15881 = w3499 & w5663;
assign w15882 = ~w15879 & ~w15880;
assign w15883 = ~w15878 & w15882;
assign w15884 = ~w15881 & w15883;
assign w15885 = a[44] & ~w15884;
assign w15886 = ~a[44] & w15884;
assign w15887 = ~w15885 & ~w15886;
assign w15888 = ~w15701 & ~w15713;
assign w15889 = ~w15685 & ~w15697;
assign w15890 = b[25] & w7586;
assign w15891 = b[27] & w7314;
assign w15892 = b[26] & w7307;
assign w15893 = w2378 & w7312;
assign w15894 = ~w15891 & ~w15892;
assign w15895 = ~w15890 & w15894;
assign w15896 = ~w15893 & w15895;
assign w15897 = a[50] & ~w15896;
assign w15898 = ~a[50] & w15896;
assign w15899 = ~w15897 & ~w15898;
assign w15900 = ~w15679 & ~w15681;
assign w15901 = b[22] & w8515;
assign w15902 = b[24] & w8202;
assign w15903 = b[23] & w8200;
assign w15904 = w1895 & w8195;
assign w15905 = ~w15902 & ~w15903;
assign w15906 = ~w15901 & w15905;
assign w15907 = ~w15904 & w15906;
assign w15908 = a[53] & ~w15907;
assign w15909 = ~a[53] & w15907;
assign w15910 = ~w15908 & ~w15909;
assign w15911 = ~w15656 & ~w15659;
assign w15912 = b[16] & w10496;
assign w15913 = b[17] & w10146;
assign w15914 = b[18] & w10148;
assign w15915 = ~w1108 & w10141;
assign w15916 = ~w15913 & ~w15914;
assign w15917 = ~w15912 & w15916;
assign w15918 = ~w15915 & w15917;
assign w15919 = a[59] & ~w15918;
assign w15920 = ~a[59] & w15918;
assign w15921 = ~w15919 & ~w15920;
assign w15922 = ~w15650 & ~w15653;
assign w15923 = b[13] & w11561;
assign w15924 = b[14] & w11194;
assign w15925 = b[15] & w11196;
assign w15926 = ~w799 & w11189;
assign w15927 = ~w15924 & ~w15925;
assign w15928 = ~w15923 & w15927;
assign w15929 = ~w15926 & w15928;
assign w15930 = a[62] & ~w15929;
assign w15931 = ~a[62] & w15929;
assign w15932 = ~w15930 & ~w15931;
assign w15933 = b[11] & w11921;
assign w15934 = b[12] & w11923;
assign w15935 = ~w15933 & ~w15934;
assign w15936 = ~a[11] & ~w15394;
assign w15937 = a[11] & w15394;
assign w15938 = ~w15936 & ~w15937;
assign w15939 = ~w15935 & w15938;
assign w15940 = w15935 & ~w15938;
assign w15941 = ~w15939 & ~w15940;
assign w15942 = ~w15932 & ~w15941;
assign w15943 = w15932 & w15941;
assign w15944 = ~w15942 & ~w15943;
assign w15945 = ~w15922 & w15944;
assign w15946 = w15922 & ~w15944;
assign w15947 = ~w15945 & ~w15946;
assign w15948 = w15921 & w15947;
assign w15949 = ~w15921 & ~w15947;
assign w15950 = ~w15948 & ~w15949;
assign w15951 = w15911 & ~w15950;
assign w15952 = ~w15911 & w15950;
assign w15953 = ~w15951 & ~w15952;
assign w15954 = b[19] & w9482;
assign w15955 = b[21] & w9160;
assign w15956 = b[20] & w9165;
assign w15957 = w1467 & w9158;
assign w15958 = ~w15955 & ~w15956;
assign w15959 = ~w15954 & w15958;
assign w15960 = ~w15957 & w15959;
assign w15961 = a[56] & ~w15960;
assign w15962 = ~a[56] & w15960;
assign w15963 = ~w15961 & ~w15962;
assign w15964 = w15953 & w15963;
assign w15965 = ~w15953 & ~w15963;
assign w15966 = ~w15964 & ~w15965;
assign w15967 = ~w15662 & ~w15676;
assign w15968 = w15966 & ~w15967;
assign w15969 = ~w15966 & w15967;
assign w15970 = ~w15968 & ~w15969;
assign w15971 = ~w15910 & ~w15970;
assign w15972 = w15910 & w15970;
assign w15973 = ~w15971 & ~w15972;
assign w15974 = ~w15900 & w15973;
assign w15975 = w15900 & ~w15973;
assign w15976 = ~w15974 & ~w15975;
assign w15977 = w15899 & w15976;
assign w15978 = ~w15899 & ~w15976;
assign w15979 = ~w15977 & ~w15978;
assign w15980 = w15889 & ~w15979;
assign w15981 = ~w15889 & w15979;
assign w15982 = ~w15980 & ~w15981;
assign w15983 = b[28] & w6732;
assign w15984 = b[30] & w6476;
assign w15985 = b[29] & w6474;
assign w15986 = ~w2908 & w6469;
assign w15987 = ~w15984 & ~w15985;
assign w15988 = ~w15983 & w15987;
assign w15989 = ~w15986 & w15988;
assign w15990 = a[47] & ~w15989;
assign w15991 = ~a[47] & w15989;
assign w15992 = ~w15990 & ~w15991;
assign w15993 = ~w15982 & ~w15992;
assign w15994 = w15982 & w15992;
assign w15995 = ~w15993 & ~w15994;
assign w15996 = w15888 & w15995;
assign w15997 = ~w15888 & ~w15995;
assign w15998 = ~w15996 & ~w15997;
assign w15999 = w15887 & ~w15998;
assign w16000 = ~w15887 & w15998;
assign w16001 = ~w15999 & ~w16000;
assign w16002 = ~w15877 & w16001;
assign w16003 = w15877 & ~w16001;
assign w16004 = ~w16002 & ~w16003;
assign w16005 = w15876 & w16004;
assign w16006 = ~w15876 & ~w16004;
assign w16007 = ~w16005 & ~w16006;
assign w16008 = w15866 & ~w16007;
assign w16009 = ~w15866 & w16007;
assign w16010 = ~w16008 & ~w16009;
assign w16011 = b[37] & w4453;
assign w16012 = b[38] & w4241;
assign w16013 = b[39] & w4243;
assign w16014 = w4236 & ~w4812;
assign w16015 = ~w16012 & ~w16013;
assign w16016 = ~w16011 & w16015;
assign w16017 = ~w16014 & w16016;
assign w16018 = a[38] & ~w16017;
assign w16019 = ~a[38] & w16017;
assign w16020 = ~w16018 & ~w16019;
assign w16021 = w16010 & w16020;
assign w16022 = ~w16010 & ~w16020;
assign w16023 = ~w16021 & ~w16022;
assign w16024 = ~w15865 & w16023;
assign w16025 = w15865 & ~w16023;
assign w16026 = ~w16024 & ~w16025;
assign w16027 = w15864 & w16026;
assign w16028 = ~w15864 & ~w16026;
assign w16029 = ~w16027 & ~w16028;
assign w16030 = w15854 & ~w16029;
assign w16031 = ~w15854 & w16029;
assign w16032 = ~w16030 & ~w16031;
assign w16033 = ~w15764 & ~w15767;
assign w16034 = b[43] & w3177;
assign w16035 = b[44] & w2973;
assign w16036 = b[45] & w2978;
assign w16037 = w2980 & w6334;
assign w16038 = ~w16035 & ~w16036;
assign w16039 = ~w16034 & w16038;
assign w16040 = ~w16037 & w16039;
assign w16041 = a[32] & ~w16040;
assign w16042 = ~a[32] & w16040;
assign w16043 = ~w16041 & ~w16042;
assign w16044 = ~w16033 & w16043;
assign w16045 = w16033 & ~w16043;
assign w16046 = ~w16044 & ~w16045;
assign w16047 = w16032 & w16046;
assign w16048 = ~w16032 & ~w16046;
assign w16049 = ~w16047 & ~w16048;
assign w16050 = ~w15781 & ~w15784;
assign w16051 = b[46] & ~w2622;
assign w16052 = b[48] & w2438;
assign w16053 = b[47] & w2436;
assign w16054 = w2432 & ~w7170;
assign w16055 = ~w16051 & ~w16052;
assign w16056 = ~w16053 & w16055;
assign w16057 = ~w16054 & w16056;
assign w16058 = a[29] & ~w16057;
assign w16059 = ~a[29] & w16057;
assign w16060 = ~w16058 & ~w16059;
assign w16061 = ~w16050 & w16060;
assign w16062 = w16050 & ~w16060;
assign w16063 = ~w16061 & ~w16062;
assign w16064 = ~w16049 & ~w16063;
assign w16065 = w16049 & w16063;
assign w16066 = ~w16064 & ~w16065;
assign w16067 = b[49] & ~w2114;
assign w16068 = b[50] & w1955;
assign w16069 = b[51] & w1957;
assign w16070 = w1951 & ~w8058;
assign w16071 = ~w16067 & ~w16068;
assign w16072 = ~w16069 & w16071;
assign w16073 = ~w16070 & w16072;
assign w16074 = a[26] & ~w16073;
assign w16075 = ~a[26] & w16073;
assign w16076 = ~w16074 & ~w16075;
assign w16077 = ~w15798 & ~w15801;
assign w16078 = w16076 & ~w16077;
assign w16079 = ~w16076 & w16077;
assign w16080 = ~w16078 & ~w16079;
assign w16081 = w16066 & w16080;
assign w16082 = ~w16066 & ~w16080;
assign w16083 = ~w16081 & ~w16082;
assign w16084 = ~w15814 & ~w15817;
assign w16085 = b[52] & ~w1676;
assign w16086 = b[53] & w1517;
assign w16087 = b[54] & w1519;
assign w16088 = w1513 & ~w8998;
assign w16089 = ~w16085 & ~w16086;
assign w16090 = ~w16087 & w16089;
assign w16091 = ~w16088 & w16090;
assign w16092 = a[23] & ~w16091;
assign w16093 = ~a[23] & w16091;
assign w16094 = ~w16092 & ~w16093;
assign w16095 = ~w16084 & w16094;
assign w16096 = w16084 & ~w16094;
assign w16097 = ~w16095 & ~w16096;
assign w16098 = ~w16083 & ~w16097;
assign w16099 = w16083 & w16097;
assign w16100 = ~w16098 & ~w16099;
assign w16101 = b[56] & w1154;
assign w16102 = b[55] & ~w1272;
assign w16103 = b[57] & w1156;
assign w16104 = w1150 & ~w9992;
assign w16105 = ~w16101 & ~w16102;
assign w16106 = ~w16103 & w16105;
assign w16107 = ~w16104 & w16106;
assign w16108 = a[20] & ~w16107;
assign w16109 = ~a[20] & w16107;
assign w16110 = ~w16108 & ~w16109;
assign w16111 = ~w15578 & ~w15820;
assign w16112 = w16110 & ~w16111;
assign w16113 = ~w16110 & w16111;
assign w16114 = ~w16112 & ~w16113;
assign w16115 = w16100 & w16114;
assign w16116 = ~w16100 & ~w16114;
assign w16117 = ~w16115 & ~w16116;
assign w16118 = (~w15566 & ~w15568) | (~w15566 & w25449) | (~w15568 & w25449);
assign w16119 = b[60] & w834;
assign w16120 = b[59] & w838;
assign w16121 = b[58] & ~w934;
assign w16122 = ~w16119 & ~w16120;
assign w16123 = ~w16121 & w16122;
assign w16124 = (w11035 & w25574) | (w11035 & w25575) | (w25574 & w25575);
assign w16125 = ~a[17] & w25732;
assign w16126 = ~w16124 & ~w16125;
assign w16127 = ~w16118 & w16126;
assign w16128 = w16118 & ~w16126;
assign w16129 = ~w16127 & ~w16128;
assign w16130 = ~w16117 & ~w16129;
assign w16131 = w16117 & w16129;
assign w16132 = ~w16130 & ~w16131;
assign w16133 = ~w15835 & ~w15838;
assign w16134 = b[62] & w573;
assign w16135 = b[63] & w575;
assign w16136 = b[61] & ~w649;
assign w16137 = w569 & w12132;
assign w16138 = ~w16134 & ~w16135;
assign w16139 = ~w16136 & w16138;
assign w16140 = ~w16137 & w16139;
assign w16141 = a[14] & ~w16140;
assign w16142 = ~a[14] & w16140;
assign w16143 = ~w16141 & ~w16142;
assign w16144 = ~w16133 & w16143;
assign w16145 = w16133 & ~w16143;
assign w16146 = ~w16144 & ~w16145;
assign w16147 = w16132 & w16146;
assign w16148 = ~w16132 & ~w16146;
assign w16149 = ~w16147 & ~w16148;
assign w16150 = ~w15853 & w16149;
assign w16151 = w15853 & ~w16149;
assign w16152 = ~w16150 & ~w16151;
assign w16153 = w15852 & ~w16152;
assign w16154 = ~w15852 & w16152;
assign w16155 = ~w16153 & ~w16154;
assign w16156 = ~w16144 & ~w16147;
assign w16157 = b[61] & w834;
assign w16158 = b[59] & ~w934;
assign w16159 = b[60] & w838;
assign w16160 = ~w16157 & ~w16158;
assign w16161 = ~w16159 & w16160;
assign w16162 = (w11400 & w25451) | (w11400 & w25452) | (w25451 & w25452);
assign w16163 = (~w11400 & w25453) | (~w11400 & w25454) | (w25453 & w25454);
assign w16164 = ~w16162 & ~w16163;
assign w16165 = ~w16112 & ~w16115;
assign w16166 = w16164 & ~w16165;
assign w16167 = ~w16164 & w16165;
assign w16168 = ~w16166 & ~w16167;
assign w16169 = b[47] & ~w2622;
assign w16170 = b[49] & w2438;
assign w16171 = b[48] & w2436;
assign w16172 = w2432 & ~w7468;
assign w16173 = ~w16169 & ~w16170;
assign w16174 = ~w16171 & w16173;
assign w16175 = ~w16172 & w16174;
assign w16176 = a[29] & ~w16175;
assign w16177 = ~a[29] & w16175;
assign w16178 = ~w16176 & ~w16177;
assign w16179 = ~w16044 & ~w16047;
assign w16180 = w16178 & ~w16179;
assign w16181 = ~w16178 & w16179;
assign w16182 = ~w16180 & ~w16181;
assign w16183 = ~w16021 & ~w16024;
assign w16184 = b[38] & w4453;
assign w16185 = b[39] & w4241;
assign w16186 = b[40] & w4243;
assign w16187 = w4236 & ~w5058;
assign w16188 = ~w16185 & ~w16186;
assign w16189 = ~w16184 & w16188;
assign w16190 = ~w16187 & w16189;
assign w16191 = a[38] & ~w16190;
assign w16192 = ~a[38] & w16190;
assign w16193 = ~w16191 & ~w16192;
assign w16194 = ~w16005 & ~w16009;
assign w16195 = b[35] & w5167;
assign w16196 = b[36] & w4918;
assign w16197 = b[37] & w4925;
assign w16198 = ~w4357 & w4923;
assign w16199 = ~w16196 & ~w16197;
assign w16200 = ~w16195 & w16199;
assign w16201 = ~w16198 & w16200;
assign w16202 = a[41] & ~w16201;
assign w16203 = ~a[41] & w16201;
assign w16204 = ~w16202 & ~w16203;
assign w16205 = ~w15999 & ~w16002;
assign w16206 = b[32] & w5939;
assign w16207 = b[34] & w5665;
assign w16208 = b[33] & w5670;
assign w16209 = ~w3710 & w5663;
assign w16210 = ~w16207 & ~w16208;
assign w16211 = ~w16206 & w16210;
assign w16212 = ~w16209 & w16211;
assign w16213 = a[44] & ~w16212;
assign w16214 = ~a[44] & w16212;
assign w16215 = ~w16213 & ~w16214;
assign w16216 = b[29] & w6732;
assign w16217 = b[31] & w6476;
assign w16218 = b[30] & w6474;
assign w16219 = ~w3112 & w6469;
assign w16220 = ~w16217 & ~w16218;
assign w16221 = ~w16216 & w16220;
assign w16222 = ~w16219 & w16221;
assign w16223 = a[47] & ~w16222;
assign w16224 = ~a[47] & w16222;
assign w16225 = ~w16223 & ~w16224;
assign w16226 = ~w15977 & ~w15981;
assign w16227 = b[26] & w7586;
assign w16228 = b[28] & w7314;
assign w16229 = b[27] & w7307;
assign w16230 = w2559 & w7312;
assign w16231 = ~w16228 & ~w16229;
assign w16232 = ~w16227 & w16231;
assign w16233 = ~w16230 & w16232;
assign w16234 = a[50] & ~w16233;
assign w16235 = ~a[50] & w16233;
assign w16236 = ~w16234 & ~w16235;
assign w16237 = b[23] & w8515;
assign w16238 = b[25] & w8202;
assign w16239 = b[24] & w8200;
assign w16240 = w2061 & w8195;
assign w16241 = ~w16238 & ~w16239;
assign w16242 = ~w16237 & w16241;
assign w16243 = ~w16240 & w16242;
assign w16244 = a[53] & ~w16243;
assign w16245 = ~a[53] & w16243;
assign w16246 = ~w16244 & ~w16245;
assign w16247 = b[20] & w9482;
assign w16248 = b[21] & w9165;
assign w16249 = b[22] & w9160;
assign w16250 = w1615 & w9158;
assign w16251 = ~w16248 & ~w16249;
assign w16252 = ~w16247 & w16251;
assign w16253 = ~w16250 & w16252;
assign w16254 = a[56] & ~w16253;
assign w16255 = ~a[56] & w16253;
assign w16256 = ~w16254 & ~w16255;
assign w16257 = b[17] & w10496;
assign w16258 = b[18] & w10146;
assign w16259 = b[19] & w10148;
assign w16260 = ~w1231 & w10141;
assign w16261 = ~w16258 & ~w16259;
assign w16262 = ~w16257 & w16261;
assign w16263 = ~w16260 & w16262;
assign w16264 = a[59] & ~w16263;
assign w16265 = ~a[59] & w16263;
assign w16266 = ~w16264 & ~w16265;
assign w16267 = ~w15943 & ~w15945;
assign w16268 = b[12] & w11921;
assign w16269 = b[13] & w11923;
assign w16270 = ~w16268 & ~w16269;
assign w16271 = ~w15936 & ~w15939;
assign w16272 = w16270 & ~w16271;
assign w16273 = ~w16270 & w16271;
assign w16274 = ~w16272 & ~w16273;
assign w16275 = b[14] & w11561;
assign w16276 = b[16] & w11196;
assign w16277 = b[15] & w11194;
assign w16278 = w905 & w11189;
assign w16279 = ~w16276 & ~w16277;
assign w16280 = ~w16275 & w16279;
assign w16281 = ~w16278 & w16280;
assign w16282 = a[62] & ~w16281;
assign w16283 = ~a[62] & w16281;
assign w16284 = ~w16282 & ~w16283;
assign w16285 = w16274 & w16284;
assign w16286 = ~w16274 & ~w16284;
assign w16287 = ~w16285 & ~w16286;
assign w16288 = ~w16267 & w16287;
assign w16289 = w16267 & ~w16287;
assign w16290 = ~w16288 & ~w16289;
assign w16291 = w16266 & w16290;
assign w16292 = ~w16266 & ~w16290;
assign w16293 = ~w16291 & ~w16292;
assign w16294 = ~w15948 & ~w15952;
assign w16295 = w16293 & ~w16294;
assign w16296 = ~w16293 & w16294;
assign w16297 = ~w16295 & ~w16296;
assign w16298 = w16256 & w16297;
assign w16299 = ~w16256 & ~w16297;
assign w16300 = ~w16298 & ~w16299;
assign w16301 = ~w15964 & ~w15968;
assign w16302 = w16300 & ~w16301;
assign w16303 = ~w16300 & w16301;
assign w16304 = ~w16302 & ~w16303;
assign w16305 = w16246 & w16304;
assign w16306 = ~w16246 & ~w16304;
assign w16307 = ~w16305 & ~w16306;
assign w16308 = ~w15972 & ~w15974;
assign w16309 = w16307 & ~w16308;
assign w16310 = ~w16307 & w16308;
assign w16311 = ~w16309 & ~w16310;
assign w16312 = ~w16236 & ~w16311;
assign w16313 = w16236 & w16311;
assign w16314 = ~w16312 & ~w16313;
assign w16315 = w16226 & ~w16314;
assign w16316 = ~w16226 & w16314;
assign w16317 = ~w16315 & ~w16316;
assign w16318 = w16225 & w16317;
assign w16319 = ~w16225 & ~w16317;
assign w16320 = ~w16318 & ~w16319;
assign w16321 = ~w15993 & ~w15996;
assign w16322 = ~w16320 & ~w16321;
assign w16323 = w16320 & w16321;
assign w16324 = ~w16322 & ~w16323;
assign w16325 = w16215 & w16324;
assign w16326 = ~w16215 & ~w16324;
assign w16327 = ~w16325 & ~w16326;
assign w16328 = w16205 & ~w16327;
assign w16329 = ~w16205 & w16327;
assign w16330 = ~w16328 & ~w16329;
assign w16331 = w16204 & w16330;
assign w16332 = ~w16204 & ~w16330;
assign w16333 = ~w16331 & ~w16332;
assign w16334 = w16194 & ~w16333;
assign w16335 = ~w16194 & w16333;
assign w16336 = ~w16334 & ~w16335;
assign w16337 = w16193 & w16336;
assign w16338 = ~w16193 & ~w16336;
assign w16339 = ~w16337 & ~w16338;
assign w16340 = w16183 & ~w16339;
assign w16341 = ~w16183 & w16339;
assign w16342 = ~w16340 & ~w16341;
assign w16343 = b[41] & w3785;
assign w16344 = b[43] & w3580;
assign w16345 = b[42] & w3578;
assign w16346 = w3573 & w5811;
assign w16347 = ~w16344 & ~w16345;
assign w16348 = ~w16343 & w16347;
assign w16349 = ~w16346 & w16348;
assign w16350 = a[35] & ~w16349;
assign w16351 = ~a[35] & w16349;
assign w16352 = ~w16350 & ~w16351;
assign w16353 = w16342 & w16352;
assign w16354 = ~w16342 & ~w16352;
assign w16355 = ~w16353 & ~w16354;
assign w16356 = ~w16027 & ~w16031;
assign w16357 = b[44] & w3177;
assign w16358 = b[46] & w2978;
assign w16359 = b[45] & w2973;
assign w16360 = w2980 & ~w6613;
assign w16361 = ~w16358 & ~w16359;
assign w16362 = ~w16357 & w16361;
assign w16363 = ~w16360 & w16362;
assign w16364 = a[32] & ~w16363;
assign w16365 = ~a[32] & w16363;
assign w16366 = ~w16364 & ~w16365;
assign w16367 = ~w16356 & w16366;
assign w16368 = w16356 & ~w16366;
assign w16369 = ~w16367 & ~w16368;
assign w16370 = w16355 & w16369;
assign w16371 = ~w16355 & ~w16369;
assign w16372 = ~w16370 & ~w16371;
assign w16373 = w16182 & w16372;
assign w16374 = ~w16182 & ~w16372;
assign w16375 = ~w16373 & ~w16374;
assign w16376 = ~w16061 & ~w16065;
assign w16377 = b[51] & w1955;
assign w16378 = b[50] & ~w2114;
assign w16379 = b[52] & w1957;
assign w16380 = w1951 & ~w8371;
assign w16381 = ~w16377 & ~w16378;
assign w16382 = ~w16379 & w16381;
assign w16383 = ~w16380 & w16382;
assign w16384 = a[26] & ~w16383;
assign w16385 = ~a[26] & w16383;
assign w16386 = ~w16384 & ~w16385;
assign w16387 = ~w16376 & w16386;
assign w16388 = w16376 & ~w16386;
assign w16389 = ~w16387 & ~w16388;
assign w16390 = ~w16375 & ~w16389;
assign w16391 = w16375 & w16389;
assign w16392 = ~w16390 & ~w16391;
assign w16393 = b[53] & ~w1676;
assign w16394 = b[55] & w1519;
assign w16395 = b[54] & w1517;
assign w16396 = w1513 & ~w9330;
assign w16397 = ~w16393 & ~w16394;
assign w16398 = ~w16395 & w16397;
assign w16399 = ~w16396 & w16398;
assign w16400 = a[23] & ~w16399;
assign w16401 = ~a[23] & w16399;
assign w16402 = ~w16400 & ~w16401;
assign w16403 = ~w16078 & ~w16081;
assign w16404 = w16402 & ~w16403;
assign w16405 = ~w16402 & w16403;
assign w16406 = ~w16404 & ~w16405;
assign w16407 = w16392 & w16406;
assign w16408 = ~w16392 & ~w16406;
assign w16409 = ~w16407 & ~w16408;
assign w16410 = ~w16095 & ~w16099;
assign w16411 = b[56] & ~w1272;
assign w16412 = b[57] & w1154;
assign w16413 = b[58] & w1156;
assign w16414 = ~w16411 & ~w16412;
assign w16415 = ~w16413 & w16414;
assign w16416 = a[20] & w25733;
assign w16417 = (w10339 & w25576) | (w10339 & w25577) | (w25576 & w25577);
assign w16418 = ~w16416 & ~w16417;
assign w16419 = ~w16410 & w16418;
assign w16420 = w16410 & ~w16418;
assign w16421 = ~w16419 & ~w16420;
assign w16422 = w16409 & w16421;
assign w16423 = ~w16409 & ~w16421;
assign w16424 = ~w16422 & ~w16423;
assign w16425 = w16168 & w16424;
assign w16426 = ~w16168 & ~w16424;
assign w16427 = ~w16425 & ~w16426;
assign w16428 = (~w16127 & ~w16129) | (~w16127 & w25578) | (~w16129 & w25578);
assign w16429 = b[62] & ~w649;
assign w16430 = b[63] & w573;
assign w16431 = ~w12153 & w25579;
assign w16432 = ~w16429 & ~w16430;
assign w16433 = ~w16431 & w16432;
assign w16434 = a[14] & ~w16433;
assign w16435 = ~a[14] & w16433;
assign w16436 = ~w16434 & ~w16435;
assign w16437 = ~w16428 & w16436;
assign w16438 = w16428 & ~w16436;
assign w16439 = ~w16437 & ~w16438;
assign w16440 = w16427 & w16439;
assign w16441 = ~w16427 & ~w16439;
assign w16442 = ~w16440 & ~w16441;
assign w16443 = w16156 & ~w16442;
assign w16444 = ~w16156 & w16442;
assign w16445 = ~w16443 & ~w16444;
assign w16446 = (w15542 & w24419) | (w15542 & w24420) | (w24419 & w24420);
assign w16447 = w16445 & w16446;
assign w16448 = ~w16445 & ~w16446;
assign w16449 = ~w16447 & ~w16448;
assign w16450 = (~w15542 & w24421) | (~w15542 & w24422) | (w24421 & w24422);
assign w16451 = ~w16437 & ~w16440;
assign w16452 = b[42] & w3785;
assign w16453 = b[44] & w3580;
assign w16454 = b[43] & w3578;
assign w16455 = w3573 & w6069;
assign w16456 = ~w16453 & ~w16454;
assign w16457 = ~w16452 & w16456;
assign w16458 = ~w16455 & w16457;
assign w16459 = a[35] & ~w16458;
assign w16460 = ~a[35] & w16458;
assign w16461 = ~w16459 & ~w16460;
assign w16462 = ~w16335 & ~w16337;
assign w16463 = b[39] & w4453;
assign w16464 = b[41] & w4243;
assign w16465 = b[40] & w4241;
assign w16466 = w4236 & w5302;
assign w16467 = ~w16464 & ~w16465;
assign w16468 = ~w16463 & w16467;
assign w16469 = ~w16466 & w16468;
assign w16470 = a[38] & ~w16469;
assign w16471 = ~a[38] & w16469;
assign w16472 = ~w16470 & ~w16471;
assign w16473 = ~w16329 & ~w16331;
assign w16474 = b[36] & w5167;
assign w16475 = b[38] & w4925;
assign w16476 = b[37] & w4918;
assign w16477 = w4582 & w4923;
assign w16478 = ~w16475 & ~w16476;
assign w16479 = ~w16474 & w16478;
assign w16480 = ~w16477 & w16479;
assign w16481 = a[41] & ~w16480;
assign w16482 = ~a[41] & w16480;
assign w16483 = ~w16481 & ~w16482;
assign w16484 = b[33] & w5939;
assign w16485 = b[35] & w5665;
assign w16486 = b[34] & w5670;
assign w16487 = w3918 & w5663;
assign w16488 = ~w16485 & ~w16486;
assign w16489 = ~w16484 & w16488;
assign w16490 = ~w16487 & w16489;
assign w16491 = a[44] & ~w16490;
assign w16492 = ~a[44] & w16490;
assign w16493 = ~w16491 & ~w16492;
assign w16494 = ~w16316 & ~w16318;
assign w16495 = b[30] & w6732;
assign w16496 = b[31] & w6474;
assign w16497 = b[32] & w6476;
assign w16498 = w3304 & w6469;
assign w16499 = ~w16496 & ~w16497;
assign w16500 = ~w16495 & w16499;
assign w16501 = ~w16498 & w16500;
assign w16502 = a[47] & ~w16501;
assign w16503 = ~a[47] & w16501;
assign w16504 = ~w16502 & ~w16503;
assign w16505 = ~w16302 & ~w16305;
assign w16506 = ~w16295 & ~w16298;
assign w16507 = b[21] & w9482;
assign w16508 = b[23] & w9160;
assign w16509 = b[22] & w9165;
assign w16510 = w1755 & w9158;
assign w16511 = ~w16508 & ~w16509;
assign w16512 = ~w16507 & w16511;
assign w16513 = ~w16510 & w16512;
assign w16514 = a[56] & ~w16513;
assign w16515 = ~a[56] & w16513;
assign w16516 = ~w16514 & ~w16515;
assign w16517 = ~w16272 & ~w16285;
assign w16518 = b[13] & w11921;
assign w16519 = b[14] & w11923;
assign w16520 = ~w16518 & ~w16519;
assign w16521 = w16270 & ~w16520;
assign w16522 = ~w16270 & w16520;
assign w16523 = ~w16521 & ~w16522;
assign w16524 = b[15] & w11561;
assign w16525 = b[16] & w11194;
assign w16526 = b[17] & w11196;
assign w16527 = w1008 & w11189;
assign w16528 = ~w16525 & ~w16526;
assign w16529 = ~w16524 & w16528;
assign w16530 = ~w16527 & w16529;
assign w16531 = a[62] & ~w16530;
assign w16532 = ~a[62] & w16530;
assign w16533 = ~w16531 & ~w16532;
assign w16534 = w16523 & w16533;
assign w16535 = ~w16523 & ~w16533;
assign w16536 = ~w16534 & ~w16535;
assign w16537 = w16517 & ~w16536;
assign w16538 = ~w16517 & w16536;
assign w16539 = ~w16537 & ~w16538;
assign w16540 = b[18] & w10496;
assign w16541 = b[19] & w10146;
assign w16542 = b[20] & w10148;
assign w16543 = w1347 & w10141;
assign w16544 = ~w16541 & ~w16542;
assign w16545 = ~w16540 & w16544;
assign w16546 = ~w16543 & w16545;
assign w16547 = a[59] & ~w16546;
assign w16548 = ~a[59] & w16546;
assign w16549 = ~w16547 & ~w16548;
assign w16550 = w16539 & w16549;
assign w16551 = ~w16539 & ~w16549;
assign w16552 = ~w16550 & ~w16551;
assign w16553 = ~w16288 & ~w16291;
assign w16554 = w16552 & ~w16553;
assign w16555 = ~w16552 & w16553;
assign w16556 = ~w16554 & ~w16555;
assign w16557 = ~w16516 & ~w16556;
assign w16558 = w16516 & w16556;
assign w16559 = ~w16557 & ~w16558;
assign w16560 = w16506 & ~w16559;
assign w16561 = ~w16506 & w16559;
assign w16562 = ~w16560 & ~w16561;
assign w16563 = b[24] & w8515;
assign w16564 = b[26] & w8202;
assign w16565 = b[25] & w8200;
assign w16566 = w2219 & w8195;
assign w16567 = ~w16564 & ~w16565;
assign w16568 = ~w16563 & w16567;
assign w16569 = ~w16566 & w16568;
assign w16570 = a[53] & ~w16569;
assign w16571 = ~a[53] & w16569;
assign w16572 = ~w16570 & ~w16571;
assign w16573 = w16562 & w16572;
assign w16574 = ~w16562 & ~w16572;
assign w16575 = ~w16573 & ~w16574;
assign w16576 = w16505 & ~w16575;
assign w16577 = ~w16505 & w16575;
assign w16578 = ~w16576 & ~w16577;
assign w16579 = b[27] & w7586;
assign w16580 = b[28] & w7307;
assign w16581 = b[29] & w7314;
assign w16582 = w2734 & w7312;
assign w16583 = ~w16580 & ~w16581;
assign w16584 = ~w16579 & w16583;
assign w16585 = ~w16582 & w16584;
assign w16586 = a[50] & ~w16585;
assign w16587 = ~a[50] & w16585;
assign w16588 = ~w16586 & ~w16587;
assign w16589 = w16578 & w16588;
assign w16590 = ~w16578 & ~w16588;
assign w16591 = ~w16589 & ~w16590;
assign w16592 = ~w16309 & ~w16313;
assign w16593 = w16591 & ~w16592;
assign w16594 = ~w16591 & w16592;
assign w16595 = ~w16593 & ~w16594;
assign w16596 = w16504 & w16595;
assign w16597 = ~w16504 & ~w16595;
assign w16598 = ~w16596 & ~w16597;
assign w16599 = ~w16494 & w16598;
assign w16600 = w16494 & ~w16598;
assign w16601 = ~w16599 & ~w16600;
assign w16602 = w16493 & w16601;
assign w16603 = ~w16493 & ~w16601;
assign w16604 = ~w16602 & ~w16603;
assign w16605 = ~w16323 & ~w16325;
assign w16606 = w16604 & ~w16605;
assign w16607 = ~w16604 & w16605;
assign w16608 = ~w16606 & ~w16607;
assign w16609 = ~w16483 & ~w16608;
assign w16610 = w16483 & w16608;
assign w16611 = ~w16609 & ~w16610;
assign w16612 = w16473 & ~w16611;
assign w16613 = ~w16473 & w16611;
assign w16614 = ~w16612 & ~w16613;
assign w16615 = w16472 & w16614;
assign w16616 = ~w16472 & ~w16614;
assign w16617 = ~w16615 & ~w16616;
assign w16618 = w16462 & ~w16617;
assign w16619 = ~w16462 & w16617;
assign w16620 = ~w16618 & ~w16619;
assign w16621 = ~w16461 & ~w16620;
assign w16622 = w16461 & w16620;
assign w16623 = ~w16621 & ~w16622;
assign w16624 = ~w16341 & ~w16353;
assign w16625 = b[45] & w3177;
assign w16626 = b[46] & w2973;
assign w16627 = b[47] & w2978;
assign w16628 = w2980 & w6889;
assign w16629 = ~w16626 & ~w16627;
assign w16630 = ~w16625 & w16629;
assign w16631 = ~w16628 & w16630;
assign w16632 = a[32] & ~w16631;
assign w16633 = ~a[32] & w16631;
assign w16634 = ~w16632 & ~w16633;
assign w16635 = ~w16624 & w16634;
assign w16636 = w16624 & ~w16634;
assign w16637 = ~w16635 & ~w16636;
assign w16638 = w16623 & w16637;
assign w16639 = ~w16623 & ~w16637;
assign w16640 = ~w16638 & ~w16639;
assign w16641 = ~w16367 & ~w16370;
assign w16642 = b[48] & ~w2622;
assign w16643 = b[49] & w2436;
assign w16644 = b[50] & w2438;
assign w16645 = w2432 & w7759;
assign w16646 = ~w16642 & ~w16643;
assign w16647 = ~w16644 & w16646;
assign w16648 = ~w16645 & w16647;
assign w16649 = a[29] & ~w16648;
assign w16650 = ~a[29] & w16648;
assign w16651 = ~w16649 & ~w16650;
assign w16652 = ~w16641 & w16651;
assign w16653 = w16641 & ~w16651;
assign w16654 = ~w16652 & ~w16653;
assign w16655 = ~w16640 & ~w16654;
assign w16656 = w16640 & w16654;
assign w16657 = ~w16655 & ~w16656;
assign w16658 = b[53] & w1957;
assign w16659 = b[51] & ~w2114;
assign w16660 = b[52] & w1955;
assign w16661 = ~w16658 & ~w16659;
assign w16662 = ~w16660 & w16661;
assign w16663 = (w16662 & ~w8683) | (w16662 & w25456) | (~w8683 & w25456);
assign w16664 = a[26] & ~w16663;
assign w16665 = ~a[26] & w16663;
assign w16666 = ~w16664 & ~w16665;
assign w16667 = ~w16180 & ~w16373;
assign w16668 = w16666 & ~w16667;
assign w16669 = ~w16666 & w16667;
assign w16670 = ~w16668 & ~w16669;
assign w16671 = w16657 & w16670;
assign w16672 = ~w16657 & ~w16670;
assign w16673 = ~w16671 & ~w16672;
assign w16674 = b[54] & ~w1676;
assign w16675 = b[56] & w1519;
assign w16676 = b[55] & w1517;
assign w16677 = w1513 & w9657;
assign w16678 = ~w16674 & ~w16675;
assign w16679 = ~w16676 & w16678;
assign w16680 = ~w16677 & w16679;
assign w16681 = a[23] & ~w16680;
assign w16682 = ~a[23] & w16680;
assign w16683 = ~w16681 & ~w16682;
assign w16684 = ~w16387 & ~w16391;
assign w16685 = w16683 & ~w16684;
assign w16686 = ~w16683 & w16684;
assign w16687 = ~w16685 & ~w16686;
assign w16688 = w16673 & w16687;
assign w16689 = ~w16673 & ~w16687;
assign w16690 = ~w16688 & ~w16689;
assign w16691 = b[59] & w1156;
assign w16692 = b[58] & w1154;
assign w16693 = b[57] & ~w1272;
assign w16694 = ~w16691 & ~w16692;
assign w16695 = ~w16693 & w16694;
assign w16696 = (w10371 & w25580) | (w10371 & w25581) | (w25580 & w25581);
assign w16697 = (~w10371 & w25582) | (~w10371 & w25583) | (w25582 & w25583);
assign w16698 = ~w16696 & ~w16697;
assign w16699 = ~w16404 & ~w16407;
assign w16700 = w16698 & ~w16699;
assign w16701 = ~w16698 & w16699;
assign w16702 = ~w16700 & ~w16701;
assign w16703 = w16690 & w16702;
assign w16704 = ~w16690 & ~w16702;
assign w16705 = ~w16703 & ~w16704;
assign w16706 = ~w16419 & ~w16422;
assign w16707 = b[60] & ~w934;
assign w16708 = b[61] & w838;
assign w16709 = b[62] & w834;
assign w16710 = ~w16707 & ~w16708;
assign w16711 = ~w16709 & w16710;
assign w16712 = (w11763 & w25458) | (w11763 & w25459) | (w25458 & w25459);
assign w16713 = (~w11763 & w25460) | (~w11763 & w25461) | (w25460 & w25461);
assign w16714 = ~w16712 & ~w16713;
assign w16715 = ~w16706 & w16714;
assign w16716 = w16706 & ~w16714;
assign w16717 = ~w16715 & ~w16716;
assign w16718 = w16705 & w16717;
assign w16719 = ~w16705 & ~w16717;
assign w16720 = ~w16718 & ~w16719;
assign w16721 = (~w16166 & ~w16168) | (~w16166 & w25584) | (~w16168 & w25584);
assign w16722 = w569 & ~w12154;
assign w16723 = w649 & ~w16722;
assign w16724 = b[63] & ~w16723;
assign w16725 = ~a[14] & ~w16724;
assign w16726 = a[14] & w16724;
assign w16727 = ~w16725 & ~w16726;
assign w16728 = ~w16721 & w16727;
assign w16729 = w16721 & ~w16727;
assign w16730 = ~w16728 & ~w16729;
assign w16731 = w16720 & w16730;
assign w16732 = ~w16720 & ~w16730;
assign w16733 = ~w16731 & ~w16732;
assign w16734 = ~w16451 & w16733;
assign w16735 = w16451 & ~w16733;
assign w16736 = ~w16734 & ~w16735;
assign w16737 = ~w16443 & w16736;
assign w16738 = ~w16450 & w16737;
assign w16739 = ~w16444 & ~w16736;
assign w16740 = ~w16447 & w16739;
assign w16741 = ~w16738 & ~w16740;
assign w16742 = b[53] & w1955;
assign w16743 = b[54] & w1957;
assign w16744 = b[52] & ~w2114;
assign w16745 = w1951 & ~w8998;
assign w16746 = ~w16742 & ~w16743;
assign w16747 = ~w16744 & w16746;
assign w16748 = ~w16745 & w16747;
assign w16749 = a[26] & ~w16748;
assign w16750 = ~a[26] & w16748;
assign w16751 = ~w16749 & ~w16750;
assign w16752 = ~w16668 & ~w16671;
assign w16753 = w16751 & ~w16752;
assign w16754 = ~w16751 & w16752;
assign w16755 = ~w16753 & ~w16754;
assign w16756 = ~w16613 & ~w16615;
assign w16757 = b[40] & w4453;
assign w16758 = b[42] & w4243;
assign w16759 = b[41] & w4241;
assign w16760 = w4236 & w5548;
assign w16761 = ~w16758 & ~w16759;
assign w16762 = ~w16757 & w16761;
assign w16763 = ~w16760 & w16762;
assign w16764 = a[38] & ~w16763;
assign w16765 = ~a[38] & w16763;
assign w16766 = ~w16764 & ~w16765;
assign w16767 = ~w16606 & ~w16610;
assign w16768 = ~w16599 & ~w16602;
assign w16769 = b[34] & w5939;
assign w16770 = b[36] & w5665;
assign w16771 = b[35] & w5670;
assign w16772 = w4129 & w5663;
assign w16773 = ~w16770 & ~w16771;
assign w16774 = ~w16769 & w16773;
assign w16775 = ~w16772 & w16774;
assign w16776 = a[44] & ~w16775;
assign w16777 = ~a[44] & w16775;
assign w16778 = ~w16776 & ~w16777;
assign w16779 = ~w16593 & ~w16596;
assign w16780 = ~w16561 & ~w16573;
assign w16781 = b[25] & w8515;
assign w16782 = b[26] & w8200;
assign w16783 = b[27] & w8202;
assign w16784 = w2378 & w8195;
assign w16785 = ~w16782 & ~w16783;
assign w16786 = ~w16781 & w16785;
assign w16787 = ~w16784 & w16786;
assign w16788 = a[53] & ~w16787;
assign w16789 = ~a[53] & w16787;
assign w16790 = ~w16788 & ~w16789;
assign w16791 = ~w16554 & ~w16558;
assign w16792 = ~w16521 & ~w16534;
assign w16793 = b[16] & w11561;
assign w16794 = b[17] & w11194;
assign w16795 = b[18] & w11196;
assign w16796 = ~w1108 & w11189;
assign w16797 = ~w16794 & ~w16795;
assign w16798 = ~w16793 & w16797;
assign w16799 = ~w16796 & w16798;
assign w16800 = a[62] & ~w16799;
assign w16801 = ~a[62] & w16799;
assign w16802 = ~w16800 & ~w16801;
assign w16803 = b[14] & w11921;
assign w16804 = b[15] & w11923;
assign w16805 = ~w16803 & ~w16804;
assign w16806 = ~a[14] & ~w16805;
assign w16807 = a[14] & w16805;
assign w16808 = ~w16806 & ~w16807;
assign w16809 = ~w16270 & w16808;
assign w16810 = w16270 & ~w16808;
assign w16811 = ~w16809 & ~w16810;
assign w16812 = w16802 & w16811;
assign w16813 = ~w16802 & ~w16811;
assign w16814 = ~w16812 & ~w16813;
assign w16815 = w16792 & ~w16814;
assign w16816 = ~w16792 & w16814;
assign w16817 = ~w16815 & ~w16816;
assign w16818 = b[19] & w10496;
assign w16819 = b[21] & w10148;
assign w16820 = b[20] & w10146;
assign w16821 = w1467 & w10141;
assign w16822 = ~w16819 & ~w16820;
assign w16823 = ~w16818 & w16822;
assign w16824 = ~w16821 & w16823;
assign w16825 = a[59] & ~w16824;
assign w16826 = ~a[59] & w16824;
assign w16827 = ~w16825 & ~w16826;
assign w16828 = w16817 & w16827;
assign w16829 = ~w16817 & ~w16827;
assign w16830 = ~w16828 & ~w16829;
assign w16831 = ~w16538 & ~w16550;
assign w16832 = ~w16830 & w16831;
assign w16833 = w16830 & ~w16831;
assign w16834 = ~w16832 & ~w16833;
assign w16835 = b[22] & w9482;
assign w16836 = b[24] & w9160;
assign w16837 = b[23] & w9165;
assign w16838 = w1895 & w9158;
assign w16839 = ~w16836 & ~w16837;
assign w16840 = ~w16835 & w16839;
assign w16841 = ~w16838 & w16840;
assign w16842 = a[56] & ~w16841;
assign w16843 = ~a[56] & w16841;
assign w16844 = ~w16842 & ~w16843;
assign w16845 = ~w16834 & ~w16844;
assign w16846 = w16834 & w16844;
assign w16847 = ~w16845 & ~w16846;
assign w16848 = w16791 & w16847;
assign w16849 = ~w16791 & ~w16847;
assign w16850 = ~w16848 & ~w16849;
assign w16851 = w16790 & ~w16850;
assign w16852 = ~w16790 & w16850;
assign w16853 = ~w16851 & ~w16852;
assign w16854 = w16780 & ~w16853;
assign w16855 = ~w16780 & w16853;
assign w16856 = ~w16854 & ~w16855;
assign w16857 = b[28] & w7586;
assign w16858 = b[29] & w7307;
assign w16859 = b[30] & w7314;
assign w16860 = ~w2908 & w7312;
assign w16861 = ~w16858 & ~w16859;
assign w16862 = ~w16857 & w16861;
assign w16863 = ~w16860 & w16862;
assign w16864 = a[50] & ~w16863;
assign w16865 = ~a[50] & w16863;
assign w16866 = ~w16864 & ~w16865;
assign w16867 = w16856 & w16866;
assign w16868 = ~w16856 & ~w16866;
assign w16869 = ~w16867 & ~w16868;
assign w16870 = ~w16577 & ~w16589;
assign w16871 = ~w16869 & w16870;
assign w16872 = w16869 & ~w16870;
assign w16873 = ~w16871 & ~w16872;
assign w16874 = b[31] & w6732;
assign w16875 = b[33] & w6476;
assign w16876 = b[32] & w6474;
assign w16877 = w3499 & w6469;
assign w16878 = ~w16875 & ~w16876;
assign w16879 = ~w16874 & w16878;
assign w16880 = ~w16877 & w16879;
assign w16881 = a[47] & ~w16880;
assign w16882 = ~a[47] & w16880;
assign w16883 = ~w16881 & ~w16882;
assign w16884 = w16873 & w16883;
assign w16885 = ~w16873 & ~w16883;
assign w16886 = ~w16884 & ~w16885;
assign w16887 = ~w16779 & w16886;
assign w16888 = w16779 & ~w16886;
assign w16889 = ~w16887 & ~w16888;
assign w16890 = w16778 & w16889;
assign w16891 = ~w16778 & ~w16889;
assign w16892 = ~w16890 & ~w16891;
assign w16893 = w16768 & ~w16892;
assign w16894 = ~w16768 & w16892;
assign w16895 = ~w16893 & ~w16894;
assign w16896 = b[37] & w5167;
assign w16897 = b[39] & w4925;
assign w16898 = b[38] & w4918;
assign w16899 = ~w4812 & w4923;
assign w16900 = ~w16897 & ~w16898;
assign w16901 = ~w16896 & w16900;
assign w16902 = ~w16899 & w16901;
assign w16903 = a[41] & ~w16902;
assign w16904 = ~a[41] & w16902;
assign w16905 = ~w16903 & ~w16904;
assign w16906 = w16895 & w16905;
assign w16907 = ~w16895 & ~w16905;
assign w16908 = ~w16906 & ~w16907;
assign w16909 = ~w16767 & w16908;
assign w16910 = w16767 & ~w16908;
assign w16911 = ~w16909 & ~w16910;
assign w16912 = w16766 & w16911;
assign w16913 = ~w16766 & ~w16911;
assign w16914 = ~w16912 & ~w16913;
assign w16915 = w16756 & ~w16914;
assign w16916 = ~w16756 & w16914;
assign w16917 = ~w16915 & ~w16916;
assign w16918 = b[43] & w3785;
assign w16919 = b[44] & w3578;
assign w16920 = b[45] & w3580;
assign w16921 = w3573 & w6334;
assign w16922 = ~w16919 & ~w16920;
assign w16923 = ~w16918 & w16922;
assign w16924 = ~w16921 & w16923;
assign w16925 = a[35] & ~w16924;
assign w16926 = ~a[35] & w16924;
assign w16927 = ~w16925 & ~w16926;
assign w16928 = w16917 & w16927;
assign w16929 = ~w16917 & ~w16927;
assign w16930 = ~w16928 & ~w16929;
assign w16931 = ~w16619 & ~w16622;
assign w16932 = ~w16930 & w16931;
assign w16933 = w16930 & ~w16931;
assign w16934 = ~w16932 & ~w16933;
assign w16935 = ~w16635 & ~w16638;
assign w16936 = b[46] & w3177;
assign w16937 = b[48] & w2978;
assign w16938 = b[47] & w2973;
assign w16939 = w2980 & ~w7170;
assign w16940 = ~w16937 & ~w16938;
assign w16941 = ~w16936 & w16940;
assign w16942 = ~w16939 & w16941;
assign w16943 = a[32] & ~w16942;
assign w16944 = ~a[32] & w16942;
assign w16945 = ~w16943 & ~w16944;
assign w16946 = ~w16935 & w16945;
assign w16947 = w16935 & ~w16945;
assign w16948 = ~w16946 & ~w16947;
assign w16949 = w16934 & w16948;
assign w16950 = ~w16934 & ~w16948;
assign w16951 = ~w16949 & ~w16950;
assign w16952 = b[51] & w2438;
assign w16953 = b[50] & w2436;
assign w16954 = b[49] & ~w2622;
assign w16955 = w2432 & ~w8058;
assign w16956 = ~w16952 & ~w16953;
assign w16957 = ~w16954 & w16956;
assign w16958 = ~w16955 & w16957;
assign w16959 = a[29] & ~w16958;
assign w16960 = ~a[29] & w16958;
assign w16961 = ~w16959 & ~w16960;
assign w16962 = ~w16652 & ~w16656;
assign w16963 = w16961 & ~w16962;
assign w16964 = ~w16961 & w16962;
assign w16965 = ~w16963 & ~w16964;
assign w16966 = w16951 & w16965;
assign w16967 = ~w16951 & ~w16965;
assign w16968 = ~w16966 & ~w16967;
assign w16969 = w16755 & w16968;
assign w16970 = ~w16755 & ~w16968;
assign w16971 = ~w16969 & ~w16970;
assign w16972 = ~w16685 & ~w16688;
assign w16973 = b[55] & ~w1676;
assign w16974 = b[57] & w1519;
assign w16975 = b[56] & w1517;
assign w16976 = w1513 & ~w9992;
assign w16977 = ~w16973 & ~w16974;
assign w16978 = ~w16975 & w16977;
assign w16979 = ~w16976 & w16978;
assign w16980 = a[23] & ~w16979;
assign w16981 = ~a[23] & w16979;
assign w16982 = ~w16980 & ~w16981;
assign w16983 = ~w16972 & w16982;
assign w16984 = w16972 & ~w16982;
assign w16985 = ~w16983 & ~w16984;
assign w16986 = ~w16971 & ~w16985;
assign w16987 = w16971 & w16985;
assign w16988 = ~w16986 & ~w16987;
assign w16989 = b[59] & w1154;
assign w16990 = b[58] & ~w1272;
assign w16991 = b[60] & w1156;
assign w16992 = w1150 & w11035;
assign w16993 = ~w16989 & ~w16990;
assign w16994 = ~w16991 & w16993;
assign w16995 = ~w16992 & w16994;
assign w16996 = a[20] & ~w16995;
assign w16997 = ~a[20] & w16995;
assign w16998 = ~w16996 & ~w16997;
assign w16999 = ~w16700 & ~w16703;
assign w17000 = w16998 & ~w16999;
assign w17001 = ~w16998 & w16999;
assign w17002 = ~w17000 & ~w17001;
assign w17003 = w16988 & w17002;
assign w17004 = ~w16988 & ~w17002;
assign w17005 = ~w17003 & ~w17004;
assign w17006 = (~w16715 & ~w16717) | (~w16715 & w25585) | (~w16717 & w25585);
assign w17007 = b[61] & ~w934;
assign w17008 = b[63] & w834;
assign w17009 = b[62] & w838;
assign w17010 = w832 & w12132;
assign w17011 = ~w17007 & ~w17008;
assign w17012 = ~w17009 & w17011;
assign w17013 = ~w17010 & w17012;
assign w17014 = a[17] & ~w17013;
assign w17015 = ~a[17] & w17013;
assign w17016 = ~w17014 & ~w17015;
assign w17017 = ~w17006 & w17016;
assign w17018 = w17006 & ~w17016;
assign w17019 = ~w17017 & ~w17018;
assign w17020 = ~w17005 & ~w17019;
assign w17021 = w17005 & w17019;
assign w17022 = ~w17020 & ~w17021;
assign w17023 = ~w16728 & ~w16731;
assign w17024 = ~w17022 & w17023;
assign w17025 = w17022 & ~w17023;
assign w17026 = ~w17024 & ~w17025;
assign w17027 = (~w16734 & w16450) | (~w16734 & w24423) | (w16450 & w24423);
assign w17028 = ~w17026 & w17027;
assign w17029 = (~w16450 & w24424) | (~w16450 & w24425) | (w24424 & w24425);
assign w17030 = ~w17028 & ~w17029;
assign w17031 = ~w17017 & ~w17021;
assign w17032 = b[61] & w1156;
assign w17033 = b[60] & w1154;
assign w17034 = b[59] & ~w1272;
assign w17035 = w1150 & w11400;
assign w17036 = ~w17032 & ~w17033;
assign w17037 = ~w17034 & w17036;
assign w17038 = ~w17035 & w17037;
assign w17039 = a[20] & ~w17038;
assign w17040 = ~a[20] & w17038;
assign w17041 = ~w17039 & ~w17040;
assign w17042 = ~w16983 & ~w16987;
assign w17043 = w17041 & ~w17042;
assign w17044 = ~w17041 & w17042;
assign w17045 = ~w17043 & ~w17044;
assign w17046 = b[44] & w3785;
assign w17047 = b[45] & w3578;
assign w17048 = b[46] & w3580;
assign w17049 = w3573 & ~w6613;
assign w17050 = ~w17047 & ~w17048;
assign w17051 = ~w17046 & w17050;
assign w17052 = ~w17049 & w17051;
assign w17053 = a[35] & ~w17052;
assign w17054 = ~a[35] & w17052;
assign w17055 = ~w17053 & ~w17054;
assign w17056 = ~w16906 & ~w16909;
assign w17057 = b[38] & w5167;
assign w17058 = b[39] & w4918;
assign w17059 = b[40] & w4925;
assign w17060 = w4923 & ~w5058;
assign w17061 = ~w17058 & ~w17059;
assign w17062 = ~w17057 & w17061;
assign w17063 = ~w17060 & w17062;
assign w17064 = a[41] & ~w17063;
assign w17065 = ~a[41] & w17063;
assign w17066 = ~w17064 & ~w17065;
assign w17067 = ~w16890 & ~w16894;
assign w17068 = b[35] & w5939;
assign w17069 = b[37] & w5665;
assign w17070 = b[36] & w5670;
assign w17071 = ~w4357 & w5663;
assign w17072 = ~w17069 & ~w17070;
assign w17073 = ~w17068 & w17072;
assign w17074 = ~w17071 & w17073;
assign w17075 = a[44] & ~w17074;
assign w17076 = ~a[44] & w17074;
assign w17077 = ~w17075 & ~w17076;
assign w17078 = ~w16884 & ~w16887;
assign w17079 = b[32] & w6732;
assign w17080 = b[34] & w6476;
assign w17081 = b[33] & w6474;
assign w17082 = ~w3710 & w6469;
assign w17083 = ~w17080 & ~w17081;
assign w17084 = ~w17079 & w17083;
assign w17085 = ~w17082 & w17084;
assign w17086 = a[47] & ~w17085;
assign w17087 = ~a[47] & w17085;
assign w17088 = ~w17086 & ~w17087;
assign w17089 = ~w16851 & ~w16855;
assign w17090 = b[26] & w8515;
assign w17091 = b[27] & w8200;
assign w17092 = b[28] & w8202;
assign w17093 = w2559 & w8195;
assign w17094 = ~w17091 & ~w17092;
assign w17095 = ~w17090 & w17094;
assign w17096 = ~w17093 & w17095;
assign w17097 = a[53] & ~w17096;
assign w17098 = ~a[53] & w17096;
assign w17099 = ~w17097 & ~w17098;
assign w17100 = b[23] & w9482;
assign w17101 = b[25] & w9160;
assign w17102 = b[24] & w9165;
assign w17103 = w2061 & w9158;
assign w17104 = ~w17101 & ~w17102;
assign w17105 = ~w17100 & w17104;
assign w17106 = ~w17103 & w17105;
assign w17107 = a[56] & ~w17106;
assign w17108 = ~a[56] & w17106;
assign w17109 = ~w17107 & ~w17108;
assign w17110 = ~w16812 & ~w16816;
assign w17111 = b[15] & w11921;
assign w17112 = b[16] & w11923;
assign w17113 = ~w17111 & ~w17112;
assign w17114 = ~w16806 & ~w16809;
assign w17115 = w17113 & ~w17114;
assign w17116 = ~w17113 & w17114;
assign w17117 = ~w17115 & ~w17116;
assign w17118 = b[17] & w11561;
assign w17119 = b[18] & w11194;
assign w17120 = b[19] & w11196;
assign w17121 = ~w1231 & w11189;
assign w17122 = ~w17119 & ~w17120;
assign w17123 = ~w17118 & w17122;
assign w17124 = ~w17121 & w17123;
assign w17125 = a[62] & ~w17124;
assign w17126 = ~a[62] & w17124;
assign w17127 = ~w17125 & ~w17126;
assign w17128 = w17117 & w17127;
assign w17129 = ~w17117 & ~w17127;
assign w17130 = ~w17128 & ~w17129;
assign w17131 = w17110 & ~w17130;
assign w17132 = ~w17110 & w17130;
assign w17133 = ~w17131 & ~w17132;
assign w17134 = b[20] & w10496;
assign w17135 = b[21] & w10146;
assign w17136 = b[22] & w10148;
assign w17137 = w1615 & w10141;
assign w17138 = ~w17135 & ~w17136;
assign w17139 = ~w17134 & w17138;
assign w17140 = ~w17137 & w17139;
assign w17141 = a[59] & ~w17140;
assign w17142 = ~a[59] & w17140;
assign w17143 = ~w17141 & ~w17142;
assign w17144 = w17133 & w17143;
assign w17145 = ~w17133 & ~w17143;
assign w17146 = ~w17144 & ~w17145;
assign w17147 = ~w16828 & ~w16833;
assign w17148 = w17146 & ~w17147;
assign w17149 = ~w17146 & w17147;
assign w17150 = ~w17148 & ~w17149;
assign w17151 = w17109 & w17150;
assign w17152 = ~w17109 & ~w17150;
assign w17153 = ~w17151 & ~w17152;
assign w17154 = ~w16845 & ~w16848;
assign w17155 = w17153 & w17154;
assign w17156 = ~w17153 & ~w17154;
assign w17157 = ~w17155 & ~w17156;
assign w17158 = w17099 & w17157;
assign w17159 = ~w17099 & ~w17157;
assign w17160 = ~w17158 & ~w17159;
assign w17161 = ~w17089 & w17160;
assign w17162 = w17089 & ~w17160;
assign w17163 = ~w17161 & ~w17162;
assign w17164 = b[29] & w7586;
assign w17165 = b[31] & w7314;
assign w17166 = b[30] & w7307;
assign w17167 = ~w3112 & w7312;
assign w17168 = ~w17165 & ~w17166;
assign w17169 = ~w17164 & w17168;
assign w17170 = ~w17167 & w17169;
assign w17171 = a[50] & ~w17170;
assign w17172 = ~a[50] & w17170;
assign w17173 = ~w17171 & ~w17172;
assign w17174 = w17163 & w17173;
assign w17175 = ~w17163 & ~w17173;
assign w17176 = ~w17174 & ~w17175;
assign w17177 = ~w16867 & ~w16872;
assign w17178 = w17176 & ~w17177;
assign w17179 = ~w17176 & w17177;
assign w17180 = ~w17178 & ~w17179;
assign w17181 = ~w17088 & ~w17180;
assign w17182 = w17088 & w17180;
assign w17183 = ~w17181 & ~w17182;
assign w17184 = w17078 & ~w17183;
assign w17185 = ~w17078 & w17183;
assign w17186 = ~w17184 & ~w17185;
assign w17187 = w17077 & w17186;
assign w17188 = ~w17077 & ~w17186;
assign w17189 = ~w17187 & ~w17188;
assign w17190 = w17067 & ~w17189;
assign w17191 = ~w17067 & w17189;
assign w17192 = ~w17190 & ~w17191;
assign w17193 = w17066 & w17192;
assign w17194 = ~w17066 & ~w17192;
assign w17195 = ~w17193 & ~w17194;
assign w17196 = w17056 & ~w17195;
assign w17197 = ~w17056 & w17195;
assign w17198 = ~w17196 & ~w17197;
assign w17199 = b[41] & w4453;
assign w17200 = b[42] & w4241;
assign w17201 = b[43] & w4243;
assign w17202 = w4236 & w5811;
assign w17203 = ~w17200 & ~w17201;
assign w17204 = ~w17199 & w17203;
assign w17205 = ~w17202 & w17204;
assign w17206 = a[38] & ~w17205;
assign w17207 = ~a[38] & w17205;
assign w17208 = ~w17206 & ~w17207;
assign w17209 = w17198 & w17208;
assign w17210 = ~w17198 & ~w17208;
assign w17211 = ~w17209 & ~w17210;
assign w17212 = ~w16912 & ~w16916;
assign w17213 = w17211 & ~w17212;
assign w17214 = ~w17211 & w17212;
assign w17215 = ~w17213 & ~w17214;
assign w17216 = w17055 & w17215;
assign w17217 = ~w17055 & ~w17215;
assign w17218 = ~w17216 & ~w17217;
assign w17219 = b[47] & w3177;
assign w17220 = b[49] & w2978;
assign w17221 = b[48] & w2973;
assign w17222 = w2980 & ~w7468;
assign w17223 = ~w17220 & ~w17221;
assign w17224 = ~w17219 & w17223;
assign w17225 = ~w17222 & w17224;
assign w17226 = a[32] & ~w17225;
assign w17227 = ~a[32] & w17225;
assign w17228 = ~w17226 & ~w17227;
assign w17229 = ~w16928 & ~w16933;
assign w17230 = w17228 & ~w17229;
assign w17231 = ~w17228 & w17229;
assign w17232 = ~w17230 & ~w17231;
assign w17233 = w17218 & w17232;
assign w17234 = ~w17218 & ~w17232;
assign w17235 = ~w17233 & ~w17234;
assign w17236 = b[51] & w2436;
assign w17237 = b[52] & w2438;
assign w17238 = b[50] & ~w2622;
assign w17239 = w2432 & ~w8371;
assign w17240 = ~w17236 & ~w17237;
assign w17241 = ~w17238 & w17240;
assign w17242 = ~w17239 & w17241;
assign w17243 = a[29] & ~w17242;
assign w17244 = ~a[29] & w17242;
assign w17245 = ~w17243 & ~w17244;
assign w17246 = ~w16946 & ~w16949;
assign w17247 = w17245 & ~w17246;
assign w17248 = ~w17245 & w17246;
assign w17249 = ~w17247 & ~w17248;
assign w17250 = ~w17235 & ~w17249;
assign w17251 = w17235 & w17249;
assign w17252 = ~w17250 & ~w17251;
assign w17253 = b[53] & ~w2114;
assign w17254 = b[55] & w1957;
assign w17255 = b[54] & w1955;
assign w17256 = w1951 & ~w9330;
assign w17257 = ~w17253 & ~w17254;
assign w17258 = ~w17255 & w17257;
assign w17259 = ~w17256 & w17258;
assign w17260 = a[26] & ~w17259;
assign w17261 = ~a[26] & w17259;
assign w17262 = ~w17260 & ~w17261;
assign w17263 = ~w16963 & ~w16966;
assign w17264 = w17262 & ~w17263;
assign w17265 = ~w17262 & w17263;
assign w17266 = ~w17264 & ~w17265;
assign w17267 = w17252 & w17266;
assign w17268 = ~w17252 & ~w17266;
assign w17269 = ~w17267 & ~w17268;
assign w17270 = ~w16753 & ~w16969;
assign w17271 = b[58] & w1519;
assign w17272 = b[56] & ~w1676;
assign w17273 = b[57] & w1517;
assign w17274 = ~w17271 & ~w17272;
assign w17275 = ~w17273 & w17274;
assign w17276 = a[23] & w25734;
assign w17277 = (w10339 & w25462) | (w10339 & w25463) | (w25462 & w25463);
assign w17278 = ~w17276 & ~w17277;
assign w17279 = ~w17270 & w17278;
assign w17280 = w17270 & ~w17278;
assign w17281 = ~w17279 & ~w17280;
assign w17282 = w17269 & w17281;
assign w17283 = ~w17269 & ~w17281;
assign w17284 = ~w17282 & ~w17283;
assign w17285 = w17045 & w17284;
assign w17286 = ~w17045 & ~w17284;
assign w17287 = ~w17285 & ~w17286;
assign w17288 = ~w17000 & ~w17003;
assign w17289 = b[62] & ~w934;
assign w17290 = b[63] & w838;
assign w17291 = w832 & w12156;
assign w17292 = ~w17289 & ~w17290;
assign w17293 = ~w17291 & w17292;
assign w17294 = a[17] & ~w17293;
assign w17295 = ~a[17] & w17293;
assign w17296 = ~w17294 & ~w17295;
assign w17297 = ~w17288 & w17296;
assign w17298 = w17288 & ~w17296;
assign w17299 = ~w17297 & ~w17298;
assign w17300 = w17287 & w17299;
assign w17301 = ~w17287 & ~w17299;
assign w17302 = ~w17300 & ~w17301;
assign w17303 = w17031 & ~w17302;
assign w17304 = ~w17031 & w17302;
assign w17305 = ~w17303 & ~w17304;
assign w17306 = (w16450 & w24426) | (w16450 & w24427) | (w24426 & w24427);
assign w17307 = w17305 & ~w17306;
assign w17308 = ~w17305 & w17306;
assign w17309 = ~w17307 & ~w17308;
assign w17310 = ~w17297 & ~w17300;
assign w17311 = ~w17197 & ~w17209;
assign w17312 = b[42] & w4453;
assign w17313 = b[44] & w4243;
assign w17314 = b[43] & w4241;
assign w17315 = w4236 & w6069;
assign w17316 = ~w17313 & ~w17314;
assign w17317 = ~w17312 & w17316;
assign w17318 = ~w17315 & w17317;
assign w17319 = a[38] & ~w17318;
assign w17320 = ~a[38] & w17318;
assign w17321 = ~w17319 & ~w17320;
assign w17322 = ~w17191 & ~w17193;
assign w17323 = b[39] & w5167;
assign w17324 = b[41] & w4925;
assign w17325 = b[40] & w4918;
assign w17326 = w4923 & w5302;
assign w17327 = ~w17324 & ~w17325;
assign w17328 = ~w17323 & w17327;
assign w17329 = ~w17326 & w17328;
assign w17330 = a[41] & ~w17329;
assign w17331 = ~a[41] & w17329;
assign w17332 = ~w17330 & ~w17331;
assign w17333 = ~w17185 & ~w17187;
assign w17334 = b[36] & w5939;
assign w17335 = b[38] & w5665;
assign w17336 = b[37] & w5670;
assign w17337 = w4582 & w5663;
assign w17338 = ~w17335 & ~w17336;
assign w17339 = ~w17334 & w17338;
assign w17340 = ~w17337 & w17339;
assign w17341 = a[44] & ~w17340;
assign w17342 = ~a[44] & w17340;
assign w17343 = ~w17341 & ~w17342;
assign w17344 = b[33] & w6732;
assign w17345 = b[34] & w6474;
assign w17346 = b[35] & w6476;
assign w17347 = w3918 & w6469;
assign w17348 = ~w17345 & ~w17346;
assign w17349 = ~w17344 & w17348;
assign w17350 = ~w17347 & w17349;
assign w17351 = a[47] & ~w17350;
assign w17352 = ~a[47] & w17350;
assign w17353 = ~w17351 & ~w17352;
assign w17354 = ~w17161 & ~w17174;
assign w17355 = b[30] & w7586;
assign w17356 = b[32] & w7314;
assign w17357 = b[31] & w7307;
assign w17358 = w3304 & w7312;
assign w17359 = ~w17356 & ~w17357;
assign w17360 = ~w17355 & w17359;
assign w17361 = ~w17358 & w17360;
assign w17362 = a[50] & ~w17361;
assign w17363 = ~a[50] & w17361;
assign w17364 = ~w17362 & ~w17363;
assign w17365 = ~w17148 & ~w17151;
assign w17366 = b[24] & w9482;
assign w17367 = b[25] & w9165;
assign w17368 = b[26] & w9160;
assign w17369 = w2219 & w9158;
assign w17370 = ~w17367 & ~w17368;
assign w17371 = ~w17366 & w17370;
assign w17372 = ~w17369 & w17371;
assign w17373 = a[56] & ~w17372;
assign w17374 = ~a[56] & w17372;
assign w17375 = ~w17373 & ~w17374;
assign w17376 = ~w17132 & ~w17144;
assign w17377 = b[21] & w10496;
assign w17378 = b[23] & w10148;
assign w17379 = b[22] & w10146;
assign w17380 = w1755 & w10141;
assign w17381 = ~w17378 & ~w17379;
assign w17382 = ~w17377 & w17381;
assign w17383 = ~w17380 & w17382;
assign w17384 = a[59] & ~w17383;
assign w17385 = ~a[59] & w17383;
assign w17386 = ~w17384 & ~w17385;
assign w17387 = ~w17115 & ~w17128;
assign w17388 = b[18] & w11561;
assign w17389 = b[19] & w11194;
assign w17390 = b[20] & w11196;
assign w17391 = w1347 & w11189;
assign w17392 = ~w17389 & ~w17390;
assign w17393 = ~w17388 & w17392;
assign w17394 = ~w17391 & w17393;
assign w17395 = a[62] & ~w17394;
assign w17396 = ~a[62] & w17394;
assign w17397 = ~w17395 & ~w17396;
assign w17398 = b[16] & w11921;
assign w17399 = b[17] & w11923;
assign w17400 = ~w17398 & ~w17399;
assign w17401 = w17113 & ~w17400;
assign w17402 = ~w17113 & w17400;
assign w17403 = ~w17401 & ~w17402;
assign w17404 = w17397 & ~w17403;
assign w17405 = ~w17397 & w17403;
assign w17406 = ~w17404 & ~w17405;
assign w17407 = ~w17387 & ~w17406;
assign w17408 = w17387 & w17406;
assign w17409 = ~w17407 & ~w17408;
assign w17410 = ~w17386 & ~w17409;
assign w17411 = w17386 & w17409;
assign w17412 = ~w17410 & ~w17411;
assign w17413 = w17376 & ~w17412;
assign w17414 = ~w17376 & w17412;
assign w17415 = ~w17413 & ~w17414;
assign w17416 = w17375 & w17415;
assign w17417 = ~w17375 & ~w17415;
assign w17418 = ~w17416 & ~w17417;
assign w17419 = w17365 & ~w17418;
assign w17420 = ~w17365 & w17418;
assign w17421 = ~w17419 & ~w17420;
assign w17422 = b[27] & w8515;
assign w17423 = b[29] & w8202;
assign w17424 = b[28] & w8200;
assign w17425 = w2734 & w8195;
assign w17426 = ~w17423 & ~w17424;
assign w17427 = ~w17422 & w17426;
assign w17428 = ~w17425 & w17427;
assign w17429 = a[53] & ~w17428;
assign w17430 = ~a[53] & w17428;
assign w17431 = ~w17429 & ~w17430;
assign w17432 = w17421 & w17431;
assign w17433 = ~w17421 & ~w17431;
assign w17434 = ~w17432 & ~w17433;
assign w17435 = ~w17155 & ~w17158;
assign w17436 = w17434 & ~w17435;
assign w17437 = ~w17434 & w17435;
assign w17438 = ~w17436 & ~w17437;
assign w17439 = w17364 & w17438;
assign w17440 = ~w17364 & ~w17438;
assign w17441 = ~w17439 & ~w17440;
assign w17442 = ~w17354 & w17441;
assign w17443 = w17354 & ~w17441;
assign w17444 = ~w17442 & ~w17443;
assign w17445 = w17353 & w17444;
assign w17446 = ~w17353 & ~w17444;
assign w17447 = ~w17445 & ~w17446;
assign w17448 = ~w17178 & ~w17182;
assign w17449 = w17447 & ~w17448;
assign w17450 = ~w17447 & w17448;
assign w17451 = ~w17449 & ~w17450;
assign w17452 = w17343 & w17451;
assign w17453 = ~w17343 & ~w17451;
assign w17454 = ~w17452 & ~w17453;
assign w17455 = ~w17333 & w17454;
assign w17456 = w17333 & ~w17454;
assign w17457 = ~w17455 & ~w17456;
assign w17458 = w17332 & w17457;
assign w17459 = ~w17332 & ~w17457;
assign w17460 = ~w17458 & ~w17459;
assign w17461 = w17322 & ~w17460;
assign w17462 = ~w17322 & w17460;
assign w17463 = ~w17461 & ~w17462;
assign w17464 = w17321 & w17463;
assign w17465 = ~w17321 & ~w17463;
assign w17466 = ~w17464 & ~w17465;
assign w17467 = w17311 & ~w17466;
assign w17468 = ~w17311 & w17466;
assign w17469 = ~w17467 & ~w17468;
assign w17470 = b[45] & w3785;
assign w17471 = b[46] & w3578;
assign w17472 = b[47] & w3580;
assign w17473 = w3573 & w6889;
assign w17474 = ~w17471 & ~w17472;
assign w17475 = ~w17470 & w17474;
assign w17476 = ~w17473 & w17475;
assign w17477 = a[35] & ~w17476;
assign w17478 = ~a[35] & w17476;
assign w17479 = ~w17477 & ~w17478;
assign w17480 = w17469 & w17479;
assign w17481 = ~w17469 & ~w17479;
assign w17482 = ~w17480 & ~w17481;
assign w17483 = b[48] & w3177;
assign w17484 = b[50] & w2978;
assign w17485 = b[49] & w2973;
assign w17486 = w2980 & w7759;
assign w17487 = ~w17484 & ~w17485;
assign w17488 = ~w17483 & w17487;
assign w17489 = ~w17486 & w17488;
assign w17490 = a[32] & ~w17489;
assign w17491 = ~a[32] & w17489;
assign w17492 = ~w17490 & ~w17491;
assign w17493 = ~w17213 & ~w17216;
assign w17494 = w17492 & ~w17493;
assign w17495 = ~w17492 & w17493;
assign w17496 = ~w17494 & ~w17495;
assign w17497 = w17482 & w17496;
assign w17498 = ~w17482 & ~w17496;
assign w17499 = ~w17497 & ~w17498;
assign w17500 = b[52] & w2436;
assign w17501 = b[51] & ~w2622;
assign w17502 = b[53] & w2438;
assign w17503 = ~w17500 & ~w17501;
assign w17504 = ~w17502 & w17503;
assign w17505 = (w17504 & ~w8683) | (w17504 & w25464) | (~w8683 & w25464);
assign w17506 = a[29] & ~w17505;
assign w17507 = ~a[29] & w17505;
assign w17508 = ~w17506 & ~w17507;
assign w17509 = ~w17230 & ~w17233;
assign w17510 = w17508 & ~w17509;
assign w17511 = ~w17508 & w17509;
assign w17512 = ~w17510 & ~w17511;
assign w17513 = ~w17499 & ~w17512;
assign w17514 = w17499 & w17512;
assign w17515 = ~w17513 & ~w17514;
assign w17516 = b[54] & ~w2114;
assign w17517 = b[56] & w1957;
assign w17518 = b[55] & w1955;
assign w17519 = ~w17516 & ~w17517;
assign w17520 = ~w17518 & w17519;
assign w17521 = (w9657 & w25319) | (w9657 & w25320) | (w25319 & w25320);
assign w17522 = ~a[26] & w25735;
assign w17523 = ~w17521 & ~w17522;
assign w17524 = ~w17247 & ~w17251;
assign w17525 = w17523 & ~w17524;
assign w17526 = ~w17523 & w17524;
assign w17527 = ~w17525 & ~w17526;
assign w17528 = w17515 & w17527;
assign w17529 = ~w17515 & ~w17527;
assign w17530 = ~w17528 & ~w17529;
assign w17531 = b[58] & w1517;
assign w17532 = b[59] & w1519;
assign w17533 = b[57] & ~w1676;
assign w17534 = ~w17531 & ~w17532;
assign w17535 = ~w17533 & w17534;
assign w17536 = (w10371 & w24868) | (w10371 & w24869) | (w24868 & w24869);
assign w17537 = (~w10371 & w24870) | (~w10371 & w24871) | (w24870 & w24871);
assign w17538 = ~w17536 & ~w17537;
assign w17539 = ~w17264 & ~w17267;
assign w17540 = w17538 & ~w17539;
assign w17541 = ~w17538 & w17539;
assign w17542 = ~w17540 & ~w17541;
assign w17543 = ~w17530 & ~w17542;
assign w17544 = w17530 & w17542;
assign w17545 = ~w17543 & ~w17544;
assign w17546 = b[62] & w1156;
assign w17547 = b[61] & w1154;
assign w17548 = b[60] & ~w1272;
assign w17549 = ~w17546 & ~w17547;
assign w17550 = ~w17548 & w17549;
assign w17551 = (w11763 & w24872) | (w11763 & w24873) | (w24872 & w24873);
assign w17552 = ~a[20] & w25736;
assign w17553 = ~w17551 & ~w17552;
assign w17554 = ~w17279 & ~w17282;
assign w17555 = w17553 & ~w17554;
assign w17556 = ~w17553 & w17554;
assign w17557 = ~w17555 & ~w17556;
assign w17558 = ~w17545 & ~w17557;
assign w17559 = w17545 & w17557;
assign w17560 = ~w17558 & ~w17559;
assign w17561 = ~w17043 & ~w17285;
assign w17562 = w832 & ~w12154;
assign w17563 = w934 & ~w17562;
assign w17564 = b[63] & ~w17563;
assign w17565 = ~a[17] & ~w17564;
assign w17566 = a[17] & w17564;
assign w17567 = ~w17565 & ~w17566;
assign w17568 = ~w17561 & w17567;
assign w17569 = w17561 & ~w17567;
assign w17570 = ~w17568 & ~w17569;
assign w17571 = w17560 & w17570;
assign w17572 = ~w17560 & ~w17570;
assign w17573 = ~w17571 & ~w17572;
assign w17574 = w17310 & ~w17573;
assign w17575 = ~w17310 & w17573;
assign w17576 = ~w17574 & ~w17575;
assign w17577 = (w16450 & w24430) | (w16450 & w24431) | (w24430 & w24431);
assign w17578 = w17576 & ~w17577;
assign w17579 = ~w17576 & w17577;
assign w17580 = ~w17578 & ~w17579;
assign w17581 = (w16450 & w24434) | (w16450 & w24435) | (w24434 & w24435);
assign w17582 = ~w17568 & ~w17571;
assign w17583 = b[54] & w2438;
assign w17584 = b[53] & w2436;
assign w17585 = b[52] & ~w2622;
assign w17586 = w2432 & ~w8998;
assign w17587 = ~w17583 & ~w17584;
assign w17588 = ~w17585 & w17587;
assign w17589 = ~w17586 & w17588;
assign w17590 = a[29] & ~w17589;
assign w17591 = ~a[29] & w17589;
assign w17592 = ~w17590 & ~w17591;
assign w17593 = ~w17510 & ~w17514;
assign w17594 = w17592 & ~w17593;
assign w17595 = ~w17592 & w17593;
assign w17596 = ~w17594 & ~w17595;
assign w17597 = ~w17455 & ~w17458;
assign w17598 = b[40] & w5167;
assign w17599 = b[41] & w4918;
assign w17600 = b[42] & w4925;
assign w17601 = w4923 & w5548;
assign w17602 = ~w17599 & ~w17600;
assign w17603 = ~w17598 & w17602;
assign w17604 = ~w17601 & w17603;
assign w17605 = a[41] & ~w17604;
assign w17606 = ~a[41] & w17604;
assign w17607 = ~w17605 & ~w17606;
assign w17608 = ~w17449 & ~w17452;
assign w17609 = ~w17442 & ~w17445;
assign w17610 = b[34] & w6732;
assign w17611 = b[36] & w6476;
assign w17612 = b[35] & w6474;
assign w17613 = w4129 & w6469;
assign w17614 = ~w17611 & ~w17612;
assign w17615 = ~w17610 & w17614;
assign w17616 = ~w17613 & w17615;
assign w17617 = a[47] & ~w17616;
assign w17618 = ~a[47] & w17616;
assign w17619 = ~w17617 & ~w17618;
assign w17620 = ~w17407 & ~w17411;
assign w17621 = b[22] & w10496;
assign w17622 = b[24] & w10148;
assign w17623 = b[23] & w10146;
assign w17624 = w1895 & w10141;
assign w17625 = ~w17622 & ~w17623;
assign w17626 = ~w17621 & w17625;
assign w17627 = ~w17624 & w17626;
assign w17628 = a[59] & ~w17627;
assign w17629 = ~a[59] & w17627;
assign w17630 = ~w17628 & ~w17629;
assign w17631 = b[19] & w11561;
assign w17632 = b[20] & w11194;
assign w17633 = b[21] & w11196;
assign w17634 = w1467 & w11189;
assign w17635 = ~w17632 & ~w17633;
assign w17636 = ~w17631 & w17635;
assign w17637 = ~w17634 & w17636;
assign w17638 = a[62] & ~w17637;
assign w17639 = ~a[62] & w17637;
assign w17640 = ~w17638 & ~w17639;
assign w17641 = b[17] & w11921;
assign w17642 = b[18] & w11923;
assign w17643 = ~w17641 & ~w17642;
assign w17644 = ~a[17] & ~w17643;
assign w17645 = a[17] & w17643;
assign w17646 = ~w17644 & ~w17645;
assign w17647 = ~w17400 & w17646;
assign w17648 = w17400 & ~w17646;
assign w17649 = ~w17647 & ~w17648;
assign w17650 = ~w17640 & ~w17649;
assign w17651 = w17640 & w17649;
assign w17652 = ~w17650 & ~w17651;
assign w17653 = ~w17401 & ~w17405;
assign w17654 = w17652 & w17653;
assign w17655 = ~w17652 & ~w17653;
assign w17656 = ~w17654 & ~w17655;
assign w17657 = w17630 & w17656;
assign w17658 = ~w17630 & ~w17656;
assign w17659 = ~w17657 & ~w17658;
assign w17660 = ~w17620 & w17659;
assign w17661 = w17620 & ~w17659;
assign w17662 = ~w17660 & ~w17661;
assign w17663 = b[25] & w9482;
assign w17664 = b[26] & w9165;
assign w17665 = b[27] & w9160;
assign w17666 = w2378 & w9158;
assign w17667 = ~w17664 & ~w17665;
assign w17668 = ~w17663 & w17667;
assign w17669 = ~w17666 & w17668;
assign w17670 = a[56] & ~w17669;
assign w17671 = ~a[56] & w17669;
assign w17672 = ~w17670 & ~w17671;
assign w17673 = w17662 & w17672;
assign w17674 = ~w17662 & ~w17672;
assign w17675 = ~w17673 & ~w17674;
assign w17676 = ~w17414 & ~w17416;
assign w17677 = ~w17675 & w17676;
assign w17678 = w17675 & ~w17676;
assign w17679 = ~w17677 & ~w17678;
assign w17680 = b[28] & w8515;
assign w17681 = b[29] & w8200;
assign w17682 = b[30] & w8202;
assign w17683 = ~w2908 & w8195;
assign w17684 = ~w17681 & ~w17682;
assign w17685 = ~w17680 & w17684;
assign w17686 = ~w17683 & w17685;
assign w17687 = a[53] & ~w17686;
assign w17688 = ~a[53] & w17686;
assign w17689 = ~w17687 & ~w17688;
assign w17690 = w17679 & w17689;
assign w17691 = ~w17679 & ~w17689;
assign w17692 = ~w17690 & ~w17691;
assign w17693 = ~w17420 & ~w17432;
assign w17694 = ~w17692 & w17693;
assign w17695 = w17692 & ~w17693;
assign w17696 = ~w17694 & ~w17695;
assign w17697 = b[31] & w7586;
assign w17698 = b[32] & w7307;
assign w17699 = b[33] & w7314;
assign w17700 = w3499 & w7312;
assign w17701 = ~w17698 & ~w17699;
assign w17702 = ~w17697 & w17701;
assign w17703 = ~w17700 & w17702;
assign w17704 = a[50] & ~w17703;
assign w17705 = ~a[50] & w17703;
assign w17706 = ~w17704 & ~w17705;
assign w17707 = ~w17436 & ~w17439;
assign w17708 = w17706 & ~w17707;
assign w17709 = ~w17706 & w17707;
assign w17710 = ~w17708 & ~w17709;
assign w17711 = w17696 & w17710;
assign w17712 = ~w17696 & ~w17710;
assign w17713 = ~w17711 & ~w17712;
assign w17714 = w17619 & w17713;
assign w17715 = ~w17619 & ~w17713;
assign w17716 = ~w17714 & ~w17715;
assign w17717 = w17609 & ~w17716;
assign w17718 = ~w17609 & w17716;
assign w17719 = ~w17717 & ~w17718;
assign w17720 = b[37] & w5939;
assign w17721 = b[39] & w5665;
assign w17722 = b[38] & w5670;
assign w17723 = ~w4812 & w5663;
assign w17724 = ~w17721 & ~w17722;
assign w17725 = ~w17720 & w17724;
assign w17726 = ~w17723 & w17725;
assign w17727 = a[44] & ~w17726;
assign w17728 = ~a[44] & w17726;
assign w17729 = ~w17727 & ~w17728;
assign w17730 = w17719 & w17729;
assign w17731 = ~w17719 & ~w17729;
assign w17732 = ~w17730 & ~w17731;
assign w17733 = ~w17608 & w17732;
assign w17734 = w17608 & ~w17732;
assign w17735 = ~w17733 & ~w17734;
assign w17736 = w17607 & w17735;
assign w17737 = ~w17607 & ~w17735;
assign w17738 = ~w17736 & ~w17737;
assign w17739 = w17597 & ~w17738;
assign w17740 = ~w17597 & w17738;
assign w17741 = ~w17739 & ~w17740;
assign w17742 = b[43] & w4453;
assign w17743 = b[45] & w4243;
assign w17744 = b[44] & w4241;
assign w17745 = w4236 & w6334;
assign w17746 = ~w17743 & ~w17744;
assign w17747 = ~w17742 & w17746;
assign w17748 = ~w17745 & w17747;
assign w17749 = a[38] & ~w17748;
assign w17750 = ~a[38] & w17748;
assign w17751 = ~w17749 & ~w17750;
assign w17752 = w17741 & w17751;
assign w17753 = ~w17741 & ~w17751;
assign w17754 = ~w17752 & ~w17753;
assign w17755 = ~w17462 & ~w17464;
assign w17756 = ~w17754 & w17755;
assign w17757 = w17754 & ~w17755;
assign w17758 = ~w17756 & ~w17757;
assign w17759 = b[46] & w3785;
assign w17760 = b[47] & w3578;
assign w17761 = b[48] & w3580;
assign w17762 = w3573 & ~w7170;
assign w17763 = ~w17760 & ~w17761;
assign w17764 = ~w17759 & w17763;
assign w17765 = ~w17762 & w17764;
assign w17766 = a[35] & ~w17765;
assign w17767 = ~a[35] & w17765;
assign w17768 = ~w17766 & ~w17767;
assign w17769 = w17758 & w17768;
assign w17770 = ~w17758 & ~w17768;
assign w17771 = ~w17769 & ~w17770;
assign w17772 = ~w17468 & ~w17480;
assign w17773 = ~w17771 & w17772;
assign w17774 = w17771 & ~w17772;
assign w17775 = ~w17773 & ~w17774;
assign w17776 = ~w17494 & ~w17497;
assign w17777 = b[49] & w3177;
assign w17778 = b[51] & w2978;
assign w17779 = b[50] & w2973;
assign w17780 = w2980 & ~w8058;
assign w17781 = ~w17778 & ~w17779;
assign w17782 = ~w17777 & w17781;
assign w17783 = ~w17780 & w17782;
assign w17784 = a[32] & ~w17783;
assign w17785 = ~a[32] & w17783;
assign w17786 = ~w17784 & ~w17785;
assign w17787 = ~w17776 & w17786;
assign w17788 = w17776 & ~w17786;
assign w17789 = ~w17787 & ~w17788;
assign w17790 = w17775 & w17789;
assign w17791 = ~w17775 & ~w17789;
assign w17792 = ~w17790 & ~w17791;
assign w17793 = w17596 & w17792;
assign w17794 = ~w17596 & ~w17792;
assign w17795 = ~w17793 & ~w17794;
assign w17796 = b[55] & ~w2114;
assign w17797 = b[56] & w1955;
assign w17798 = b[57] & w1957;
assign w17799 = w1951 & ~w9992;
assign w17800 = ~w17796 & ~w17797;
assign w17801 = ~w17798 & w17800;
assign w17802 = ~w17799 & w17801;
assign w17803 = a[26] & ~w17802;
assign w17804 = ~a[26] & w17802;
assign w17805 = ~w17803 & ~w17804;
assign w17806 = ~w17525 & ~w17528;
assign w17807 = w17805 & ~w17806;
assign w17808 = ~w17805 & w17806;
assign w17809 = ~w17807 & ~w17808;
assign w17810 = ~w17795 & ~w17809;
assign w17811 = w17795 & w17809;
assign w17812 = ~w17810 & ~w17811;
assign w17813 = b[59] & w1517;
assign w17814 = b[58] & ~w1676;
assign w17815 = b[60] & w1519;
assign w17816 = ~w17813 & ~w17814;
assign w17817 = ~w17815 & w17816;
assign w17818 = (w11035 & w25209) | (w11035 & w25210) | (w25209 & w25210);
assign w17819 = ~a[23] & w25737;
assign w17820 = ~w17818 & ~w17819;
assign w17821 = (~w17540 & ~w17542) | (~w17540 & w25023) | (~w17542 & w25023);
assign w17822 = w17820 & ~w17821;
assign w17823 = ~w17820 & w17821;
assign w17824 = ~w17822 & ~w17823;
assign w17825 = w17812 & w17824;
assign w17826 = ~w17812 & ~w17824;
assign w17827 = ~w17825 & ~w17826;
assign w17828 = (~w17555 & ~w17557) | (~w17555 & w25024) | (~w17557 & w25024);
assign w17829 = b[63] & w1156;
assign w17830 = b[62] & w1154;
assign w17831 = b[61] & ~w1272;
assign w17832 = ~w17829 & ~w17830;
assign w17833 = ~w17831 & w17832;
assign w17834 = (w17833 & ~w12132) | (w17833 & w25465) | (~w12132 & w25465);
assign w17835 = a[20] & ~w17834;
assign w17836 = ~a[20] & w17834;
assign w17837 = ~w17835 & ~w17836;
assign w17838 = ~w17828 & w17837;
assign w17839 = w17828 & ~w17837;
assign w17840 = ~w17838 & ~w17839;
assign w17841 = w17827 & w17840;
assign w17842 = ~w17827 & ~w17840;
assign w17843 = ~w17841 & ~w17842;
assign w17844 = ~w17582 & w17843;
assign w17845 = w17582 & ~w17843;
assign w17846 = ~w17844 & ~w17845;
assign w17847 = w17581 & ~w17846;
assign w17848 = ~w17581 & w17846;
assign w17849 = ~w17847 & ~w17848;
assign w17850 = (~w17838 & ~w17840) | (~w17838 & w25466) | (~w17840 & w25466);
assign w17851 = b[56] & ~w2114;
assign w17852 = b[58] & w1957;
assign w17853 = b[57] & w1955;
assign w17854 = ~w17851 & ~w17852;
assign w17855 = ~w17853 & w17854;
assign w17856 = a[26] & w25738;
assign w17857 = (w10339 & w25467) | (w10339 & w25468) | (w25467 & w25468);
assign w17858 = ~w17856 & ~w17857;
assign w17859 = ~w17594 & ~w17793;
assign w17860 = w17858 & ~w17859;
assign w17861 = ~w17858 & w17859;
assign w17862 = ~w17860 & ~w17861;
assign w17863 = b[47] & w3785;
assign w17864 = b[49] & w3580;
assign w17865 = b[48] & w3578;
assign w17866 = w3573 & ~w7468;
assign w17867 = ~w17864 & ~w17865;
assign w17868 = ~w17863 & w17867;
assign w17869 = ~w17866 & w17868;
assign w17870 = a[35] & ~w17869;
assign w17871 = ~a[35] & w17869;
assign w17872 = ~w17870 & ~w17871;
assign w17873 = b[44] & w4453;
assign w17874 = b[46] & w4243;
assign w17875 = b[45] & w4241;
assign w17876 = w4236 & ~w6613;
assign w17877 = ~w17874 & ~w17875;
assign w17878 = ~w17873 & w17877;
assign w17879 = ~w17876 & w17878;
assign w17880 = a[38] & ~w17879;
assign w17881 = ~a[38] & w17879;
assign w17882 = ~w17880 & ~w17881;
assign w17883 = ~w17730 & ~w17733;
assign w17884 = b[38] & w5939;
assign w17885 = b[40] & w5665;
assign w17886 = b[39] & w5670;
assign w17887 = ~w5058 & w5663;
assign w17888 = ~w17885 & ~w17886;
assign w17889 = ~w17884 & w17888;
assign w17890 = ~w17887 & w17889;
assign w17891 = a[44] & ~w17890;
assign w17892 = ~a[44] & w17890;
assign w17893 = ~w17891 & ~w17892;
assign w17894 = ~w17714 & ~w17718;
assign w17895 = b[35] & w6732;
assign w17896 = b[37] & w6476;
assign w17897 = b[36] & w6474;
assign w17898 = ~w4357 & w6469;
assign w17899 = ~w17896 & ~w17897;
assign w17900 = ~w17895 & w17899;
assign w17901 = ~w17898 & w17900;
assign w17902 = a[47] & ~w17901;
assign w17903 = ~a[47] & w17901;
assign w17904 = ~w17902 & ~w17903;
assign w17905 = b[32] & w7586;
assign w17906 = b[34] & w7314;
assign w17907 = b[33] & w7307;
assign w17908 = ~w3710 & w7312;
assign w17909 = ~w17906 & ~w17907;
assign w17910 = ~w17905 & w17909;
assign w17911 = ~w17908 & w17910;
assign w17912 = a[50] & ~w17911;
assign w17913 = ~a[50] & w17911;
assign w17914 = ~w17912 & ~w17913;
assign w17915 = ~w17673 & ~w17678;
assign w17916 = b[26] & w9482;
assign w17917 = b[28] & w9160;
assign w17918 = b[27] & w9165;
assign w17919 = w2559 & w9158;
assign w17920 = ~w17917 & ~w17918;
assign w17921 = ~w17916 & w17920;
assign w17922 = ~w17919 & w17921;
assign w17923 = a[56] & ~w17922;
assign w17924 = ~a[56] & w17922;
assign w17925 = ~w17923 & ~w17924;
assign w17926 = ~w17657 & ~w17660;
assign w17927 = b[18] & w11921;
assign w17928 = b[19] & w11923;
assign w17929 = ~w17927 & ~w17928;
assign w17930 = ~w17644 & ~w17647;
assign w17931 = w17929 & ~w17930;
assign w17932 = ~w17929 & w17930;
assign w17933 = ~w17931 & ~w17932;
assign w17934 = b[20] & w11561;
assign w17935 = b[21] & w11194;
assign w17936 = b[22] & w11196;
assign w17937 = w1615 & w11189;
assign w17938 = ~w17935 & ~w17936;
assign w17939 = ~w17934 & w17938;
assign w17940 = ~w17937 & w17939;
assign w17941 = a[62] & ~w17940;
assign w17942 = ~a[62] & w17940;
assign w17943 = ~w17941 & ~w17942;
assign w17944 = ~w17933 & ~w17943;
assign w17945 = w17933 & w17943;
assign w17946 = ~w17944 & ~w17945;
assign w17947 = ~w17651 & ~w17654;
assign w17948 = w17946 & ~w17947;
assign w17949 = ~w17946 & w17947;
assign w17950 = ~w17948 & ~w17949;
assign w17951 = b[23] & w10496;
assign w17952 = b[24] & w10146;
assign w17953 = b[25] & w10148;
assign w17954 = w2061 & w10141;
assign w17955 = ~w17952 & ~w17953;
assign w17956 = ~w17951 & w17955;
assign w17957 = ~w17954 & w17956;
assign w17958 = a[59] & ~w17957;
assign w17959 = ~a[59] & w17957;
assign w17960 = ~w17958 & ~w17959;
assign w17961 = w17950 & w17960;
assign w17962 = ~w17950 & ~w17960;
assign w17963 = ~w17961 & ~w17962;
assign w17964 = ~w17926 & w17963;
assign w17965 = w17926 & ~w17963;
assign w17966 = ~w17964 & ~w17965;
assign w17967 = w17925 & w17966;
assign w17968 = ~w17925 & ~w17966;
assign w17969 = ~w17967 & ~w17968;
assign w17970 = ~w17915 & w17969;
assign w17971 = w17915 & ~w17969;
assign w17972 = ~w17970 & ~w17971;
assign w17973 = b[29] & w8515;
assign w17974 = b[30] & w8200;
assign w17975 = b[31] & w8202;
assign w17976 = ~w3112 & w8195;
assign w17977 = ~w17974 & ~w17975;
assign w17978 = ~w17973 & w17977;
assign w17979 = ~w17976 & w17978;
assign w17980 = a[53] & ~w17979;
assign w17981 = ~a[53] & w17979;
assign w17982 = ~w17980 & ~w17981;
assign w17983 = w17972 & w17982;
assign w17984 = ~w17972 & ~w17982;
assign w17985 = ~w17983 & ~w17984;
assign w17986 = ~w17690 & ~w17695;
assign w17987 = w17985 & ~w17986;
assign w17988 = ~w17985 & w17986;
assign w17989 = ~w17987 & ~w17988;
assign w17990 = w17914 & w17989;
assign w17991 = ~w17914 & ~w17989;
assign w17992 = ~w17990 & ~w17991;
assign w17993 = ~w17708 & ~w17711;
assign w17994 = w17992 & ~w17993;
assign w17995 = ~w17992 & w17993;
assign w17996 = ~w17994 & ~w17995;
assign w17997 = ~w17904 & ~w17996;
assign w17998 = w17904 & w17996;
assign w17999 = ~w17997 & ~w17998;
assign w18000 = w17894 & ~w17999;
assign w18001 = ~w17894 & w17999;
assign w18002 = ~w18000 & ~w18001;
assign w18003 = w17893 & w18002;
assign w18004 = ~w17893 & ~w18002;
assign w18005 = ~w18003 & ~w18004;
assign w18006 = w17883 & ~w18005;
assign w18007 = ~w17883 & w18005;
assign w18008 = ~w18006 & ~w18007;
assign w18009 = b[41] & w5167;
assign w18010 = b[42] & w4918;
assign w18011 = b[43] & w4925;
assign w18012 = w4923 & w5811;
assign w18013 = ~w18010 & ~w18011;
assign w18014 = ~w18009 & w18013;
assign w18015 = ~w18012 & w18014;
assign w18016 = a[41] & ~w18015;
assign w18017 = ~a[41] & w18015;
assign w18018 = ~w18016 & ~w18017;
assign w18019 = w18008 & w18018;
assign w18020 = ~w18008 & ~w18018;
assign w18021 = ~w18019 & ~w18020;
assign w18022 = ~w17736 & ~w17740;
assign w18023 = w18021 & ~w18022;
assign w18024 = ~w18021 & w18022;
assign w18025 = ~w18023 & ~w18024;
assign w18026 = w17882 & w18025;
assign w18027 = ~w17882 & ~w18025;
assign w18028 = ~w18026 & ~w18027;
assign w18029 = ~w17752 & ~w17757;
assign w18030 = w18028 & ~w18029;
assign w18031 = ~w18028 & w18029;
assign w18032 = ~w18030 & ~w18031;
assign w18033 = w17872 & w18032;
assign w18034 = ~w17872 & ~w18032;
assign w18035 = ~w18033 & ~w18034;
assign w18036 = b[50] & w3177;
assign w18037 = b[51] & w2973;
assign w18038 = b[52] & w2978;
assign w18039 = w2980 & ~w8371;
assign w18040 = ~w18037 & ~w18038;
assign w18041 = ~w18036 & w18040;
assign w18042 = ~w18039 & w18041;
assign w18043 = a[32] & ~w18042;
assign w18044 = ~a[32] & w18042;
assign w18045 = ~w18043 & ~w18044;
assign w18046 = ~w17769 & ~w17774;
assign w18047 = w18045 & ~w18046;
assign w18048 = ~w18045 & w18046;
assign w18049 = ~w18047 & ~w18048;
assign w18050 = w18035 & w18049;
assign w18051 = ~w18035 & ~w18049;
assign w18052 = ~w18050 & ~w18051;
assign w18053 = b[53] & ~w2622;
assign w18054 = b[54] & w2436;
assign w18055 = b[55] & w2438;
assign w18056 = w2432 & ~w9330;
assign w18057 = ~w18053 & ~w18054;
assign w18058 = ~w18055 & w18057;
assign w18059 = ~w18056 & w18058;
assign w18060 = a[29] & ~w18059;
assign w18061 = ~a[29] & w18059;
assign w18062 = ~w18060 & ~w18061;
assign w18063 = ~w17787 & ~w17790;
assign w18064 = w18062 & ~w18063;
assign w18065 = ~w18062 & w18063;
assign w18066 = ~w18064 & ~w18065;
assign w18067 = w18052 & w18066;
assign w18068 = ~w18052 & ~w18066;
assign w18069 = ~w18067 & ~w18068;
assign w18070 = w17862 & w18069;
assign w18071 = ~w17862 & ~w18069;
assign w18072 = ~w18070 & ~w18071;
assign w18073 = b[61] & w1519;
assign w18074 = b[59] & ~w1676;
assign w18075 = b[60] & w1517;
assign w18076 = ~w18073 & ~w18074;
assign w18077 = ~w18075 & w18076;
assign w18078 = (w11400 & w24874) | (w11400 & w24875) | (w24874 & w24875);
assign w18079 = (~w11400 & w24876) | (~w11400 & w24877) | (w24876 & w24877);
assign w18080 = ~w18078 & ~w18079;
assign w18081 = ~w17807 & ~w17811;
assign w18082 = w18080 & ~w18081;
assign w18083 = ~w18080 & w18081;
assign w18084 = ~w18082 & ~w18083;
assign w18085 = w18072 & w18084;
assign w18086 = ~w18072 & ~w18084;
assign w18087 = ~w18085 & ~w18086;
assign w18088 = (~w17822 & ~w17824) | (~w17822 & w25211) | (~w17824 & w25211);
assign w18089 = b[63] & w1154;
assign w18090 = b[62] & ~w1272;
assign w18091 = ~w12153 & w24720;
assign w18092 = ~w18089 & ~w18090;
assign w18093 = (a[20] & w18091) | (a[20] & w25025) | (w18091 & w25025);
assign w18094 = ~w18091 & w25026;
assign w18095 = ~w18093 & ~w18094;
assign w18096 = ~w18088 & w18095;
assign w18097 = w18088 & ~w18095;
assign w18098 = ~w18096 & ~w18097;
assign w18099 = w18087 & w18098;
assign w18100 = ~w18087 & ~w18098;
assign w18101 = ~w18099 & ~w18100;
assign w18102 = w17850 & ~w18101;
assign w18103 = ~w17850 & w18101;
assign w18104 = ~w18102 & ~w18103;
assign w18105 = ~w17845 & w25739;
assign w18106 = w18104 & w18105;
assign w18107 = ~w18104 & ~w18105;
assign w18108 = ~w18106 & ~w18107;
assign w18109 = (w16450 & w24440) | (w16450 & w24441) | (w24440 & w24441);
assign w18110 = (~w18096 & ~w18098) | (~w18096 & w25322) | (~w18098 & w25322);
assign w18111 = (~w18082 & ~w18084) | (~w18082 & w25027) | (~w18084 & w25027);
assign w18112 = w1150 & ~w12154;
assign w18113 = w1272 & ~w18112;
assign w18114 = b[63] & ~w18113;
assign w18115 = ~a[20] & ~w18114;
assign w18116 = a[20] & w18114;
assign w18117 = ~w18115 & ~w18116;
assign w18118 = ~w18111 & w18117;
assign w18119 = w18111 & ~w18117;
assign w18120 = ~w18118 & ~w18119;
assign w18121 = b[58] & w1955;
assign w18122 = b[57] & ~w2114;
assign w18123 = b[59] & w1957;
assign w18124 = ~w18121 & ~w18122;
assign w18125 = ~w18123 & w18124;
assign w18126 = (w10371 & w25212) | (w10371 & w25213) | (w25212 & w25213);
assign w18127 = (~w10371 & w25214) | (~w10371 & w25215) | (w25214 & w25215);
assign w18128 = ~w18126 & ~w18127;
assign w18129 = ~w18064 & ~w18067;
assign w18130 = w18128 & ~w18129;
assign w18131 = ~w18128 & w18129;
assign w18132 = ~w18130 & ~w18131;
assign w18133 = b[54] & ~w2622;
assign w18134 = b[56] & w2438;
assign w18135 = b[55] & w2436;
assign w18136 = ~w18133 & ~w18134;
assign w18137 = ~w18135 & w18136;
assign w18138 = (w18137 & ~w9657) | (w18137 & w25586) | (~w9657 & w25586);
assign w18139 = a[29] & ~w18138;
assign w18140 = ~a[29] & w18138;
assign w18141 = ~w18139 & ~w18140;
assign w18142 = ~w18047 & ~w18050;
assign w18143 = w18141 & ~w18142;
assign w18144 = ~w18141 & w18142;
assign w18145 = ~w18143 & ~w18144;
assign w18146 = b[48] & w3785;
assign w18147 = b[49] & w3578;
assign w18148 = b[50] & w3580;
assign w18149 = w3573 & w7759;
assign w18150 = ~w18147 & ~w18148;
assign w18151 = ~w18146 & w18150;
assign w18152 = ~w18149 & w18151;
assign w18153 = a[35] & ~w18152;
assign w18154 = ~a[35] & w18152;
assign w18155 = ~w18153 & ~w18154;
assign w18156 = ~w18007 & ~w18019;
assign w18157 = b[42] & w5167;
assign w18158 = b[43] & w4918;
assign w18159 = b[44] & w4925;
assign w18160 = w4923 & w6069;
assign w18161 = ~w18158 & ~w18159;
assign w18162 = ~w18157 & w18161;
assign w18163 = ~w18160 & w18162;
assign w18164 = a[41] & ~w18163;
assign w18165 = ~a[41] & w18163;
assign w18166 = ~w18164 & ~w18165;
assign w18167 = ~w18001 & ~w18003;
assign w18168 = b[39] & w5939;
assign w18169 = b[41] & w5665;
assign w18170 = b[40] & w5670;
assign w18171 = w5302 & w5663;
assign w18172 = ~w18169 & ~w18170;
assign w18173 = ~w18168 & w18172;
assign w18174 = ~w18171 & w18173;
assign w18175 = a[44] & ~w18174;
assign w18176 = ~a[44] & w18174;
assign w18177 = ~w18175 & ~w18176;
assign w18178 = ~w17994 & ~w17998;
assign w18179 = b[36] & w6732;
assign w18180 = b[38] & w6476;
assign w18181 = b[37] & w6474;
assign w18182 = w4582 & w6469;
assign w18183 = ~w18180 & ~w18181;
assign w18184 = ~w18179 & w18183;
assign w18185 = ~w18182 & w18184;
assign w18186 = a[47] & ~w18185;
assign w18187 = ~a[47] & w18185;
assign w18188 = ~w18186 & ~w18187;
assign w18189 = ~w17987 & ~w17990;
assign w18190 = b[33] & w7586;
assign w18191 = b[35] & w7314;
assign w18192 = b[34] & w7307;
assign w18193 = w3918 & w7312;
assign w18194 = ~w18191 & ~w18192;
assign w18195 = ~w18190 & w18194;
assign w18196 = ~w18193 & w18195;
assign w18197 = a[50] & ~w18196;
assign w18198 = ~a[50] & w18196;
assign w18199 = ~w18197 & ~w18198;
assign w18200 = ~w17970 & ~w17983;
assign w18201 = b[30] & w8515;
assign w18202 = b[31] & w8200;
assign w18203 = b[32] & w8202;
assign w18204 = w3304 & w8195;
assign w18205 = ~w18202 & ~w18203;
assign w18206 = ~w18201 & w18205;
assign w18207 = ~w18204 & w18206;
assign w18208 = a[53] & ~w18207;
assign w18209 = ~a[53] & w18207;
assign w18210 = ~w18208 & ~w18209;
assign w18211 = ~w17948 & ~w17961;
assign w18212 = b[24] & w10496;
assign w18213 = b[25] & w10146;
assign w18214 = b[26] & w10148;
assign w18215 = w2219 & w10141;
assign w18216 = ~w18213 & ~w18214;
assign w18217 = ~w18212 & w18216;
assign w18218 = ~w18215 & w18217;
assign w18219 = a[59] & ~w18218;
assign w18220 = ~a[59] & w18218;
assign w18221 = ~w18219 & ~w18220;
assign w18222 = ~w17931 & ~w17945;
assign w18223 = b[19] & w11921;
assign w18224 = b[20] & w11923;
assign w18225 = ~w18223 & ~w18224;
assign w18226 = w17929 & ~w18225;
assign w18227 = ~w17929 & w18225;
assign w18228 = ~w18226 & ~w18227;
assign w18229 = b[21] & w11561;
assign w18230 = b[23] & w11196;
assign w18231 = b[22] & w11194;
assign w18232 = w1755 & w11189;
assign w18233 = ~w18230 & ~w18231;
assign w18234 = ~w18229 & w18233;
assign w18235 = ~w18232 & w18234;
assign w18236 = a[62] & ~w18235;
assign w18237 = ~a[62] & w18235;
assign w18238 = ~w18236 & ~w18237;
assign w18239 = w18228 & w18238;
assign w18240 = ~w18228 & ~w18238;
assign w18241 = ~w18239 & ~w18240;
assign w18242 = w18222 & ~w18241;
assign w18243 = ~w18222 & w18241;
assign w18244 = ~w18242 & ~w18243;
assign w18245 = w18221 & w18244;
assign w18246 = ~w18221 & ~w18244;
assign w18247 = ~w18245 & ~w18246;
assign w18248 = w18211 & ~w18247;
assign w18249 = ~w18211 & w18247;
assign w18250 = ~w18248 & ~w18249;
assign w18251 = b[27] & w9482;
assign w18252 = b[29] & w9160;
assign w18253 = b[28] & w9165;
assign w18254 = w2734 & w9158;
assign w18255 = ~w18252 & ~w18253;
assign w18256 = ~w18251 & w18255;
assign w18257 = ~w18254 & w18256;
assign w18258 = a[56] & ~w18257;
assign w18259 = ~a[56] & w18257;
assign w18260 = ~w18258 & ~w18259;
assign w18261 = w18250 & w18260;
assign w18262 = ~w18250 & ~w18260;
assign w18263 = ~w18261 & ~w18262;
assign w18264 = ~w17964 & ~w17967;
assign w18265 = w18263 & ~w18264;
assign w18266 = ~w18263 & w18264;
assign w18267 = ~w18265 & ~w18266;
assign w18268 = w18210 & w18267;
assign w18269 = ~w18210 & ~w18267;
assign w18270 = ~w18268 & ~w18269;
assign w18271 = ~w18200 & w18270;
assign w18272 = w18200 & ~w18270;
assign w18273 = ~w18271 & ~w18272;
assign w18274 = w18199 & w18273;
assign w18275 = ~w18199 & ~w18273;
assign w18276 = ~w18274 & ~w18275;
assign w18277 = w18189 & ~w18276;
assign w18278 = ~w18189 & w18276;
assign w18279 = ~w18277 & ~w18278;
assign w18280 = w18188 & w18279;
assign w18281 = ~w18188 & ~w18279;
assign w18282 = ~w18280 & ~w18281;
assign w18283 = w18178 & ~w18282;
assign w18284 = ~w18178 & w18282;
assign w18285 = ~w18283 & ~w18284;
assign w18286 = w18177 & w18285;
assign w18287 = ~w18177 & ~w18285;
assign w18288 = ~w18286 & ~w18287;
assign w18289 = w18167 & ~w18288;
assign w18290 = ~w18167 & w18288;
assign w18291 = ~w18289 & ~w18290;
assign w18292 = w18166 & w18291;
assign w18293 = ~w18166 & ~w18291;
assign w18294 = ~w18292 & ~w18293;
assign w18295 = w18156 & ~w18294;
assign w18296 = ~w18156 & w18294;
assign w18297 = ~w18295 & ~w18296;
assign w18298 = b[45] & w4453;
assign w18299 = b[46] & w4241;
assign w18300 = b[47] & w4243;
assign w18301 = w4236 & w6889;
assign w18302 = ~w18299 & ~w18300;
assign w18303 = ~w18298 & w18302;
assign w18304 = ~w18301 & w18303;
assign w18305 = a[38] & ~w18304;
assign w18306 = ~a[38] & w18304;
assign w18307 = ~w18305 & ~w18306;
assign w18308 = w18297 & w18307;
assign w18309 = ~w18297 & ~w18307;
assign w18310 = ~w18308 & ~w18309;
assign w18311 = ~w18023 & ~w18026;
assign w18312 = w18310 & ~w18311;
assign w18313 = ~w18310 & w18311;
assign w18314 = ~w18312 & ~w18313;
assign w18315 = w18155 & w18314;
assign w18316 = ~w18155 & ~w18314;
assign w18317 = ~w18315 & ~w18316;
assign w18318 = b[51] & w3177;
assign w18319 = b[53] & w2978;
assign w18320 = b[52] & w2973;
assign w18321 = w2980 & w8683;
assign w18322 = ~w18319 & ~w18320;
assign w18323 = ~w18318 & w18322;
assign w18324 = ~w18321 & w18323;
assign w18325 = a[32] & ~w18324;
assign w18326 = ~a[32] & w18324;
assign w18327 = ~w18325 & ~w18326;
assign w18328 = ~w18030 & ~w18033;
assign w18329 = w18327 & ~w18328;
assign w18330 = ~w18327 & w18328;
assign w18331 = ~w18329 & ~w18330;
assign w18332 = w18317 & w18331;
assign w18333 = ~w18317 & ~w18331;
assign w18334 = ~w18332 & ~w18333;
assign w18335 = w18145 & w18334;
assign w18336 = ~w18145 & ~w18334;
assign w18337 = ~w18335 & ~w18336;
assign w18338 = w18132 & w18337;
assign w18339 = ~w18132 & ~w18337;
assign w18340 = ~w18338 & ~w18339;
assign w18341 = b[60] & ~w1676;
assign w18342 = b[62] & w1519;
assign w18343 = b[61] & w1517;
assign w18344 = ~w18341 & ~w18342;
assign w18345 = ~w18343 & w18344;
assign w18346 = (w11763 & w24878) | (w11763 & w24879) | (w24878 & w24879);
assign w18347 = (~w11763 & w24880) | (~w11763 & w24881) | (w24880 & w24881);
assign w18348 = ~w18346 & ~w18347;
assign w18349 = ~w17860 & ~w18070;
assign w18350 = w18348 & ~w18349;
assign w18351 = ~w18348 & w18349;
assign w18352 = ~w18350 & ~w18351;
assign w18353 = w18340 & w18352;
assign w18354 = ~w18340 & ~w18352;
assign w18355 = ~w18353 & ~w18354;
assign w18356 = w18120 & w18355;
assign w18357 = ~w18120 & ~w18355;
assign w18358 = ~w18356 & ~w18357;
assign w18359 = ~w18110 & w18358;
assign w18360 = w18110 & ~w18358;
assign w18361 = ~w18359 & ~w18360;
assign w18362 = ~w18102 & w18361;
assign w18363 = ~w18109 & w18362;
assign w18364 = ~w18103 & ~w18361;
assign w18365 = ~w18106 & w18364;
assign w18366 = ~w18363 & ~w18365;
assign w18367 = b[52] & w3177;
assign w18368 = b[54] & w2978;
assign w18369 = b[53] & w2973;
assign w18370 = w2980 & ~w8998;
assign w18371 = ~w18368 & ~w18369;
assign w18372 = ~w18367 & w18371;
assign w18373 = ~w18370 & w18372;
assign w18374 = a[32] & ~w18373;
assign w18375 = ~a[32] & w18373;
assign w18376 = ~w18374 & ~w18375;
assign w18377 = ~w18329 & ~w18332;
assign w18378 = w18376 & ~w18377;
assign w18379 = ~w18376 & w18377;
assign w18380 = ~w18378 & ~w18379;
assign w18381 = ~w18312 & ~w18315;
assign w18382 = ~w18271 & ~w18274;
assign w18383 = b[34] & w7586;
assign w18384 = b[35] & w7307;
assign w18385 = b[36] & w7314;
assign w18386 = w4129 & w7312;
assign w18387 = ~w18384 & ~w18385;
assign w18388 = ~w18383 & w18387;
assign w18389 = ~w18386 & w18388;
assign w18390 = a[50] & ~w18389;
assign w18391 = ~a[50] & w18389;
assign w18392 = ~w18390 & ~w18391;
assign w18393 = ~w18243 & ~w18245;
assign w18394 = b[25] & w10496;
assign w18395 = b[26] & w10146;
assign w18396 = b[27] & w10148;
assign w18397 = w2378 & w10141;
assign w18398 = ~w18395 & ~w18396;
assign w18399 = ~w18394 & w18398;
assign w18400 = ~w18397 & w18399;
assign w18401 = a[59] & ~w18400;
assign w18402 = ~a[59] & w18400;
assign w18403 = ~w18401 & ~w18402;
assign w18404 = b[20] & w11921;
assign w18405 = b[21] & w11923;
assign w18406 = ~w18404 & ~w18405;
assign w18407 = ~a[20] & ~w18406;
assign w18408 = a[20] & w18406;
assign w18409 = ~w18407 & ~w18408;
assign w18410 = ~w18225 & w18409;
assign w18411 = w18225 & ~w18409;
assign w18412 = ~w18410 & ~w18411;
assign w18413 = b[22] & w11561;
assign w18414 = b[24] & w11196;
assign w18415 = b[23] & w11194;
assign w18416 = w1895 & w11189;
assign w18417 = ~w18414 & ~w18415;
assign w18418 = ~w18413 & w18417;
assign w18419 = ~w18416 & w18418;
assign w18420 = a[62] & ~w18419;
assign w18421 = ~a[62] & w18419;
assign w18422 = ~w18420 & ~w18421;
assign w18423 = w18412 & w18422;
assign w18424 = ~w18412 & ~w18422;
assign w18425 = ~w18423 & ~w18424;
assign w18426 = ~w18227 & ~w18239;
assign w18427 = w18425 & ~w18426;
assign w18428 = ~w18425 & w18426;
assign w18429 = ~w18427 & ~w18428;
assign w18430 = w18403 & w18429;
assign w18431 = ~w18403 & ~w18429;
assign w18432 = ~w18430 & ~w18431;
assign w18433 = w18393 & ~w18432;
assign w18434 = ~w18393 & w18432;
assign w18435 = ~w18433 & ~w18434;
assign w18436 = b[28] & w9482;
assign w18437 = b[29] & w9165;
assign w18438 = b[30] & w9160;
assign w18439 = ~w2908 & w9158;
assign w18440 = ~w18437 & ~w18438;
assign w18441 = ~w18436 & w18440;
assign w18442 = ~w18439 & w18441;
assign w18443 = a[56] & ~w18442;
assign w18444 = ~a[56] & w18442;
assign w18445 = ~w18443 & ~w18444;
assign w18446 = w18435 & w18445;
assign w18447 = ~w18435 & ~w18445;
assign w18448 = ~w18446 & ~w18447;
assign w18449 = ~w18249 & ~w18261;
assign w18450 = ~w18448 & w18449;
assign w18451 = w18448 & ~w18449;
assign w18452 = ~w18450 & ~w18451;
assign w18453 = b[31] & w8515;
assign w18454 = b[32] & w8200;
assign w18455 = b[33] & w8202;
assign w18456 = w3499 & w8195;
assign w18457 = ~w18454 & ~w18455;
assign w18458 = ~w18453 & w18457;
assign w18459 = ~w18456 & w18458;
assign w18460 = a[53] & ~w18459;
assign w18461 = ~a[53] & w18459;
assign w18462 = ~w18460 & ~w18461;
assign w18463 = ~w18265 & ~w18268;
assign w18464 = w18462 & ~w18463;
assign w18465 = ~w18462 & w18463;
assign w18466 = ~w18464 & ~w18465;
assign w18467 = w18452 & w18466;
assign w18468 = ~w18452 & ~w18466;
assign w18469 = ~w18467 & ~w18468;
assign w18470 = w18392 & w18469;
assign w18471 = ~w18392 & ~w18469;
assign w18472 = ~w18470 & ~w18471;
assign w18473 = w18382 & ~w18472;
assign w18474 = ~w18382 & w18472;
assign w18475 = ~w18473 & ~w18474;
assign w18476 = b[37] & w6732;
assign w18477 = b[38] & w6474;
assign w18478 = b[39] & w6476;
assign w18479 = ~w4812 & w6469;
assign w18480 = ~w18477 & ~w18478;
assign w18481 = ~w18476 & w18480;
assign w18482 = ~w18479 & w18481;
assign w18483 = a[47] & ~w18482;
assign w18484 = ~a[47] & w18482;
assign w18485 = ~w18483 & ~w18484;
assign w18486 = w18475 & w18485;
assign w18487 = ~w18475 & ~w18485;
assign w18488 = ~w18486 & ~w18487;
assign w18489 = ~w18278 & ~w18280;
assign w18490 = ~w18488 & w18489;
assign w18491 = w18488 & ~w18489;
assign w18492 = ~w18490 & ~w18491;
assign w18493 = b[40] & w5939;
assign w18494 = b[41] & w5670;
assign w18495 = b[42] & w5665;
assign w18496 = w5548 & w5663;
assign w18497 = ~w18494 & ~w18495;
assign w18498 = ~w18493 & w18497;
assign w18499 = ~w18496 & w18498;
assign w18500 = a[44] & ~w18499;
assign w18501 = ~a[44] & w18499;
assign w18502 = ~w18500 & ~w18501;
assign w18503 = w18492 & w18502;
assign w18504 = ~w18492 & ~w18502;
assign w18505 = ~w18503 & ~w18504;
assign w18506 = ~w18284 & ~w18286;
assign w18507 = ~w18505 & w18506;
assign w18508 = w18505 & ~w18506;
assign w18509 = ~w18507 & ~w18508;
assign w18510 = b[43] & w5167;
assign w18511 = b[45] & w4925;
assign w18512 = b[44] & w4918;
assign w18513 = w4923 & w6334;
assign w18514 = ~w18511 & ~w18512;
assign w18515 = ~w18510 & w18514;
assign w18516 = ~w18513 & w18515;
assign w18517 = a[41] & ~w18516;
assign w18518 = ~a[41] & w18516;
assign w18519 = ~w18517 & ~w18518;
assign w18520 = w18509 & w18519;
assign w18521 = ~w18509 & ~w18519;
assign w18522 = ~w18520 & ~w18521;
assign w18523 = ~w18290 & ~w18292;
assign w18524 = ~w18522 & w18523;
assign w18525 = w18522 & ~w18523;
assign w18526 = ~w18524 & ~w18525;
assign w18527 = b[46] & w4453;
assign w18528 = b[47] & w4241;
assign w18529 = b[48] & w4243;
assign w18530 = w4236 & ~w7170;
assign w18531 = ~w18528 & ~w18529;
assign w18532 = ~w18527 & w18531;
assign w18533 = ~w18530 & w18532;
assign w18534 = a[38] & ~w18533;
assign w18535 = ~a[38] & w18533;
assign w18536 = ~w18534 & ~w18535;
assign w18537 = w18526 & w18536;
assign w18538 = ~w18526 & ~w18536;
assign w18539 = ~w18537 & ~w18538;
assign w18540 = ~w18296 & ~w18308;
assign w18541 = ~w18539 & w18540;
assign w18542 = w18539 & ~w18540;
assign w18543 = ~w18541 & ~w18542;
assign w18544 = b[49] & w3785;
assign w18545 = b[51] & w3580;
assign w18546 = b[50] & w3578;
assign w18547 = w3573 & ~w8058;
assign w18548 = ~w18545 & ~w18546;
assign w18549 = ~w18544 & w18548;
assign w18550 = ~w18547 & w18549;
assign w18551 = a[35] & ~w18550;
assign w18552 = ~a[35] & w18550;
assign w18553 = ~w18551 & ~w18552;
assign w18554 = ~w18543 & ~w18553;
assign w18555 = w18543 & w18553;
assign w18556 = ~w18554 & ~w18555;
assign w18557 = w18381 & w18556;
assign w18558 = ~w18381 & ~w18556;
assign w18559 = ~w18557 & ~w18558;
assign w18560 = w18380 & ~w18559;
assign w18561 = ~w18380 & w18559;
assign w18562 = ~w18560 & ~w18561;
assign w18563 = ~w18143 & ~w18335;
assign w18564 = b[56] & w2436;
assign w18565 = b[57] & w2438;
assign w18566 = b[55] & ~w2622;
assign w18567 = w2432 & ~w9992;
assign w18568 = ~w18564 & ~w18565;
assign w18569 = ~w18566 & w18568;
assign w18570 = ~w18567 & w18569;
assign w18571 = a[29] & ~w18570;
assign w18572 = ~a[29] & w18570;
assign w18573 = ~w18571 & ~w18572;
assign w18574 = ~w18563 & w18573;
assign w18575 = w18563 & ~w18573;
assign w18576 = ~w18574 & ~w18575;
assign w18577 = ~w18562 & ~w18576;
assign w18578 = w18562 & w18576;
assign w18579 = ~w18577 & ~w18578;
assign w18580 = b[59] & w1955;
assign w18581 = b[58] & ~w2114;
assign w18582 = b[60] & w1957;
assign w18583 = ~w18580 & ~w18581;
assign w18584 = ~w18582 & w18583;
assign w18585 = (w11035 & w25469) | (w11035 & w25470) | (w25469 & w25470);
assign w18586 = ~a[26] & w25740;
assign w18587 = ~w18585 & ~w18586;
assign w18588 = (~w18130 & ~w18132) | (~w18130 & w25324) | (~w18132 & w25324);
assign w18589 = w18587 & ~w18588;
assign w18590 = ~w18587 & w18588;
assign w18591 = ~w18589 & ~w18590;
assign w18592 = w18579 & w18591;
assign w18593 = ~w18579 & ~w18591;
assign w18594 = ~w18592 & ~w18593;
assign w18595 = (~w18350 & ~w18352) | (~w18350 & w25029) | (~w18352 & w25029);
assign w18596 = b[61] & ~w1676;
assign w18597 = b[62] & w1517;
assign w18598 = b[63] & w1519;
assign w18599 = ~w18596 & ~w18597;
assign w18600 = ~w18598 & w18599;
assign w18601 = (w18600 & ~w12132) | (w18600 & w25471) | (~w12132 & w25471);
assign w18602 = a[23] & ~w18601;
assign w18603 = ~a[23] & w18601;
assign w18604 = ~w18602 & ~w18603;
assign w18605 = ~w18595 & w18604;
assign w18606 = w18595 & ~w18604;
assign w18607 = ~w18605 & ~w18606;
assign w18608 = ~w18594 & ~w18607;
assign w18609 = w18594 & w18607;
assign w18610 = ~w18608 & ~w18609;
assign w18611 = (~w18118 & ~w18120) | (~w18118 & w25472) | (~w18120 & w25472);
assign w18612 = ~w18610 & w18611;
assign w18613 = w18610 & ~w18611;
assign w18614 = ~w18612 & ~w18613;
assign w18615 = (~w18359 & w18109) | (~w18359 & w24442) | (w18109 & w24442);
assign w18616 = ~w18614 & w18615;
assign w18617 = w18614 & ~w18615;
assign w18618 = ~w18616 & ~w18617;
assign w18619 = (~w18605 & ~w18607) | (~w18605 & w25587) | (~w18607 & w25587);
assign w18620 = b[61] & w1957;
assign w18621 = b[60] & w1955;
assign w18622 = b[59] & ~w2114;
assign w18623 = ~w18620 & ~w18621;
assign w18624 = ~w18622 & w18623;
assign w18625 = (w11400 & w25588) | (w11400 & w25589) | (w25588 & w25589);
assign w18626 = (~w11400 & w25590) | (~w11400 & w25591) | (w25590 & w25591);
assign w18627 = ~w18625 & ~w18626;
assign w18628 = ~w18574 & ~w18578;
assign w18629 = w18627 & ~w18628;
assign w18630 = ~w18627 & w18628;
assign w18631 = ~w18629 & ~w18630;
assign w18632 = b[50] & w3785;
assign w18633 = b[51] & w3578;
assign w18634 = b[52] & w3580;
assign w18635 = w3573 & ~w8371;
assign w18636 = ~w18633 & ~w18634;
assign w18637 = ~w18632 & w18636;
assign w18638 = ~w18635 & w18637;
assign w18639 = a[35] & ~w18638;
assign w18640 = ~a[35] & w18638;
assign w18641 = ~w18639 & ~w18640;
assign w18642 = b[47] & w4453;
assign w18643 = b[49] & w4243;
assign w18644 = b[48] & w4241;
assign w18645 = w4236 & ~w7468;
assign w18646 = ~w18643 & ~w18644;
assign w18647 = ~w18642 & w18646;
assign w18648 = ~w18645 & w18647;
assign w18649 = a[38] & ~w18648;
assign w18650 = ~a[38] & w18648;
assign w18651 = ~w18649 & ~w18650;
assign w18652 = b[44] & w5167;
assign w18653 = b[46] & w4925;
assign w18654 = b[45] & w4918;
assign w18655 = w4923 & ~w6613;
assign w18656 = ~w18653 & ~w18654;
assign w18657 = ~w18652 & w18656;
assign w18658 = ~w18655 & w18657;
assign w18659 = a[41] & ~w18658;
assign w18660 = ~a[41] & w18658;
assign w18661 = ~w18659 & ~w18660;
assign w18662 = ~w18486 & ~w18491;
assign w18663 = b[38] & w6732;
assign w18664 = b[39] & w6474;
assign w18665 = b[40] & w6476;
assign w18666 = ~w5058 & w6469;
assign w18667 = ~w18664 & ~w18665;
assign w18668 = ~w18663 & w18667;
assign w18669 = ~w18666 & w18668;
assign w18670 = a[47] & ~w18669;
assign w18671 = ~a[47] & w18669;
assign w18672 = ~w18670 & ~w18671;
assign w18673 = ~w18470 & ~w18474;
assign w18674 = b[35] & w7586;
assign w18675 = b[37] & w7314;
assign w18676 = b[36] & w7307;
assign w18677 = ~w4357 & w7312;
assign w18678 = ~w18675 & ~w18676;
assign w18679 = ~w18674 & w18678;
assign w18680 = ~w18677 & w18679;
assign w18681 = a[50] & ~w18680;
assign w18682 = ~a[50] & w18680;
assign w18683 = ~w18681 & ~w18682;
assign w18684 = b[32] & w8515;
assign w18685 = b[33] & w8200;
assign w18686 = b[34] & w8202;
assign w18687 = ~w3710 & w8195;
assign w18688 = ~w18685 & ~w18686;
assign w18689 = ~w18684 & w18688;
assign w18690 = ~w18687 & w18689;
assign w18691 = a[53] & ~w18690;
assign w18692 = ~a[53] & w18690;
assign w18693 = ~w18691 & ~w18692;
assign w18694 = ~w18430 & ~w18434;
assign w18695 = b[26] & w10496;
assign w18696 = b[28] & w10148;
assign w18697 = b[27] & w10146;
assign w18698 = w2559 & w10141;
assign w18699 = ~w18696 & ~w18697;
assign w18700 = ~w18695 & w18699;
assign w18701 = ~w18698 & w18700;
assign w18702 = a[59] & ~w18701;
assign w18703 = ~a[59] & w18701;
assign w18704 = ~w18702 & ~w18703;
assign w18705 = ~w18423 & ~w18427;
assign w18706 = b[21] & w11921;
assign w18707 = b[22] & w11923;
assign w18708 = ~w18706 & ~w18707;
assign w18709 = ~w18407 & ~w18410;
assign w18710 = w18708 & ~w18709;
assign w18711 = ~w18708 & w18709;
assign w18712 = ~w18710 & ~w18711;
assign w18713 = b[23] & w11561;
assign w18714 = b[24] & w11194;
assign w18715 = b[25] & w11196;
assign w18716 = w2061 & w11189;
assign w18717 = ~w18714 & ~w18715;
assign w18718 = ~w18713 & w18717;
assign w18719 = ~w18716 & w18718;
assign w18720 = a[62] & ~w18719;
assign w18721 = ~a[62] & w18719;
assign w18722 = ~w18720 & ~w18721;
assign w18723 = w18712 & w18722;
assign w18724 = ~w18712 & ~w18722;
assign w18725 = ~w18723 & ~w18724;
assign w18726 = w18705 & ~w18725;
assign w18727 = ~w18705 & w18725;
assign w18728 = ~w18726 & ~w18727;
assign w18729 = w18704 & w18728;
assign w18730 = ~w18704 & ~w18728;
assign w18731 = ~w18729 & ~w18730;
assign w18732 = w18694 & ~w18731;
assign w18733 = ~w18694 & w18731;
assign w18734 = ~w18732 & ~w18733;
assign w18735 = b[29] & w9482;
assign w18736 = b[30] & w9165;
assign w18737 = b[31] & w9160;
assign w18738 = ~w3112 & w9158;
assign w18739 = ~w18736 & ~w18737;
assign w18740 = ~w18735 & w18739;
assign w18741 = ~w18738 & w18740;
assign w18742 = a[56] & ~w18741;
assign w18743 = ~a[56] & w18741;
assign w18744 = ~w18742 & ~w18743;
assign w18745 = w18734 & w18744;
assign w18746 = ~w18734 & ~w18744;
assign w18747 = ~w18745 & ~w18746;
assign w18748 = ~w18446 & ~w18451;
assign w18749 = w18747 & ~w18748;
assign w18750 = ~w18747 & w18748;
assign w18751 = ~w18749 & ~w18750;
assign w18752 = w18693 & w18751;
assign w18753 = ~w18693 & ~w18751;
assign w18754 = ~w18752 & ~w18753;
assign w18755 = ~w18464 & ~w18467;
assign w18756 = w18754 & ~w18755;
assign w18757 = ~w18754 & w18755;
assign w18758 = ~w18756 & ~w18757;
assign w18759 = ~w18683 & ~w18758;
assign w18760 = w18683 & w18758;
assign w18761 = ~w18759 & ~w18760;
assign w18762 = w18673 & ~w18761;
assign w18763 = ~w18673 & w18761;
assign w18764 = ~w18762 & ~w18763;
assign w18765 = w18672 & w18764;
assign w18766 = ~w18672 & ~w18764;
assign w18767 = ~w18765 & ~w18766;
assign w18768 = w18662 & ~w18767;
assign w18769 = ~w18662 & w18767;
assign w18770 = ~w18768 & ~w18769;
assign w18771 = b[41] & w5939;
assign w18772 = b[43] & w5665;
assign w18773 = b[42] & w5670;
assign w18774 = w5663 & w5811;
assign w18775 = ~w18772 & ~w18773;
assign w18776 = ~w18771 & w18775;
assign w18777 = ~w18774 & w18776;
assign w18778 = a[44] & ~w18777;
assign w18779 = ~a[44] & w18777;
assign w18780 = ~w18778 & ~w18779;
assign w18781 = w18770 & w18780;
assign w18782 = ~w18770 & ~w18780;
assign w18783 = ~w18781 & ~w18782;
assign w18784 = ~w18503 & ~w18508;
assign w18785 = w18783 & ~w18784;
assign w18786 = ~w18783 & w18784;
assign w18787 = ~w18785 & ~w18786;
assign w18788 = w18661 & w18787;
assign w18789 = ~w18661 & ~w18787;
assign w18790 = ~w18788 & ~w18789;
assign w18791 = ~w18520 & ~w18525;
assign w18792 = w18790 & ~w18791;
assign w18793 = ~w18790 & w18791;
assign w18794 = ~w18792 & ~w18793;
assign w18795 = w18651 & w18794;
assign w18796 = ~w18651 & ~w18794;
assign w18797 = ~w18795 & ~w18796;
assign w18798 = ~w18537 & ~w18542;
assign w18799 = w18797 & ~w18798;
assign w18800 = ~w18797 & w18798;
assign w18801 = ~w18799 & ~w18800;
assign w18802 = w18641 & w18801;
assign w18803 = ~w18641 & ~w18801;
assign w18804 = ~w18802 & ~w18803;
assign w18805 = b[53] & w3177;
assign w18806 = b[54] & w2973;
assign w18807 = b[55] & w2978;
assign w18808 = w2980 & ~w9330;
assign w18809 = ~w18806 & ~w18807;
assign w18810 = ~w18805 & w18809;
assign w18811 = ~w18808 & w18810;
assign w18812 = a[32] & ~w18811;
assign w18813 = ~a[32] & w18811;
assign w18814 = ~w18812 & ~w18813;
assign w18815 = ~w18554 & ~w18557;
assign w18816 = w18814 & w18815;
assign w18817 = ~w18814 & ~w18815;
assign w18818 = ~w18816 & ~w18817;
assign w18819 = w18804 & w18818;
assign w18820 = ~w18804 & ~w18818;
assign w18821 = ~w18819 & ~w18820;
assign w18822 = ~w18378 & ~w18560;
assign w18823 = b[58] & w2438;
assign w18824 = b[56] & ~w2622;
assign w18825 = b[57] & w2436;
assign w18826 = w2432 & ~w10339;
assign w18827 = ~w18823 & ~w18824;
assign w18828 = ~w18825 & w18827;
assign w18829 = ~w18826 & w18828;
assign w18830 = a[29] & ~w18829;
assign w18831 = ~a[29] & w18829;
assign w18832 = ~w18830 & ~w18831;
assign w18833 = ~w18822 & w18832;
assign w18834 = w18822 & ~w18832;
assign w18835 = ~w18833 & ~w18834;
assign w18836 = w18821 & w18835;
assign w18837 = ~w18821 & ~w18835;
assign w18838 = ~w18836 & ~w18837;
assign w18839 = w18631 & w18838;
assign w18840 = ~w18631 & ~w18838;
assign w18841 = ~w18839 & ~w18840;
assign w18842 = (~w18589 & ~w18591) | (~w18589 & w25474) | (~w18591 & w25474);
assign w18843 = b[62] & ~w1676;
assign w18844 = b[63] & w1517;
assign w18845 = ~w12153 & w25475;
assign w18846 = ~w18843 & ~w18844;
assign w18847 = (a[23] & w18845) | (a[23] & w25592) | (w18845 & w25592);
assign w18848 = ~w18845 & w25593;
assign w18849 = ~w18847 & ~w18848;
assign w18850 = ~w18842 & w18849;
assign w18851 = w18842 & ~w18849;
assign w18852 = ~w18850 & ~w18851;
assign w18853 = w18841 & w18852;
assign w18854 = ~w18841 & ~w18852;
assign w18855 = ~w18853 & ~w18854;
assign w18856 = w18619 & ~w18855;
assign w18857 = ~w18619 & w18855;
assign w18858 = ~w18856 & ~w18857;
assign w18859 = (w18109 & w24443) | (w18109 & w24444) | (w24443 & w24444);
assign w18860 = w18858 & ~w18859;
assign w18861 = ~w18858 & w18859;
assign w18862 = ~w18860 & ~w18861;
assign w18863 = ~w18850 & ~w18853;
assign w18864 = b[62] & w1957;
assign w18865 = b[60] & ~w2114;
assign w18866 = b[61] & w1955;
assign w18867 = w1951 & w11763;
assign w18868 = ~w18864 & ~w18865;
assign w18869 = ~w18866 & w18868;
assign w18870 = ~w18867 & w18869;
assign w18871 = a[26] & ~w18870;
assign w18872 = ~a[26] & w18870;
assign w18873 = ~w18871 & ~w18872;
assign w18874 = ~w18833 & ~w18836;
assign w18875 = w18873 & ~w18874;
assign w18876 = ~w18873 & w18874;
assign w18877 = ~w18875 & ~w18876;
assign w18878 = b[54] & w3177;
assign w18879 = b[56] & w2978;
assign w18880 = b[55] & w2973;
assign w18881 = w2980 & w9657;
assign w18882 = ~w18879 & ~w18880;
assign w18883 = ~w18878 & w18882;
assign w18884 = ~w18881 & w18883;
assign w18885 = a[32] & ~w18884;
assign w18886 = ~a[32] & w18884;
assign w18887 = ~w18885 & ~w18886;
assign w18888 = ~w18799 & ~w18802;
assign w18889 = w18887 & ~w18888;
assign w18890 = ~w18887 & w18888;
assign w18891 = ~w18889 & ~w18890;
assign w18892 = b[51] & w3785;
assign w18893 = b[52] & w3578;
assign w18894 = b[53] & w3580;
assign w18895 = w3573 & w8683;
assign w18896 = ~w18893 & ~w18894;
assign w18897 = ~w18892 & w18896;
assign w18898 = ~w18895 & w18897;
assign w18899 = a[35] & ~w18898;
assign w18900 = ~a[35] & w18898;
assign w18901 = ~w18899 & ~w18900;
assign w18902 = ~w18792 & ~w18795;
assign w18903 = b[48] & w4453;
assign w18904 = b[50] & w4243;
assign w18905 = b[49] & w4241;
assign w18906 = w4236 & w7759;
assign w18907 = ~w18904 & ~w18905;
assign w18908 = ~w18903 & w18907;
assign w18909 = ~w18906 & w18908;
assign w18910 = a[38] & ~w18909;
assign w18911 = ~a[38] & w18909;
assign w18912 = ~w18910 & ~w18911;
assign w18913 = ~w18769 & ~w18781;
assign w18914 = b[42] & w5939;
assign w18915 = b[43] & w5670;
assign w18916 = b[44] & w5665;
assign w18917 = w5663 & w6069;
assign w18918 = ~w18915 & ~w18916;
assign w18919 = ~w18914 & w18918;
assign w18920 = ~w18917 & w18919;
assign w18921 = a[44] & ~w18920;
assign w18922 = ~a[44] & w18920;
assign w18923 = ~w18921 & ~w18922;
assign w18924 = ~w18763 & ~w18765;
assign w18925 = b[39] & w6732;
assign w18926 = b[41] & w6476;
assign w18927 = b[40] & w6474;
assign w18928 = w5302 & w6469;
assign w18929 = ~w18926 & ~w18927;
assign w18930 = ~w18925 & w18929;
assign w18931 = ~w18928 & w18930;
assign w18932 = a[47] & ~w18931;
assign w18933 = ~a[47] & w18931;
assign w18934 = ~w18932 & ~w18933;
assign w18935 = ~w18749 & ~w18752;
assign w18936 = b[33] & w8515;
assign w18937 = b[35] & w8202;
assign w18938 = b[34] & w8200;
assign w18939 = w3918 & w8195;
assign w18940 = ~w18937 & ~w18938;
assign w18941 = ~w18936 & w18940;
assign w18942 = ~w18939 & w18941;
assign w18943 = a[53] & ~w18942;
assign w18944 = ~a[53] & w18942;
assign w18945 = ~w18943 & ~w18944;
assign w18946 = ~w18733 & ~w18745;
assign w18947 = b[30] & w9482;
assign w18948 = b[31] & w9165;
assign w18949 = b[32] & w9160;
assign w18950 = w3304 & w9158;
assign w18951 = ~w18948 & ~w18949;
assign w18952 = ~w18947 & w18951;
assign w18953 = ~w18950 & w18952;
assign w18954 = a[56] & ~w18953;
assign w18955 = ~a[56] & w18953;
assign w18956 = ~w18954 & ~w18955;
assign w18957 = ~w18710 & ~w18723;
assign w18958 = b[22] & w11921;
assign w18959 = b[23] & w11923;
assign w18960 = ~w18958 & ~w18959;
assign w18961 = w18708 & ~w18960;
assign w18962 = ~w18708 & w18960;
assign w18963 = ~w18961 & ~w18962;
assign w18964 = b[24] & w11561;
assign w18965 = b[26] & w11196;
assign w18966 = b[25] & w11194;
assign w18967 = w2219 & w11189;
assign w18968 = ~w18965 & ~w18966;
assign w18969 = ~w18964 & w18968;
assign w18970 = ~w18967 & w18969;
assign w18971 = a[62] & ~w18970;
assign w18972 = ~a[62] & w18970;
assign w18973 = ~w18971 & ~w18972;
assign w18974 = w18963 & w18973;
assign w18975 = ~w18963 & ~w18973;
assign w18976 = ~w18974 & ~w18975;
assign w18977 = w18957 & ~w18976;
assign w18978 = ~w18957 & w18976;
assign w18979 = ~w18977 & ~w18978;
assign w18980 = b[27] & w10496;
assign w18981 = b[29] & w10148;
assign w18982 = b[28] & w10146;
assign w18983 = w2734 & w10141;
assign w18984 = ~w18981 & ~w18982;
assign w18985 = ~w18980 & w18984;
assign w18986 = ~w18983 & w18985;
assign w18987 = a[59] & ~w18986;
assign w18988 = ~a[59] & w18986;
assign w18989 = ~w18987 & ~w18988;
assign w18990 = w18979 & w18989;
assign w18991 = ~w18979 & ~w18989;
assign w18992 = ~w18990 & ~w18991;
assign w18993 = ~w18727 & ~w18729;
assign w18994 = w18992 & ~w18993;
assign w18995 = ~w18992 & w18993;
assign w18996 = ~w18994 & ~w18995;
assign w18997 = ~w18956 & ~w18996;
assign w18998 = w18956 & w18996;
assign w18999 = ~w18997 & ~w18998;
assign w19000 = w18946 & ~w18999;
assign w19001 = ~w18946 & w18999;
assign w19002 = ~w19000 & ~w19001;
assign w19003 = w18945 & w19002;
assign w19004 = ~w18945 & ~w19002;
assign w19005 = ~w19003 & ~w19004;
assign w19006 = w18935 & ~w19005;
assign w19007 = ~w18935 & w19005;
assign w19008 = ~w19006 & ~w19007;
assign w19009 = b[36] & w7586;
assign w19010 = b[38] & w7314;
assign w19011 = b[37] & w7307;
assign w19012 = w4582 & w7312;
assign w19013 = ~w19010 & ~w19011;
assign w19014 = ~w19009 & w19013;
assign w19015 = ~w19012 & w19014;
assign w19016 = a[50] & ~w19015;
assign w19017 = ~a[50] & w19015;
assign w19018 = ~w19016 & ~w19017;
assign w19019 = w19008 & w19018;
assign w19020 = ~w19008 & ~w19018;
assign w19021 = ~w19019 & ~w19020;
assign w19022 = ~w18756 & ~w18760;
assign w19023 = w19021 & ~w19022;
assign w19024 = ~w19021 & w19022;
assign w19025 = ~w19023 & ~w19024;
assign w19026 = w18934 & w19025;
assign w19027 = ~w18934 & ~w19025;
assign w19028 = ~w19026 & ~w19027;
assign w19029 = ~w18924 & w19028;
assign w19030 = w18924 & ~w19028;
assign w19031 = ~w19029 & ~w19030;
assign w19032 = w18923 & w19031;
assign w19033 = ~w18923 & ~w19031;
assign w19034 = ~w19032 & ~w19033;
assign w19035 = w18913 & ~w19034;
assign w19036 = ~w18913 & w19034;
assign w19037 = ~w19035 & ~w19036;
assign w19038 = b[45] & w5167;
assign w19039 = b[47] & w4925;
assign w19040 = b[46] & w4918;
assign w19041 = w4923 & w6889;
assign w19042 = ~w19039 & ~w19040;
assign w19043 = ~w19038 & w19042;
assign w19044 = ~w19041 & w19043;
assign w19045 = a[41] & ~w19044;
assign w19046 = ~a[41] & w19044;
assign w19047 = ~w19045 & ~w19046;
assign w19048 = w19037 & w19047;
assign w19049 = ~w19037 & ~w19047;
assign w19050 = ~w19048 & ~w19049;
assign w19051 = ~w18785 & ~w18788;
assign w19052 = w19050 & ~w19051;
assign w19053 = ~w19050 & w19051;
assign w19054 = ~w19052 & ~w19053;
assign w19055 = ~w18912 & ~w19054;
assign w19056 = w18912 & w19054;
assign w19057 = ~w19055 & ~w19056;
assign w19058 = w18902 & ~w19057;
assign w19059 = ~w18902 & w19057;
assign w19060 = ~w19058 & ~w19059;
assign w19061 = w18901 & w19060;
assign w19062 = ~w18901 & ~w19060;
assign w19063 = ~w19061 & ~w19062;
assign w19064 = w18891 & w19063;
assign w19065 = ~w18891 & ~w19063;
assign w19066 = ~w19064 & ~w19065;
assign w19067 = b[57] & ~w2622;
assign w19068 = b[58] & w2436;
assign w19069 = b[59] & w2438;
assign w19070 = w2432 & w10371;
assign w19071 = ~w19067 & ~w19068;
assign w19072 = ~w19069 & w19071;
assign w19073 = ~w19070 & w19072;
assign w19074 = a[29] & ~w19073;
assign w19075 = ~a[29] & w19073;
assign w19076 = ~w19074 & ~w19075;
assign w19077 = ~w18816 & ~w18819;
assign w19078 = w19076 & ~w19077;
assign w19079 = ~w19076 & w19077;
assign w19080 = ~w19078 & ~w19079;
assign w19081 = w19066 & w19080;
assign w19082 = ~w19066 & ~w19080;
assign w19083 = ~w19081 & ~w19082;
assign w19084 = w18877 & w19083;
assign w19085 = ~w18877 & ~w19083;
assign w19086 = ~w19084 & ~w19085;
assign w19087 = ~w18629 & ~w18839;
assign w19088 = w1513 & ~w12154;
assign w19089 = w1676 & ~w19088;
assign w19090 = b[63] & ~w19089;
assign w19091 = ~a[23] & ~w19090;
assign w19092 = a[23] & w19090;
assign w19093 = ~w19091 & ~w19092;
assign w19094 = ~w19087 & w19093;
assign w19095 = w19087 & ~w19093;
assign w19096 = ~w19094 & ~w19095;
assign w19097 = w19086 & w19096;
assign w19098 = ~w19086 & ~w19096;
assign w19099 = ~w19097 & ~w19098;
assign w19100 = ~w18863 & w19099;
assign w19101 = w18863 & ~w19099;
assign w19102 = ~w19100 & ~w19101;
assign w19103 = (w18109 & w24445) | (w18109 & w24446) | (w24445 & w24446);
assign w19104 = w19102 & ~w19103;
assign w19105 = ~w19102 & w19103;
assign w19106 = ~w19104 & ~w19105;
assign w19107 = (w18109 & w24447) | (w18109 & w24448) | (w24447 & w24448);
assign w19108 = ~w19094 & ~w19097;
assign w19109 = ~w19059 & ~w19061;
assign w19110 = b[52] & w3785;
assign w19111 = b[54] & w3580;
assign w19112 = b[53] & w3578;
assign w19113 = w3573 & ~w8998;
assign w19114 = ~w19111 & ~w19112;
assign w19115 = ~w19110 & w19114;
assign w19116 = ~w19113 & w19115;
assign w19117 = a[35] & ~w19116;
assign w19118 = ~a[35] & w19116;
assign w19119 = ~w19117 & ~w19118;
assign w19120 = ~w19052 & ~w19056;
assign w19121 = ~w19029 & ~w19032;
assign w19122 = b[43] & w5939;
assign w19123 = b[44] & w5670;
assign w19124 = b[45] & w5665;
assign w19125 = w5663 & w6334;
assign w19126 = ~w19123 & ~w19124;
assign w19127 = ~w19122 & w19126;
assign w19128 = ~w19125 & w19127;
assign w19129 = a[44] & ~w19128;
assign w19130 = ~a[44] & w19128;
assign w19131 = ~w19129 & ~w19130;
assign w19132 = ~w19023 & ~w19026;
assign w19133 = ~w18978 & ~w18990;
assign w19134 = b[28] & w10496;
assign w19135 = b[29] & w10146;
assign w19136 = b[30] & w10148;
assign w19137 = ~w2908 & w10141;
assign w19138 = ~w19135 & ~w19136;
assign w19139 = ~w19134 & w19138;
assign w19140 = ~w19137 & w19139;
assign w19141 = a[59] & ~w19140;
assign w19142 = ~a[59] & w19140;
assign w19143 = ~w19141 & ~w19142;
assign w19144 = ~w18962 & ~w18974;
assign w19145 = b[23] & w11921;
assign w19146 = b[24] & w11923;
assign w19147 = ~w19145 & ~w19146;
assign w19148 = ~a[23] & ~w19147;
assign w19149 = a[23] & w19147;
assign w19150 = ~w19148 & ~w19149;
assign w19151 = ~w18960 & w19150;
assign w19152 = w18960 & ~w19150;
assign w19153 = ~w19151 & ~w19152;
assign w19154 = b[25] & w11561;
assign w19155 = b[26] & w11194;
assign w19156 = b[27] & w11196;
assign w19157 = w2378 & w11189;
assign w19158 = ~w19155 & ~w19156;
assign w19159 = ~w19154 & w19158;
assign w19160 = ~w19157 & w19159;
assign w19161 = a[62] & ~w19160;
assign w19162 = ~a[62] & w19160;
assign w19163 = ~w19161 & ~w19162;
assign w19164 = w19153 & w19163;
assign w19165 = ~w19153 & ~w19163;
assign w19166 = ~w19164 & ~w19165;
assign w19167 = ~w19144 & w19166;
assign w19168 = w19144 & ~w19166;
assign w19169 = ~w19167 & ~w19168;
assign w19170 = w19143 & w19169;
assign w19171 = ~w19143 & ~w19169;
assign w19172 = ~w19170 & ~w19171;
assign w19173 = w19133 & ~w19172;
assign w19174 = ~w19133 & w19172;
assign w19175 = ~w19173 & ~w19174;
assign w19176 = b[31] & w9482;
assign w19177 = b[33] & w9160;
assign w19178 = b[32] & w9165;
assign w19179 = w3499 & w9158;
assign w19180 = ~w19177 & ~w19178;
assign w19181 = ~w19176 & w19180;
assign w19182 = ~w19179 & w19181;
assign w19183 = a[56] & ~w19182;
assign w19184 = ~a[56] & w19182;
assign w19185 = ~w19183 & ~w19184;
assign w19186 = ~w18994 & ~w18998;
assign w19187 = w19185 & ~w19186;
assign w19188 = ~w19185 & w19186;
assign w19189 = ~w19187 & ~w19188;
assign w19190 = w19175 & w19189;
assign w19191 = ~w19175 & ~w19189;
assign w19192 = ~w19190 & ~w19191;
assign w19193 = b[34] & w8515;
assign w19194 = b[36] & w8202;
assign w19195 = b[35] & w8200;
assign w19196 = w4129 & w8195;
assign w19197 = ~w19194 & ~w19195;
assign w19198 = ~w19193 & w19197;
assign w19199 = ~w19196 & w19198;
assign w19200 = a[53] & ~w19199;
assign w19201 = ~a[53] & w19199;
assign w19202 = ~w19200 & ~w19201;
assign w19203 = w19192 & w19202;
assign w19204 = ~w19192 & ~w19202;
assign w19205 = ~w19203 & ~w19204;
assign w19206 = ~w19001 & ~w19003;
assign w19207 = ~w19205 & w19206;
assign w19208 = w19205 & ~w19206;
assign w19209 = ~w19207 & ~w19208;
assign w19210 = b[37] & w7586;
assign w19211 = b[38] & w7307;
assign w19212 = b[39] & w7314;
assign w19213 = ~w4812 & w7312;
assign w19214 = ~w19211 & ~w19212;
assign w19215 = ~w19210 & w19214;
assign w19216 = ~w19213 & w19215;
assign w19217 = a[50] & ~w19216;
assign w19218 = ~a[50] & w19216;
assign w19219 = ~w19217 & ~w19218;
assign w19220 = w19209 & w19219;
assign w19221 = ~w19209 & ~w19219;
assign w19222 = ~w19220 & ~w19221;
assign w19223 = ~w19007 & ~w19019;
assign w19224 = ~w19222 & w19223;
assign w19225 = w19222 & ~w19223;
assign w19226 = ~w19224 & ~w19225;
assign w19227 = b[40] & w6732;
assign w19228 = b[41] & w6474;
assign w19229 = b[42] & w6476;
assign w19230 = w5548 & w6469;
assign w19231 = ~w19228 & ~w19229;
assign w19232 = ~w19227 & w19231;
assign w19233 = ~w19230 & w19232;
assign w19234 = a[47] & ~w19233;
assign w19235 = ~a[47] & w19233;
assign w19236 = ~w19234 & ~w19235;
assign w19237 = w19226 & w19236;
assign w19238 = ~w19226 & ~w19236;
assign w19239 = ~w19237 & ~w19238;
assign w19240 = ~w19132 & w19239;
assign w19241 = w19132 & ~w19239;
assign w19242 = ~w19240 & ~w19241;
assign w19243 = w19131 & w19242;
assign w19244 = ~w19131 & ~w19242;
assign w19245 = ~w19243 & ~w19244;
assign w19246 = w19121 & ~w19245;
assign w19247 = ~w19121 & w19245;
assign w19248 = ~w19246 & ~w19247;
assign w19249 = b[46] & w5167;
assign w19250 = b[47] & w4918;
assign w19251 = b[48] & w4925;
assign w19252 = w4923 & ~w7170;
assign w19253 = ~w19250 & ~w19251;
assign w19254 = ~w19249 & w19253;
assign w19255 = ~w19252 & w19254;
assign w19256 = a[41] & ~w19255;
assign w19257 = ~a[41] & w19255;
assign w19258 = ~w19256 & ~w19257;
assign w19259 = w19248 & w19258;
assign w19260 = ~w19248 & ~w19258;
assign w19261 = ~w19259 & ~w19260;
assign w19262 = ~w19036 & ~w19048;
assign w19263 = ~w19261 & w19262;
assign w19264 = w19261 & ~w19262;
assign w19265 = ~w19263 & ~w19264;
assign w19266 = b[49] & w4453;
assign w19267 = b[51] & w4243;
assign w19268 = b[50] & w4241;
assign w19269 = w4236 & ~w8058;
assign w19270 = ~w19267 & ~w19268;
assign w19271 = ~w19266 & w19270;
assign w19272 = ~w19269 & w19271;
assign w19273 = a[38] & ~w19272;
assign w19274 = ~a[38] & w19272;
assign w19275 = ~w19273 & ~w19274;
assign w19276 = ~w19265 & ~w19275;
assign w19277 = w19265 & w19275;
assign w19278 = ~w19276 & ~w19277;
assign w19279 = w19120 & w19278;
assign w19280 = ~w19120 & ~w19278;
assign w19281 = ~w19279 & ~w19280;
assign w19282 = w19119 & ~w19281;
assign w19283 = ~w19119 & w19281;
assign w19284 = ~w19282 & ~w19283;
assign w19285 = ~w19109 & w19284;
assign w19286 = w19109 & ~w19284;
assign w19287 = ~w19285 & ~w19286;
assign w19288 = b[55] & w3177;
assign w19289 = b[57] & w2978;
assign w19290 = b[56] & w2973;
assign w19291 = w2980 & ~w9992;
assign w19292 = ~w19289 & ~w19290;
assign w19293 = ~w19288 & w19292;
assign w19294 = ~w19291 & w19293;
assign w19295 = a[32] & ~w19294;
assign w19296 = ~a[32] & w19294;
assign w19297 = ~w19295 & ~w19296;
assign w19298 = ~w18889 & ~w19064;
assign w19299 = w19297 & ~w19298;
assign w19300 = ~w19297 & w19298;
assign w19301 = ~w19299 & ~w19300;
assign w19302 = w19287 & w19301;
assign w19303 = ~w19287 & ~w19301;
assign w19304 = ~w19302 & ~w19303;
assign w19305 = ~w19078 & ~w19081;
assign w19306 = b[58] & ~w2622;
assign w19307 = b[60] & w2438;
assign w19308 = b[59] & w2436;
assign w19309 = w2432 & w11035;
assign w19310 = ~w19306 & ~w19307;
assign w19311 = ~w19308 & w19310;
assign w19312 = ~w19309 & w19311;
assign w19313 = a[29] & ~w19312;
assign w19314 = ~a[29] & w19312;
assign w19315 = ~w19313 & ~w19314;
assign w19316 = ~w19305 & w19315;
assign w19317 = w19305 & ~w19315;
assign w19318 = ~w19316 & ~w19317;
assign w19319 = ~w19304 & ~w19318;
assign w19320 = w19304 & w19318;
assign w19321 = ~w19319 & ~w19320;
assign w19322 = ~w18875 & ~w19084;
assign w19323 = b[62] & w1955;
assign w19324 = b[61] & ~w2114;
assign w19325 = b[63] & w1957;
assign w19326 = w1951 & w12132;
assign w19327 = ~w19323 & ~w19324;
assign w19328 = ~w19325 & w19327;
assign w19329 = ~w19326 & w19328;
assign w19330 = a[26] & ~w19329;
assign w19331 = ~a[26] & w19329;
assign w19332 = ~w19330 & ~w19331;
assign w19333 = ~w19322 & w19332;
assign w19334 = w19322 & ~w19332;
assign w19335 = ~w19333 & ~w19334;
assign w19336 = w19321 & w19335;
assign w19337 = ~w19321 & ~w19335;
assign w19338 = ~w19336 & ~w19337;
assign w19339 = ~w19108 & w19338;
assign w19340 = w19108 & ~w19338;
assign w19341 = ~w19339 & ~w19340;
assign w19342 = ~w19107 & ~w19341;
assign w19343 = (w18109 & w24449) | (w18109 & w24450) | (w24449 & w24450);
assign w19344 = ~w19342 & ~w19343;
assign w19345 = ~w19333 & ~w19336;
assign w19346 = b[53] & w3785;
assign w19347 = b[54] & w3578;
assign w19348 = b[55] & w3580;
assign w19349 = w3573 & ~w9330;
assign w19350 = ~w19347 & ~w19348;
assign w19351 = ~w19346 & w19350;
assign w19352 = ~w19349 & w19351;
assign w19353 = a[35] & ~w19352;
assign w19354 = ~a[35] & w19352;
assign w19355 = ~w19353 & ~w19354;
assign w19356 = b[50] & w4453;
assign w19357 = b[51] & w4241;
assign w19358 = b[52] & w4243;
assign w19359 = w4236 & ~w8371;
assign w19360 = ~w19357 & ~w19358;
assign w19361 = ~w19356 & w19360;
assign w19362 = ~w19359 & w19361;
assign w19363 = a[38] & ~w19362;
assign w19364 = ~a[38] & w19362;
assign w19365 = ~w19363 & ~w19364;
assign w19366 = b[47] & w5167;
assign w19367 = b[48] & w4918;
assign w19368 = b[49] & w4925;
assign w19369 = w4923 & ~w7468;
assign w19370 = ~w19367 & ~w19368;
assign w19371 = ~w19366 & w19370;
assign w19372 = ~w19369 & w19371;
assign w19373 = a[41] & ~w19372;
assign w19374 = ~a[41] & w19372;
assign w19375 = ~w19373 & ~w19374;
assign w19376 = b[44] & w5939;
assign w19377 = b[45] & w5670;
assign w19378 = b[46] & w5665;
assign w19379 = w5663 & ~w6613;
assign w19380 = ~w19377 & ~w19378;
assign w19381 = ~w19376 & w19380;
assign w19382 = ~w19379 & w19381;
assign w19383 = a[44] & ~w19382;
assign w19384 = ~a[44] & w19382;
assign w19385 = ~w19383 & ~w19384;
assign w19386 = ~w19220 & ~w19225;
assign w19387 = b[38] & w7586;
assign w19388 = b[40] & w7314;
assign w19389 = b[39] & w7307;
assign w19390 = ~w5058 & w7312;
assign w19391 = ~w19388 & ~w19389;
assign w19392 = ~w19387 & w19391;
assign w19393 = ~w19390 & w19392;
assign w19394 = a[50] & ~w19393;
assign w19395 = ~a[50] & w19393;
assign w19396 = ~w19394 & ~w19395;
assign w19397 = ~w19203 & ~w19208;
assign w19398 = b[35] & w8515;
assign w19399 = b[36] & w8200;
assign w19400 = b[37] & w8202;
assign w19401 = ~w4357 & w8195;
assign w19402 = ~w19399 & ~w19400;
assign w19403 = ~w19398 & w19402;
assign w19404 = ~w19401 & w19403;
assign w19405 = a[53] & ~w19404;
assign w19406 = ~a[53] & w19404;
assign w19407 = ~w19405 & ~w19406;
assign w19408 = b[32] & w9482;
assign w19409 = b[33] & w9165;
assign w19410 = b[34] & w9160;
assign w19411 = ~w3710 & w9158;
assign w19412 = ~w19409 & ~w19410;
assign w19413 = ~w19408 & w19412;
assign w19414 = ~w19411 & w19413;
assign w19415 = a[56] & ~w19414;
assign w19416 = ~a[56] & w19414;
assign w19417 = ~w19415 & ~w19416;
assign w19418 = ~w19164 & ~w19167;
assign w19419 = b[24] & w11921;
assign w19420 = b[25] & w11923;
assign w19421 = ~w19419 & ~w19420;
assign w19422 = ~w19148 & ~w19151;
assign w19423 = w19421 & ~w19422;
assign w19424 = ~w19421 & w19422;
assign w19425 = ~w19423 & ~w19424;
assign w19426 = b[26] & w11561;
assign w19427 = b[27] & w11194;
assign w19428 = b[28] & w11196;
assign w19429 = w2559 & w11189;
assign w19430 = ~w19427 & ~w19428;
assign w19431 = ~w19426 & w19430;
assign w19432 = ~w19429 & w19431;
assign w19433 = a[62] & ~w19432;
assign w19434 = ~a[62] & w19432;
assign w19435 = ~w19433 & ~w19434;
assign w19436 = w19425 & w19435;
assign w19437 = ~w19425 & ~w19435;
assign w19438 = ~w19436 & ~w19437;
assign w19439 = w19418 & ~w19438;
assign w19440 = ~w19418 & w19438;
assign w19441 = ~w19439 & ~w19440;
assign w19442 = b[29] & w10496;
assign w19443 = b[30] & w10146;
assign w19444 = b[31] & w10148;
assign w19445 = ~w3112 & w10141;
assign w19446 = ~w19443 & ~w19444;
assign w19447 = ~w19442 & w19446;
assign w19448 = ~w19445 & w19447;
assign w19449 = a[59] & ~w19448;
assign w19450 = ~a[59] & w19448;
assign w19451 = ~w19449 & ~w19450;
assign w19452 = w19441 & w19451;
assign w19453 = ~w19441 & ~w19451;
assign w19454 = ~w19452 & ~w19453;
assign w19455 = ~w19170 & ~w19174;
assign w19456 = w19454 & ~w19455;
assign w19457 = ~w19454 & w19455;
assign w19458 = ~w19456 & ~w19457;
assign w19459 = w19417 & w19458;
assign w19460 = ~w19417 & ~w19458;
assign w19461 = ~w19459 & ~w19460;
assign w19462 = ~w19187 & ~w19190;
assign w19463 = w19461 & ~w19462;
assign w19464 = ~w19461 & w19462;
assign w19465 = ~w19463 & ~w19464;
assign w19466 = ~w19407 & ~w19465;
assign w19467 = w19407 & w19465;
assign w19468 = ~w19466 & ~w19467;
assign w19469 = w19397 & ~w19468;
assign w19470 = ~w19397 & w19468;
assign w19471 = ~w19469 & ~w19470;
assign w19472 = w19396 & w19471;
assign w19473 = ~w19396 & ~w19471;
assign w19474 = ~w19472 & ~w19473;
assign w19475 = w19386 & ~w19474;
assign w19476 = ~w19386 & w19474;
assign w19477 = ~w19475 & ~w19476;
assign w19478 = b[41] & w6732;
assign w19479 = b[42] & w6474;
assign w19480 = b[43] & w6476;
assign w19481 = w5811 & w6469;
assign w19482 = ~w19479 & ~w19480;
assign w19483 = ~w19478 & w19482;
assign w19484 = ~w19481 & w19483;
assign w19485 = a[47] & ~w19484;
assign w19486 = ~a[47] & w19484;
assign w19487 = ~w19485 & ~w19486;
assign w19488 = w19477 & w19487;
assign w19489 = ~w19477 & ~w19487;
assign w19490 = ~w19488 & ~w19489;
assign w19491 = ~w19237 & ~w19240;
assign w19492 = w19490 & ~w19491;
assign w19493 = ~w19490 & w19491;
assign w19494 = ~w19492 & ~w19493;
assign w19495 = w19385 & w19494;
assign w19496 = ~w19385 & ~w19494;
assign w19497 = ~w19495 & ~w19496;
assign w19498 = ~w19243 & ~w19247;
assign w19499 = w19497 & ~w19498;
assign w19500 = ~w19497 & w19498;
assign w19501 = ~w19499 & ~w19500;
assign w19502 = w19375 & w19501;
assign w19503 = ~w19375 & ~w19501;
assign w19504 = ~w19502 & ~w19503;
assign w19505 = ~w19259 & ~w19264;
assign w19506 = w19504 & ~w19505;
assign w19507 = ~w19504 & w19505;
assign w19508 = ~w19506 & ~w19507;
assign w19509 = w19365 & w19508;
assign w19510 = ~w19365 & ~w19508;
assign w19511 = ~w19509 & ~w19510;
assign w19512 = ~w19276 & ~w19279;
assign w19513 = w19511 & w19512;
assign w19514 = ~w19511 & ~w19512;
assign w19515 = ~w19513 & ~w19514;
assign w19516 = w19355 & w19515;
assign w19517 = ~w19355 & ~w19515;
assign w19518 = ~w19516 & ~w19517;
assign w19519 = ~w19282 & ~w19285;
assign w19520 = b[56] & w3177;
assign w19521 = b[57] & w2973;
assign w19522 = b[58] & w2978;
assign w19523 = w2980 & ~w10339;
assign w19524 = ~w19521 & ~w19522;
assign w19525 = ~w19520 & w19524;
assign w19526 = ~w19523 & w19525;
assign w19527 = a[32] & ~w19526;
assign w19528 = ~a[32] & w19526;
assign w19529 = ~w19527 & ~w19528;
assign w19530 = ~w19519 & w19529;
assign w19531 = w19519 & ~w19529;
assign w19532 = ~w19530 & ~w19531;
assign w19533 = w19518 & w19532;
assign w19534 = ~w19518 & ~w19532;
assign w19535 = ~w19533 & ~w19534;
assign w19536 = b[59] & ~w2622;
assign w19537 = b[61] & w2438;
assign w19538 = b[60] & w2436;
assign w19539 = w2432 & w11400;
assign w19540 = ~w19536 & ~w19537;
assign w19541 = ~w19538 & w19540;
assign w19542 = ~w19539 & w19541;
assign w19543 = a[29] & ~w19542;
assign w19544 = ~a[29] & w19542;
assign w19545 = ~w19543 & ~w19544;
assign w19546 = ~w19299 & ~w19302;
assign w19547 = w19545 & ~w19546;
assign w19548 = ~w19545 & w19546;
assign w19549 = ~w19547 & ~w19548;
assign w19550 = ~w19535 & ~w19549;
assign w19551 = w19535 & w19549;
assign w19552 = ~w19550 & ~w19551;
assign w19553 = ~w19316 & ~w19320;
assign w19554 = b[62] & ~w2114;
assign w19555 = b[63] & w1955;
assign w19556 = w1951 & w12156;
assign w19557 = ~w19554 & ~w19555;
assign w19558 = ~w19556 & w19557;
assign w19559 = a[26] & ~w19558;
assign w19560 = ~a[26] & w19558;
assign w19561 = ~w19559 & ~w19560;
assign w19562 = ~w19553 & w19561;
assign w19563 = w19553 & ~w19561;
assign w19564 = ~w19562 & ~w19563;
assign w19565 = w19552 & w19564;
assign w19566 = ~w19552 & ~w19564;
assign w19567 = ~w19565 & ~w19566;
assign w19568 = w19345 & ~w19567;
assign w19569 = ~w19345 & w19567;
assign w19570 = ~w19568 & ~w19569;
assign w19571 = (~w18109 & w24451) | (~w18109 & w24452) | (w24451 & w24452);
assign w19572 = w19570 & w19571;
assign w19573 = ~w19570 & ~w19571;
assign w19574 = ~w19572 & ~w19573;
assign w19575 = ~w19562 & ~w19565;
assign w19576 = b[54] & w3785;
assign w19577 = b[55] & w3578;
assign w19578 = b[56] & w3580;
assign w19579 = w3573 & w9657;
assign w19580 = ~w19577 & ~w19578;
assign w19581 = ~w19576 & w19580;
assign w19582 = ~w19579 & w19581;
assign w19583 = a[35] & ~w19582;
assign w19584 = ~a[35] & w19582;
assign w19585 = ~w19583 & ~w19584;
assign w19586 = ~w19506 & ~w19509;
assign w19587 = b[51] & w4453;
assign w19588 = b[53] & w4243;
assign w19589 = b[52] & w4241;
assign w19590 = w4236 & w8683;
assign w19591 = ~w19588 & ~w19589;
assign w19592 = ~w19587 & w19591;
assign w19593 = ~w19590 & w19592;
assign w19594 = a[38] & ~w19593;
assign w19595 = ~a[38] & w19593;
assign w19596 = ~w19594 & ~w19595;
assign w19597 = ~w19499 & ~w19502;
assign w19598 = b[48] & w5167;
assign w19599 = b[49] & w4918;
assign w19600 = b[50] & w4925;
assign w19601 = w4923 & w7759;
assign w19602 = ~w19599 & ~w19600;
assign w19603 = ~w19598 & w19602;
assign w19604 = ~w19601 & w19603;
assign w19605 = a[41] & ~w19604;
assign w19606 = ~a[41] & w19604;
assign w19607 = ~w19605 & ~w19606;
assign w19608 = ~w19476 & ~w19488;
assign w19609 = b[42] & w6732;
assign w19610 = b[43] & w6474;
assign w19611 = b[44] & w6476;
assign w19612 = w6069 & w6469;
assign w19613 = ~w19610 & ~w19611;
assign w19614 = ~w19609 & w19613;
assign w19615 = ~w19612 & w19614;
assign w19616 = a[47] & ~w19615;
assign w19617 = ~a[47] & w19615;
assign w19618 = ~w19616 & ~w19617;
assign w19619 = ~w19470 & ~w19472;
assign w19620 = b[39] & w7586;
assign w19621 = b[40] & w7307;
assign w19622 = b[41] & w7314;
assign w19623 = w5302 & w7312;
assign w19624 = ~w19621 & ~w19622;
assign w19625 = ~w19620 & w19624;
assign w19626 = ~w19623 & w19625;
assign w19627 = a[50] & ~w19626;
assign w19628 = ~a[50] & w19626;
assign w19629 = ~w19627 & ~w19628;
assign w19630 = ~w19456 & ~w19459;
assign w19631 = b[33] & w9482;
assign w19632 = b[35] & w9160;
assign w19633 = b[34] & w9165;
assign w19634 = w3918 & w9158;
assign w19635 = ~w19632 & ~w19633;
assign w19636 = ~w19631 & w19635;
assign w19637 = ~w19634 & w19636;
assign w19638 = a[56] & ~w19637;
assign w19639 = ~a[56] & w19637;
assign w19640 = ~w19638 & ~w19639;
assign w19641 = ~w19440 & ~w19452;
assign w19642 = b[30] & w10496;
assign w19643 = b[31] & w10146;
assign w19644 = b[32] & w10148;
assign w19645 = w3304 & w10141;
assign w19646 = ~w19643 & ~w19644;
assign w19647 = ~w19642 & w19646;
assign w19648 = ~w19645 & w19647;
assign w19649 = a[59] & ~w19648;
assign w19650 = ~a[59] & w19648;
assign w19651 = ~w19649 & ~w19650;
assign w19652 = ~w19423 & ~w19436;
assign w19653 = b[25] & w11921;
assign w19654 = b[26] & w11923;
assign w19655 = ~w19653 & ~w19654;
assign w19656 = w19421 & ~w19655;
assign w19657 = ~w19421 & w19655;
assign w19658 = ~w19656 & ~w19657;
assign w19659 = b[27] & w11561;
assign w19660 = b[29] & w11196;
assign w19661 = b[28] & w11194;
assign w19662 = w2734 & w11189;
assign w19663 = ~w19660 & ~w19661;
assign w19664 = ~w19659 & w19663;
assign w19665 = ~w19662 & w19664;
assign w19666 = a[62] & ~w19665;
assign w19667 = ~a[62] & w19665;
assign w19668 = ~w19666 & ~w19667;
assign w19669 = w19658 & w19668;
assign w19670 = ~w19658 & ~w19668;
assign w19671 = ~w19669 & ~w19670;
assign w19672 = w19652 & ~w19671;
assign w19673 = ~w19652 & w19671;
assign w19674 = ~w19672 & ~w19673;
assign w19675 = w19651 & w19674;
assign w19676 = ~w19651 & ~w19674;
assign w19677 = ~w19675 & ~w19676;
assign w19678 = w19641 & ~w19677;
assign w19679 = ~w19641 & w19677;
assign w19680 = ~w19678 & ~w19679;
assign w19681 = w19640 & w19680;
assign w19682 = ~w19640 & ~w19680;
assign w19683 = ~w19681 & ~w19682;
assign w19684 = w19630 & ~w19683;
assign w19685 = ~w19630 & w19683;
assign w19686 = ~w19684 & ~w19685;
assign w19687 = b[36] & w8515;
assign w19688 = b[37] & w8200;
assign w19689 = b[38] & w8202;
assign w19690 = w4582 & w8195;
assign w19691 = ~w19688 & ~w19689;
assign w19692 = ~w19687 & w19691;
assign w19693 = ~w19690 & w19692;
assign w19694 = a[53] & ~w19693;
assign w19695 = ~a[53] & w19693;
assign w19696 = ~w19694 & ~w19695;
assign w19697 = w19686 & w19696;
assign w19698 = ~w19686 & ~w19696;
assign w19699 = ~w19697 & ~w19698;
assign w19700 = ~w19463 & ~w19467;
assign w19701 = w19699 & ~w19700;
assign w19702 = ~w19699 & w19700;
assign w19703 = ~w19701 & ~w19702;
assign w19704 = w19629 & w19703;
assign w19705 = ~w19629 & ~w19703;
assign w19706 = ~w19704 & ~w19705;
assign w19707 = ~w19619 & w19706;
assign w19708 = w19619 & ~w19706;
assign w19709 = ~w19707 & ~w19708;
assign w19710 = w19618 & w19709;
assign w19711 = ~w19618 & ~w19709;
assign w19712 = ~w19710 & ~w19711;
assign w19713 = w19608 & ~w19712;
assign w19714 = ~w19608 & w19712;
assign w19715 = ~w19713 & ~w19714;
assign w19716 = b[45] & w5939;
assign w19717 = b[47] & w5665;
assign w19718 = b[46] & w5670;
assign w19719 = w5663 & w6889;
assign w19720 = ~w19717 & ~w19718;
assign w19721 = ~w19716 & w19720;
assign w19722 = ~w19719 & w19721;
assign w19723 = a[44] & ~w19722;
assign w19724 = ~a[44] & w19722;
assign w19725 = ~w19723 & ~w19724;
assign w19726 = w19715 & w19725;
assign w19727 = ~w19715 & ~w19725;
assign w19728 = ~w19726 & ~w19727;
assign w19729 = ~w19492 & ~w19495;
assign w19730 = w19728 & ~w19729;
assign w19731 = ~w19728 & w19729;
assign w19732 = ~w19730 & ~w19731;
assign w19733 = ~w19607 & ~w19732;
assign w19734 = w19607 & w19732;
assign w19735 = ~w19733 & ~w19734;
assign w19736 = w19597 & ~w19735;
assign w19737 = ~w19597 & w19735;
assign w19738 = ~w19736 & ~w19737;
assign w19739 = w19596 & w19738;
assign w19740 = ~w19596 & ~w19738;
assign w19741 = ~w19739 & ~w19740;
assign w19742 = w19586 & ~w19741;
assign w19743 = ~w19586 & w19741;
assign w19744 = ~w19742 & ~w19743;
assign w19745 = ~w19585 & ~w19744;
assign w19746 = w19585 & w19744;
assign w19747 = ~w19745 & ~w19746;
assign w19748 = b[57] & w3177;
assign w19749 = b[58] & w2973;
assign w19750 = b[59] & w2978;
assign w19751 = w2980 & w10371;
assign w19752 = ~w19749 & ~w19750;
assign w19753 = ~w19748 & w19752;
assign w19754 = ~w19751 & w19753;
assign w19755 = a[32] & ~w19754;
assign w19756 = ~a[32] & w19754;
assign w19757 = ~w19755 & ~w19756;
assign w19758 = ~w19513 & ~w19516;
assign w19759 = w19757 & ~w19758;
assign w19760 = ~w19757 & w19758;
assign w19761 = ~w19759 & ~w19760;
assign w19762 = w19747 & w19761;
assign w19763 = ~w19747 & ~w19761;
assign w19764 = ~w19762 & ~w19763;
assign w19765 = b[60] & ~w2622;
assign w19766 = b[61] & w2436;
assign w19767 = b[62] & w2438;
assign w19768 = w2432 & w11763;
assign w19769 = ~w19765 & ~w19766;
assign w19770 = ~w19767 & w19769;
assign w19771 = ~w19768 & w19770;
assign w19772 = a[29] & ~w19771;
assign w19773 = ~a[29] & w19771;
assign w19774 = ~w19772 & ~w19773;
assign w19775 = ~w19530 & ~w19533;
assign w19776 = w19774 & ~w19775;
assign w19777 = ~w19774 & w19775;
assign w19778 = ~w19776 & ~w19777;
assign w19779 = ~w19764 & ~w19778;
assign w19780 = w19764 & w19778;
assign w19781 = ~w19779 & ~w19780;
assign w19782 = ~w19547 & ~w19551;
assign w19783 = w1951 & ~w12154;
assign w19784 = w2114 & ~w19783;
assign w19785 = b[63] & ~w19784;
assign w19786 = ~a[26] & ~w19785;
assign w19787 = a[26] & w19785;
assign w19788 = ~w19786 & ~w19787;
assign w19789 = ~w19782 & w19788;
assign w19790 = w19782 & ~w19788;
assign w19791 = ~w19789 & ~w19790;
assign w19792 = w19781 & w19791;
assign w19793 = ~w19781 & ~w19791;
assign w19794 = ~w19792 & ~w19793;
assign w19795 = ~w19575 & w19794;
assign w19796 = w19575 & ~w19794;
assign w19797 = ~w19795 & ~w19796;
assign w19798 = (w18109 & w24455) | (w18109 & w24456) | (w24455 & w24456);
assign w19799 = w19797 & ~w19798;
assign w19800 = ~w19797 & w19798;
assign w19801 = ~w19799 & ~w19800;
assign w19802 = ~w19789 & ~w19792;
assign w19803 = ~w19776 & ~w19780;
assign w19804 = b[61] & ~w2622;
assign w19805 = b[63] & w2438;
assign w19806 = b[62] & w2436;
assign w19807 = w2432 & w12132;
assign w19808 = ~w19804 & ~w19805;
assign w19809 = ~w19806 & w19808;
assign w19810 = ~w19807 & w19809;
assign w19811 = a[29] & ~w19810;
assign w19812 = ~a[29] & w19810;
assign w19813 = ~w19811 & ~w19812;
assign w19814 = ~w19803 & w19813;
assign w19815 = w19803 & ~w19813;
assign w19816 = ~w19814 & ~w19815;
assign w19817 = ~w19737 & ~w19739;
assign w19818 = b[52] & w4453;
assign w19819 = b[54] & w4243;
assign w19820 = b[53] & w4241;
assign w19821 = w4236 & ~w8998;
assign w19822 = ~w19819 & ~w19820;
assign w19823 = ~w19818 & w19822;
assign w19824 = ~w19821 & w19823;
assign w19825 = a[38] & ~w19824;
assign w19826 = ~a[38] & w19824;
assign w19827 = ~w19825 & ~w19826;
assign w19828 = ~w19730 & ~w19734;
assign w19829 = ~w19707 & ~w19710;
assign w19830 = b[43] & w6732;
assign w19831 = b[44] & w6474;
assign w19832 = b[45] & w6476;
assign w19833 = w6334 & w6469;
assign w19834 = ~w19831 & ~w19832;
assign w19835 = ~w19830 & w19834;
assign w19836 = ~w19833 & w19835;
assign w19837 = a[47] & ~w19836;
assign w19838 = ~a[47] & w19836;
assign w19839 = ~w19837 & ~w19838;
assign w19840 = ~w19701 & ~w19704;
assign w19841 = ~w19657 & ~w19669;
assign w19842 = b[26] & w11921;
assign w19843 = b[27] & w11923;
assign w19844 = ~w19842 & ~w19843;
assign w19845 = ~a[26] & ~w19844;
assign w19846 = a[26] & w19844;
assign w19847 = ~w19845 & ~w19846;
assign w19848 = ~w19655 & w19847;
assign w19849 = w19655 & ~w19847;
assign w19850 = ~w19848 & ~w19849;
assign w19851 = w19841 & ~w19850;
assign w19852 = ~w19841 & w19850;
assign w19853 = ~w19851 & ~w19852;
assign w19854 = b[28] & w11561;
assign w19855 = b[30] & w11196;
assign w19856 = b[29] & w11194;
assign w19857 = ~w2908 & w11189;
assign w19858 = ~w19855 & ~w19856;
assign w19859 = ~w19854 & w19858;
assign w19860 = ~w19857 & w19859;
assign w19861 = a[62] & ~w19860;
assign w19862 = ~a[62] & w19860;
assign w19863 = ~w19861 & ~w19862;
assign w19864 = w19853 & w19863;
assign w19865 = ~w19853 & ~w19863;
assign w19866 = ~w19864 & ~w19865;
assign w19867 = b[31] & w10496;
assign w19868 = b[33] & w10148;
assign w19869 = b[32] & w10146;
assign w19870 = w3499 & w10141;
assign w19871 = ~w19868 & ~w19869;
assign w19872 = ~w19867 & w19871;
assign w19873 = ~w19870 & w19872;
assign w19874 = a[59] & ~w19873;
assign w19875 = ~a[59] & w19873;
assign w19876 = ~w19874 & ~w19875;
assign w19877 = ~w19673 & ~w19675;
assign w19878 = w19876 & ~w19877;
assign w19879 = ~w19876 & w19877;
assign w19880 = ~w19878 & ~w19879;
assign w19881 = ~w19866 & ~w19880;
assign w19882 = w19866 & w19880;
assign w19883 = ~w19881 & ~w19882;
assign w19884 = b[34] & w9482;
assign w19885 = b[36] & w9160;
assign w19886 = b[35] & w9165;
assign w19887 = w4129 & w9158;
assign w19888 = ~w19885 & ~w19886;
assign w19889 = ~w19884 & w19888;
assign w19890 = ~w19887 & w19889;
assign w19891 = a[56] & ~w19890;
assign w19892 = ~a[56] & w19890;
assign w19893 = ~w19891 & ~w19892;
assign w19894 = w19883 & w19893;
assign w19895 = ~w19883 & ~w19893;
assign w19896 = ~w19894 & ~w19895;
assign w19897 = ~w19679 & ~w19681;
assign w19898 = ~w19896 & w19897;
assign w19899 = w19896 & ~w19897;
assign w19900 = ~w19898 & ~w19899;
assign w19901 = b[37] & w8515;
assign w19902 = b[38] & w8200;
assign w19903 = b[39] & w8202;
assign w19904 = ~w4812 & w8195;
assign w19905 = ~w19902 & ~w19903;
assign w19906 = ~w19901 & w19905;
assign w19907 = ~w19904 & w19906;
assign w19908 = a[53] & ~w19907;
assign w19909 = ~a[53] & w19907;
assign w19910 = ~w19908 & ~w19909;
assign w19911 = w19900 & w19910;
assign w19912 = ~w19900 & ~w19910;
assign w19913 = ~w19911 & ~w19912;
assign w19914 = ~w19685 & ~w19697;
assign w19915 = ~w19913 & w19914;
assign w19916 = w19913 & ~w19914;
assign w19917 = ~w19915 & ~w19916;
assign w19918 = b[40] & w7586;
assign w19919 = b[41] & w7307;
assign w19920 = b[42] & w7314;
assign w19921 = w5548 & w7312;
assign w19922 = ~w19919 & ~w19920;
assign w19923 = ~w19918 & w19922;
assign w19924 = ~w19921 & w19923;
assign w19925 = a[50] & ~w19924;
assign w19926 = ~a[50] & w19924;
assign w19927 = ~w19925 & ~w19926;
assign w19928 = w19917 & w19927;
assign w19929 = ~w19917 & ~w19927;
assign w19930 = ~w19928 & ~w19929;
assign w19931 = ~w19840 & w19930;
assign w19932 = w19840 & ~w19930;
assign w19933 = ~w19931 & ~w19932;
assign w19934 = w19839 & w19933;
assign w19935 = ~w19839 & ~w19933;
assign w19936 = ~w19934 & ~w19935;
assign w19937 = w19829 & ~w19936;
assign w19938 = ~w19829 & w19936;
assign w19939 = ~w19937 & ~w19938;
assign w19940 = b[46] & w5939;
assign w19941 = b[47] & w5670;
assign w19942 = b[48] & w5665;
assign w19943 = w5663 & ~w7170;
assign w19944 = ~w19941 & ~w19942;
assign w19945 = ~w19940 & w19944;
assign w19946 = ~w19943 & w19945;
assign w19947 = a[44] & ~w19946;
assign w19948 = ~a[44] & w19946;
assign w19949 = ~w19947 & ~w19948;
assign w19950 = w19939 & w19949;
assign w19951 = ~w19939 & ~w19949;
assign w19952 = ~w19950 & ~w19951;
assign w19953 = ~w19714 & ~w19726;
assign w19954 = ~w19952 & w19953;
assign w19955 = w19952 & ~w19953;
assign w19956 = ~w19954 & ~w19955;
assign w19957 = b[49] & w5167;
assign w19958 = b[50] & w4918;
assign w19959 = b[51] & w4925;
assign w19960 = w4923 & ~w8058;
assign w19961 = ~w19958 & ~w19959;
assign w19962 = ~w19957 & w19961;
assign w19963 = ~w19960 & w19962;
assign w19964 = a[41] & ~w19963;
assign w19965 = ~a[41] & w19963;
assign w19966 = ~w19964 & ~w19965;
assign w19967 = ~w19956 & ~w19966;
assign w19968 = w19956 & w19966;
assign w19969 = ~w19967 & ~w19968;
assign w19970 = w19828 & w19969;
assign w19971 = ~w19828 & ~w19969;
assign w19972 = ~w19970 & ~w19971;
assign w19973 = w19827 & ~w19972;
assign w19974 = ~w19827 & w19972;
assign w19975 = ~w19973 & ~w19974;
assign w19976 = ~w19817 & w19975;
assign w19977 = w19817 & ~w19975;
assign w19978 = ~w19976 & ~w19977;
assign w19979 = b[55] & w3785;
assign w19980 = b[56] & w3578;
assign w19981 = b[57] & w3580;
assign w19982 = w3573 & ~w9992;
assign w19983 = ~w19980 & ~w19981;
assign w19984 = ~w19979 & w19983;
assign w19985 = ~w19982 & w19984;
assign w19986 = a[35] & ~w19985;
assign w19987 = ~a[35] & w19985;
assign w19988 = ~w19986 & ~w19987;
assign w19989 = w19978 & w19988;
assign w19990 = ~w19978 & ~w19988;
assign w19991 = ~w19989 & ~w19990;
assign w19992 = ~w19743 & ~w19746;
assign w19993 = ~w19991 & w19992;
assign w19994 = w19991 & ~w19992;
assign w19995 = ~w19993 & ~w19994;
assign w19996 = b[58] & w3177;
assign w19997 = b[60] & w2978;
assign w19998 = b[59] & w2973;
assign w19999 = w2980 & w11035;
assign w20000 = ~w19997 & ~w19998;
assign w20001 = ~w19996 & w20000;
assign w20002 = ~w19999 & w20001;
assign w20003 = a[32] & ~w20002;
assign w20004 = ~a[32] & w20002;
assign w20005 = ~w20003 & ~w20004;
assign w20006 = ~w19759 & ~w19762;
assign w20007 = w20005 & ~w20006;
assign w20008 = ~w20005 & w20006;
assign w20009 = ~w20007 & ~w20008;
assign w20010 = w19995 & w20009;
assign w20011 = ~w19995 & ~w20009;
assign w20012 = ~w20010 & ~w20011;
assign w20013 = w19816 & w20012;
assign w20014 = ~w19816 & ~w20012;
assign w20015 = ~w20013 & ~w20014;
assign w20016 = w19802 & ~w20015;
assign w20017 = ~w19802 & w20015;
assign w20018 = ~w20016 & ~w20017;
assign w20019 = (w18109 & w24459) | (w18109 & w24460) | (w24459 & w24460);
assign w20020 = ~w20018 & w20019;
assign w20021 = (~w16450 & w25671) | (~w16450 & w25672) | (w25671 & w25672);
assign w20022 = ~w20020 & ~w20021;
assign w20023 = ~w19814 & ~w20013;
assign w20024 = ~w19973 & ~w19976;
assign w20025 = b[53] & w4453;
assign w20026 = b[54] & w4241;
assign w20027 = b[55] & w4243;
assign w20028 = w4236 & ~w9330;
assign w20029 = ~w20026 & ~w20027;
assign w20030 = ~w20025 & w20029;
assign w20031 = ~w20028 & w20030;
assign w20032 = a[38] & ~w20031;
assign w20033 = ~a[38] & w20031;
assign w20034 = ~w20032 & ~w20033;
assign w20035 = b[50] & w5167;
assign w20036 = b[52] & w4925;
assign w20037 = b[51] & w4918;
assign w20038 = w4923 & ~w8371;
assign w20039 = ~w20036 & ~w20037;
assign w20040 = ~w20035 & w20039;
assign w20041 = ~w20038 & w20040;
assign w20042 = a[41] & ~w20041;
assign w20043 = ~a[41] & w20041;
assign w20044 = ~w20042 & ~w20043;
assign w20045 = b[47] & w5939;
assign w20046 = b[48] & w5670;
assign w20047 = b[49] & w5665;
assign w20048 = w5663 & ~w7468;
assign w20049 = ~w20046 & ~w20047;
assign w20050 = ~w20045 & w20049;
assign w20051 = ~w20048 & w20050;
assign w20052 = a[44] & ~w20051;
assign w20053 = ~a[44] & w20051;
assign w20054 = ~w20052 & ~w20053;
assign w20055 = b[44] & w6732;
assign w20056 = b[45] & w6474;
assign w20057 = b[46] & w6476;
assign w20058 = w6469 & ~w6613;
assign w20059 = ~w20056 & ~w20057;
assign w20060 = ~w20055 & w20059;
assign w20061 = ~w20058 & w20060;
assign w20062 = a[47] & ~w20061;
assign w20063 = ~a[47] & w20061;
assign w20064 = ~w20062 & ~w20063;
assign w20065 = ~w19911 & ~w19916;
assign w20066 = b[38] & w8515;
assign w20067 = b[40] & w8202;
assign w20068 = b[39] & w8200;
assign w20069 = ~w5058 & w8195;
assign w20070 = ~w20067 & ~w20068;
assign w20071 = ~w20066 & w20070;
assign w20072 = ~w20069 & w20071;
assign w20073 = a[53] & ~w20072;
assign w20074 = ~a[53] & w20072;
assign w20075 = ~w20073 & ~w20074;
assign w20076 = ~w19894 & ~w19899;
assign w20077 = b[35] & w9482;
assign w20078 = b[36] & w9165;
assign w20079 = b[37] & w9160;
assign w20080 = ~w4357 & w9158;
assign w20081 = ~w20078 & ~w20079;
assign w20082 = ~w20077 & w20081;
assign w20083 = ~w20080 & w20082;
assign w20084 = a[56] & ~w20083;
assign w20085 = ~a[56] & w20083;
assign w20086 = ~w20084 & ~w20085;
assign w20087 = b[27] & w11921;
assign w20088 = b[28] & w11923;
assign w20089 = ~w20087 & ~w20088;
assign w20090 = ~w19845 & ~w19848;
assign w20091 = w20089 & ~w20090;
assign w20092 = ~w20089 & w20090;
assign w20093 = ~w20091 & ~w20092;
assign w20094 = b[29] & w11561;
assign w20095 = b[31] & w11196;
assign w20096 = b[30] & w11194;
assign w20097 = ~w3112 & w11189;
assign w20098 = ~w20095 & ~w20096;
assign w20099 = ~w20094 & w20098;
assign w20100 = ~w20097 & w20099;
assign w20101 = a[62] & ~w20100;
assign w20102 = ~a[62] & w20100;
assign w20103 = ~w20101 & ~w20102;
assign w20104 = ~w20093 & ~w20103;
assign w20105 = w20093 & w20103;
assign w20106 = ~w20104 & ~w20105;
assign w20107 = ~w19852 & ~w19864;
assign w20108 = w20106 & ~w20107;
assign w20109 = ~w20106 & w20107;
assign w20110 = ~w20108 & ~w20109;
assign w20111 = b[32] & w10496;
assign w20112 = b[33] & w10146;
assign w20113 = b[34] & w10148;
assign w20114 = ~w3710 & w10141;
assign w20115 = ~w20112 & ~w20113;
assign w20116 = ~w20111 & w20115;
assign w20117 = ~w20114 & w20116;
assign w20118 = a[59] & ~w20117;
assign w20119 = ~a[59] & w20117;
assign w20120 = ~w20118 & ~w20119;
assign w20121 = w20110 & w20120;
assign w20122 = ~w20110 & ~w20120;
assign w20123 = ~w20121 & ~w20122;
assign w20124 = ~w19878 & ~w19882;
assign w20125 = w20123 & ~w20124;
assign w20126 = ~w20123 & w20124;
assign w20127 = ~w20125 & ~w20126;
assign w20128 = w20086 & w20127;
assign w20129 = ~w20086 & ~w20127;
assign w20130 = ~w20128 & ~w20129;
assign w20131 = ~w20076 & w20130;
assign w20132 = w20076 & ~w20130;
assign w20133 = ~w20131 & ~w20132;
assign w20134 = w20075 & w20133;
assign w20135 = ~w20075 & ~w20133;
assign w20136 = ~w20134 & ~w20135;
assign w20137 = w20065 & ~w20136;
assign w20138 = ~w20065 & w20136;
assign w20139 = ~w20137 & ~w20138;
assign w20140 = b[41] & w7586;
assign w20141 = b[42] & w7307;
assign w20142 = b[43] & w7314;
assign w20143 = w5811 & w7312;
assign w20144 = ~w20141 & ~w20142;
assign w20145 = ~w20140 & w20144;
assign w20146 = ~w20143 & w20145;
assign w20147 = a[50] & ~w20146;
assign w20148 = ~a[50] & w20146;
assign w20149 = ~w20147 & ~w20148;
assign w20150 = w20139 & w20149;
assign w20151 = ~w20139 & ~w20149;
assign w20152 = ~w20150 & ~w20151;
assign w20153 = ~w19928 & ~w19931;
assign w20154 = w20152 & ~w20153;
assign w20155 = ~w20152 & w20153;
assign w20156 = ~w20154 & ~w20155;
assign w20157 = w20064 & w20156;
assign w20158 = ~w20064 & ~w20156;
assign w20159 = ~w20157 & ~w20158;
assign w20160 = ~w19934 & ~w19938;
assign w20161 = w20159 & ~w20160;
assign w20162 = ~w20159 & w20160;
assign w20163 = ~w20161 & ~w20162;
assign w20164 = w20054 & w20163;
assign w20165 = ~w20054 & ~w20163;
assign w20166 = ~w20164 & ~w20165;
assign w20167 = ~w19950 & ~w19955;
assign w20168 = w20166 & ~w20167;
assign w20169 = ~w20166 & w20167;
assign w20170 = ~w20168 & ~w20169;
assign w20171 = w20044 & w20170;
assign w20172 = ~w20044 & ~w20170;
assign w20173 = ~w20171 & ~w20172;
assign w20174 = ~w19967 & ~w19970;
assign w20175 = w20173 & w20174;
assign w20176 = ~w20173 & ~w20174;
assign w20177 = ~w20175 & ~w20176;
assign w20178 = w20034 & w20177;
assign w20179 = ~w20034 & ~w20177;
assign w20180 = ~w20178 & ~w20179;
assign w20181 = w20024 & ~w20180;
assign w20182 = ~w20024 & w20180;
assign w20183 = ~w20181 & ~w20182;
assign w20184 = b[56] & w3785;
assign w20185 = b[57] & w3578;
assign w20186 = b[58] & w3580;
assign w20187 = w3573 & ~w10339;
assign w20188 = ~w20185 & ~w20186;
assign w20189 = ~w20184 & w20188;
assign w20190 = ~w20187 & w20189;
assign w20191 = a[35] & ~w20190;
assign w20192 = ~a[35] & w20190;
assign w20193 = ~w20191 & ~w20192;
assign w20194 = w20183 & w20193;
assign w20195 = ~w20183 & ~w20193;
assign w20196 = ~w20194 & ~w20195;
assign w20197 = b[59] & w3177;
assign w20198 = b[61] & w2978;
assign w20199 = b[60] & w2973;
assign w20200 = w2980 & w11400;
assign w20201 = ~w20198 & ~w20199;
assign w20202 = ~w20197 & w20201;
assign w20203 = ~w20200 & w20202;
assign w20204 = a[32] & ~w20203;
assign w20205 = ~a[32] & w20203;
assign w20206 = ~w20204 & ~w20205;
assign w20207 = ~w19989 & ~w19994;
assign w20208 = w20206 & ~w20207;
assign w20209 = ~w20206 & w20207;
assign w20210 = ~w20208 & ~w20209;
assign w20211 = w20196 & w20210;
assign w20212 = ~w20196 & ~w20210;
assign w20213 = ~w20211 & ~w20212;
assign w20214 = ~w20007 & ~w20010;
assign w20215 = b[63] & w2436;
assign w20216 = b[62] & ~w2622;
assign w20217 = w2432 & w12156;
assign w20218 = ~w20215 & ~w20216;
assign w20219 = ~w20217 & w20218;
assign w20220 = a[29] & ~w20219;
assign w20221 = ~a[29] & w20219;
assign w20222 = ~w20220 & ~w20221;
assign w20223 = ~w20214 & w20222;
assign w20224 = w20214 & ~w20222;
assign w20225 = ~w20223 & ~w20224;
assign w20226 = w20213 & w20225;
assign w20227 = ~w20213 & ~w20225;
assign w20228 = ~w20226 & ~w20227;
assign w20229 = w20023 & ~w20228;
assign w20230 = ~w20023 & w20228;
assign w20231 = ~w20229 & ~w20230;
assign w20232 = ~w20017 & ~w20021;
assign w20233 = (w20231 & w20021) | (w20231 & w24463) | (w20021 & w24463);
assign w20234 = ~w20231 & w20232;
assign w20235 = ~w20233 & ~w20234;
assign w20236 = ~w20223 & ~w20226;
assign w20237 = ~w20175 & ~w20178;
assign w20238 = b[54] & w4453;
assign w20239 = b[55] & w4241;
assign w20240 = b[56] & w4243;
assign w20241 = ~w20239 & ~w20240;
assign w20242 = ~w20238 & w20241;
assign w20243 = (w20242 & ~w9657) | (w20242 & w25594) | (~w9657 & w25594);
assign w20244 = a[38] & ~w20243;
assign w20245 = ~a[38] & w20243;
assign w20246 = ~w20244 & ~w20245;
assign w20247 = ~w20168 & ~w20171;
assign w20248 = b[51] & w5167;
assign w20249 = b[53] & w4925;
assign w20250 = b[52] & w4918;
assign w20251 = w4923 & w8683;
assign w20252 = ~w20249 & ~w20250;
assign w20253 = ~w20248 & w20252;
assign w20254 = ~w20251 & w20253;
assign w20255 = a[41] & ~w20254;
assign w20256 = ~a[41] & w20254;
assign w20257 = ~w20255 & ~w20256;
assign w20258 = ~w20161 & ~w20164;
assign w20259 = b[48] & w5939;
assign w20260 = b[49] & w5670;
assign w20261 = b[50] & w5665;
assign w20262 = w5663 & w7759;
assign w20263 = ~w20260 & ~w20261;
assign w20264 = ~w20259 & w20263;
assign w20265 = ~w20262 & w20264;
assign w20266 = a[44] & ~w20265;
assign w20267 = ~a[44] & w20265;
assign w20268 = ~w20266 & ~w20267;
assign w20269 = ~w20138 & ~w20150;
assign w20270 = b[42] & w7586;
assign w20271 = b[44] & w7314;
assign w20272 = b[43] & w7307;
assign w20273 = w6069 & w7312;
assign w20274 = ~w20271 & ~w20272;
assign w20275 = ~w20270 & w20274;
assign w20276 = ~w20273 & w20275;
assign w20277 = a[50] & ~w20276;
assign w20278 = ~a[50] & w20276;
assign w20279 = ~w20277 & ~w20278;
assign w20280 = ~w20131 & ~w20134;
assign w20281 = b[39] & w8515;
assign w20282 = b[40] & w8200;
assign w20283 = b[41] & w8202;
assign w20284 = w5302 & w8195;
assign w20285 = ~w20282 & ~w20283;
assign w20286 = ~w20281 & w20285;
assign w20287 = ~w20284 & w20286;
assign w20288 = a[53] & ~w20287;
assign w20289 = ~a[53] & w20287;
assign w20290 = ~w20288 & ~w20289;
assign w20291 = ~w20108 & ~w20121;
assign w20292 = b[33] & w10496;
assign w20293 = b[34] & w10146;
assign w20294 = b[35] & w10148;
assign w20295 = w3918 & w10141;
assign w20296 = ~w20293 & ~w20294;
assign w20297 = ~w20292 & w20296;
assign w20298 = ~w20295 & w20297;
assign w20299 = a[59] & ~w20298;
assign w20300 = ~a[59] & w20298;
assign w20301 = ~w20299 & ~w20300;
assign w20302 = b[30] & w11561;
assign w20303 = b[32] & w11196;
assign w20304 = b[31] & w11194;
assign w20305 = w3304 & w11189;
assign w20306 = ~w20303 & ~w20304;
assign w20307 = ~w20302 & w20306;
assign w20308 = ~w20305 & w20307;
assign w20309 = a[62] & ~w20308;
assign w20310 = ~a[62] & w20308;
assign w20311 = ~w20309 & ~w20310;
assign w20312 = ~w20091 & ~w20105;
assign w20313 = b[28] & w11921;
assign w20314 = b[29] & w11923;
assign w20315 = ~w20313 & ~w20314;
assign w20316 = w20089 & ~w20315;
assign w20317 = ~w20089 & w20315;
assign w20318 = ~w20316 & ~w20317;
assign w20319 = w20312 & w20318;
assign w20320 = ~w20312 & ~w20318;
assign w20321 = ~w20319 & ~w20320;
assign w20322 = w20311 & ~w20321;
assign w20323 = ~w20311 & w20321;
assign w20324 = ~w20322 & ~w20323;
assign w20325 = w20301 & w20324;
assign w20326 = ~w20301 & ~w20324;
assign w20327 = ~w20325 & ~w20326;
assign w20328 = w20291 & ~w20327;
assign w20329 = ~w20291 & w20327;
assign w20330 = ~w20328 & ~w20329;
assign w20331 = b[36] & w9482;
assign w20332 = b[38] & w9160;
assign w20333 = b[37] & w9165;
assign w20334 = w4582 & w9158;
assign w20335 = ~w20332 & ~w20333;
assign w20336 = ~w20331 & w20335;
assign w20337 = ~w20334 & w20336;
assign w20338 = a[56] & ~w20337;
assign w20339 = ~a[56] & w20337;
assign w20340 = ~w20338 & ~w20339;
assign w20341 = w20330 & w20340;
assign w20342 = ~w20330 & ~w20340;
assign w20343 = ~w20341 & ~w20342;
assign w20344 = ~w20125 & ~w20128;
assign w20345 = w20343 & ~w20344;
assign w20346 = ~w20343 & w20344;
assign w20347 = ~w20345 & ~w20346;
assign w20348 = w20290 & w20347;
assign w20349 = ~w20290 & ~w20347;
assign w20350 = ~w20348 & ~w20349;
assign w20351 = ~w20280 & w20350;
assign w20352 = w20280 & ~w20350;
assign w20353 = ~w20351 & ~w20352;
assign w20354 = w20279 & w20353;
assign w20355 = ~w20279 & ~w20353;
assign w20356 = ~w20354 & ~w20355;
assign w20357 = w20269 & ~w20356;
assign w20358 = ~w20269 & w20356;
assign w20359 = ~w20357 & ~w20358;
assign w20360 = b[45] & w6732;
assign w20361 = b[47] & w6476;
assign w20362 = b[46] & w6474;
assign w20363 = w6469 & w6889;
assign w20364 = ~w20361 & ~w20362;
assign w20365 = ~w20360 & w20364;
assign w20366 = ~w20363 & w20365;
assign w20367 = a[47] & ~w20366;
assign w20368 = ~a[47] & w20366;
assign w20369 = ~w20367 & ~w20368;
assign w20370 = w20359 & w20369;
assign w20371 = ~w20359 & ~w20369;
assign w20372 = ~w20370 & ~w20371;
assign w20373 = ~w20154 & ~w20157;
assign w20374 = w20372 & ~w20373;
assign w20375 = ~w20372 & w20373;
assign w20376 = ~w20374 & ~w20375;
assign w20377 = ~w20268 & ~w20376;
assign w20378 = w20268 & w20376;
assign w20379 = ~w20377 & ~w20378;
assign w20380 = w20258 & ~w20379;
assign w20381 = ~w20258 & w20379;
assign w20382 = ~w20380 & ~w20381;
assign w20383 = w20257 & w20382;
assign w20384 = ~w20257 & ~w20382;
assign w20385 = ~w20383 & ~w20384;
assign w20386 = w20247 & ~w20385;
assign w20387 = ~w20247 & w20385;
assign w20388 = ~w20386 & ~w20387;
assign w20389 = w20246 & w20388;
assign w20390 = ~w20246 & ~w20388;
assign w20391 = ~w20389 & ~w20390;
assign w20392 = w20237 & ~w20391;
assign w20393 = ~w20237 & w20391;
assign w20394 = ~w20392 & ~w20393;
assign w20395 = b[57] & w3785;
assign w20396 = b[58] & w3578;
assign w20397 = b[59] & w3580;
assign w20398 = ~w20396 & ~w20397;
assign w20399 = ~w20395 & w20398;
assign w20400 = (w10371 & w25476) | (w10371 & w25477) | (w25476 & w25477);
assign w20401 = ~a[35] & w25741;
assign w20402 = ~w20400 & ~w20401;
assign w20403 = w20394 & w20402;
assign w20404 = ~w20394 & ~w20402;
assign w20405 = ~w20403 & ~w20404;
assign w20406 = b[60] & w3177;
assign w20407 = b[61] & w2973;
assign w20408 = b[62] & w2978;
assign w20409 = ~w20407 & ~w20408;
assign w20410 = ~w20406 & w20409;
assign w20411 = (w11763 & w24882) | (w11763 & w24883) | (w24882 & w24883);
assign w20412 = (~w11763 & w24884) | (~w11763 & w24885) | (w24884 & w24885);
assign w20413 = ~w20411 & ~w20412;
assign w20414 = ~w20182 & ~w20194;
assign w20415 = w20413 & ~w20414;
assign w20416 = ~w20413 & w20414;
assign w20417 = ~w20415 & ~w20416;
assign w20418 = ~w20405 & ~w20417;
assign w20419 = w20405 & w20417;
assign w20420 = ~w20418 & ~w20419;
assign w20421 = ~w20208 & ~w20211;
assign w20422 = w2432 & ~w12154;
assign w20423 = w2622 & ~w20422;
assign w20424 = b[63] & ~w20423;
assign w20425 = ~a[29] & ~w20424;
assign w20426 = a[29] & w20424;
assign w20427 = ~w20425 & ~w20426;
assign w20428 = ~w20421 & w20427;
assign w20429 = w20421 & ~w20427;
assign w20430 = ~w20428 & ~w20429;
assign w20431 = w20420 & w20430;
assign w20432 = ~w20420 & ~w20430;
assign w20433 = ~w20431 & ~w20432;
assign w20434 = w20236 & ~w20433;
assign w20435 = ~w20236 & w20433;
assign w20436 = ~w20434 & ~w20435;
assign w20437 = (~w20021 & w24464) | (~w20021 & w24465) | (w24464 & w24465);
assign w20438 = (w20021 & w24466) | (w20021 & w24467) | (w24466 & w24467);
assign w20439 = ~w20436 & w20437;
assign w20440 = ~w20438 & ~w20439;
assign w20441 = (~w20021 & w24468) | (~w20021 & w24469) | (w24468 & w24469);
assign w20442 = ~w20428 & ~w20431;
assign w20443 = ~w20381 & ~w20383;
assign w20444 = b[52] & w5167;
assign w20445 = b[53] & w4918;
assign w20446 = b[54] & w4925;
assign w20447 = ~w20445 & ~w20446;
assign w20448 = ~w20444 & w20447;
assign w20449 = a[41] & w25742;
assign w20450 = (w8998 & w25595) | (w8998 & w25596) | (w25595 & w25596);
assign w20451 = ~w20449 & ~w20450;
assign w20452 = ~w20374 & ~w20378;
assign w20453 = ~w20351 & ~w20354;
assign w20454 = b[43] & w7586;
assign w20455 = b[45] & w7314;
assign w20456 = b[44] & w7307;
assign w20457 = w6334 & w7312;
assign w20458 = ~w20455 & ~w20456;
assign w20459 = ~w20454 & w20458;
assign w20460 = ~w20457 & w20459;
assign w20461 = a[50] & ~w20460;
assign w20462 = ~a[50] & w20460;
assign w20463 = ~w20461 & ~w20462;
assign w20464 = ~w20345 & ~w20348;
assign w20465 = ~w20322 & ~w20325;
assign w20466 = b[34] & w10496;
assign w20467 = b[36] & w10148;
assign w20468 = b[35] & w10146;
assign w20469 = w4129 & w10141;
assign w20470 = ~w20467 & ~w20468;
assign w20471 = ~w20466 & w20470;
assign w20472 = ~w20469 & w20471;
assign w20473 = a[59] & ~w20472;
assign w20474 = ~a[59] & w20472;
assign w20475 = ~w20473 & ~w20474;
assign w20476 = b[31] & w11561;
assign w20477 = b[33] & w11196;
assign w20478 = b[32] & w11194;
assign w20479 = w3499 & w11189;
assign w20480 = ~w20477 & ~w20478;
assign w20481 = ~w20476 & w20480;
assign w20482 = ~w20479 & w20481;
assign w20483 = a[62] & ~w20482;
assign w20484 = ~a[62] & w20482;
assign w20485 = ~w20483 & ~w20484;
assign w20486 = b[29] & w11921;
assign w20487 = b[30] & w11923;
assign w20488 = ~w20486 & ~w20487;
assign w20489 = ~a[29] & ~w20488;
assign w20490 = a[29] & w20488;
assign w20491 = ~w20489 & ~w20490;
assign w20492 = w20315 & ~w20491;
assign w20493 = ~w20315 & w20491;
assign w20494 = ~w20492 & ~w20493;
assign w20495 = ~w20316 & ~w20319;
assign w20496 = w20494 & w20495;
assign w20497 = ~w20494 & ~w20495;
assign w20498 = ~w20496 & ~w20497;
assign w20499 = w20485 & w20498;
assign w20500 = ~w20485 & ~w20498;
assign w20501 = ~w20499 & ~w20500;
assign w20502 = w20475 & w20501;
assign w20503 = ~w20475 & ~w20501;
assign w20504 = ~w20502 & ~w20503;
assign w20505 = ~w20465 & w20504;
assign w20506 = w20465 & ~w20504;
assign w20507 = ~w20505 & ~w20506;
assign w20508 = b[37] & w9482;
assign w20509 = b[38] & w9165;
assign w20510 = b[39] & w9160;
assign w20511 = ~w4812 & w9158;
assign w20512 = ~w20509 & ~w20510;
assign w20513 = ~w20508 & w20512;
assign w20514 = ~w20511 & w20513;
assign w20515 = a[56] & ~w20514;
assign w20516 = ~a[56] & w20514;
assign w20517 = ~w20515 & ~w20516;
assign w20518 = w20507 & w20517;
assign w20519 = ~w20507 & ~w20517;
assign w20520 = ~w20518 & ~w20519;
assign w20521 = ~w20329 & ~w20341;
assign w20522 = ~w20520 & w20521;
assign w20523 = w20520 & ~w20521;
assign w20524 = ~w20522 & ~w20523;
assign w20525 = b[40] & w8515;
assign w20526 = b[42] & w8202;
assign w20527 = b[41] & w8200;
assign w20528 = w5548 & w8195;
assign w20529 = ~w20526 & ~w20527;
assign w20530 = ~w20525 & w20529;
assign w20531 = ~w20528 & w20530;
assign w20532 = a[53] & ~w20531;
assign w20533 = ~a[53] & w20531;
assign w20534 = ~w20532 & ~w20533;
assign w20535 = w20524 & w20534;
assign w20536 = ~w20524 & ~w20534;
assign w20537 = ~w20535 & ~w20536;
assign w20538 = ~w20464 & w20537;
assign w20539 = w20464 & ~w20537;
assign w20540 = ~w20538 & ~w20539;
assign w20541 = w20463 & w20540;
assign w20542 = ~w20463 & ~w20540;
assign w20543 = ~w20541 & ~w20542;
assign w20544 = w20453 & ~w20543;
assign w20545 = ~w20453 & w20543;
assign w20546 = ~w20544 & ~w20545;
assign w20547 = b[46] & w6732;
assign w20548 = b[48] & w6476;
assign w20549 = b[47] & w6474;
assign w20550 = ~w20548 & ~w20549;
assign w20551 = ~w20547 & w20550;
assign w20552 = (w20551 & w7170) | (w20551 & w25597) | (w7170 & w25597);
assign w20553 = a[47] & ~w20552;
assign w20554 = ~a[47] & w20552;
assign w20555 = ~w20553 & ~w20554;
assign w20556 = w20546 & w20555;
assign w20557 = ~w20546 & ~w20555;
assign w20558 = ~w20556 & ~w20557;
assign w20559 = ~w20358 & ~w20370;
assign w20560 = ~w20558 & w20559;
assign w20561 = w20558 & ~w20559;
assign w20562 = ~w20560 & ~w20561;
assign w20563 = b[49] & w5939;
assign w20564 = b[51] & w5665;
assign w20565 = b[50] & w5670;
assign w20566 = ~w20564 & ~w20565;
assign w20567 = ~w20563 & w20566;
assign w20568 = (w20567 & w8058) | (w20567 & w25598) | (w8058 & w25598);
assign w20569 = a[44] & ~w20568;
assign w20570 = ~a[44] & w20568;
assign w20571 = ~w20569 & ~w20570;
assign w20572 = ~w20562 & ~w20571;
assign w20573 = w20562 & w20571;
assign w20574 = ~w20572 & ~w20573;
assign w20575 = w20452 & w20574;
assign w20576 = ~w20452 & ~w20574;
assign w20577 = ~w20575 & ~w20576;
assign w20578 = w20451 & ~w20577;
assign w20579 = ~w20451 & w20577;
assign w20580 = ~w20578 & ~w20579;
assign w20581 = ~w20443 & w20580;
assign w20582 = w20443 & ~w20580;
assign w20583 = ~w20581 & ~w20582;
assign w20584 = b[55] & w4453;
assign w20585 = b[57] & w4243;
assign w20586 = b[56] & w4241;
assign w20587 = ~w20585 & ~w20586;
assign w20588 = ~w20584 & w20587;
assign w20589 = a[38] & w25743;
assign w20590 = (w9992 & w25479) | (w9992 & w25480) | (w25479 & w25480);
assign w20591 = ~w20589 & ~w20590;
assign w20592 = w20583 & w20591;
assign w20593 = ~w20583 & ~w20591;
assign w20594 = ~w20592 & ~w20593;
assign w20595 = ~w20387 & ~w20389;
assign w20596 = ~w20594 & w20595;
assign w20597 = w20594 & ~w20595;
assign w20598 = ~w20596 & ~w20597;
assign w20599 = b[58] & w3785;
assign w20600 = b[59] & w3578;
assign w20601 = b[60] & w3580;
assign w20602 = ~w20600 & ~w20601;
assign w20603 = ~w20599 & w20602;
assign w20604 = (w11035 & w25216) | (w11035 & w25217) | (w25216 & w25217);
assign w20605 = (~w11035 & w25218) | (~w11035 & w25219) | (w25218 & w25219);
assign w20606 = ~w20604 & ~w20605;
assign w20607 = w20598 & w20606;
assign w20608 = ~w20598 & ~w20606;
assign w20609 = ~w20607 & ~w20608;
assign w20610 = ~w20393 & ~w20403;
assign w20611 = ~w20609 & w20610;
assign w20612 = w20609 & ~w20610;
assign w20613 = ~w20611 & ~w20612;
assign w20614 = (~w20415 & ~w20417) | (~w20415 & w25031) | (~w20417 & w25031);
assign w20615 = b[61] & w3177;
assign w20616 = b[63] & w2978;
assign w20617 = b[62] & w2973;
assign w20618 = ~w20616 & ~w20617;
assign w20619 = ~w20615 & w20618;
assign w20620 = (w20619 & ~w12132) | (w20619 & w25481) | (~w12132 & w25481);
assign w20621 = a[32] & ~w20620;
assign w20622 = ~a[32] & w20620;
assign w20623 = ~w20621 & ~w20622;
assign w20624 = ~w20614 & w20623;
assign w20625 = w20614 & ~w20623;
assign w20626 = ~w20624 & ~w20625;
assign w20627 = ~w20613 & ~w20626;
assign w20628 = w20613 & w20626;
assign w20629 = ~w20627 & ~w20628;
assign w20630 = ~w20442 & w20629;
assign w20631 = w20442 & ~w20629;
assign w20632 = ~w20630 & ~w20631;
assign w20633 = w20441 & ~w20632;
assign w20634 = ~w20441 & w20632;
assign w20635 = ~w20633 & ~w20634;
assign w20636 = (~w20624 & ~w20626) | (~w20624 & w25482) | (~w20626 & w25482);
assign w20637 = b[59] & w3785;
assign w20638 = b[60] & w3578;
assign w20639 = b[61] & w3580;
assign w20640 = ~w20638 & ~w20639;
assign w20641 = ~w20637 & w20640;
assign w20642 = (w11400 & w25327) | (w11400 & w25328) | (w25327 & w25328);
assign w20643 = (~w11400 & w25329) | (~w11400 & w25330) | (w25329 & w25330);
assign w20644 = ~w20642 & ~w20643;
assign w20645 = ~w20578 & ~w20581;
assign w20646 = b[53] & w5167;
assign w20647 = b[54] & w4918;
assign w20648 = b[55] & w4925;
assign w20649 = ~w20647 & ~w20648;
assign w20650 = ~w20646 & w20649;
assign w20651 = (w20650 & w9330) | (w20650 & w25599) | (w9330 & w25599);
assign w20652 = a[41] & ~w20651;
assign w20653 = ~a[41] & w20651;
assign w20654 = ~w20652 & ~w20653;
assign w20655 = b[50] & w5939;
assign w20656 = b[52] & w5665;
assign w20657 = b[51] & w5670;
assign w20658 = ~w20656 & ~w20657;
assign w20659 = ~w20655 & w20658;
assign w20660 = (w20659 & w8371) | (w20659 & w25600) | (w8371 & w25600);
assign w20661 = a[44] & ~w20660;
assign w20662 = ~a[44] & w20660;
assign w20663 = ~w20661 & ~w20662;
assign w20664 = b[47] & w6732;
assign w20665 = b[49] & w6476;
assign w20666 = b[48] & w6474;
assign w20667 = ~w20665 & ~w20666;
assign w20668 = ~w20664 & w20667;
assign w20669 = (w20668 & w7468) | (w20668 & w25601) | (w7468 & w25601);
assign w20670 = a[47] & ~w20669;
assign w20671 = ~a[47] & w20669;
assign w20672 = ~w20670 & ~w20671;
assign w20673 = b[44] & w7586;
assign w20674 = b[46] & w7314;
assign w20675 = b[45] & w7307;
assign w20676 = ~w6613 & w7312;
assign w20677 = ~w20674 & ~w20675;
assign w20678 = ~w20673 & w20677;
assign w20679 = ~w20676 & w20678;
assign w20680 = a[50] & ~w20679;
assign w20681 = ~a[50] & w20679;
assign w20682 = ~w20680 & ~w20681;
assign w20683 = ~w20518 & ~w20523;
assign w20684 = b[38] & w9482;
assign w20685 = b[40] & w9160;
assign w20686 = b[39] & w9165;
assign w20687 = ~w5058 & w9158;
assign w20688 = ~w20685 & ~w20686;
assign w20689 = ~w20684 & w20688;
assign w20690 = ~w20687 & w20689;
assign w20691 = a[56] & ~w20690;
assign w20692 = ~a[56] & w20690;
assign w20693 = ~w20691 & ~w20692;
assign w20694 = ~w20502 & ~w20505;
assign w20695 = b[35] & w10496;
assign w20696 = b[37] & w10148;
assign w20697 = b[36] & w10146;
assign w20698 = ~w4357 & w10141;
assign w20699 = ~w20696 & ~w20697;
assign w20700 = ~w20695 & w20699;
assign w20701 = ~w20698 & w20700;
assign w20702 = a[59] & ~w20701;
assign w20703 = ~a[59] & w20701;
assign w20704 = ~w20702 & ~w20703;
assign w20705 = ~w20496 & ~w20499;
assign w20706 = b[30] & w11921;
assign w20707 = b[31] & w11923;
assign w20708 = ~w20706 & ~w20707;
assign w20709 = ~w20489 & ~w20493;
assign w20710 = w20708 & ~w20709;
assign w20711 = ~w20708 & w20709;
assign w20712 = ~w20710 & ~w20711;
assign w20713 = b[32] & w11561;
assign w20714 = b[34] & w11196;
assign w20715 = b[33] & w11194;
assign w20716 = ~w3710 & w11189;
assign w20717 = ~w20714 & ~w20715;
assign w20718 = ~w20713 & w20717;
assign w20719 = ~w20716 & w20718;
assign w20720 = a[62] & ~w20719;
assign w20721 = ~a[62] & w20719;
assign w20722 = ~w20720 & ~w20721;
assign w20723 = ~w20712 & ~w20722;
assign w20724 = w20712 & w20722;
assign w20725 = ~w20723 & ~w20724;
assign w20726 = w20705 & ~w20725;
assign w20727 = ~w20705 & w20725;
assign w20728 = ~w20726 & ~w20727;
assign w20729 = w20704 & w20728;
assign w20730 = ~w20704 & ~w20728;
assign w20731 = ~w20729 & ~w20730;
assign w20732 = w20694 & ~w20731;
assign w20733 = ~w20694 & w20731;
assign w20734 = ~w20732 & ~w20733;
assign w20735 = w20693 & w20734;
assign w20736 = ~w20693 & ~w20734;
assign w20737 = ~w20735 & ~w20736;
assign w20738 = w20683 & ~w20737;
assign w20739 = ~w20683 & w20737;
assign w20740 = ~w20738 & ~w20739;
assign w20741 = b[41] & w8515;
assign w20742 = b[42] & w8200;
assign w20743 = b[43] & w8202;
assign w20744 = w5811 & w8195;
assign w20745 = ~w20742 & ~w20743;
assign w20746 = ~w20741 & w20745;
assign w20747 = ~w20744 & w20746;
assign w20748 = a[53] & ~w20747;
assign w20749 = ~a[53] & w20747;
assign w20750 = ~w20748 & ~w20749;
assign w20751 = w20740 & w20750;
assign w20752 = ~w20740 & ~w20750;
assign w20753 = ~w20751 & ~w20752;
assign w20754 = ~w20535 & ~w20538;
assign w20755 = w20753 & ~w20754;
assign w20756 = ~w20753 & w20754;
assign w20757 = ~w20755 & ~w20756;
assign w20758 = w20682 & w20757;
assign w20759 = ~w20682 & ~w20757;
assign w20760 = ~w20758 & ~w20759;
assign w20761 = ~w20541 & ~w20545;
assign w20762 = w20760 & ~w20761;
assign w20763 = ~w20760 & w20761;
assign w20764 = ~w20762 & ~w20763;
assign w20765 = w20672 & w20764;
assign w20766 = ~w20672 & ~w20764;
assign w20767 = ~w20765 & ~w20766;
assign w20768 = ~w20556 & ~w20561;
assign w20769 = w20767 & ~w20768;
assign w20770 = ~w20767 & w20768;
assign w20771 = ~w20769 & ~w20770;
assign w20772 = w20663 & w20771;
assign w20773 = ~w20663 & ~w20771;
assign w20774 = ~w20772 & ~w20773;
assign w20775 = ~w20572 & ~w20575;
assign w20776 = w20774 & w20775;
assign w20777 = ~w20774 & ~w20775;
assign w20778 = ~w20776 & ~w20777;
assign w20779 = w20654 & w20778;
assign w20780 = ~w20654 & ~w20778;
assign w20781 = ~w20779 & ~w20780;
assign w20782 = w20645 & ~w20781;
assign w20783 = ~w20645 & w20781;
assign w20784 = ~w20782 & ~w20783;
assign w20785 = b[56] & w4453;
assign w20786 = b[57] & w4241;
assign w20787 = b[58] & w4243;
assign w20788 = ~w20786 & ~w20787;
assign w20789 = ~w20785 & w20788;
assign w20790 = (~w10339 & w25483) | (~w10339 & w25484) | (w25483 & w25484);
assign w20791 = (w10339 & w25485) | (w10339 & w25486) | (w25485 & w25486);
assign w20792 = ~w20790 & ~w20791;
assign w20793 = w20784 & w20792;
assign w20794 = ~w20784 & ~w20792;
assign w20795 = ~w20793 & ~w20794;
assign w20796 = (~w20592 & ~w20594) | (~w20592 & w25602) | (~w20594 & w25602);
assign w20797 = w20795 & ~w20796;
assign w20798 = ~w20795 & w20796;
assign w20799 = ~w20797 & ~w20798;
assign w20800 = w20644 & w20799;
assign w20801 = ~w20644 & ~w20799;
assign w20802 = ~w20800 & ~w20801;
assign w20803 = (~w20607 & ~w20609) | (~w20607 & w25332) | (~w20609 & w25332);
assign w20804 = b[62] & w3177;
assign w20805 = b[63] & w2973;
assign w20806 = ~w12153 & w24723;
assign w20807 = ~w20804 & ~w20805;
assign w20808 = ~w20806 & w25033;
assign w20809 = (a[32] & w20806) | (a[32] & w25034) | (w20806 & w25034);
assign w20810 = ~w20808 & ~w20809;
assign w20811 = ~w20803 & w20810;
assign w20812 = w20803 & ~w20810;
assign w20813 = ~w20811 & ~w20812;
assign w20814 = w20802 & w20813;
assign w20815 = ~w20802 & ~w20813;
assign w20816 = ~w20814 & ~w20815;
assign w20817 = ~w20636 & w20816;
assign w20818 = w20636 & ~w20816;
assign w20819 = ~w20817 & ~w20818;
assign w20820 = (~w18109 & w24724) | (~w18109 & w24725) | (w24724 & w24725);
assign w20821 = w20819 & w20820;
assign w20822 = ~w20819 & ~w20820;
assign w20823 = ~w20821 & ~w20822;
assign w20824 = (~w20811 & ~w20813) | (~w20811 & w25487) | (~w20813 & w25487);
assign w20825 = b[60] & w3785;
assign w20826 = b[61] & w3578;
assign w20827 = b[62] & w3580;
assign w20828 = ~w20826 & ~w20827;
assign w20829 = ~w20825 & w20828;
assign w20830 = (w11763 & w25488) | (w11763 & w25489) | (w25488 & w25489);
assign w20831 = (~w11763 & w25490) | (~w11763 & w25491) | (w25490 & w25491);
assign w20832 = ~w20830 & ~w20831;
assign w20833 = ~w20776 & ~w20779;
assign w20834 = b[54] & w5167;
assign w20835 = b[55] & w4918;
assign w20836 = b[56] & w4925;
assign w20837 = ~w20835 & ~w20836;
assign w20838 = ~w20834 & w20837;
assign w20839 = (w20838 & ~w9657) | (w20838 & w25492) | (~w9657 & w25492);
assign w20840 = a[41] & ~w20839;
assign w20841 = ~a[41] & w20839;
assign w20842 = ~w20840 & ~w20841;
assign w20843 = ~w20769 & ~w20772;
assign w20844 = b[51] & w5939;
assign w20845 = b[53] & w5665;
assign w20846 = b[52] & w5670;
assign w20847 = w5663 & w8683;
assign w20848 = ~w20845 & ~w20846;
assign w20849 = ~w20844 & w20848;
assign w20850 = ~w20847 & w20849;
assign w20851 = a[44] & ~w20850;
assign w20852 = ~a[44] & w20850;
assign w20853 = ~w20851 & ~w20852;
assign w20854 = ~w20762 & ~w20765;
assign w20855 = b[48] & w6732;
assign w20856 = b[50] & w6476;
assign w20857 = b[49] & w6474;
assign w20858 = w6469 & w7759;
assign w20859 = ~w20856 & ~w20857;
assign w20860 = ~w20855 & w20859;
assign w20861 = ~w20858 & w20860;
assign w20862 = a[47] & ~w20861;
assign w20863 = ~a[47] & w20861;
assign w20864 = ~w20862 & ~w20863;
assign w20865 = ~w20739 & ~w20751;
assign w20866 = b[42] & w8515;
assign w20867 = b[44] & w8202;
assign w20868 = b[43] & w8200;
assign w20869 = w6069 & w8195;
assign w20870 = ~w20867 & ~w20868;
assign w20871 = ~w20866 & w20870;
assign w20872 = ~w20869 & w20871;
assign w20873 = a[53] & ~w20872;
assign w20874 = ~a[53] & w20872;
assign w20875 = ~w20873 & ~w20874;
assign w20876 = ~w20733 & ~w20735;
assign w20877 = b[39] & w9482;
assign w20878 = b[40] & w9165;
assign w20879 = b[41] & w9160;
assign w20880 = w5302 & w9158;
assign w20881 = ~w20878 & ~w20879;
assign w20882 = ~w20877 & w20881;
assign w20883 = ~w20880 & w20882;
assign w20884 = a[56] & ~w20883;
assign w20885 = ~a[56] & w20883;
assign w20886 = ~w20884 & ~w20885;
assign w20887 = ~w20727 & ~w20729;
assign w20888 = b[36] & w10496;
assign w20889 = b[38] & w10148;
assign w20890 = b[37] & w10146;
assign w20891 = w4582 & w10141;
assign w20892 = ~w20889 & ~w20890;
assign w20893 = ~w20888 & w20892;
assign w20894 = ~w20891 & w20893;
assign w20895 = a[59] & ~w20894;
assign w20896 = ~a[59] & w20894;
assign w20897 = ~w20895 & ~w20896;
assign w20898 = b[33] & w11561;
assign w20899 = b[35] & w11196;
assign w20900 = b[34] & w11194;
assign w20901 = w3918 & w11189;
assign w20902 = ~w20899 & ~w20900;
assign w20903 = ~w20898 & w20902;
assign w20904 = ~w20901 & w20903;
assign w20905 = a[62] & ~w20904;
assign w20906 = ~a[62] & w20904;
assign w20907 = ~w20905 & ~w20906;
assign w20908 = ~w20710 & ~w20724;
assign w20909 = b[31] & w11921;
assign w20910 = b[32] & w11923;
assign w20911 = ~w20909 & ~w20910;
assign w20912 = w20708 & ~w20911;
assign w20913 = ~w20708 & w20911;
assign w20914 = ~w20912 & ~w20913;
assign w20915 = w20908 & w20914;
assign w20916 = ~w20908 & ~w20914;
assign w20917 = ~w20915 & ~w20916;
assign w20918 = w20907 & ~w20917;
assign w20919 = ~w20907 & w20917;
assign w20920 = ~w20918 & ~w20919;
assign w20921 = w20897 & w20920;
assign w20922 = ~w20897 & ~w20920;
assign w20923 = ~w20921 & ~w20922;
assign w20924 = ~w20887 & w20923;
assign w20925 = w20887 & ~w20923;
assign w20926 = ~w20924 & ~w20925;
assign w20927 = w20886 & w20926;
assign w20928 = ~w20886 & ~w20926;
assign w20929 = ~w20927 & ~w20928;
assign w20930 = w20876 & ~w20929;
assign w20931 = ~w20876 & w20929;
assign w20932 = ~w20930 & ~w20931;
assign w20933 = w20875 & w20932;
assign w20934 = ~w20875 & ~w20932;
assign w20935 = ~w20933 & ~w20934;
assign w20936 = w20865 & ~w20935;
assign w20937 = ~w20865 & w20935;
assign w20938 = ~w20936 & ~w20937;
assign w20939 = b[45] & w7586;
assign w20940 = b[47] & w7314;
assign w20941 = b[46] & w7307;
assign w20942 = w6889 & w7312;
assign w20943 = ~w20940 & ~w20941;
assign w20944 = ~w20939 & w20943;
assign w20945 = ~w20942 & w20944;
assign w20946 = a[50] & ~w20945;
assign w20947 = ~a[50] & w20945;
assign w20948 = ~w20946 & ~w20947;
assign w20949 = w20938 & w20948;
assign w20950 = ~w20938 & ~w20948;
assign w20951 = ~w20949 & ~w20950;
assign w20952 = ~w20755 & ~w20758;
assign w20953 = w20951 & ~w20952;
assign w20954 = ~w20951 & w20952;
assign w20955 = ~w20953 & ~w20954;
assign w20956 = ~w20864 & ~w20955;
assign w20957 = w20864 & w20955;
assign w20958 = ~w20956 & ~w20957;
assign w20959 = w20854 & ~w20958;
assign w20960 = ~w20854 & w20958;
assign w20961 = ~w20959 & ~w20960;
assign w20962 = w20853 & w20961;
assign w20963 = ~w20853 & ~w20961;
assign w20964 = ~w20962 & ~w20963;
assign w20965 = w20843 & ~w20964;
assign w20966 = ~w20843 & w20964;
assign w20967 = ~w20965 & ~w20966;
assign w20968 = w20842 & w20967;
assign w20969 = ~w20842 & ~w20967;
assign w20970 = ~w20968 & ~w20969;
assign w20971 = w20833 & ~w20970;
assign w20972 = ~w20833 & w20970;
assign w20973 = ~w20971 & ~w20972;
assign w20974 = b[57] & w4453;
assign w20975 = b[58] & w4241;
assign w20976 = b[59] & w4243;
assign w20977 = ~w20975 & ~w20976;
assign w20978 = ~w20974 & w20977;
assign w20979 = (w10371 & w25333) | (w10371 & w25334) | (w25333 & w25334);
assign w20980 = (~w10371 & w25335) | (~w10371 & w25336) | (w25335 & w25336);
assign w20981 = ~w20979 & ~w20980;
assign w20982 = w20973 & w20981;
assign w20983 = ~w20973 & ~w20981;
assign w20984 = ~w20982 & ~w20983;
assign w20985 = ~w20783 & ~w20793;
assign w20986 = w20984 & ~w20985;
assign w20987 = ~w20984 & w20985;
assign w20988 = ~w20986 & ~w20987;
assign w20989 = w20832 & w20988;
assign w20990 = ~w20832 & ~w20988;
assign w20991 = ~w20989 & ~w20990;
assign w20992 = (~w20797 & ~w20644) | (~w20797 & w25493) | (~w20644 & w25493);
assign w20993 = (w25495 & w25494) | (w25495 & ~w11757) | (w25494 & ~w11757);
assign w20994 = ~w3177 & ~w20993;
assign w20995 = b[63] & ~w20994;
assign w20996 = ~a[32] & ~w20995;
assign w20997 = a[32] & w20995;
assign w20998 = ~w20996 & ~w20997;
assign w20999 = ~w20992 & w20998;
assign w21000 = w20992 & ~w20998;
assign w21001 = ~w20999 & ~w21000;
assign w21002 = w20991 & w21001;
assign w21003 = ~w20991 & ~w21001;
assign w21004 = ~w21002 & ~w21003;
assign w21005 = ~w20824 & w21004;
assign w21006 = w20824 & ~w21004;
assign w21007 = ~w21005 & ~w21006;
assign w21008 = (w18109 & w25673) | (w18109 & w25674) | (w25673 & w25674);
assign w21009 = (w20820 & w24475) | (w20820 & w24476) | (w24475 & w24476);
assign w21010 = ~w21007 & w21008;
assign w21011 = ~w21009 & ~w21010;
assign w21012 = (w18109 & w25675) | (w18109 & w25676) | (w25675 & w25676);
assign w21013 = ~w20999 & ~w21002;
assign w21014 = ~w20960 & ~w20962;
assign w21015 = b[52] & w5939;
assign w21016 = b[54] & w5665;
assign w21017 = b[53] & w5670;
assign w21018 = w5663 & ~w8998;
assign w21019 = ~w21016 & ~w21017;
assign w21020 = ~w21015 & w21019;
assign w21021 = ~w21018 & w21020;
assign w21022 = a[44] & ~w21021;
assign w21023 = ~a[44] & w21021;
assign w21024 = ~w21022 & ~w21023;
assign w21025 = ~w20953 & ~w20957;
assign w21026 = ~w20918 & ~w20921;
assign w21027 = b[37] & w10496;
assign w21028 = b[39] & w10148;
assign w21029 = b[38] & w10146;
assign w21030 = ~w4812 & w10141;
assign w21031 = ~w21028 & ~w21029;
assign w21032 = ~w21027 & w21031;
assign w21033 = ~w21030 & w21032;
assign w21034 = a[59] & ~w21033;
assign w21035 = ~a[59] & w21033;
assign w21036 = ~w21034 & ~w21035;
assign w21037 = b[34] & w11561;
assign w21038 = b[36] & w11196;
assign w21039 = b[35] & w11194;
assign w21040 = w4129 & w11189;
assign w21041 = ~w21038 & ~w21039;
assign w21042 = ~w21037 & w21041;
assign w21043 = ~w21040 & w21042;
assign w21044 = a[62] & ~w21043;
assign w21045 = ~a[62] & w21043;
assign w21046 = ~w21044 & ~w21045;
assign w21047 = b[32] & w11921;
assign w21048 = b[33] & w11923;
assign w21049 = ~w21047 & ~w21048;
assign w21050 = ~a[32] & ~w21049;
assign w21051 = a[32] & w21049;
assign w21052 = ~w21050 & ~w21051;
assign w21053 = w20911 & ~w21052;
assign w21054 = ~w20911 & w21052;
assign w21055 = ~w21053 & ~w21054;
assign w21056 = ~w20912 & ~w20915;
assign w21057 = w21055 & w21056;
assign w21058 = ~w21055 & ~w21056;
assign w21059 = ~w21057 & ~w21058;
assign w21060 = w21046 & w21059;
assign w21061 = ~w21046 & ~w21059;
assign w21062 = ~w21060 & ~w21061;
assign w21063 = w21036 & w21062;
assign w21064 = ~w21036 & ~w21062;
assign w21065 = ~w21063 & ~w21064;
assign w21066 = ~w21026 & w21065;
assign w21067 = w21026 & ~w21065;
assign w21068 = ~w21066 & ~w21067;
assign w21069 = b[40] & w9482;
assign w21070 = b[42] & w9160;
assign w21071 = b[41] & w9165;
assign w21072 = w5548 & w9158;
assign w21073 = ~w21070 & ~w21071;
assign w21074 = ~w21069 & w21073;
assign w21075 = ~w21072 & w21074;
assign w21076 = a[56] & ~w21075;
assign w21077 = ~a[56] & w21075;
assign w21078 = ~w21076 & ~w21077;
assign w21079 = w21068 & w21078;
assign w21080 = ~w21068 & ~w21078;
assign w21081 = ~w21079 & ~w21080;
assign w21082 = ~w20924 & ~w20927;
assign w21083 = ~w21081 & w21082;
assign w21084 = w21081 & ~w21082;
assign w21085 = ~w21083 & ~w21084;
assign w21086 = b[43] & w8515;
assign w21087 = b[44] & w8200;
assign w21088 = b[45] & w8202;
assign w21089 = w6334 & w8195;
assign w21090 = ~w21087 & ~w21088;
assign w21091 = ~w21086 & w21090;
assign w21092 = ~w21089 & w21091;
assign w21093 = a[53] & ~w21092;
assign w21094 = ~a[53] & w21092;
assign w21095 = ~w21093 & ~w21094;
assign w21096 = w21085 & w21095;
assign w21097 = ~w21085 & ~w21095;
assign w21098 = ~w21096 & ~w21097;
assign w21099 = ~w20931 & ~w20933;
assign w21100 = ~w21098 & w21099;
assign w21101 = w21098 & ~w21099;
assign w21102 = ~w21100 & ~w21101;
assign w21103 = b[46] & w7586;
assign w21104 = b[47] & w7307;
assign w21105 = b[48] & w7314;
assign w21106 = ~w7170 & w7312;
assign w21107 = ~w21104 & ~w21105;
assign w21108 = ~w21103 & w21107;
assign w21109 = ~w21106 & w21108;
assign w21110 = a[50] & ~w21109;
assign w21111 = ~a[50] & w21109;
assign w21112 = ~w21110 & ~w21111;
assign w21113 = w21102 & w21112;
assign w21114 = ~w21102 & ~w21112;
assign w21115 = ~w21113 & ~w21114;
assign w21116 = ~w20937 & ~w20949;
assign w21117 = ~w21115 & w21116;
assign w21118 = w21115 & ~w21116;
assign w21119 = ~w21117 & ~w21118;
assign w21120 = b[49] & w6732;
assign w21121 = b[51] & w6476;
assign w21122 = b[50] & w6474;
assign w21123 = w6469 & ~w8058;
assign w21124 = ~w21121 & ~w21122;
assign w21125 = ~w21120 & w21124;
assign w21126 = ~w21123 & w21125;
assign w21127 = a[47] & ~w21126;
assign w21128 = ~a[47] & w21126;
assign w21129 = ~w21127 & ~w21128;
assign w21130 = ~w21119 & ~w21129;
assign w21131 = w21119 & w21129;
assign w21132 = ~w21130 & ~w21131;
assign w21133 = w21025 & w21132;
assign w21134 = ~w21025 & ~w21132;
assign w21135 = ~w21133 & ~w21134;
assign w21136 = w21024 & ~w21135;
assign w21137 = ~w21024 & w21135;
assign w21138 = ~w21136 & ~w21137;
assign w21139 = ~w21014 & w21138;
assign w21140 = w21014 & ~w21138;
assign w21141 = ~w21139 & ~w21140;
assign w21142 = b[55] & w5167;
assign w21143 = b[56] & w4918;
assign w21144 = b[57] & w4925;
assign w21145 = w4923 & ~w9992;
assign w21146 = ~w21143 & ~w21144;
assign w21147 = ~w21142 & w21146;
assign w21148 = ~w21145 & w21147;
assign w21149 = a[41] & ~w21148;
assign w21150 = ~a[41] & w21148;
assign w21151 = ~w21149 & ~w21150;
assign w21152 = w21141 & w21151;
assign w21153 = ~w21141 & ~w21151;
assign w21154 = ~w21152 & ~w21153;
assign w21155 = ~w20966 & ~w20968;
assign w21156 = ~w21154 & w21155;
assign w21157 = w21154 & ~w21155;
assign w21158 = ~w21156 & ~w21157;
assign w21159 = b[58] & w4453;
assign w21160 = b[59] & w4241;
assign w21161 = b[60] & w4243;
assign w21162 = ~w21160 & ~w21161;
assign w21163 = ~w21159 & w21162;
assign w21164 = (w11035 & w25603) | (w11035 & w25604) | (w25603 & w25604);
assign w21165 = ~a[38] & w25744;
assign w21166 = ~w21164 & ~w21165;
assign w21167 = w21158 & w21166;
assign w21168 = ~w21158 & ~w21166;
assign w21169 = ~w21167 & ~w21168;
assign w21170 = ~w20972 & ~w20982;
assign w21171 = ~w21169 & w21170;
assign w21172 = w21169 & ~w21170;
assign w21173 = ~w21171 & ~w21172;
assign w21174 = (~w20986 & ~w20988) | (~w20986 & w25497) | (~w20988 & w25497);
assign w21175 = b[61] & w3785;
assign w21176 = b[62] & w3578;
assign w21177 = b[63] & w3580;
assign w21178 = ~w21176 & ~w21177;
assign w21179 = ~w21175 & w21178;
assign w21180 = (w12132 & w25605) | (w12132 & w25606) | (w25605 & w25606);
assign w21181 = ~a[35] & w25745;
assign w21182 = ~w21180 & ~w21181;
assign w21183 = ~w21174 & w21182;
assign w21184 = w21174 & ~w21182;
assign w21185 = ~w21183 & ~w21184;
assign w21186 = ~w21173 & ~w21185;
assign w21187 = w21173 & w21185;
assign w21188 = ~w21186 & ~w21187;
assign w21189 = ~w21013 & w21188;
assign w21190 = w21013 & ~w21188;
assign w21191 = ~w21189 & ~w21190;
assign w21192 = ~w21012 & ~w21191;
assign w21193 = (~w20820 & w24479) | (~w20820 & w24480) | (w24479 & w24480);
assign w21194 = ~w21192 & ~w21193;
assign w21195 = ~w21183 & ~w21187;
assign w21196 = b[59] & w4453;
assign w21197 = b[60] & w4241;
assign w21198 = b[61] & w4243;
assign w21199 = w4236 & w11400;
assign w21200 = ~w21197 & ~w21198;
assign w21201 = ~w21196 & w21200;
assign w21202 = ~w21199 & w21201;
assign w21203 = a[38] & ~w21202;
assign w21204 = ~a[38] & w21202;
assign w21205 = ~w21203 & ~w21204;
assign w21206 = ~w21136 & ~w21139;
assign w21207 = b[53] & w5939;
assign w21208 = b[55] & w5665;
assign w21209 = b[54] & w5670;
assign w21210 = w5663 & ~w9330;
assign w21211 = ~w21208 & ~w21209;
assign w21212 = ~w21207 & w21211;
assign w21213 = ~w21210 & w21212;
assign w21214 = a[44] & ~w21213;
assign w21215 = ~a[44] & w21213;
assign w21216 = ~w21214 & ~w21215;
assign w21217 = b[50] & w6732;
assign w21218 = b[51] & w6474;
assign w21219 = b[52] & w6476;
assign w21220 = w6469 & ~w8371;
assign w21221 = ~w21218 & ~w21219;
assign w21222 = ~w21217 & w21221;
assign w21223 = ~w21220 & w21222;
assign w21224 = a[47] & ~w21223;
assign w21225 = ~a[47] & w21223;
assign w21226 = ~w21224 & ~w21225;
assign w21227 = b[47] & w7586;
assign w21228 = b[48] & w7307;
assign w21229 = b[49] & w7314;
assign w21230 = w7312 & ~w7468;
assign w21231 = ~w21228 & ~w21229;
assign w21232 = ~w21227 & w21231;
assign w21233 = ~w21230 & w21232;
assign w21234 = a[50] & ~w21233;
assign w21235 = ~a[50] & w21233;
assign w21236 = ~w21234 & ~w21235;
assign w21237 = b[44] & w8515;
assign w21238 = b[46] & w8202;
assign w21239 = b[45] & w8200;
assign w21240 = ~w6613 & w8195;
assign w21241 = ~w21238 & ~w21239;
assign w21242 = ~w21237 & w21241;
assign w21243 = ~w21240 & w21242;
assign w21244 = a[53] & ~w21243;
assign w21245 = ~a[53] & w21243;
assign w21246 = ~w21244 & ~w21245;
assign w21247 = ~w21063 & ~w21066;
assign w21248 = b[38] & w10496;
assign w21249 = b[39] & w10146;
assign w21250 = b[40] & w10148;
assign w21251 = ~w5058 & w10141;
assign w21252 = ~w21249 & ~w21250;
assign w21253 = ~w21248 & w21252;
assign w21254 = ~w21251 & w21253;
assign w21255 = a[59] & ~w21254;
assign w21256 = ~a[59] & w21254;
assign w21257 = ~w21255 & ~w21256;
assign w21258 = ~w21057 & ~w21060;
assign w21259 = b[33] & w11921;
assign w21260 = b[34] & w11923;
assign w21261 = ~w21259 & ~w21260;
assign w21262 = ~w21050 & ~w21054;
assign w21263 = w21261 & ~w21262;
assign w21264 = ~w21261 & w21262;
assign w21265 = ~w21263 & ~w21264;
assign w21266 = b[35] & w11561;
assign w21267 = b[37] & w11196;
assign w21268 = b[36] & w11194;
assign w21269 = ~w4357 & w11189;
assign w21270 = ~w21267 & ~w21268;
assign w21271 = ~w21266 & w21270;
assign w21272 = ~w21269 & w21271;
assign w21273 = a[62] & ~w21272;
assign w21274 = ~a[62] & w21272;
assign w21275 = ~w21273 & ~w21274;
assign w21276 = ~w21265 & ~w21275;
assign w21277 = w21265 & w21275;
assign w21278 = ~w21276 & ~w21277;
assign w21279 = w21258 & ~w21278;
assign w21280 = ~w21258 & w21278;
assign w21281 = ~w21279 & ~w21280;
assign w21282 = w21257 & w21281;
assign w21283 = ~w21257 & ~w21281;
assign w21284 = ~w21282 & ~w21283;
assign w21285 = w21247 & ~w21284;
assign w21286 = ~w21247 & w21284;
assign w21287 = ~w21285 & ~w21286;
assign w21288 = b[41] & w9482;
assign w21289 = b[43] & w9160;
assign w21290 = b[42] & w9165;
assign w21291 = w5811 & w9158;
assign w21292 = ~w21289 & ~w21290;
assign w21293 = ~w21288 & w21292;
assign w21294 = ~w21291 & w21293;
assign w21295 = a[56] & ~w21294;
assign w21296 = ~a[56] & w21294;
assign w21297 = ~w21295 & ~w21296;
assign w21298 = w21287 & w21297;
assign w21299 = ~w21287 & ~w21297;
assign w21300 = ~w21298 & ~w21299;
assign w21301 = ~w21079 & ~w21084;
assign w21302 = w21300 & ~w21301;
assign w21303 = ~w21300 & w21301;
assign w21304 = ~w21302 & ~w21303;
assign w21305 = w21246 & w21304;
assign w21306 = ~w21246 & ~w21304;
assign w21307 = ~w21305 & ~w21306;
assign w21308 = ~w21096 & ~w21101;
assign w21309 = w21307 & ~w21308;
assign w21310 = ~w21307 & w21308;
assign w21311 = ~w21309 & ~w21310;
assign w21312 = w21236 & w21311;
assign w21313 = ~w21236 & ~w21311;
assign w21314 = ~w21312 & ~w21313;
assign w21315 = ~w21113 & ~w21118;
assign w21316 = w21314 & ~w21315;
assign w21317 = ~w21314 & w21315;
assign w21318 = ~w21316 & ~w21317;
assign w21319 = w21226 & w21318;
assign w21320 = ~w21226 & ~w21318;
assign w21321 = ~w21319 & ~w21320;
assign w21322 = ~w21130 & ~w21133;
assign w21323 = w21321 & w21322;
assign w21324 = ~w21321 & ~w21322;
assign w21325 = ~w21323 & ~w21324;
assign w21326 = w21216 & w21325;
assign w21327 = ~w21216 & ~w21325;
assign w21328 = ~w21326 & ~w21327;
assign w21329 = w21206 & ~w21328;
assign w21330 = ~w21206 & w21328;
assign w21331 = ~w21329 & ~w21330;
assign w21332 = b[56] & w5167;
assign w21333 = b[58] & w4925;
assign w21334 = b[57] & w4918;
assign w21335 = w4923 & ~w10339;
assign w21336 = ~w21333 & ~w21334;
assign w21337 = ~w21332 & w21336;
assign w21338 = ~w21335 & w21337;
assign w21339 = a[41] & ~w21338;
assign w21340 = ~a[41] & w21338;
assign w21341 = ~w21339 & ~w21340;
assign w21342 = w21331 & w21341;
assign w21343 = ~w21331 & ~w21341;
assign w21344 = ~w21342 & ~w21343;
assign w21345 = ~w21152 & ~w21157;
assign w21346 = w21344 & ~w21345;
assign w21347 = ~w21344 & w21345;
assign w21348 = ~w21346 & ~w21347;
assign w21349 = w21205 & w21348;
assign w21350 = ~w21205 & ~w21348;
assign w21351 = ~w21349 & ~w21350;
assign w21352 = ~w21167 & ~w21172;
assign w21353 = b[62] & w3785;
assign w21354 = b[63] & w3578;
assign w21355 = w3573 & w12156;
assign w21356 = ~w21353 & ~w21354;
assign w21357 = ~w21355 & w21356;
assign w21358 = a[35] & ~w21357;
assign w21359 = ~a[35] & w21357;
assign w21360 = ~w21358 & ~w21359;
assign w21361 = ~w21352 & w21360;
assign w21362 = w21352 & ~w21360;
assign w21363 = ~w21361 & ~w21362;
assign w21364 = w21351 & w21363;
assign w21365 = ~w21351 & ~w21363;
assign w21366 = ~w21364 & ~w21365;
assign w21367 = ~w21195 & w21366;
assign w21368 = w21195 & ~w21366;
assign w21369 = ~w21367 & ~w21368;
assign w21370 = (~w18109 & w25677) | (~w18109 & w25678) | (w25677 & w25678);
assign w21371 = (w20820 & w24483) | (w20820 & w24484) | (w24483 & w24484);
assign w21372 = ~w21369 & ~w21370;
assign w21373 = ~w21371 & ~w21372;
assign w21374 = ~w21361 & ~w21364;
assign w21375 = b[60] & w4453;
assign w21376 = b[62] & w4243;
assign w21377 = b[61] & w4241;
assign w21378 = w4236 & w11763;
assign w21379 = ~w21376 & ~w21377;
assign w21380 = ~w21375 & w21379;
assign w21381 = ~w21378 & w21380;
assign w21382 = a[38] & ~w21381;
assign w21383 = ~a[38] & w21381;
assign w21384 = ~w21382 & ~w21383;
assign w21385 = ~w21323 & ~w21326;
assign w21386 = b[54] & w5939;
assign w21387 = b[56] & w5665;
assign w21388 = b[55] & w5670;
assign w21389 = w5663 & w9657;
assign w21390 = ~w21387 & ~w21388;
assign w21391 = ~w21386 & w21390;
assign w21392 = ~w21389 & w21391;
assign w21393 = a[44] & ~w21392;
assign w21394 = ~a[44] & w21392;
assign w21395 = ~w21393 & ~w21394;
assign w21396 = ~w21316 & ~w21319;
assign w21397 = b[51] & w6732;
assign w21398 = b[53] & w6476;
assign w21399 = b[52] & w6474;
assign w21400 = w6469 & w8683;
assign w21401 = ~w21398 & ~w21399;
assign w21402 = ~w21397 & w21401;
assign w21403 = ~w21400 & w21402;
assign w21404 = a[47] & ~w21403;
assign w21405 = ~a[47] & w21403;
assign w21406 = ~w21404 & ~w21405;
assign w21407 = ~w21309 & ~w21312;
assign w21408 = b[48] & w7586;
assign w21409 = b[49] & w7307;
assign w21410 = b[50] & w7314;
assign w21411 = w7312 & w7759;
assign w21412 = ~w21409 & ~w21410;
assign w21413 = ~w21408 & w21412;
assign w21414 = ~w21411 & w21413;
assign w21415 = a[50] & ~w21414;
assign w21416 = ~a[50] & w21414;
assign w21417 = ~w21415 & ~w21416;
assign w21418 = ~w21286 & ~w21298;
assign w21419 = b[42] & w9482;
assign w21420 = b[44] & w9160;
assign w21421 = b[43] & w9165;
assign w21422 = w6069 & w9158;
assign w21423 = ~w21420 & ~w21421;
assign w21424 = ~w21419 & w21423;
assign w21425 = ~w21422 & w21424;
assign w21426 = a[56] & ~w21425;
assign w21427 = ~a[56] & w21425;
assign w21428 = ~w21426 & ~w21427;
assign w21429 = ~w21280 & ~w21282;
assign w21430 = b[39] & w10496;
assign w21431 = b[40] & w10146;
assign w21432 = b[41] & w10148;
assign w21433 = w5302 & w10141;
assign w21434 = ~w21431 & ~w21432;
assign w21435 = ~w21430 & w21434;
assign w21436 = ~w21433 & w21435;
assign w21437 = a[59] & ~w21436;
assign w21438 = ~a[59] & w21436;
assign w21439 = ~w21437 & ~w21438;
assign w21440 = b[36] & w11561;
assign w21441 = b[37] & w11194;
assign w21442 = b[38] & w11196;
assign w21443 = w4582 & w11189;
assign w21444 = ~w21441 & ~w21442;
assign w21445 = ~w21440 & w21444;
assign w21446 = ~w21443 & w21445;
assign w21447 = a[62] & ~w21446;
assign w21448 = ~a[62] & w21446;
assign w21449 = ~w21447 & ~w21448;
assign w21450 = ~w21263 & ~w21277;
assign w21451 = b[34] & w11921;
assign w21452 = b[35] & w11923;
assign w21453 = ~w21451 & ~w21452;
assign w21454 = w21261 & ~w21453;
assign w21455 = ~w21261 & w21453;
assign w21456 = ~w21454 & ~w21455;
assign w21457 = w21450 & w21456;
assign w21458 = ~w21450 & ~w21456;
assign w21459 = ~w21457 & ~w21458;
assign w21460 = w21449 & ~w21459;
assign w21461 = ~w21449 & w21459;
assign w21462 = ~w21460 & ~w21461;
assign w21463 = w21439 & w21462;
assign w21464 = ~w21439 & ~w21462;
assign w21465 = ~w21463 & ~w21464;
assign w21466 = ~w21429 & w21465;
assign w21467 = w21429 & ~w21465;
assign w21468 = ~w21466 & ~w21467;
assign w21469 = w21428 & w21468;
assign w21470 = ~w21428 & ~w21468;
assign w21471 = ~w21469 & ~w21470;
assign w21472 = w21418 & ~w21471;
assign w21473 = ~w21418 & w21471;
assign w21474 = ~w21472 & ~w21473;
assign w21475 = b[45] & w8515;
assign w21476 = b[47] & w8202;
assign w21477 = b[46] & w8200;
assign w21478 = w6889 & w8195;
assign w21479 = ~w21476 & ~w21477;
assign w21480 = ~w21475 & w21479;
assign w21481 = ~w21478 & w21480;
assign w21482 = a[53] & ~w21481;
assign w21483 = ~a[53] & w21481;
assign w21484 = ~w21482 & ~w21483;
assign w21485 = w21474 & w21484;
assign w21486 = ~w21474 & ~w21484;
assign w21487 = ~w21485 & ~w21486;
assign w21488 = ~w21302 & ~w21305;
assign w21489 = w21487 & ~w21488;
assign w21490 = ~w21487 & w21488;
assign w21491 = ~w21489 & ~w21490;
assign w21492 = ~w21417 & ~w21491;
assign w21493 = w21417 & w21491;
assign w21494 = ~w21492 & ~w21493;
assign w21495 = w21407 & ~w21494;
assign w21496 = ~w21407 & w21494;
assign w21497 = ~w21495 & ~w21496;
assign w21498 = w21406 & w21497;
assign w21499 = ~w21406 & ~w21497;
assign w21500 = ~w21498 & ~w21499;
assign w21501 = w21396 & ~w21500;
assign w21502 = ~w21396 & w21500;
assign w21503 = ~w21501 & ~w21502;
assign w21504 = w21395 & w21503;
assign w21505 = ~w21395 & ~w21503;
assign w21506 = ~w21504 & ~w21505;
assign w21507 = w21385 & ~w21506;
assign w21508 = ~w21385 & w21506;
assign w21509 = ~w21507 & ~w21508;
assign w21510 = b[57] & w5167;
assign w21511 = b[59] & w4925;
assign w21512 = b[58] & w4918;
assign w21513 = w4923 & w10371;
assign w21514 = ~w21511 & ~w21512;
assign w21515 = ~w21510 & w21514;
assign w21516 = ~w21513 & w21515;
assign w21517 = a[41] & ~w21516;
assign w21518 = ~a[41] & w21516;
assign w21519 = ~w21517 & ~w21518;
assign w21520 = w21509 & w21519;
assign w21521 = ~w21509 & ~w21519;
assign w21522 = ~w21520 & ~w21521;
assign w21523 = ~w21330 & ~w21342;
assign w21524 = w21522 & ~w21523;
assign w21525 = ~w21522 & w21523;
assign w21526 = ~w21524 & ~w21525;
assign w21527 = w21384 & w21526;
assign w21528 = ~w21384 & ~w21526;
assign w21529 = ~w21527 & ~w21528;
assign w21530 = ~w21346 & ~w21349;
assign w21531 = w3573 & ~w12154;
assign w21532 = ~w3785 & ~w21531;
assign w21533 = b[63] & ~w21532;
assign w21534 = ~a[35] & ~w21533;
assign w21535 = a[35] & w21533;
assign w21536 = ~w21534 & ~w21535;
assign w21537 = ~w21530 & w21536;
assign w21538 = w21530 & ~w21536;
assign w21539 = ~w21537 & ~w21538;
assign w21540 = w21529 & w21539;
assign w21541 = ~w21529 & ~w21539;
assign w21542 = ~w21540 & ~w21541;
assign w21543 = ~w21374 & w21542;
assign w21544 = w21374 & ~w21542;
assign w21545 = ~w21543 & ~w21544;
assign w21546 = (w18109 & w25679) | (w18109 & w25680) | (w25679 & w25680);
assign w21547 = (w20820 & w24487) | (w20820 & w24488) | (w24487 & w24488);
assign w21548 = ~w21545 & w21546;
assign w21549 = ~w21547 & ~w21548;
assign w21550 = (w18109 & w25681) | (w18109 & w25682) | (w25681 & w25682);
assign w21551 = ~w21496 & ~w21498;
assign w21552 = b[52] & w6732;
assign w21553 = b[53] & w6474;
assign w21554 = b[54] & w6476;
assign w21555 = w6469 & ~w8998;
assign w21556 = ~w21553 & ~w21554;
assign w21557 = ~w21552 & w21556;
assign w21558 = ~w21555 & w21557;
assign w21559 = a[47] & ~w21558;
assign w21560 = ~a[47] & w21558;
assign w21561 = ~w21559 & ~w21560;
assign w21562 = ~w21489 & ~w21493;
assign w21563 = ~w21466 & ~w21469;
assign w21564 = b[43] & w9482;
assign w21565 = b[45] & w9160;
assign w21566 = b[44] & w9165;
assign w21567 = w6334 & w9158;
assign w21568 = ~w21565 & ~w21566;
assign w21569 = ~w21564 & w21568;
assign w21570 = ~w21567 & w21569;
assign w21571 = a[56] & ~w21570;
assign w21572 = ~a[56] & w21570;
assign w21573 = ~w21571 & ~w21572;
assign w21574 = b[35] & w11921;
assign w21575 = b[36] & w11923;
assign w21576 = ~w21574 & ~w21575;
assign w21577 = ~a[35] & ~w21453;
assign w21578 = a[35] & w21453;
assign w21579 = ~w21577 & ~w21578;
assign w21580 = ~w21576 & w21579;
assign w21581 = w21576 & ~w21579;
assign w21582 = ~w21580 & ~w21581;
assign w21583 = ~w21454 & ~w21457;
assign w21584 = ~w21582 & ~w21583;
assign w21585 = w21582 & w21583;
assign w21586 = ~w21584 & ~w21585;
assign w21587 = b[37] & w11561;
assign w21588 = b[39] & w11196;
assign w21589 = b[38] & w11194;
assign w21590 = ~w4812 & w11189;
assign w21591 = ~w21588 & ~w21589;
assign w21592 = ~w21587 & w21591;
assign w21593 = ~w21590 & w21592;
assign w21594 = a[62] & ~w21593;
assign w21595 = ~a[62] & w21593;
assign w21596 = ~w21594 & ~w21595;
assign w21597 = ~w21586 & ~w21596;
assign w21598 = w21586 & w21596;
assign w21599 = ~w21597 & ~w21598;
assign w21600 = b[40] & w10496;
assign w21601 = b[42] & w10148;
assign w21602 = b[41] & w10146;
assign w21603 = w5548 & w10141;
assign w21604 = ~w21601 & ~w21602;
assign w21605 = ~w21600 & w21604;
assign w21606 = ~w21603 & w21605;
assign w21607 = a[59] & ~w21606;
assign w21608 = ~a[59] & w21606;
assign w21609 = ~w21607 & ~w21608;
assign w21610 = w21599 & w21609;
assign w21611 = ~w21599 & ~w21609;
assign w21612 = ~w21610 & ~w21611;
assign w21613 = ~w21460 & ~w21463;
assign w21614 = w21612 & ~w21613;
assign w21615 = ~w21612 & w21613;
assign w21616 = ~w21614 & ~w21615;
assign w21617 = w21573 & w21616;
assign w21618 = ~w21573 & ~w21616;
assign w21619 = ~w21617 & ~w21618;
assign w21620 = w21563 & ~w21619;
assign w21621 = ~w21563 & w21619;
assign w21622 = ~w21620 & ~w21621;
assign w21623 = b[46] & w8515;
assign w21624 = b[48] & w8202;
assign w21625 = b[47] & w8200;
assign w21626 = ~w7170 & w8195;
assign w21627 = ~w21624 & ~w21625;
assign w21628 = ~w21623 & w21627;
assign w21629 = ~w21626 & w21628;
assign w21630 = a[53] & ~w21629;
assign w21631 = ~a[53] & w21629;
assign w21632 = ~w21630 & ~w21631;
assign w21633 = w21622 & w21632;
assign w21634 = ~w21622 & ~w21632;
assign w21635 = ~w21633 & ~w21634;
assign w21636 = ~w21473 & ~w21485;
assign w21637 = ~w21635 & w21636;
assign w21638 = w21635 & ~w21636;
assign w21639 = ~w21637 & ~w21638;
assign w21640 = b[49] & w7586;
assign w21641 = b[51] & w7314;
assign w21642 = b[50] & w7307;
assign w21643 = w7312 & ~w8058;
assign w21644 = ~w21641 & ~w21642;
assign w21645 = ~w21640 & w21644;
assign w21646 = ~w21643 & w21645;
assign w21647 = a[50] & ~w21646;
assign w21648 = ~a[50] & w21646;
assign w21649 = ~w21647 & ~w21648;
assign w21650 = w21639 & w21649;
assign w21651 = ~w21639 & ~w21649;
assign w21652 = ~w21650 & ~w21651;
assign w21653 = ~w21562 & w21652;
assign w21654 = w21562 & ~w21652;
assign w21655 = ~w21653 & ~w21654;
assign w21656 = ~w21561 & ~w21655;
assign w21657 = w21561 & w21655;
assign w21658 = ~w21656 & ~w21657;
assign w21659 = ~w21551 & w21658;
assign w21660 = w21551 & ~w21658;
assign w21661 = ~w21659 & ~w21660;
assign w21662 = b[55] & w5939;
assign w21663 = b[56] & w5670;
assign w21664 = b[57] & w5665;
assign w21665 = ~w21663 & ~w21664;
assign w21666 = ~w21662 & w21665;
assign w21667 = (w21666 & w9992) | (w21666 & w25337) | (w9992 & w25337);
assign w21668 = a[44] & ~w21667;
assign w21669 = ~a[44] & w21667;
assign w21670 = ~w21668 & ~w21669;
assign w21671 = w21661 & w21670;
assign w21672 = ~w21661 & ~w21670;
assign w21673 = ~w21671 & ~w21672;
assign w21674 = ~w21502 & ~w21504;
assign w21675 = ~w21673 & w21674;
assign w21676 = w21673 & ~w21674;
assign w21677 = ~w21675 & ~w21676;
assign w21678 = b[58] & w5167;
assign w21679 = b[59] & w4918;
assign w21680 = b[60] & w4925;
assign w21681 = w4923 & w11035;
assign w21682 = ~w21679 & ~w21680;
assign w21683 = ~w21678 & w21682;
assign w21684 = ~w21681 & w21683;
assign w21685 = a[41] & ~w21684;
assign w21686 = ~a[41] & w21684;
assign w21687 = ~w21685 & ~w21686;
assign w21688 = w21677 & w21687;
assign w21689 = ~w21677 & ~w21687;
assign w21690 = ~w21688 & ~w21689;
assign w21691 = ~w21508 & ~w21520;
assign w21692 = ~w21690 & w21691;
assign w21693 = w21690 & ~w21691;
assign w21694 = ~w21692 & ~w21693;
assign w21695 = b[61] & w4453;
assign w21696 = b[62] & w4241;
assign w21697 = b[63] & w4243;
assign w21698 = w4236 & w12132;
assign w21699 = ~w21696 & ~w21697;
assign w21700 = ~w21695 & w21699;
assign w21701 = ~w21698 & w21700;
assign w21702 = a[38] & ~w21701;
assign w21703 = ~a[38] & w21701;
assign w21704 = ~w21702 & ~w21703;
assign w21705 = w21694 & w21704;
assign w21706 = ~w21694 & ~w21704;
assign w21707 = ~w21705 & ~w21706;
assign w21708 = ~w21524 & ~w21527;
assign w21709 = ~w21707 & w21708;
assign w21710 = w21707 & ~w21708;
assign w21711 = ~w21709 & ~w21710;
assign w21712 = ~w21537 & ~w21540;
assign w21713 = w21711 & ~w21712;
assign w21714 = ~w21711 & w21712;
assign w21715 = ~w21713 & ~w21714;
assign w21716 = ~w21550 & ~w21715;
assign w21717 = w21715 & w25746;
assign w21718 = ~w21716 & ~w21717;
assign w21719 = ~w21705 & ~w21710;
assign w21720 = b[59] & w5167;
assign w21721 = b[61] & w4925;
assign w21722 = b[60] & w4918;
assign w21723 = ~w21721 & ~w21722;
assign w21724 = ~w21720 & w21723;
assign w21725 = (w11400 & w25338) | (w11400 & w25339) | (w25338 & w25339);
assign w21726 = ~a[41] & w25747;
assign w21727 = ~w21725 & ~w21726;
assign w21728 = b[56] & w5939;
assign w21729 = b[57] & w5670;
assign w21730 = b[58] & w5665;
assign w21731 = ~w21729 & ~w21730;
assign w21732 = ~w21728 & w21731;
assign w21733 = (w21732 & w10339) | (w21732 & w25340) | (w10339 & w25340);
assign w21734 = a[44] & ~w21733;
assign w21735 = ~a[44] & w21733;
assign w21736 = ~w21734 & ~w21735;
assign w21737 = ~w21657 & ~w21659;
assign w21738 = b[53] & w6732;
assign w21739 = b[54] & w6474;
assign w21740 = b[55] & w6476;
assign w21741 = w6469 & ~w9330;
assign w21742 = ~w21739 & ~w21740;
assign w21743 = ~w21738 & w21742;
assign w21744 = ~w21741 & w21743;
assign w21745 = a[47] & ~w21744;
assign w21746 = ~a[47] & w21744;
assign w21747 = ~w21745 & ~w21746;
assign w21748 = b[50] & w7586;
assign w21749 = b[51] & w7307;
assign w21750 = b[52] & w7314;
assign w21751 = w7312 & ~w8371;
assign w21752 = ~w21749 & ~w21750;
assign w21753 = ~w21748 & w21752;
assign w21754 = ~w21751 & w21753;
assign w21755 = a[50] & ~w21754;
assign w21756 = ~a[50] & w21754;
assign w21757 = ~w21755 & ~w21756;
assign w21758 = b[47] & w8515;
assign w21759 = b[48] & w8200;
assign w21760 = b[49] & w8202;
assign w21761 = ~w7468 & w8195;
assign w21762 = ~w21759 & ~w21760;
assign w21763 = ~w21758 & w21762;
assign w21764 = ~w21761 & w21763;
assign w21765 = a[53] & ~w21764;
assign w21766 = ~a[53] & w21764;
assign w21767 = ~w21765 & ~w21766;
assign w21768 = b[44] & w9482;
assign w21769 = b[46] & w9160;
assign w21770 = b[45] & w9165;
assign w21771 = ~w6613 & w9158;
assign w21772 = ~w21769 & ~w21770;
assign w21773 = ~w21768 & w21772;
assign w21774 = ~w21771 & w21773;
assign w21775 = a[56] & ~w21774;
assign w21776 = ~a[56] & w21774;
assign w21777 = ~w21775 & ~w21776;
assign w21778 = b[41] & w10496;
assign w21779 = b[42] & w10146;
assign w21780 = b[43] & w10148;
assign w21781 = w5811 & w10141;
assign w21782 = ~w21779 & ~w21780;
assign w21783 = ~w21778 & w21782;
assign w21784 = ~w21781 & w21783;
assign w21785 = a[59] & ~w21784;
assign w21786 = ~a[59] & w21784;
assign w21787 = ~w21785 & ~w21786;
assign w21788 = ~w21585 & ~w21598;
assign w21789 = b[38] & w11561;
assign w21790 = b[40] & w11196;
assign w21791 = b[39] & w11194;
assign w21792 = ~w5058 & w11189;
assign w21793 = ~w21790 & ~w21791;
assign w21794 = ~w21789 & w21793;
assign w21795 = ~w21792 & w21794;
assign w21796 = a[62] & ~w21795;
assign w21797 = ~a[62] & w21795;
assign w21798 = ~w21796 & ~w21797;
assign w21799 = b[36] & w11921;
assign w21800 = b[37] & w11923;
assign w21801 = ~w21799 & ~w21800;
assign w21802 = ~w21577 & ~w21580;
assign w21803 = w21801 & ~w21802;
assign w21804 = ~w21801 & w21802;
assign w21805 = ~w21803 & ~w21804;
assign w21806 = w21798 & w21805;
assign w21807 = ~w21798 & ~w21805;
assign w21808 = ~w21806 & ~w21807;
assign w21809 = ~w21788 & w21808;
assign w21810 = w21788 & ~w21808;
assign w21811 = ~w21809 & ~w21810;
assign w21812 = w21787 & w21811;
assign w21813 = ~w21787 & ~w21811;
assign w21814 = ~w21812 & ~w21813;
assign w21815 = ~w21610 & ~w21614;
assign w21816 = w21814 & ~w21815;
assign w21817 = ~w21814 & w21815;
assign w21818 = ~w21816 & ~w21817;
assign w21819 = w21777 & w21818;
assign w21820 = ~w21777 & ~w21818;
assign w21821 = ~w21819 & ~w21820;
assign w21822 = ~w21617 & ~w21621;
assign w21823 = w21821 & ~w21822;
assign w21824 = ~w21821 & w21822;
assign w21825 = ~w21823 & ~w21824;
assign w21826 = w21767 & w21825;
assign w21827 = ~w21767 & ~w21825;
assign w21828 = ~w21826 & ~w21827;
assign w21829 = ~w21633 & ~w21638;
assign w21830 = w21828 & ~w21829;
assign w21831 = ~w21828 & w21829;
assign w21832 = ~w21830 & ~w21831;
assign w21833 = w21757 & w21832;
assign w21834 = ~w21757 & ~w21832;
assign w21835 = ~w21833 & ~w21834;
assign w21836 = ~w21650 & ~w21653;
assign w21837 = w21835 & ~w21836;
assign w21838 = ~w21835 & w21836;
assign w21839 = ~w21837 & ~w21838;
assign w21840 = w21747 & w21839;
assign w21841 = ~w21747 & ~w21839;
assign w21842 = ~w21840 & ~w21841;
assign w21843 = ~w21737 & w21842;
assign w21844 = w21737 & ~w21842;
assign w21845 = ~w21843 & ~w21844;
assign w21846 = w21736 & w21845;
assign w21847 = ~w21736 & ~w21845;
assign w21848 = ~w21846 & ~w21847;
assign w21849 = ~w21671 & ~w21676;
assign w21850 = w21848 & ~w21849;
assign w21851 = ~w21848 & w21849;
assign w21852 = ~w21850 & ~w21851;
assign w21853 = w21727 & w21852;
assign w21854 = ~w21727 & ~w21852;
assign w21855 = ~w21853 & ~w21854;
assign w21856 = ~w21688 & ~w21693;
assign w21857 = b[62] & w4453;
assign w21858 = b[63] & w4241;
assign w21859 = w4236 & w12156;
assign w21860 = ~w21857 & ~w21858;
assign w21861 = ~w21859 & w21860;
assign w21862 = ~a[38] & w21861;
assign w21863 = a[38] & ~w21861;
assign w21864 = ~w21862 & ~w21863;
assign w21865 = ~w21856 & w21864;
assign w21866 = w21856 & ~w21864;
assign w21867 = ~w21865 & ~w21866;
assign w21868 = w21855 & w21867;
assign w21869 = ~w21855 & ~w21867;
assign w21870 = ~w21868 & ~w21869;
assign w21871 = w21719 & ~w21870;
assign w21872 = ~w21719 & w21870;
assign w21873 = ~w21871 & ~w21872;
assign w21874 = (~w18109 & w25683) | (~w18109 & w25684) | (w25683 & w25684);
assign w21875 = (w20820 & w24495) | (w20820 & w24496) | (w24495 & w24496);
assign w21876 = ~w21873 & ~w21874;
assign w21877 = ~w21875 & ~w21876;
assign w21878 = ~w21865 & ~w21868;
assign w21879 = b[60] & w5167;
assign w21880 = b[62] & w4925;
assign w21881 = b[61] & w4918;
assign w21882 = ~w21880 & ~w21881;
assign w21883 = ~w21879 & w21882;
assign w21884 = (w21883 & ~w11763) | (w21883 & w25499) | (~w11763 & w25499);
assign w21885 = a[41] & ~w21884;
assign w21886 = ~a[41] & w21884;
assign w21887 = ~w21885 & ~w21886;
assign w21888 = ~w21837 & ~w21840;
assign w21889 = b[54] & w6732;
assign w21890 = b[55] & w6474;
assign w21891 = b[56] & w6476;
assign w21892 = ~w21890 & ~w21891;
assign w21893 = ~w21889 & w21892;
assign w21894 = (w21893 & ~w9657) | (w21893 & w25607) | (~w9657 & w25607);
assign w21895 = a[47] & ~w21894;
assign w21896 = ~a[47] & w21894;
assign w21897 = ~w21895 & ~w21896;
assign w21898 = ~w21830 & ~w21833;
assign w21899 = b[51] & w7586;
assign w21900 = b[53] & w7314;
assign w21901 = b[52] & w7307;
assign w21902 = w7312 & w8683;
assign w21903 = ~w21900 & ~w21901;
assign w21904 = ~w21899 & w21903;
assign w21905 = ~w21902 & w21904;
assign w21906 = a[50] & ~w21905;
assign w21907 = ~a[50] & w21905;
assign w21908 = ~w21906 & ~w21907;
assign w21909 = ~w21823 & ~w21826;
assign w21910 = b[45] & w9482;
assign w21911 = b[47] & w9160;
assign w21912 = b[46] & w9165;
assign w21913 = w6889 & w9158;
assign w21914 = ~w21911 & ~w21912;
assign w21915 = ~w21910 & w21914;
assign w21916 = ~w21913 & w21915;
assign w21917 = a[56] & ~w21916;
assign w21918 = ~a[56] & w21916;
assign w21919 = ~w21917 & ~w21918;
assign w21920 = ~w21809 & ~w21812;
assign w21921 = b[42] & w10496;
assign w21922 = b[44] & w10148;
assign w21923 = b[43] & w10146;
assign w21924 = w6069 & w10141;
assign w21925 = ~w21922 & ~w21923;
assign w21926 = ~w21921 & w21925;
assign w21927 = ~w21924 & w21926;
assign w21928 = a[59] & ~w21927;
assign w21929 = ~a[59] & w21927;
assign w21930 = ~w21928 & ~w21929;
assign w21931 = b[39] & w11561;
assign w21932 = b[41] & w11196;
assign w21933 = b[40] & w11194;
assign w21934 = w5302 & w11189;
assign w21935 = ~w21932 & ~w21933;
assign w21936 = ~w21931 & w21935;
assign w21937 = ~w21934 & w21936;
assign w21938 = a[62] & ~w21937;
assign w21939 = ~a[62] & w21937;
assign w21940 = ~w21938 & ~w21939;
assign w21941 = ~w21803 & ~w21806;
assign w21942 = b[37] & w11921;
assign w21943 = b[38] & w11923;
assign w21944 = ~w21942 & ~w21943;
assign w21945 = w21801 & ~w21944;
assign w21946 = ~w21801 & w21944;
assign w21947 = ~w21945 & ~w21946;
assign w21948 = ~w21941 & w21947;
assign w21949 = w21941 & ~w21947;
assign w21950 = ~w21948 & ~w21949;
assign w21951 = w21940 & w21950;
assign w21952 = ~w21940 & ~w21950;
assign w21953 = ~w21951 & ~w21952;
assign w21954 = w21930 & w21953;
assign w21955 = ~w21930 & ~w21953;
assign w21956 = ~w21954 & ~w21955;
assign w21957 = ~w21920 & w21956;
assign w21958 = w21920 & ~w21956;
assign w21959 = ~w21957 & ~w21958;
assign w21960 = w21919 & w21959;
assign w21961 = ~w21919 & ~w21959;
assign w21962 = ~w21960 & ~w21961;
assign w21963 = ~w21816 & ~w21819;
assign w21964 = w21962 & ~w21963;
assign w21965 = ~w21962 & w21963;
assign w21966 = ~w21964 & ~w21965;
assign w21967 = b[48] & w8515;
assign w21968 = b[50] & w8202;
assign w21969 = b[49] & w8200;
assign w21970 = w7759 & w8195;
assign w21971 = ~w21968 & ~w21969;
assign w21972 = ~w21967 & w21971;
assign w21973 = ~w21970 & w21972;
assign w21974 = a[53] & ~w21973;
assign w21975 = ~a[53] & w21973;
assign w21976 = ~w21974 & ~w21975;
assign w21977 = ~w21966 & ~w21976;
assign w21978 = w21966 & w21976;
assign w21979 = ~w21977 & ~w21978;
assign w21980 = w21909 & ~w21979;
assign w21981 = ~w21909 & w21979;
assign w21982 = ~w21980 & ~w21981;
assign w21983 = w21908 & w21982;
assign w21984 = ~w21908 & ~w21982;
assign w21985 = ~w21983 & ~w21984;
assign w21986 = w21898 & ~w21985;
assign w21987 = ~w21898 & w21985;
assign w21988 = ~w21986 & ~w21987;
assign w21989 = w21897 & w21988;
assign w21990 = ~w21897 & ~w21988;
assign w21991 = ~w21989 & ~w21990;
assign w21992 = w21888 & ~w21991;
assign w21993 = ~w21888 & w21991;
assign w21994 = ~w21992 & ~w21993;
assign w21995 = b[57] & w5939;
assign w21996 = b[59] & w5665;
assign w21997 = b[58] & w5670;
assign w21998 = ~w21996 & ~w21997;
assign w21999 = ~w21995 & w21998;
assign w22000 = (w10371 & w25500) | (w10371 & w25501) | (w25500 & w25501);
assign w22001 = ~a[44] & w25748;
assign w22002 = ~w22000 & ~w22001;
assign w22003 = w21994 & w22002;
assign w22004 = ~w21994 & ~w22002;
assign w22005 = ~w22003 & ~w22004;
assign w22006 = ~w21843 & ~w21846;
assign w22007 = w22005 & ~w22006;
assign w22008 = ~w22005 & w22006;
assign w22009 = ~w22007 & ~w22008;
assign w22010 = w21887 & w22009;
assign w22011 = ~w21887 & ~w22009;
assign w22012 = ~w22010 & ~w22011;
assign w22013 = ~w21850 & ~w21853;
assign w22014 = w4236 & ~w12154;
assign w22015 = ~w4453 & ~w22014;
assign w22016 = b[63] & ~w22015;
assign w22017 = ~a[38] & ~w22016;
assign w22018 = a[38] & w22016;
assign w22019 = ~w22017 & ~w22018;
assign w22020 = ~w22013 & w22019;
assign w22021 = w22013 & ~w22019;
assign w22022 = ~w22020 & ~w22021;
assign w22023 = w22012 & w22022;
assign w22024 = ~w22012 & ~w22022;
assign w22025 = ~w22023 & ~w22024;
assign w22026 = ~w21878 & w22025;
assign w22027 = w21878 & ~w22025;
assign w22028 = ~w22026 & ~w22027;
assign w22029 = (w18109 & w25685) | (w18109 & w25686) | (w25685 & w25686);
assign w22030 = (w20820 & w24499) | (w20820 & w24500) | (w24499 & w24500);
assign w22031 = ~w22028 & w22029;
assign w22032 = ~w22030 & ~w22031;
assign w22033 = (w18109 & w25687) | (w18109 & w25688) | (w25687 & w25688);
assign w22034 = ~w21981 & ~w21983;
assign w22035 = b[52] & w7586;
assign w22036 = b[54] & w7314;
assign w22037 = b[53] & w7307;
assign w22038 = ~w22036 & ~w22037;
assign w22039 = ~w22035 & w22038;
assign w22040 = a[50] & w25749;
assign w22041 = (w8998 & w25608) | (w8998 & w25609) | (w25608 & w25609);
assign w22042 = ~w22040 & ~w22041;
assign w22043 = ~w21964 & ~w21978;
assign w22044 = ~w21957 & ~w21960;
assign w22045 = b[46] & w9482;
assign w22046 = b[48] & w9160;
assign w22047 = b[47] & w9165;
assign w22048 = ~w22046 & ~w22047;
assign w22049 = ~w22045 & w22048;
assign w22050 = (w22049 & w7170) | (w22049 & w25610) | (w7170 & w25610);
assign w22051 = a[56] & ~w22050;
assign w22052 = ~a[56] & w22050;
assign w22053 = ~w22051 & ~w22052;
assign w22054 = ~w21951 & ~w21954;
assign w22055 = ~w21945 & ~w21948;
assign w22056 = b[38] & w11921;
assign w22057 = b[39] & w11923;
assign w22058 = ~w22056 & ~w22057;
assign w22059 = ~a[38] & ~w21801;
assign w22060 = a[38] & w21801;
assign w22061 = ~w22059 & ~w22060;
assign w22062 = ~w22058 & w22061;
assign w22063 = w22058 & ~w22061;
assign w22064 = ~w22062 & ~w22063;
assign w22065 = w22055 & ~w22064;
assign w22066 = ~w22055 & w22064;
assign w22067 = ~w22065 & ~w22066;
assign w22068 = b[40] & w11561;
assign w22069 = b[41] & w11194;
assign w22070 = b[42] & w11196;
assign w22071 = w5548 & w11189;
assign w22072 = ~w22069 & ~w22070;
assign w22073 = ~w22068 & w22072;
assign w22074 = ~w22071 & w22073;
assign w22075 = a[62] & ~w22074;
assign w22076 = ~a[62] & w22074;
assign w22077 = ~w22075 & ~w22076;
assign w22078 = w22067 & w22077;
assign w22079 = ~w22067 & ~w22077;
assign w22080 = ~w22078 & ~w22079;
assign w22081 = b[43] & w10496;
assign w22082 = b[44] & w10146;
assign w22083 = b[45] & w10148;
assign w22084 = w6334 & w10141;
assign w22085 = ~w22082 & ~w22083;
assign w22086 = ~w22081 & w22085;
assign w22087 = ~w22084 & w22086;
assign w22088 = a[59] & ~w22087;
assign w22089 = ~a[59] & w22087;
assign w22090 = ~w22088 & ~w22089;
assign w22091 = w22080 & w22090;
assign w22092 = ~w22080 & ~w22090;
assign w22093 = ~w22091 & ~w22092;
assign w22094 = ~w22054 & w22093;
assign w22095 = w22054 & ~w22093;
assign w22096 = ~w22094 & ~w22095;
assign w22097 = w22053 & w22096;
assign w22098 = ~w22053 & ~w22096;
assign w22099 = ~w22097 & ~w22098;
assign w22100 = w22044 & ~w22099;
assign w22101 = ~w22044 & w22099;
assign w22102 = ~w22100 & ~w22101;
assign w22103 = b[49] & w8515;
assign w22104 = b[50] & w8200;
assign w22105 = b[51] & w8202;
assign w22106 = ~w22104 & ~w22105;
assign w22107 = ~w22103 & w22106;
assign w22108 = (w22107 & w8058) | (w22107 & w25611) | (w8058 & w25611);
assign w22109 = a[53] & ~w22108;
assign w22110 = ~a[53] & w22108;
assign w22111 = ~w22109 & ~w22110;
assign w22112 = w22102 & w22111;
assign w22113 = ~w22102 & ~w22111;
assign w22114 = ~w22112 & ~w22113;
assign w22115 = ~w22043 & w22114;
assign w22116 = w22043 & ~w22114;
assign w22117 = ~w22115 & ~w22116;
assign w22118 = ~w22042 & ~w22117;
assign w22119 = w22042 & w22117;
assign w22120 = ~w22118 & ~w22119;
assign w22121 = ~w22034 & w22120;
assign w22122 = w22034 & ~w22120;
assign w22123 = ~w22121 & ~w22122;
assign w22124 = b[55] & w6732;
assign w22125 = b[56] & w6474;
assign w22126 = b[57] & w6476;
assign w22127 = ~w22125 & ~w22126;
assign w22128 = ~w22124 & w22127;
assign w22129 = a[47] & w25750;
assign w22130 = (w9992 & w25503) | (w9992 & w25504) | (w25503 & w25504);
assign w22131 = ~w22129 & ~w22130;
assign w22132 = w22123 & w22131;
assign w22133 = ~w22123 & ~w22131;
assign w22134 = ~w22132 & ~w22133;
assign w22135 = ~w21987 & ~w21989;
assign w22136 = ~w22134 & w22135;
assign w22137 = w22134 & ~w22135;
assign w22138 = ~w22136 & ~w22137;
assign w22139 = b[58] & w5939;
assign w22140 = b[59] & w5670;
assign w22141 = b[60] & w5665;
assign w22142 = ~w22140 & ~w22141;
assign w22143 = ~w22139 & w22142;
assign w22144 = (w11035 & w25221) | (w11035 & w25222) | (w25221 & w25222);
assign w22145 = (~w11035 & w25223) | (~w11035 & w25224) | (w25223 & w25224);
assign w22146 = ~w22144 & ~w22145;
assign w22147 = w22138 & w22146;
assign w22148 = ~w22138 & ~w22146;
assign w22149 = ~w22147 & ~w22148;
assign w22150 = ~w21993 & ~w22003;
assign w22151 = ~w22149 & w22150;
assign w22152 = w22149 & ~w22150;
assign w22153 = ~w22151 & ~w22152;
assign w22154 = b[61] & w5167;
assign w22155 = b[63] & w4925;
assign w22156 = b[62] & w4918;
assign w22157 = ~w22155 & ~w22156;
assign w22158 = ~w22154 & w22157;
assign w22159 = (w22158 & ~w12132) | (w22158 & w25038) | (~w12132 & w25038);
assign w22160 = a[41] & ~w22159;
assign w22161 = ~a[41] & w22159;
assign w22162 = ~w22160 & ~w22161;
assign w22163 = w22153 & w22162;
assign w22164 = ~w22153 & ~w22162;
assign w22165 = ~w22163 & ~w22164;
assign w22166 = ~w22007 & ~w22010;
assign w22167 = ~w22165 & w22166;
assign w22168 = w22165 & ~w22166;
assign w22169 = ~w22167 & ~w22168;
assign w22170 = ~w22020 & ~w22023;
assign w22171 = w22169 & ~w22170;
assign w22172 = ~w22169 & w22170;
assign w22173 = ~w22171 & ~w22172;
assign w22174 = ~w22033 & ~w22173;
assign w22175 = (w18109 & w25689) | (w18109 & w25690) | (w25689 & w25690);
assign w22176 = ~w22174 & ~w22175;
assign w22177 = (~w22163 & ~w22165) | (~w22163 & w25343) | (~w22165 & w25343);
assign w22178 = b[59] & w5939;
assign w22179 = b[61] & w5665;
assign w22180 = b[60] & w5670;
assign w22181 = ~w22179 & ~w22180;
assign w22182 = ~w22178 & w22181;
assign w22183 = (w11400 & w25344) | (w11400 & w25345) | (w25344 & w25345);
assign w22184 = (~w11400 & w25346) | (~w11400 & w25347) | (w25346 & w25347);
assign w22185 = ~w22183 & ~w22184;
assign w22186 = b[56] & w6732;
assign w22187 = b[57] & w6474;
assign w22188 = b[58] & w6476;
assign w22189 = ~w22187 & ~w22188;
assign w22190 = ~w22186 & w22189;
assign w22191 = (~w10339 & w25505) | (~w10339 & w25506) | (w25505 & w25506);
assign w22192 = (w10339 & w25507) | (w10339 & w25508) | (w25507 & w25508);
assign w22193 = ~w22191 & ~w22192;
assign w22194 = ~w22119 & ~w22121;
assign w22195 = b[53] & w7586;
assign w22196 = b[55] & w7314;
assign w22197 = b[54] & w7307;
assign w22198 = ~w22196 & ~w22197;
assign w22199 = ~w22195 & w22198;
assign w22200 = (w22199 & w9330) | (w22199 & w25612) | (w9330 & w25612);
assign w22201 = a[50] & ~w22200;
assign w22202 = ~a[50] & w22200;
assign w22203 = ~w22201 & ~w22202;
assign w22204 = b[50] & w8515;
assign w22205 = b[51] & w8200;
assign w22206 = b[52] & w8202;
assign w22207 = ~w22205 & ~w22206;
assign w22208 = ~w22204 & w22207;
assign w22209 = (w22208 & w8371) | (w22208 & w25613) | (w8371 & w25613);
assign w22210 = a[53] & ~w22209;
assign w22211 = ~a[53] & w22209;
assign w22212 = ~w22210 & ~w22211;
assign w22213 = b[47] & w9482;
assign w22214 = b[49] & w9160;
assign w22215 = b[48] & w9165;
assign w22216 = ~w22214 & ~w22215;
assign w22217 = ~w22213 & w22216;
assign w22218 = (w22217 & w7468) | (w22217 & w25614) | (w7468 & w25614);
assign w22219 = a[56] & ~w22218;
assign w22220 = ~a[56] & w22218;
assign w22221 = ~w22219 & ~w22220;
assign w22222 = ~w22066 & ~w22078;
assign w22223 = b[39] & w11921;
assign w22224 = b[40] & w11923;
assign w22225 = ~w22223 & ~w22224;
assign w22226 = ~w22059 & ~w22062;
assign w22227 = w22225 & ~w22226;
assign w22228 = ~w22225 & w22226;
assign w22229 = ~w22227 & ~w22228;
assign w22230 = b[41] & w11561;
assign w22231 = b[42] & w11194;
assign w22232 = b[43] & w11196;
assign w22233 = w5811 & w11189;
assign w22234 = ~w22231 & ~w22232;
assign w22235 = ~w22230 & w22234;
assign w22236 = ~w22233 & w22235;
assign w22237 = a[62] & ~w22236;
assign w22238 = ~a[62] & w22236;
assign w22239 = ~w22237 & ~w22238;
assign w22240 = w22229 & w22239;
assign w22241 = ~w22229 & ~w22239;
assign w22242 = ~w22240 & ~w22241;
assign w22243 = w22222 & ~w22242;
assign w22244 = ~w22222 & w22242;
assign w22245 = ~w22243 & ~w22244;
assign w22246 = b[44] & w10496;
assign w22247 = b[46] & w10148;
assign w22248 = b[45] & w10146;
assign w22249 = ~w6613 & w10141;
assign w22250 = ~w22247 & ~w22248;
assign w22251 = ~w22246 & w22250;
assign w22252 = ~w22249 & w22251;
assign w22253 = a[59] & ~w22252;
assign w22254 = ~a[59] & w22252;
assign w22255 = ~w22253 & ~w22254;
assign w22256 = w22245 & w22255;
assign w22257 = ~w22245 & ~w22255;
assign w22258 = ~w22256 & ~w22257;
assign w22259 = ~w22091 & ~w22094;
assign w22260 = w22258 & ~w22259;
assign w22261 = ~w22258 & w22259;
assign w22262 = ~w22260 & ~w22261;
assign w22263 = w22221 & w22262;
assign w22264 = ~w22221 & ~w22262;
assign w22265 = ~w22263 & ~w22264;
assign w22266 = ~w22097 & ~w22101;
assign w22267 = w22265 & ~w22266;
assign w22268 = ~w22265 & w22266;
assign w22269 = ~w22267 & ~w22268;
assign w22270 = w22212 & w22269;
assign w22271 = ~w22212 & ~w22269;
assign w22272 = ~w22270 & ~w22271;
assign w22273 = ~w22112 & ~w22115;
assign w22274 = w22272 & ~w22273;
assign w22275 = ~w22272 & w22273;
assign w22276 = ~w22274 & ~w22275;
assign w22277 = w22203 & w22276;
assign w22278 = ~w22203 & ~w22276;
assign w22279 = ~w22277 & ~w22278;
assign w22280 = ~w22194 & w22279;
assign w22281 = w22194 & ~w22279;
assign w22282 = ~w22280 & ~w22281;
assign w22283 = w22193 & w22282;
assign w22284 = ~w22193 & ~w22282;
assign w22285 = ~w22283 & ~w22284;
assign w22286 = (~w22132 & ~w22134) | (~w22132 & w25615) | (~w22134 & w25615);
assign w22287 = w22285 & ~w22286;
assign w22288 = ~w22285 & w22286;
assign w22289 = ~w22287 & ~w22288;
assign w22290 = w22185 & w22289;
assign w22291 = ~w22185 & ~w22289;
assign w22292 = ~w22290 & ~w22291;
assign w22293 = (~w22147 & ~w22149) | (~w22147 & w25349) | (~w22149 & w25349);
assign w22294 = b[62] & w5167;
assign w22295 = b[63] & w4918;
assign w22296 = ~w12153 & w24726;
assign w22297 = ~w22294 & ~w22295;
assign w22298 = ~w22296 & w25040;
assign w22299 = (a[41] & w22296) | (a[41] & w25041) | (w22296 & w25041);
assign w22300 = ~w22298 & ~w22299;
assign w22301 = ~w22293 & w22300;
assign w22302 = w22293 & ~w22300;
assign w22303 = ~w22301 & ~w22302;
assign w22304 = w22292 & w22303;
assign w22305 = ~w22292 & ~w22303;
assign w22306 = ~w22304 & ~w22305;
assign w22307 = w22177 & ~w22306;
assign w22308 = ~w22177 & w22306;
assign w22309 = ~w22307 & ~w22308;
assign w22310 = ~w22175 & w24505;
assign w22311 = (~w20820 & w25691) | (~w20820 & w25692) | (w25691 & w25692);
assign w22312 = ~w22310 & ~w22311;
assign w22313 = (~w22301 & ~w22303) | (~w22301 & w25509) | (~w22303 & w25509);
assign w22314 = b[60] & w5939;
assign w22315 = b[61] & w5670;
assign w22316 = b[62] & w5665;
assign w22317 = ~w22315 & ~w22316;
assign w22318 = ~w22314 & w22317;
assign w22319 = (w11763 & w25616) | (w11763 & w25617) | (w25616 & w25617);
assign w22320 = ~a[44] & w25751;
assign w22321 = ~w22319 & ~w22320;
assign w22322 = ~w22274 & ~w22277;
assign w22323 = b[54] & w7586;
assign w22324 = b[56] & w7314;
assign w22325 = b[55] & w7307;
assign w22326 = ~w22324 & ~w22325;
assign w22327 = ~w22323 & w22326;
assign w22328 = (w22327 & ~w9657) | (w22327 & w25618) | (~w9657 & w25618);
assign w22329 = a[50] & ~w22328;
assign w22330 = ~a[50] & w22328;
assign w22331 = ~w22329 & ~w22330;
assign w22332 = ~w22267 & ~w22270;
assign w22333 = b[51] & w8515;
assign w22334 = b[53] & w8202;
assign w22335 = b[52] & w8200;
assign w22336 = w8195 & w8683;
assign w22337 = ~w22334 & ~w22335;
assign w22338 = ~w22333 & w22337;
assign w22339 = ~w22336 & w22338;
assign w22340 = a[53] & ~w22339;
assign w22341 = ~a[53] & w22339;
assign w22342 = ~w22340 & ~w22341;
assign w22343 = ~w22260 & ~w22263;
assign w22344 = ~w22244 & ~w22256;
assign w22345 = b[45] & w10496;
assign w22346 = b[47] & w10148;
assign w22347 = b[46] & w10146;
assign w22348 = w6889 & w10141;
assign w22349 = ~w22346 & ~w22347;
assign w22350 = ~w22345 & w22349;
assign w22351 = ~w22348 & w22350;
assign w22352 = a[59] & ~w22351;
assign w22353 = ~a[59] & w22351;
assign w22354 = ~w22352 & ~w22353;
assign w22355 = b[42] & w11561;
assign w22356 = b[44] & w11196;
assign w22357 = b[43] & w11194;
assign w22358 = w6069 & w11189;
assign w22359 = ~w22356 & ~w22357;
assign w22360 = ~w22355 & w22359;
assign w22361 = ~w22358 & w22360;
assign w22362 = a[62] & ~w22361;
assign w22363 = ~a[62] & w22361;
assign w22364 = ~w22362 & ~w22363;
assign w22365 = ~w22227 & ~w22240;
assign w22366 = b[40] & w11921;
assign w22367 = b[41] & w11923;
assign w22368 = ~w22366 & ~w22367;
assign w22369 = w22225 & ~w22368;
assign w22370 = ~w22225 & w22368;
assign w22371 = ~w22369 & ~w22370;
assign w22372 = ~w22365 & w22371;
assign w22373 = w22365 & ~w22371;
assign w22374 = ~w22372 & ~w22373;
assign w22375 = w22364 & w22374;
assign w22376 = ~w22364 & ~w22374;
assign w22377 = ~w22375 & ~w22376;
assign w22378 = w22354 & w22377;
assign w22379 = ~w22354 & ~w22377;
assign w22380 = ~w22378 & ~w22379;
assign w22381 = w22344 & ~w22380;
assign w22382 = ~w22344 & w22380;
assign w22383 = ~w22381 & ~w22382;
assign w22384 = b[48] & w9482;
assign w22385 = b[49] & w9165;
assign w22386 = b[50] & w9160;
assign w22387 = w7759 & w9158;
assign w22388 = ~w22385 & ~w22386;
assign w22389 = ~w22384 & w22388;
assign w22390 = ~w22387 & w22389;
assign w22391 = a[56] & ~w22390;
assign w22392 = ~a[56] & w22390;
assign w22393 = ~w22391 & ~w22392;
assign w22394 = ~w22383 & ~w22393;
assign w22395 = w22383 & w22393;
assign w22396 = ~w22394 & ~w22395;
assign w22397 = w22343 & ~w22396;
assign w22398 = ~w22343 & w22396;
assign w22399 = ~w22397 & ~w22398;
assign w22400 = w22342 & w22399;
assign w22401 = ~w22342 & ~w22399;
assign w22402 = ~w22400 & ~w22401;
assign w22403 = w22332 & ~w22402;
assign w22404 = ~w22332 & w22402;
assign w22405 = ~w22403 & ~w22404;
assign w22406 = w22331 & w22405;
assign w22407 = ~w22331 & ~w22405;
assign w22408 = ~w22406 & ~w22407;
assign w22409 = w22322 & ~w22408;
assign w22410 = ~w22322 & w22408;
assign w22411 = ~w22409 & ~w22410;
assign w22412 = b[57] & w6732;
assign w22413 = b[59] & w6476;
assign w22414 = b[58] & w6474;
assign w22415 = ~w22413 & ~w22414;
assign w22416 = ~w22412 & w22415;
assign w22417 = (w10371 & w25511) | (w10371 & w25512) | (w25511 & w25512);
assign w22418 = (~w10371 & w25513) | (~w10371 & w25514) | (w25513 & w25514);
assign w22419 = ~w22417 & ~w22418;
assign w22420 = w22411 & w22419;
assign w22421 = ~w22411 & ~w22419;
assign w22422 = ~w22420 & ~w22421;
assign w22423 = ~w22280 & ~w22283;
assign w22424 = w22422 & ~w22423;
assign w22425 = ~w22422 & w22423;
assign w22426 = ~w22424 & ~w22425;
assign w22427 = w22321 & w22426;
assign w22428 = ~w22321 & ~w22426;
assign w22429 = ~w22427 & ~w22428;
assign w22430 = (~w22287 & ~w22185) | (~w22287 & w25515) | (~w22185 & w25515);
assign w22431 = (w25517 & w25516) | (w25517 & ~w11757) | (w25516 & ~w11757);
assign w22432 = ~w5167 & ~w22431;
assign w22433 = b[63] & ~w22432;
assign w22434 = ~a[41] & ~w22433;
assign w22435 = a[41] & w22433;
assign w22436 = ~w22434 & ~w22435;
assign w22437 = ~w22430 & w22436;
assign w22438 = w22430 & ~w22436;
assign w22439 = ~w22437 & ~w22438;
assign w22440 = w22429 & w22439;
assign w22441 = ~w22429 & ~w22439;
assign w22442 = ~w22440 & ~w22441;
assign w22443 = ~w22313 & w22442;
assign w22444 = w22313 & ~w22442;
assign w22445 = ~w22443 & ~w22444;
assign w22446 = (~w22175 & w24507) | (~w22175 & w24508) | (w24507 & w24508);
assign w22447 = (~w20820 & w25693) | (~w20820 & w25694) | (w25693 & w25694);
assign w22448 = ~w22446 & ~w22447;
assign w22449 = ~w22404 & ~w22406;
assign w22450 = b[55] & w7586;
assign w22451 = b[57] & w7314;
assign w22452 = b[56] & w7307;
assign w22453 = ~w22451 & ~w22452;
assign w22454 = ~w22450 & w22453;
assign w22455 = (w22454 & w9992) | (w22454 & w25619) | (w9992 & w25619);
assign w22456 = a[50] & ~w22455;
assign w22457 = ~a[50] & w22455;
assign w22458 = ~w22456 & ~w22457;
assign w22459 = ~w22398 & ~w22400;
assign w22460 = b[52] & w8515;
assign w22461 = b[53] & w8200;
assign w22462 = b[54] & w8202;
assign w22463 = w8195 & ~w8998;
assign w22464 = ~w22461 & ~w22462;
assign w22465 = ~w22460 & w22464;
assign w22466 = ~w22463 & w22465;
assign w22467 = a[53] & ~w22466;
assign w22468 = ~a[53] & w22466;
assign w22469 = ~w22467 & ~w22468;
assign w22470 = ~w22382 & ~w22395;
assign w22471 = b[49] & w9482;
assign w22472 = b[51] & w9160;
assign w22473 = b[50] & w9165;
assign w22474 = ~w8058 & w9158;
assign w22475 = ~w22472 & ~w22473;
assign w22476 = ~w22471 & w22475;
assign w22477 = ~w22474 & w22476;
assign w22478 = a[56] & ~w22477;
assign w22479 = ~a[56] & w22477;
assign w22480 = ~w22478 & ~w22479;
assign w22481 = b[41] & w11921;
assign w22482 = b[42] & w11923;
assign w22483 = ~w22481 & ~w22482;
assign w22484 = ~a[41] & ~w22225;
assign w22485 = a[41] & w22225;
assign w22486 = ~w22484 & ~w22485;
assign w22487 = w22483 & ~w22486;
assign w22488 = ~w22483 & w22486;
assign w22489 = ~w22487 & ~w22488;
assign w22490 = b[43] & w11561;
assign w22491 = b[45] & w11196;
assign w22492 = b[44] & w11194;
assign w22493 = w6334 & w11189;
assign w22494 = ~w22491 & ~w22492;
assign w22495 = ~w22490 & w22494;
assign w22496 = ~w22493 & w22495;
assign w22497 = a[62] & ~w22496;
assign w22498 = ~a[62] & w22496;
assign w22499 = ~w22497 & ~w22498;
assign w22500 = w22489 & w22499;
assign w22501 = ~w22489 & ~w22499;
assign w22502 = ~w22500 & ~w22501;
assign w22503 = ~w22369 & ~w22372;
assign w22504 = ~w22502 & w22503;
assign w22505 = w22502 & ~w22503;
assign w22506 = ~w22504 & ~w22505;
assign w22507 = b[46] & w10496;
assign w22508 = b[48] & w10148;
assign w22509 = b[47] & w10146;
assign w22510 = ~w7170 & w10141;
assign w22511 = ~w22508 & ~w22509;
assign w22512 = ~w22507 & w22511;
assign w22513 = ~w22510 & w22512;
assign w22514 = a[59] & ~w22513;
assign w22515 = ~a[59] & w22513;
assign w22516 = ~w22514 & ~w22515;
assign w22517 = w22506 & w22516;
assign w22518 = ~w22506 & ~w22516;
assign w22519 = ~w22517 & ~w22518;
assign w22520 = ~w22375 & ~w22378;
assign w22521 = w22519 & ~w22520;
assign w22522 = ~w22519 & w22520;
assign w22523 = ~w22521 & ~w22522;
assign w22524 = ~w22480 & ~w22523;
assign w22525 = w22480 & w22523;
assign w22526 = ~w22524 & ~w22525;
assign w22527 = ~w22470 & w22526;
assign w22528 = w22470 & ~w22526;
assign w22529 = ~w22527 & ~w22528;
assign w22530 = w22469 & w22529;
assign w22531 = ~w22469 & ~w22529;
assign w22532 = ~w22530 & ~w22531;
assign w22533 = ~w22459 & w22532;
assign w22534 = w22459 & ~w22532;
assign w22535 = ~w22533 & ~w22534;
assign w22536 = ~w22458 & ~w22535;
assign w22537 = w22458 & w22535;
assign w22538 = ~w22536 & ~w22537;
assign w22539 = ~w22449 & w22538;
assign w22540 = w22449 & ~w22538;
assign w22541 = ~w22539 & ~w22540;
assign w22542 = b[58] & w6732;
assign w22543 = b[59] & w6474;
assign w22544 = b[60] & w6476;
assign w22545 = ~w22543 & ~w22544;
assign w22546 = ~w22542 & w22545;
assign w22547 = (w11035 & w25518) | (w11035 & w25519) | (w25518 & w25519);
assign w22548 = (~w11035 & w25520) | (~w11035 & w25521) | (w25520 & w25521);
assign w22549 = ~w22547 & ~w22548;
assign w22550 = w22541 & w22549;
assign w22551 = ~w22541 & ~w22549;
assign w22552 = ~w22550 & ~w22551;
assign w22553 = ~w22410 & ~w22420;
assign w22554 = ~w22552 & w22553;
assign w22555 = w22552 & ~w22553;
assign w22556 = ~w22554 & ~w22555;
assign w22557 = b[61] & w5939;
assign w22558 = b[63] & w5665;
assign w22559 = b[62] & w5670;
assign w22560 = ~w22558 & ~w22559;
assign w22561 = ~w22557 & w22560;
assign w22562 = (w22561 & ~w12132) | (w22561 & w25620) | (~w12132 & w25620);
assign w22563 = a[44] & ~w22562;
assign w22564 = ~a[44] & w22562;
assign w22565 = ~w22563 & ~w22564;
assign w22566 = w22556 & w22565;
assign w22567 = ~w22556 & ~w22565;
assign w22568 = ~w22566 & ~w22567;
assign w22569 = ~w22424 & ~w22427;
assign w22570 = ~w22568 & w22569;
assign w22571 = w22568 & ~w22569;
assign w22572 = ~w22570 & ~w22571;
assign w22573 = ~w22437 & ~w22440;
assign w22574 = w22572 & ~w22573;
assign w22575 = ~w22572 & w22573;
assign w22576 = ~w22574 & ~w22575;
assign w22577 = (w20820 & w25695) | (w20820 & w25696) | (w25695 & w25696);
assign w22578 = (w22175 & w24511) | (w22175 & w24512) | (w24511 & w24512);
assign w22579 = ~w22577 & ~w22578;
assign w22580 = b[59] & w6732;
assign w22581 = b[60] & w6474;
assign w22582 = b[61] & w6476;
assign w22583 = w6469 & w11400;
assign w22584 = ~w22581 & ~w22582;
assign w22585 = ~w22580 & w22584;
assign w22586 = ~w22583 & w22585;
assign w22587 = a[47] & ~w22586;
assign w22588 = ~a[47] & w22586;
assign w22589 = ~w22587 & ~w22588;
assign w22590 = ~w22537 & ~w22539;
assign w22591 = b[56] & w7586;
assign w22592 = b[57] & w7307;
assign w22593 = b[58] & w7314;
assign w22594 = w7312 & ~w10339;
assign w22595 = ~w22592 & ~w22593;
assign w22596 = ~w22591 & w22595;
assign w22597 = ~w22594 & w22596;
assign w22598 = a[50] & ~w22597;
assign w22599 = ~a[50] & w22597;
assign w22600 = ~w22598 & ~w22599;
assign w22601 = ~w22530 & ~w22533;
assign w22602 = b[53] & w8515;
assign w22603 = b[55] & w8202;
assign w22604 = b[54] & w8200;
assign w22605 = w8195 & ~w9330;
assign w22606 = ~w22603 & ~w22604;
assign w22607 = ~w22602 & w22606;
assign w22608 = ~w22605 & w22607;
assign w22609 = a[53] & ~w22608;
assign w22610 = ~a[53] & w22608;
assign w22611 = ~w22609 & ~w22610;
assign w22612 = b[50] & w9482;
assign w22613 = b[52] & w9160;
assign w22614 = b[51] & w9165;
assign w22615 = ~w8371 & w9158;
assign w22616 = ~w22613 & ~w22614;
assign w22617 = ~w22612 & w22616;
assign w22618 = ~w22615 & w22617;
assign w22619 = a[56] & ~w22618;
assign w22620 = ~a[56] & w22618;
assign w22621 = ~w22619 & ~w22620;
assign w22622 = ~w22500 & ~w22505;
assign w22623 = b[42] & w11921;
assign w22624 = b[43] & w11923;
assign w22625 = ~w22623 & ~w22624;
assign w22626 = ~w22484 & ~w22488;
assign w22627 = w22625 & ~w22626;
assign w22628 = ~w22625 & w22626;
assign w22629 = ~w22627 & ~w22628;
assign w22630 = b[44] & w11561;
assign w22631 = b[45] & w11194;
assign w22632 = b[46] & w11196;
assign w22633 = ~w6613 & w11189;
assign w22634 = ~w22631 & ~w22632;
assign w22635 = ~w22630 & w22634;
assign w22636 = ~w22633 & w22635;
assign w22637 = a[62] & ~w22636;
assign w22638 = ~a[62] & w22636;
assign w22639 = ~w22637 & ~w22638;
assign w22640 = w22629 & w22639;
assign w22641 = ~w22629 & ~w22639;
assign w22642 = ~w22640 & ~w22641;
assign w22643 = w22622 & ~w22642;
assign w22644 = ~w22622 & w22642;
assign w22645 = ~w22643 & ~w22644;
assign w22646 = b[47] & w10496;
assign w22647 = b[49] & w10148;
assign w22648 = b[48] & w10146;
assign w22649 = ~w7468 & w10141;
assign w22650 = ~w22647 & ~w22648;
assign w22651 = ~w22646 & w22650;
assign w22652 = ~w22649 & w22651;
assign w22653 = a[59] & ~w22652;
assign w22654 = ~a[59] & w22652;
assign w22655 = ~w22653 & ~w22654;
assign w22656 = w22645 & w22655;
assign w22657 = ~w22645 & ~w22655;
assign w22658 = ~w22656 & ~w22657;
assign w22659 = ~w22517 & ~w22521;
assign w22660 = w22658 & ~w22659;
assign w22661 = ~w22658 & w22659;
assign w22662 = ~w22660 & ~w22661;
assign w22663 = w22621 & w22662;
assign w22664 = ~w22621 & ~w22662;
assign w22665 = ~w22663 & ~w22664;
assign w22666 = ~w22525 & ~w22527;
assign w22667 = w22665 & ~w22666;
assign w22668 = ~w22665 & w22666;
assign w22669 = ~w22667 & ~w22668;
assign w22670 = w22611 & w22669;
assign w22671 = ~w22611 & ~w22669;
assign w22672 = ~w22670 & ~w22671;
assign w22673 = ~w22601 & w22672;
assign w22674 = w22601 & ~w22672;
assign w22675 = ~w22673 & ~w22674;
assign w22676 = w22600 & w22675;
assign w22677 = ~w22600 & ~w22675;
assign w22678 = ~w22676 & ~w22677;
assign w22679 = w22590 & ~w22678;
assign w22680 = ~w22590 & w22678;
assign w22681 = ~w22679 & ~w22680;
assign w22682 = w22589 & w22681;
assign w22683 = ~w22589 & ~w22681;
assign w22684 = ~w22682 & ~w22683;
assign w22685 = (~w22550 & ~w22552) | (~w22550 & w25621) | (~w22552 & w25621);
assign w22686 = b[62] & w5939;
assign w22687 = b[63] & w5670;
assign w22688 = ~w12153 & w25522;
assign w22689 = ~w22686 & ~w22687;
assign w22690 = ~w22688 & w25622;
assign w22691 = (a[44] & w22688) | (a[44] & w25623) | (w22688 & w25623);
assign w22692 = ~w22690 & ~w22691;
assign w22693 = ~w22685 & w22692;
assign w22694 = w22685 & ~w22692;
assign w22695 = ~w22693 & ~w22694;
assign w22696 = w22684 & w22695;
assign w22697 = ~w22684 & ~w22695;
assign w22698 = ~w22696 & ~w22697;
assign w22699 = (~w22566 & ~w22568) | (~w22566 & w25624) | (~w22568 & w25624);
assign w22700 = ~w22698 & w22699;
assign w22701 = w22698 & ~w22699;
assign w22702 = ~w22700 & ~w22701;
assign w22703 = (~w22175 & w24515) | (~w22175 & w24516) | (w24515 & w24516);
assign w22704 = (~w20820 & w25697) | (~w20820 & w25698) | (w25697 & w25698);
assign w22705 = ~w22703 & ~w22704;
assign w22706 = ~w22693 & ~w22696;
assign w22707 = ~w22680 & ~w22682;
assign w22708 = w5663 & ~w12154;
assign w22709 = ~w5939 & ~w22708;
assign w22710 = b[63] & ~w22709;
assign w22711 = ~a[44] & ~w22710;
assign w22712 = a[44] & w22710;
assign w22713 = ~w22711 & ~w22712;
assign w22714 = ~w22707 & w22713;
assign w22715 = w22707 & ~w22713;
assign w22716 = ~w22714 & ~w22715;
assign w22717 = b[60] & w6732;
assign w22718 = b[62] & w6476;
assign w22719 = b[61] & w6474;
assign w22720 = w6469 & w11763;
assign w22721 = ~w22718 & ~w22719;
assign w22722 = ~w22717 & w22721;
assign w22723 = ~w22720 & w22722;
assign w22724 = a[47] & ~w22723;
assign w22725 = ~a[47] & w22723;
assign w22726 = ~w22724 & ~w22725;
assign w22727 = ~w22667 & ~w22670;
assign w22728 = b[54] & w8515;
assign w22729 = b[56] & w8202;
assign w22730 = b[55] & w8200;
assign w22731 = w8195 & w9657;
assign w22732 = ~w22729 & ~w22730;
assign w22733 = ~w22728 & w22732;
assign w22734 = ~w22731 & w22733;
assign w22735 = a[53] & ~w22734;
assign w22736 = ~a[53] & w22734;
assign w22737 = ~w22735 & ~w22736;
assign w22738 = ~w22660 & ~w22663;
assign w22739 = b[51] & w9482;
assign w22740 = b[53] & w9160;
assign w22741 = b[52] & w9165;
assign w22742 = w8683 & w9158;
assign w22743 = ~w22740 & ~w22741;
assign w22744 = ~w22739 & w22743;
assign w22745 = ~w22742 & w22744;
assign w22746 = a[56] & ~w22745;
assign w22747 = ~a[56] & w22745;
assign w22748 = ~w22746 & ~w22747;
assign w22749 = ~w22644 & ~w22656;
assign w22750 = ~w22627 & ~w22640;
assign w22751 = b[43] & w11921;
assign w22752 = b[44] & w11923;
assign w22753 = ~w22751 & ~w22752;
assign w22754 = w22625 & ~w22753;
assign w22755 = ~w22625 & w22753;
assign w22756 = ~w22754 & ~w22755;
assign w22757 = b[45] & w11561;
assign w22758 = b[47] & w11196;
assign w22759 = b[46] & w11194;
assign w22760 = w6889 & w11189;
assign w22761 = ~w22758 & ~w22759;
assign w22762 = ~w22757 & w22761;
assign w22763 = ~w22760 & w22762;
assign w22764 = a[62] & ~w22763;
assign w22765 = ~a[62] & w22763;
assign w22766 = ~w22764 & ~w22765;
assign w22767 = w22756 & w22766;
assign w22768 = ~w22756 & ~w22766;
assign w22769 = ~w22767 & ~w22768;
assign w22770 = w22750 & ~w22769;
assign w22771 = ~w22750 & w22769;
assign w22772 = ~w22770 & ~w22771;
assign w22773 = b[48] & w10496;
assign w22774 = b[49] & w10146;
assign w22775 = b[50] & w10148;
assign w22776 = w7759 & w10141;
assign w22777 = ~w22774 & ~w22775;
assign w22778 = ~w22773 & w22777;
assign w22779 = ~w22776 & w22778;
assign w22780 = a[59] & ~w22779;
assign w22781 = ~a[59] & w22779;
assign w22782 = ~w22780 & ~w22781;
assign w22783 = w22772 & w22782;
assign w22784 = ~w22772 & ~w22782;
assign w22785 = ~w22783 & ~w22784;
assign w22786 = w22749 & ~w22785;
assign w22787 = ~w22749 & w22785;
assign w22788 = ~w22786 & ~w22787;
assign w22789 = w22748 & w22788;
assign w22790 = ~w22748 & ~w22788;
assign w22791 = ~w22789 & ~w22790;
assign w22792 = w22738 & ~w22791;
assign w22793 = ~w22738 & w22791;
assign w22794 = ~w22792 & ~w22793;
assign w22795 = w22737 & w22794;
assign w22796 = ~w22737 & ~w22794;
assign w22797 = ~w22795 & ~w22796;
assign w22798 = w22727 & ~w22797;
assign w22799 = ~w22727 & w22797;
assign w22800 = ~w22798 & ~w22799;
assign w22801 = b[57] & w7586;
assign w22802 = b[59] & w7314;
assign w22803 = b[58] & w7307;
assign w22804 = w7312 & w10371;
assign w22805 = ~w22802 & ~w22803;
assign w22806 = ~w22801 & w22805;
assign w22807 = ~w22804 & w22806;
assign w22808 = a[50] & ~w22807;
assign w22809 = ~a[50] & w22807;
assign w22810 = ~w22808 & ~w22809;
assign w22811 = w22800 & w22810;
assign w22812 = ~w22800 & ~w22810;
assign w22813 = ~w22811 & ~w22812;
assign w22814 = ~w22673 & ~w22676;
assign w22815 = w22813 & ~w22814;
assign w22816 = ~w22813 & w22814;
assign w22817 = ~w22815 & ~w22816;
assign w22818 = w22726 & w22817;
assign w22819 = ~w22726 & ~w22817;
assign w22820 = ~w22818 & ~w22819;
assign w22821 = w22716 & w22820;
assign w22822 = ~w22716 & ~w22820;
assign w22823 = ~w22821 & ~w22822;
assign w22824 = ~w22706 & w22823;
assign w22825 = w22706 & ~w22823;
assign w22826 = ~w22824 & ~w22825;
assign w22827 = (~w22175 & w24519) | (~w22175 & w24520) | (w24519 & w24520);
assign w22828 = (~w20820 & w25699) | (~w20820 & w25700) | (w25699 & w25700);
assign w22829 = ~w22827 & ~w22828;
assign w22830 = ~w22799 & ~w22811;
assign w22831 = b[58] & w7586;
assign w22832 = b[60] & w7314;
assign w22833 = b[59] & w7307;
assign w22834 = w7312 & w11035;
assign w22835 = ~w22832 & ~w22833;
assign w22836 = ~w22831 & w22835;
assign w22837 = ~w22834 & w22836;
assign w22838 = a[50] & ~w22837;
assign w22839 = ~a[50] & w22837;
assign w22840 = ~w22838 & ~w22839;
assign w22841 = ~w22793 & ~w22795;
assign w22842 = b[55] & w8515;
assign w22843 = b[56] & w8200;
assign w22844 = b[57] & w8202;
assign w22845 = w8195 & ~w9992;
assign w22846 = ~w22843 & ~w22844;
assign w22847 = ~w22842 & w22846;
assign w22848 = ~w22845 & w22847;
assign w22849 = a[53] & ~w22848;
assign w22850 = ~a[53] & w22848;
assign w22851 = ~w22849 & ~w22850;
assign w22852 = ~w22787 & ~w22789;
assign w22853 = b[52] & w9482;
assign w22854 = b[54] & w9160;
assign w22855 = b[53] & w9165;
assign w22856 = ~w8998 & w9158;
assign w22857 = ~w22854 & ~w22855;
assign w22858 = ~w22853 & w22857;
assign w22859 = ~w22856 & w22858;
assign w22860 = a[56] & ~w22859;
assign w22861 = ~a[56] & w22859;
assign w22862 = ~w22860 & ~w22861;
assign w22863 = ~w22771 & ~w22783;
assign w22864 = b[49] & w10496;
assign w22865 = b[50] & w10146;
assign w22866 = b[51] & w10148;
assign w22867 = ~w8058 & w10141;
assign w22868 = ~w22865 & ~w22866;
assign w22869 = ~w22864 & w22868;
assign w22870 = ~w22867 & w22869;
assign w22871 = a[59] & ~w22870;
assign w22872 = ~a[59] & w22870;
assign w22873 = ~w22871 & ~w22872;
assign w22874 = b[46] & w11561;
assign w22875 = b[47] & w11194;
assign w22876 = b[48] & w11196;
assign w22877 = ~w7170 & w11189;
assign w22878 = ~w22875 & ~w22876;
assign w22879 = ~w22874 & w22878;
assign w22880 = ~w22877 & w22879;
assign w22881 = a[62] & ~w22880;
assign w22882 = ~a[62] & w22880;
assign w22883 = ~w22881 & ~w22882;
assign w22884 = ~w22754 & ~w22767;
assign w22885 = b[44] & w11921;
assign w22886 = b[45] & w11923;
assign w22887 = ~w22885 & ~w22886;
assign w22888 = ~a[44] & ~w22887;
assign w22889 = a[44] & w22887;
assign w22890 = ~w22888 & ~w22889;
assign w22891 = w22625 & ~w22890;
assign w22892 = ~w22625 & w22890;
assign w22893 = ~w22891 & ~w22892;
assign w22894 = ~w22884 & w22893;
assign w22895 = w22884 & ~w22893;
assign w22896 = ~w22894 & ~w22895;
assign w22897 = w22883 & w22896;
assign w22898 = ~w22883 & ~w22896;
assign w22899 = ~w22897 & ~w22898;
assign w22900 = w22873 & w22899;
assign w22901 = ~w22873 & ~w22899;
assign w22902 = ~w22900 & ~w22901;
assign w22903 = ~w22863 & w22902;
assign w22904 = w22863 & ~w22902;
assign w22905 = ~w22903 & ~w22904;
assign w22906 = ~w22862 & ~w22905;
assign w22907 = w22862 & w22905;
assign w22908 = ~w22906 & ~w22907;
assign w22909 = ~w22852 & w22908;
assign w22910 = w22852 & ~w22908;
assign w22911 = ~w22909 & ~w22910;
assign w22912 = ~w22851 & ~w22911;
assign w22913 = w22851 & w22911;
assign w22914 = ~w22912 & ~w22913;
assign w22915 = ~w22841 & w22914;
assign w22916 = w22841 & ~w22914;
assign w22917 = ~w22915 & ~w22916;
assign w22918 = ~w22840 & ~w22917;
assign w22919 = w22840 & w22917;
assign w22920 = ~w22918 & ~w22919;
assign w22921 = ~w22830 & w22920;
assign w22922 = w22830 & ~w22920;
assign w22923 = ~w22921 & ~w22922;
assign w22924 = b[61] & w6732;
assign w22925 = b[62] & w6474;
assign w22926 = b[63] & w6476;
assign w22927 = w6469 & w12132;
assign w22928 = ~w22925 & ~w22926;
assign w22929 = ~w22924 & w22928;
assign w22930 = ~w22927 & w22929;
assign w22931 = a[47] & ~w22930;
assign w22932 = ~a[47] & w22930;
assign w22933 = ~w22931 & ~w22932;
assign w22934 = w22923 & w22933;
assign w22935 = ~w22923 & ~w22933;
assign w22936 = ~w22934 & ~w22935;
assign w22937 = ~w22815 & ~w22818;
assign w22938 = ~w22936 & w22937;
assign w22939 = w22936 & ~w22937;
assign w22940 = ~w22938 & ~w22939;
assign w22941 = ~w22714 & ~w22821;
assign w22942 = w22940 & ~w22941;
assign w22943 = ~w22940 & w22941;
assign w22944 = ~w22942 & ~w22943;
assign w22945 = (w20820 & w25701) | (w20820 & w25702) | (w25701 & w25702);
assign w22946 = (w22175 & w24523) | (w22175 & w24524) | (w24523 & w24524);
assign w22947 = ~w22945 & ~w22946;
assign w22948 = b[59] & w7586;
assign w22949 = b[60] & w7307;
assign w22950 = b[61] & w7314;
assign w22951 = w7312 & w11400;
assign w22952 = ~w22949 & ~w22950;
assign w22953 = ~w22948 & w22952;
assign w22954 = ~w22951 & w22953;
assign w22955 = a[50] & ~w22954;
assign w22956 = ~a[50] & w22954;
assign w22957 = ~w22955 & ~w22956;
assign w22958 = ~w22913 & ~w22915;
assign w22959 = b[56] & w8515;
assign w22960 = b[58] & w8202;
assign w22961 = b[57] & w8200;
assign w22962 = w8195 & ~w10339;
assign w22963 = ~w22960 & ~w22961;
assign w22964 = ~w22959 & w22963;
assign w22965 = ~w22962 & w22964;
assign w22966 = a[53] & ~w22965;
assign w22967 = ~a[53] & w22965;
assign w22968 = ~w22966 & ~w22967;
assign w22969 = ~w22907 & ~w22909;
assign w22970 = ~w22900 & ~w22903;
assign w22971 = b[50] & w10496;
assign w22972 = b[52] & w10148;
assign w22973 = b[51] & w10146;
assign w22974 = ~w8371 & w10141;
assign w22975 = ~w22972 & ~w22973;
assign w22976 = ~w22971 & w22975;
assign w22977 = ~w22974 & w22976;
assign w22978 = a[59] & ~w22977;
assign w22979 = ~a[59] & w22977;
assign w22980 = ~w22978 & ~w22979;
assign w22981 = ~w22894 & ~w22897;
assign w22982 = b[45] & w11921;
assign w22983 = b[46] & w11923;
assign w22984 = ~w22982 & ~w22983;
assign w22985 = ~w22888 & ~w22892;
assign w22986 = w22984 & ~w22985;
assign w22987 = ~w22984 & w22985;
assign w22988 = ~w22986 & ~w22987;
assign w22989 = b[47] & w11561;
assign w22990 = b[48] & w11194;
assign w22991 = b[49] & w11196;
assign w22992 = ~w22990 & ~w22991;
assign w22993 = ~w22989 & w22992;
assign w22994 = (w22993 & w7468) | (w22993 & w25364) | (w7468 & w25364);
assign w22995 = a[62] & ~w22994;
assign w22996 = ~a[62] & w22994;
assign w22997 = ~w22995 & ~w22996;
assign w22998 = ~w22988 & ~w22997;
assign w22999 = w22988 & w22997;
assign w23000 = ~w22998 & ~w22999;
assign w23001 = w22981 & ~w23000;
assign w23002 = ~w22981 & w23000;
assign w23003 = ~w23001 & ~w23002;
assign w23004 = w22980 & w23003;
assign w23005 = ~w22980 & ~w23003;
assign w23006 = ~w23004 & ~w23005;
assign w23007 = w22970 & ~w23006;
assign w23008 = ~w22970 & w23006;
assign w23009 = ~w23007 & ~w23008;
assign w23010 = b[53] & w9482;
assign w23011 = b[55] & w9160;
assign w23012 = b[54] & w9165;
assign w23013 = w9158 & ~w9330;
assign w23014 = ~w23011 & ~w23012;
assign w23015 = ~w23010 & w23014;
assign w23016 = ~w23013 & w23015;
assign w23017 = a[56] & ~w23016;
assign w23018 = ~a[56] & w23016;
assign w23019 = ~w23017 & ~w23018;
assign w23020 = w23009 & w23019;
assign w23021 = ~w23009 & ~w23019;
assign w23022 = ~w23020 & ~w23021;
assign w23023 = ~w22969 & w23022;
assign w23024 = w22969 & ~w23022;
assign w23025 = ~w23023 & ~w23024;
assign w23026 = w22968 & w23025;
assign w23027 = ~w22968 & ~w23025;
assign w23028 = ~w23026 & ~w23027;
assign w23029 = w22958 & ~w23028;
assign w23030 = ~w22958 & w23028;
assign w23031 = ~w23029 & ~w23030;
assign w23032 = w22957 & w23031;
assign w23033 = ~w22957 & ~w23031;
assign w23034 = ~w23032 & ~w23033;
assign w23035 = ~w22919 & ~w22921;
assign w23036 = b[62] & w6732;
assign w23037 = b[63] & w6474;
assign w23038 = w6469 & w12156;
assign w23039 = ~w23036 & ~w23037;
assign w23040 = ~w23038 & w23039;
assign w23041 = a[47] & w23040;
assign w23042 = ~a[47] & ~w23040;
assign w23043 = ~w23041 & ~w23042;
assign w23044 = ~w23035 & ~w23043;
assign w23045 = w23035 & w23043;
assign w23046 = ~w23044 & ~w23045;
assign w23047 = w23034 & w23046;
assign w23048 = ~w23034 & ~w23046;
assign w23049 = ~w23047 & ~w23048;
assign w23050 = ~w22934 & ~w22939;
assign w23051 = ~w23049 & w23050;
assign w23052 = w23049 & ~w23050;
assign w23053 = ~w23051 & ~w23052;
assign w23054 = (~w20820 & w25703) | (~w20820 & w25704) | (w25703 & w25704);
assign w23055 = (~w22175 & w24527) | (~w22175 & w24528) | (w24527 & w24528);
assign w23056 = ~w23054 & ~w23055;
assign w23057 = b[60] & w7586;
assign w23058 = b[61] & w7307;
assign w23059 = b[62] & w7314;
assign w23060 = ~w23058 & ~w23059;
assign w23061 = ~w23057 & w23060;
assign w23062 = (w23061 & ~w11763) | (w23061 & w25042) | (~w11763 & w25042);
assign w23063 = a[50] & ~w23062;
assign w23064 = ~a[50] & w23062;
assign w23065 = ~w23063 & ~w23064;
assign w23066 = ~w23008 & ~w23020;
assign w23067 = b[54] & w9482;
assign w23068 = b[55] & w9165;
assign w23069 = b[56] & w9160;
assign w23070 = ~w23068 & ~w23069;
assign w23071 = ~w23067 & w23070;
assign w23072 = (w23071 & ~w9657) | (w23071 & w25367) | (~w9657 & w25367);
assign w23073 = a[56] & ~w23072;
assign w23074 = ~a[56] & w23072;
assign w23075 = ~w23073 & ~w23074;
assign w23076 = ~w23002 & ~w23004;
assign w23077 = b[51] & w10496;
assign w23078 = b[52] & w10146;
assign w23079 = b[53] & w10148;
assign w23080 = w8683 & w10141;
assign w23081 = ~w23078 & ~w23079;
assign w23082 = ~w23077 & w23081;
assign w23083 = ~w23080 & w23082;
assign w23084 = a[59] & ~w23083;
assign w23085 = ~a[59] & w23083;
assign w23086 = ~w23084 & ~w23085;
assign w23087 = b[48] & w11561;
assign w23088 = b[50] & w11196;
assign w23089 = b[49] & w11194;
assign w23090 = w7759 & w11189;
assign w23091 = ~w23088 & ~w23089;
assign w23092 = ~w23087 & w23091;
assign w23093 = ~w23090 & w23092;
assign w23094 = a[62] & ~w23093;
assign w23095 = ~a[62] & w23093;
assign w23096 = ~w23094 & ~w23095;
assign w23097 = ~w22986 & ~w22999;
assign w23098 = b[46] & w11921;
assign w23099 = b[47] & w11923;
assign w23100 = ~w23098 & ~w23099;
assign w23101 = w22984 & ~w23100;
assign w23102 = ~w22984 & w23100;
assign w23103 = ~w23101 & ~w23102;
assign w23104 = w23097 & w23103;
assign w23105 = ~w23097 & ~w23103;
assign w23106 = ~w23104 & ~w23105;
assign w23107 = w23096 & ~w23106;
assign w23108 = ~w23096 & w23106;
assign w23109 = ~w23107 & ~w23108;
assign w23110 = w23086 & w23109;
assign w23111 = ~w23086 & ~w23109;
assign w23112 = ~w23110 & ~w23111;
assign w23113 = w23076 & ~w23112;
assign w23114 = ~w23076 & w23112;
assign w23115 = ~w23113 & ~w23114;
assign w23116 = w23075 & w23115;
assign w23117 = ~w23075 & ~w23115;
assign w23118 = ~w23116 & ~w23117;
assign w23119 = w23066 & ~w23118;
assign w23120 = ~w23066 & w23118;
assign w23121 = ~w23119 & ~w23120;
assign w23122 = b[57] & w8515;
assign w23123 = b[59] & w8202;
assign w23124 = b[58] & w8200;
assign w23125 = ~w23123 & ~w23124;
assign w23126 = ~w23122 & w23125;
assign w23127 = (w10371 & w25368) | (w10371 & w25369) | (w25368 & w25369);
assign w23128 = ~a[53] & w25752;
assign w23129 = ~w23127 & ~w23128;
assign w23130 = w23121 & w23129;
assign w23131 = ~w23121 & ~w23129;
assign w23132 = ~w23130 & ~w23131;
assign w23133 = ~w23023 & ~w23026;
assign w23134 = w23132 & ~w23133;
assign w23135 = ~w23132 & w23133;
assign w23136 = ~w23134 & ~w23135;
assign w23137 = w23065 & w23136;
assign w23138 = ~w23065 & ~w23136;
assign w23139 = ~w23137 & ~w23138;
assign w23140 = ~w23030 & ~w23032;
assign w23141 = w6469 & ~w12154;
assign w23142 = ~w6732 & ~w23141;
assign w23143 = b[63] & ~w23142;
assign w23144 = a[47] & ~w23143;
assign w23145 = ~a[47] & w23143;
assign w23146 = ~w23144 & ~w23145;
assign w23147 = ~w23140 & ~w23146;
assign w23148 = w23140 & w23146;
assign w23149 = ~w23147 & ~w23148;
assign w23150 = ~w23139 & ~w23149;
assign w23151 = w23139 & w23149;
assign w23152 = ~w23150 & ~w23151;
assign w23153 = ~w23044 & ~w23047;
assign w23154 = ~w23152 & w23153;
assign w23155 = w23152 & ~w23153;
assign w23156 = ~w23154 & ~w23155;
assign w23157 = (~w22175 & w24531) | (~w22175 & w24532) | (w24531 & w24532);
assign w23158 = (~w20820 & w25705) | (~w20820 & w25706) | (w25705 & w25706);
assign w23159 = ~w23157 & ~w23158;
assign w23160 = ~w23120 & ~w23130;
assign w23161 = b[58] & w8515;
assign w23162 = b[60] & w8202;
assign w23163 = b[59] & w8200;
assign w23164 = ~w23162 & ~w23163;
assign w23165 = ~w23161 & w23164;
assign w23166 = (w11035 & w24886) | (w11035 & w24887) | (w24886 & w24887);
assign w23167 = (~w11035 & w24888) | (~w11035 & w24889) | (w24888 & w24889);
assign w23168 = ~w23166 & ~w23167;
assign w23169 = ~w23114 & ~w23116;
assign w23170 = b[55] & w9482;
assign w23171 = b[57] & w9160;
assign w23172 = b[56] & w9165;
assign w23173 = ~w23171 & ~w23172;
assign w23174 = ~w23170 & w23173;
assign w23175 = a[56] & w25753;
assign w23176 = (w9992 & w25225) | (w9992 & w25226) | (w25225 & w25226);
assign w23177 = ~w23175 & ~w23176;
assign w23178 = ~w23107 & ~w23110;
assign w23179 = b[52] & w10496;
assign w23180 = b[53] & w10146;
assign w23181 = b[54] & w10148;
assign w23182 = ~w23180 & ~w23181;
assign w23183 = ~w23179 & w23182;
assign w23184 = a[59] & w25754;
assign w23185 = (w8998 & w25372) | (w8998 & w25373) | (w25372 & w25373);
assign w23186 = ~w23184 & ~w23185;
assign w23187 = b[49] & w11561;
assign w23188 = b[50] & w11194;
assign w23189 = b[51] & w11196;
assign w23190 = ~w23188 & ~w23189;
assign w23191 = ~w23187 & w23190;
assign w23192 = (w23191 & w8058) | (w23191 & w25374) | (w8058 & w25374);
assign w23193 = a[62] & ~w23192;
assign w23194 = ~a[62] & w23192;
assign w23195 = ~w23193 & ~w23194;
assign w23196 = b[47] & w11921;
assign w23197 = b[48] & w11923;
assign w23198 = ~w23196 & ~w23197;
assign w23199 = ~a[47] & ~w23100;
assign w23200 = a[47] & w23100;
assign w23201 = ~w23199 & ~w23200;
assign w23202 = ~w23198 & w23201;
assign w23203 = w23198 & ~w23201;
assign w23204 = ~w23202 & ~w23203;
assign w23205 = ~w23195 & ~w23204;
assign w23206 = w23195 & w23204;
assign w23207 = ~w23205 & ~w23206;
assign w23208 = ~w23101 & ~w23104;
assign w23209 = w23207 & w23208;
assign w23210 = ~w23207 & ~w23208;
assign w23211 = ~w23209 & ~w23210;
assign w23212 = w23186 & w23211;
assign w23213 = ~w23186 & ~w23211;
assign w23214 = ~w23212 & ~w23213;
assign w23215 = ~w23178 & w23214;
assign w23216 = w23178 & ~w23214;
assign w23217 = ~w23215 & ~w23216;
assign w23218 = ~w23177 & ~w23217;
assign w23219 = w23177 & w23217;
assign w23220 = ~w23218 & ~w23219;
assign w23221 = ~w23169 & w23220;
assign w23222 = w23169 & ~w23220;
assign w23223 = ~w23221 & ~w23222;
assign w23224 = ~w23168 & ~w23223;
assign w23225 = w23168 & w23223;
assign w23226 = ~w23224 & ~w23225;
assign w23227 = ~w23160 & w23226;
assign w23228 = w23160 & ~w23226;
assign w23229 = ~w23227 & ~w23228;
assign w23230 = b[61] & w7586;
assign w23231 = b[62] & w7307;
assign w23232 = b[63] & w7314;
assign w23233 = ~w23231 & ~w23232;
assign w23234 = ~w23230 & w23233;
assign w23235 = (w12132 & w25045) | (w12132 & w25046) | (w25045 & w25046);
assign w23236 = ~a[50] & w25755;
assign w23237 = ~w23235 & ~w23236;
assign w23238 = w23229 & w23237;
assign w23239 = ~w23229 & ~w23237;
assign w23240 = ~w23238 & ~w23239;
assign w23241 = ~w23134 & ~w23137;
assign w23242 = ~w23240 & w23241;
assign w23243 = w23240 & ~w23241;
assign w23244 = ~w23242 & ~w23243;
assign w23245 = ~w23147 & ~w23151;
assign w23246 = ~w23244 & w23245;
assign w23247 = w23244 & ~w23245;
assign w23248 = ~w23246 & ~w23247;
assign w23249 = (~w20820 & w25707) | (~w20820 & w25708) | (w25707 & w25708);
assign w23250 = (~w22175 & w24535) | (~w22175 & w24536) | (w24535 & w24536);
assign w23251 = ~w23249 & ~w23250;
assign w23252 = (~w23225 & ~w23226) | (~w23225 & w25047) | (~w23226 & w25047);
assign w23253 = b[59] & w8515;
assign w23254 = b[60] & w8200;
assign w23255 = b[61] & w8202;
assign w23256 = ~w23254 & ~w23255;
assign w23257 = ~w23253 & w23256;
assign w23258 = (w11400 & w24890) | (w11400 & w24891) | (w24890 & w24891);
assign w23259 = (~w11400 & w24892) | (~w11400 & w24893) | (w24892 & w24893);
assign w23260 = ~w23258 & ~w23259;
assign w23261 = (~w23219 & ~w23220) | (~w23219 & w25377) | (~w23220 & w25377);
assign w23262 = b[56] & w9482;
assign w23263 = b[57] & w9165;
assign w23264 = b[58] & w9160;
assign w23265 = ~w23263 & ~w23264;
assign w23266 = ~w23262 & w23265;
assign w23267 = (~w10339 & w25228) | (~w10339 & w25229) | (w25228 & w25229);
assign w23268 = (w10339 & w25230) | (w10339 & w25231) | (w25230 & w25231);
assign w23269 = ~w23267 & ~w23268;
assign w23270 = ~w23212 & ~w23215;
assign w23271 = b[53] & w10496;
assign w23272 = b[55] & w10148;
assign w23273 = b[54] & w10146;
assign w23274 = ~w23272 & ~w23273;
assign w23275 = ~w23271 & w23274;
assign w23276 = (w23275 & w9330) | (w23275 & w25378) | (w9330 & w25378);
assign w23277 = a[59] & ~w23276;
assign w23278 = ~a[59] & w23276;
assign w23279 = ~w23277 & ~w23278;
assign w23280 = ~w23206 & ~w23209;
assign w23281 = b[48] & w11921;
assign w23282 = b[49] & w11923;
assign w23283 = ~w23281 & ~w23282;
assign w23284 = ~w23199 & ~w23202;
assign w23285 = w23283 & ~w23284;
assign w23286 = ~w23283 & w23284;
assign w23287 = ~w23285 & ~w23286;
assign w23288 = b[50] & w11561;
assign w23289 = b[51] & w11194;
assign w23290 = b[52] & w11196;
assign w23291 = ~w23289 & ~w23290;
assign w23292 = ~w23288 & w23291;
assign w23293 = (w23292 & w8371) | (w23292 & w25379) | (w8371 & w25379);
assign w23294 = a[62] & ~w23293;
assign w23295 = ~a[62] & w23293;
assign w23296 = ~w23294 & ~w23295;
assign w23297 = w23287 & w23296;
assign w23298 = ~w23287 & ~w23296;
assign w23299 = ~w23297 & ~w23298;
assign w23300 = w23280 & ~w23299;
assign w23301 = ~w23280 & w23299;
assign w23302 = ~w23300 & ~w23301;
assign w23303 = w23279 & w23302;
assign w23304 = ~w23279 & ~w23302;
assign w23305 = ~w23303 & ~w23304;
assign w23306 = w23270 & ~w23305;
assign w23307 = ~w23270 & w23305;
assign w23308 = ~w23306 & ~w23307;
assign w23309 = w23269 & w23308;
assign w23310 = ~w23269 & ~w23308;
assign w23311 = ~w23309 & ~w23310;
assign w23312 = w23261 & ~w23311;
assign w23313 = ~w23261 & w23311;
assign w23314 = ~w23312 & ~w23313;
assign w23315 = w23260 & w23314;
assign w23316 = ~w23260 & ~w23314;
assign w23317 = ~w23315 & ~w23316;
assign w23318 = w23252 & ~w23317;
assign w23319 = ~w23252 & w23317;
assign w23320 = ~w23318 & ~w23319;
assign w23321 = b[62] & w7586;
assign w23322 = b[63] & w7307;
assign w23323 = ~w12153 & w24730;
assign w23324 = ~w23321 & ~w23322;
assign w23325 = (a[50] & w23323) | (a[50] & w25049) | (w23323 & w25049);
assign w23326 = ~w23323 & w25050;
assign w23327 = ~w23325 & ~w23326;
assign w23328 = w23320 & w23327;
assign w23329 = ~w23320 & ~w23327;
assign w23330 = ~w23328 & ~w23329;
assign w23331 = (~w23238 & ~w23240) | (~w23238 & w25232) | (~w23240 & w25232);
assign w23332 = ~w23330 & w23331;
assign w23333 = w23330 & ~w23331;
assign w23334 = ~w23332 & ~w23333;
assign w23335 = (~w20820 & w25644) | (~w20820 & w25645) | (w25644 & w25645);
assign w23336 = (w22175 & w25380) | (w22175 & w25381) | (w25380 & w25381);
assign w23337 = (~w22175 & w25382) | (~w22175 & w25383) | (w25382 & w25383);
assign w23338 = ~w23336 & ~w23337;
assign w23339 = b[60] & w8515;
assign w23340 = b[62] & w8202;
assign w23341 = b[61] & w8200;
assign w23342 = ~w23340 & ~w23341;
assign w23343 = ~w23339 & w23342;
assign w23344 = (w11763 & w25051) | (w11763 & w25052) | (w25051 & w25052);
assign w23345 = ~a[53] & w25756;
assign w23346 = ~w23344 & ~w23345;
assign w23347 = ~w23301 & ~w23303;
assign w23348 = b[54] & w10496;
assign w23349 = b[56] & w10148;
assign w23350 = b[55] & w10146;
assign w23351 = ~w23349 & ~w23350;
assign w23352 = ~w23348 & w23351;
assign w23353 = (w23352 & ~w9657) | (w23352 & w25384) | (~w9657 & w25384);
assign w23354 = a[59] & ~w23353;
assign w23355 = ~a[59] & w23353;
assign w23356 = ~w23354 & ~w23355;
assign w23357 = ~w23285 & ~w23297;
assign w23358 = b[51] & w11561;
assign w23359 = b[53] & w11196;
assign w23360 = b[52] & w11194;
assign w23361 = ~w23359 & ~w23360;
assign w23362 = ~w23358 & w23361;
assign w23363 = (w23362 & ~w8683) | (w23362 & w25523) | (~w8683 & w25523);
assign w23364 = a[62] & ~w23363;
assign w23365 = ~a[62] & w23363;
assign w23366 = ~w23364 & ~w23365;
assign w23367 = b[49] & w11921;
assign w23368 = b[50] & w11923;
assign w23369 = ~w23367 & ~w23368;
assign w23370 = w23283 & ~w23369;
assign w23371 = ~w23283 & w23369;
assign w23372 = ~w23370 & ~w23371;
assign w23373 = w23366 & w23372;
assign w23374 = ~w23366 & ~w23372;
assign w23375 = ~w23373 & ~w23374;
assign w23376 = ~w23357 & w23375;
assign w23377 = w23357 & ~w23375;
assign w23378 = ~w23376 & ~w23377;
assign w23379 = ~w23356 & ~w23378;
assign w23380 = w23356 & w23378;
assign w23381 = ~w23379 & ~w23380;
assign w23382 = w23347 & ~w23381;
assign w23383 = ~w23347 & w23381;
assign w23384 = ~w23382 & ~w23383;
assign w23385 = b[57] & w9482;
assign w23386 = b[58] & w9165;
assign w23387 = b[59] & w9160;
assign w23388 = ~w23386 & ~w23387;
assign w23389 = ~w23385 & w23388;
assign w23390 = (w10371 & w25233) | (w10371 & w25234) | (w25233 & w25234);
assign w23391 = (~w10371 & w25235) | (~w10371 & w25236) | (w25235 & w25236);
assign w23392 = ~w23390 & ~w23391;
assign w23393 = w23384 & w23392;
assign w23394 = ~w23384 & ~w23392;
assign w23395 = ~w23393 & ~w23394;
assign w23396 = ~w23307 & ~w23309;
assign w23397 = w23395 & ~w23396;
assign w23398 = ~w23395 & w23396;
assign w23399 = ~w23397 & ~w23398;
assign w23400 = w23346 & w23399;
assign w23401 = ~w23346 & ~w23399;
assign w23402 = ~w23400 & ~w23401;
assign w23403 = (~w23313 & ~w23260) | (~w23313 & w25054) | (~w23260 & w25054);
assign w23404 = (w11757 & w25055) | (w11757 & w25056) | (w25055 & w25056);
assign w23405 = b[63] & ~w23404;
assign w23406 = a[50] & ~w23405;
assign w23407 = ~a[50] & w23405;
assign w23408 = ~w23406 & ~w23407;
assign w23409 = ~w23403 & ~w23408;
assign w23410 = w23403 & w23408;
assign w23411 = ~w23409 & ~w23410;
assign w23412 = ~w23402 & ~w23411;
assign w23413 = w23402 & w23411;
assign w23414 = ~w23412 & ~w23413;
assign w23415 = (~w23319 & ~w23320) | (~w23319 & w25057) | (~w23320 & w25057);
assign w23416 = ~w23414 & w23415;
assign w23417 = w23414 & ~w23415;
assign w23418 = ~w23416 & ~w23417;
assign w23419 = (~w22175 & w25385) | (~w22175 & w25386) | (w25385 & w25386);
assign w23420 = (w22175 & w25646) | (w22175 & w25647) | (w25646 & w25647);
assign w23421 = ~w23419 & ~w23420;
assign w23422 = ~w23383 & ~w23393;
assign w23423 = b[58] & w9482;
assign w23424 = b[60] & w9160;
assign w23425 = b[59] & w9165;
assign w23426 = ~w23424 & ~w23425;
assign w23427 = ~w23423 & w23426;
assign w23428 = (w11035 & w25237) | (w11035 & w25238) | (w25237 & w25238);
assign w23429 = (~w11035 & w25239) | (~w11035 & w25240) | (w25239 & w25240);
assign w23430 = ~w23428 & ~w23429;
assign w23431 = ~w23376 & ~w23380;
assign w23432 = b[55] & w10496;
assign w23433 = b[57] & w10148;
assign w23434 = b[56] & w10146;
assign w23435 = ~w23433 & ~w23434;
assign w23436 = ~w23432 & w23435;
assign w23437 = (~w9992 & w25524) | (~w9992 & w25525) | (w25524 & w25525);
assign w23438 = (w9992 & w25526) | (w9992 & w25527) | (w25526 & w25527);
assign w23439 = ~w23437 & ~w23438;
assign w23440 = b[52] & w11561;
assign w23441 = b[54] & w11196;
assign w23442 = b[53] & w11194;
assign w23443 = ~w8998 & w11189;
assign w23444 = ~w23441 & ~w23442;
assign w23445 = ~w23440 & w23444;
assign w23446 = ~w23443 & w23445;
assign w23447 = a[62] & ~w23446;
assign w23448 = ~a[62] & w23446;
assign w23449 = ~w23447 & ~w23448;
assign w23450 = ~w23370 & ~w23373;
assign w23451 = b[50] & w11921;
assign w23452 = b[51] & w11923;
assign w23453 = ~w23451 & ~w23452;
assign w23454 = ~a[50] & ~w23453;
assign w23455 = a[50] & w23453;
assign w23456 = ~w23454 & ~w23455;
assign w23457 = ~w23283 & w23456;
assign w23458 = w23283 & ~w23456;
assign w23459 = ~w23457 & ~w23458;
assign w23460 = ~w23450 & w23459;
assign w23461 = w23450 & ~w23459;
assign w23462 = ~w23460 & ~w23461;
assign w23463 = w23449 & w23462;
assign w23464 = ~w23449 & ~w23462;
assign w23465 = ~w23463 & ~w23464;
assign w23466 = w23439 & w23465;
assign w23467 = ~w23439 & ~w23465;
assign w23468 = ~w23466 & ~w23467;
assign w23469 = ~w23431 & w23468;
assign w23470 = w23431 & ~w23468;
assign w23471 = ~w23469 & ~w23470;
assign w23472 = ~w23430 & ~w23471;
assign w23473 = w23430 & w23471;
assign w23474 = ~w23472 & ~w23473;
assign w23475 = ~w23422 & w23474;
assign w23476 = w23422 & ~w23474;
assign w23477 = ~w23475 & ~w23476;
assign w23478 = b[61] & w8515;
assign w23479 = b[63] & w8202;
assign w23480 = b[62] & w8200;
assign w23481 = ~w23479 & ~w23480;
assign w23482 = ~w23478 & w23481;
assign w23483 = (w23482 & ~w12132) | (w23482 & w25061) | (~w12132 & w25061);
assign w23484 = a[53] & ~w23483;
assign w23485 = ~a[53] & w23483;
assign w23486 = ~w23484 & ~w23485;
assign w23487 = w23477 & w23486;
assign w23488 = ~w23477 & ~w23486;
assign w23489 = ~w23487 & ~w23488;
assign w23490 = ~w23397 & ~w23400;
assign w23491 = ~w23489 & w23490;
assign w23492 = w23489 & ~w23490;
assign w23493 = ~w23491 & ~w23492;
assign w23494 = ~w23409 & ~w23413;
assign w23495 = ~w23493 & w23494;
assign w23496 = w23493 & ~w23494;
assign w23497 = ~w23495 & ~w23496;
assign w23498 = (~w22175 & w25648) | (~w22175 & w25649) | (w25648 & w25649);
assign w23499 = (w22175 & w25388) | (w22175 & w25389) | (w25388 & w25389);
assign w23500 = ~w23498 & ~w23499;
assign w23501 = (~w23473 & ~w23474) | (~w23473 & w25390) | (~w23474 & w25390);
assign w23502 = b[59] & w9482;
assign w23503 = b[61] & w9160;
assign w23504 = b[60] & w9165;
assign w23505 = ~w23503 & ~w23504;
assign w23506 = ~w23502 & w23505;
assign w23507 = (w11400 & w25391) | (w11400 & w25392) | (w25391 & w25392);
assign w23508 = (~w11400 & w25393) | (~w11400 & w25394) | (w25393 & w25394);
assign w23509 = ~w23507 & ~w23508;
assign w23510 = ~w23466 & ~w23469;
assign w23511 = b[56] & w10496;
assign w23512 = b[57] & w10146;
assign w23513 = b[58] & w10148;
assign w23514 = ~w23512 & ~w23513;
assign w23515 = ~w23511 & w23514;
assign w23516 = (~w10339 & w25528) | (~w10339 & w25529) | (w25528 & w25529);
assign w23517 = (w10339 & w25530) | (w10339 & w25531) | (w25530 & w25531);
assign w23518 = ~w23516 & ~w23517;
assign w23519 = ~w23460 & ~w23463;
assign w23520 = b[51] & w11921;
assign w23521 = b[52] & w11923;
assign w23522 = ~w23520 & ~w23521;
assign w23523 = ~w23454 & ~w23457;
assign w23524 = w23522 & ~w23523;
assign w23525 = ~w23522 & w23523;
assign w23526 = ~w23524 & ~w23525;
assign w23527 = b[53] & w11561;
assign w23528 = b[55] & w11196;
assign w23529 = b[54] & w11194;
assign w23530 = ~w9330 & w11189;
assign w23531 = ~w23528 & ~w23529;
assign w23532 = ~w23527 & w23531;
assign w23533 = ~w23530 & w23532;
assign w23534 = a[62] & ~w23533;
assign w23535 = ~a[62] & w23533;
assign w23536 = ~w23534 & ~w23535;
assign w23537 = ~w23526 & ~w23536;
assign w23538 = w23526 & w23536;
assign w23539 = ~w23537 & ~w23538;
assign w23540 = w23519 & ~w23539;
assign w23541 = ~w23519 & w23539;
assign w23542 = ~w23540 & ~w23541;
assign w23543 = w23518 & w23542;
assign w23544 = ~w23518 & ~w23542;
assign w23545 = ~w23543 & ~w23544;
assign w23546 = w23510 & ~w23545;
assign w23547 = ~w23510 & w23545;
assign w23548 = ~w23546 & ~w23547;
assign w23549 = w23509 & w23548;
assign w23550 = ~w23509 & ~w23548;
assign w23551 = ~w23549 & ~w23550;
assign w23552 = w23501 & ~w23551;
assign w23553 = ~w23501 & w23551;
assign w23554 = ~w23552 & ~w23553;
assign w23555 = b[62] & w8515;
assign w23556 = b[63] & w8200;
assign w23557 = ~w12153 & w25532;
assign w23558 = ~w23555 & ~w23556;
assign w23559 = ~w23557 & w23558;
assign w23560 = ~a[53] & w23559;
assign w23561 = a[53] & ~w23559;
assign w23562 = ~w23560 & ~w23561;
assign w23563 = w23554 & w23562;
assign w23564 = ~w23554 & ~w23562;
assign w23565 = ~w23563 & ~w23564;
assign w23566 = (~w23487 & ~w23489) | (~w23487 & w25396) | (~w23489 & w25396);
assign w23567 = ~w23565 & w23566;
assign w23568 = w23565 & ~w23566;
assign w23569 = ~w23567 & ~w23568;
assign w23570 = (~w22175 & w25397) | (~w22175 & w25398) | (w25397 & w25398);
assign w23571 = (w22175 & w25650) | (w22175 & w25651) | (w25650 & w25651);
assign w23572 = ~w23570 & ~w23571;
assign w23573 = ~w23541 & ~w23543;
assign w23574 = b[57] & w10496;
assign w23575 = b[58] & w10146;
assign w23576 = b[59] & w10148;
assign w23577 = ~w23575 & ~w23576;
assign w23578 = ~w23574 & w23577;
assign w23579 = (w10371 & w25625) | (w10371 & w25626) | (w25625 & w25626);
assign w23580 = (~w10371 & w25627) | (~w10371 & w25628) | (w25627 & w25628);
assign w23581 = ~w23579 & ~w23580;
assign w23582 = b[54] & w11561;
assign w23583 = b[56] & w11196;
assign w23584 = b[55] & w11194;
assign w23585 = w9657 & w11189;
assign w23586 = ~w23583 & ~w23584;
assign w23587 = ~w23582 & w23586;
assign w23588 = ~w23585 & w23587;
assign w23589 = a[62] & ~w23588;
assign w23590 = ~a[62] & w23588;
assign w23591 = ~w23589 & ~w23590;
assign w23592 = ~w23524 & ~w23538;
assign w23593 = b[52] & w11921;
assign w23594 = b[53] & w11923;
assign w23595 = ~w23593 & ~w23594;
assign w23596 = w23522 & ~w23595;
assign w23597 = ~w23522 & w23595;
assign w23598 = ~w23596 & ~w23597;
assign w23599 = w23592 & w23598;
assign w23600 = ~w23592 & ~w23598;
assign w23601 = ~w23599 & ~w23600;
assign w23602 = w23591 & ~w23601;
assign w23603 = ~w23591 & w23601;
assign w23604 = ~w23602 & ~w23603;
assign w23605 = w23581 & w23604;
assign w23606 = ~w23581 & ~w23604;
assign w23607 = ~w23605 & ~w23606;
assign w23608 = w23573 & ~w23607;
assign w23609 = ~w23573 & w23607;
assign w23610 = ~w23608 & ~w23609;
assign w23611 = b[60] & w9482;
assign w23612 = b[62] & w9160;
assign w23613 = b[61] & w9165;
assign w23614 = ~w23612 & ~w23613;
assign w23615 = ~w23611 & w23614;
assign w23616 = (w23615 & ~w11763) | (w23615 & w25629) | (~w11763 & w25629);
assign w23617 = a[56] & ~w23616;
assign w23618 = ~a[56] & w23616;
assign w23619 = ~w23617 & ~w23618;
assign w23620 = w23610 & w23619;
assign w23621 = ~w23610 & ~w23619;
assign w23622 = ~w23620 & ~w23621;
assign w23623 = (~w23547 & ~w23509) | (~w23547 & w25630) | (~w23509 & w25630);
assign w23624 = (~w11757 & w25631) | (~w11757 & w25632) | (w25631 & w25632);
assign w23625 = ~w8515 & ~w23624;
assign w23626 = b[63] & ~w23625;
assign w23627 = a[53] & ~w23626;
assign w23628 = ~a[53] & w23626;
assign w23629 = ~w23627 & ~w23628;
assign w23630 = ~w23623 & ~w23629;
assign w23631 = w23623 & w23629;
assign w23632 = ~w23630 & ~w23631;
assign w23633 = ~w23622 & ~w23632;
assign w23634 = w23622 & w23632;
assign w23635 = ~w23633 & ~w23634;
assign w23636 = (~w23553 & ~w23554) | (~w23553 & w25633) | (~w23554 & w25633);
assign w23637 = ~w23635 & w23636;
assign w23638 = w23635 & ~w23636;
assign w23639 = ~w23637 & ~w23638;
assign w23640 = (~w22175 & w25399) | (~w22175 & w25400) | (w25399 & w25400);
assign w23641 = (w22175 & w25652) | (w22175 & w25653) | (w25652 & w25653);
assign w23642 = ~w23640 & ~w23641;
assign w23643 = ~w23630 & ~w23634;
assign w23644 = ~w23609 & ~w23620;
assign w23645 = b[61] & w9482;
assign w23646 = b[62] & w9165;
assign w23647 = b[63] & w9160;
assign w23648 = w9158 & w12132;
assign w23649 = ~w23646 & ~w23647;
assign w23650 = ~w23645 & w23649;
assign w23651 = ~w23648 & w23650;
assign w23652 = a[56] & ~w23651;
assign w23653 = ~a[56] & w23651;
assign w23654 = ~w23652 & ~w23653;
assign w23655 = ~w23644 & w23654;
assign w23656 = w23644 & ~w23654;
assign w23657 = ~w23655 & ~w23656;
assign w23658 = ~w23602 & ~w23605;
assign w23659 = b[58] & w10496;
assign w23660 = b[59] & w10146;
assign w23661 = b[60] & w10148;
assign w23662 = w10141 & w11035;
assign w23663 = ~w23660 & ~w23661;
assign w23664 = ~w23659 & w23663;
assign w23665 = ~w23662 & w23664;
assign w23666 = a[59] & ~w23665;
assign w23667 = ~a[59] & w23665;
assign w23668 = ~w23666 & ~w23667;
assign w23669 = b[53] & w11921;
assign w23670 = b[54] & w11923;
assign w23671 = ~w23669 & ~w23670;
assign w23672 = ~a[53] & ~w23595;
assign w23673 = a[53] & w23595;
assign w23674 = ~w23672 & ~w23673;
assign w23675 = w23671 & ~w23674;
assign w23676 = ~w23671 & w23674;
assign w23677 = ~w23675 & ~w23676;
assign w23678 = b[55] & w11561;
assign w23679 = b[56] & w11194;
assign w23680 = b[57] & w11196;
assign w23681 = ~w9992 & w11189;
assign w23682 = ~w23679 & ~w23680;
assign w23683 = ~w23678 & w23682;
assign w23684 = ~w23681 & w23683;
assign w23685 = a[62] & ~w23684;
assign w23686 = ~a[62] & w23684;
assign w23687 = ~w23685 & ~w23686;
assign w23688 = w23677 & w23687;
assign w23689 = ~w23677 & ~w23687;
assign w23690 = ~w23688 & ~w23689;
assign w23691 = ~w23596 & ~w23599;
assign w23692 = w23690 & w23691;
assign w23693 = ~w23690 & ~w23691;
assign w23694 = ~w23692 & ~w23693;
assign w23695 = ~w23668 & ~w23694;
assign w23696 = w23668 & w23694;
assign w23697 = ~w23695 & ~w23696;
assign w23698 = ~w23658 & w23697;
assign w23699 = w23658 & ~w23697;
assign w23700 = ~w23698 & ~w23699;
assign w23701 = w23657 & w23700;
assign w23702 = ~w23657 & ~w23700;
assign w23703 = ~w23701 & ~w23702;
assign w23704 = ~w23643 & w23703;
assign w23705 = w23643 & ~w23703;
assign w23706 = ~w23704 & ~w23705;
assign w23707 = (w22175 & w25401) | (w22175 & w25402) | (w25401 & w25402);
assign w23708 = (~w22175 & w25654) | (~w22175 & w25655) | (w25654 & w25655);
assign w23709 = ~w23707 & ~w23708;
assign w23710 = ~w23696 & ~w23698;
assign w23711 = b[59] & w10496;
assign w23712 = b[61] & w10148;
assign w23713 = b[60] & w10146;
assign w23714 = w10141 & w11400;
assign w23715 = ~w23712 & ~w23713;
assign w23716 = ~w23711 & w23715;
assign w23717 = ~w23714 & w23716;
assign w23718 = a[59] & ~w23717;
assign w23719 = ~a[59] & w23717;
assign w23720 = ~w23718 & ~w23719;
assign w23721 = ~w23688 & ~w23692;
assign w23722 = b[54] & w11921;
assign w23723 = b[55] & w11923;
assign w23724 = ~w23722 & ~w23723;
assign w23725 = ~w23672 & ~w23676;
assign w23726 = w23724 & ~w23725;
assign w23727 = ~w23724 & w23725;
assign w23728 = ~w23726 & ~w23727;
assign w23729 = b[56] & w11561;
assign w23730 = b[58] & w11196;
assign w23731 = b[57] & w11194;
assign w23732 = ~w10339 & w11189;
assign w23733 = ~w23730 & ~w23731;
assign w23734 = ~w23729 & w23733;
assign w23735 = ~w23732 & w23734;
assign w23736 = a[62] & ~w23735;
assign w23737 = ~a[62] & w23735;
assign w23738 = ~w23736 & ~w23737;
assign w23739 = w23728 & w23738;
assign w23740 = ~w23728 & ~w23738;
assign w23741 = ~w23739 & ~w23740;
assign w23742 = w23721 & ~w23741;
assign w23743 = ~w23721 & w23741;
assign w23744 = ~w23742 & ~w23743;
assign w23745 = w23720 & w23744;
assign w23746 = ~w23720 & ~w23744;
assign w23747 = ~w23745 & ~w23746;
assign w23748 = w23710 & ~w23747;
assign w23749 = ~w23710 & w23747;
assign w23750 = ~w23748 & ~w23749;
assign w23751 = b[62] & w9482;
assign w23752 = b[63] & w9165;
assign w23753 = w9158 & w12156;
assign w23754 = ~w23751 & ~w23752;
assign w23755 = ~w23753 & w23754;
assign w23756 = a[56] & w23755;
assign w23757 = ~a[56] & ~w23755;
assign w23758 = ~w23756 & ~w23757;
assign w23759 = w23750 & ~w23758;
assign w23760 = ~w23750 & w23758;
assign w23761 = ~w23759 & ~w23760;
assign w23762 = ~w23655 & ~w23701;
assign w23763 = w23761 & ~w23762;
assign w23764 = ~w23761 & w23762;
assign w23765 = ~w23763 & ~w23764;
assign w23766 = (~w22175 & w25403) | (~w22175 & w25404) | (w25403 & w25404);
assign w23767 = (w22175 & w25656) | (w22175 & w25657) | (w25656 & w25657);
assign w23768 = ~w23766 & ~w23767;
assign w23769 = b[60] & w10496;
assign w23770 = b[61] & w10146;
assign w23771 = b[62] & w10148;
assign w23772 = w10141 & w11763;
assign w23773 = ~w23770 & ~w23771;
assign w23774 = ~w23769 & w23773;
assign w23775 = ~w23772 & w23774;
assign w23776 = a[59] & ~w23775;
assign w23777 = ~a[59] & w23775;
assign w23778 = ~w23776 & ~w23777;
assign w23779 = ~w23726 & ~w23739;
assign w23780 = b[57] & w11561;
assign w23781 = b[58] & w11194;
assign w23782 = b[59] & w11196;
assign w23783 = w10371 & w11189;
assign w23784 = ~w23781 & ~w23782;
assign w23785 = ~w23780 & w23784;
assign w23786 = ~w23783 & w23785;
assign w23787 = a[62] & ~w23786;
assign w23788 = ~a[62] & w23786;
assign w23789 = ~w23787 & ~w23788;
assign w23790 = b[55] & w11921;
assign w23791 = b[56] & w11923;
assign w23792 = ~w23790 & ~w23791;
assign w23793 = w23724 & ~w23792;
assign w23794 = ~w23724 & w23792;
assign w23795 = ~w23793 & ~w23794;
assign w23796 = w23789 & w23795;
assign w23797 = ~w23789 & ~w23795;
assign w23798 = ~w23796 & ~w23797;
assign w23799 = ~w23779 & w23798;
assign w23800 = w23779 & ~w23798;
assign w23801 = ~w23799 & ~w23800;
assign w23802 = w23778 & w23801;
assign w23803 = ~w23778 & ~w23801;
assign w23804 = ~w23802 & ~w23803;
assign w23805 = ~w23743 & ~w23745;
assign w23806 = w9158 & ~w12154;
assign w23807 = ~w9482 & ~w23806;
assign w23808 = b[63] & ~w23807;
assign w23809 = a[56] & ~w23808;
assign w23810 = ~a[56] & w23808;
assign w23811 = ~w23809 & ~w23810;
assign w23812 = ~w23805 & ~w23811;
assign w23813 = w23805 & w23811;
assign w23814 = ~w23812 & ~w23813;
assign w23815 = ~w23804 & ~w23814;
assign w23816 = w23804 & w23814;
assign w23817 = ~w23815 & ~w23816;
assign w23818 = ~w23749 & ~w23759;
assign w23819 = ~w23817 & w23818;
assign w23820 = w23817 & ~w23818;
assign w23821 = ~w23819 & ~w23820;
assign w23822 = (~w22175 & w25405) | (~w22175 & w25406) | (w25405 & w25406);
assign w23823 = (w22175 & w25658) | (w22175 & w25659) | (w25658 & w25659);
assign w23824 = ~w23822 & ~w23823;
assign w23825 = b[58] & w11561;
assign w23826 = b[60] & w11196;
assign w23827 = b[59] & w11194;
assign w23828 = w11035 & w11189;
assign w23829 = ~w23826 & ~w23827;
assign w23830 = ~w23825 & w23829;
assign w23831 = ~w23828 & w23830;
assign w23832 = a[62] & ~w23831;
assign w23833 = ~a[62] & w23831;
assign w23834 = ~w23832 & ~w23833;
assign w23835 = ~w23793 & ~w23796;
assign w23836 = b[56] & w11921;
assign w23837 = b[57] & w11923;
assign w23838 = ~w23836 & ~w23837;
assign w23839 = ~a[56] & ~w23838;
assign w23840 = a[56] & w23838;
assign w23841 = ~w23839 & ~w23840;
assign w23842 = ~w23724 & w23841;
assign w23843 = w23724 & ~w23841;
assign w23844 = ~w23842 & ~w23843;
assign w23845 = ~w23835 & w23844;
assign w23846 = w23835 & ~w23844;
assign w23847 = ~w23845 & ~w23846;
assign w23848 = w23834 & w23847;
assign w23849 = ~w23834 & ~w23847;
assign w23850 = ~w23848 & ~w23849;
assign w23851 = ~w23799 & ~w23802;
assign w23852 = b[61] & w10496;
assign w23853 = b[62] & w10146;
assign w23854 = b[63] & w10148;
assign w23855 = w10141 & w12132;
assign w23856 = ~w23853 & ~w23854;
assign w23857 = ~w23852 & w23856;
assign w23858 = ~w23855 & w23857;
assign w23859 = a[59] & ~w23858;
assign w23860 = ~a[59] & w23858;
assign w23861 = ~w23859 & ~w23860;
assign w23862 = ~w23851 & w23861;
assign w23863 = w23851 & ~w23861;
assign w23864 = ~w23862 & ~w23863;
assign w23865 = ~w23850 & ~w23864;
assign w23866 = w23850 & w23864;
assign w23867 = ~w23865 & ~w23866;
assign w23868 = ~w23812 & ~w23816;
assign w23869 = ~w23867 & w23868;
assign w23870 = w23867 & ~w23868;
assign w23871 = ~w23869 & ~w23870;
assign w23872 = (w22175 & w25660) | (w22175 & w25661) | (w25660 & w25661);
assign w23873 = (~w22175 & w25407) | (~w22175 & w25408) | (w25407 & w25408);
assign w23874 = ~w23872 & ~w23873;
assign w23875 = ~w23845 & ~w23848;
assign w23876 = b[57] & w11921;
assign w23877 = b[58] & w11923;
assign w23878 = ~w23876 & ~w23877;
assign w23879 = ~w23839 & ~w23842;
assign w23880 = w23878 & ~w23879;
assign w23881 = ~w23878 & w23879;
assign w23882 = ~w23880 & ~w23881;
assign w23883 = b[59] & w11561;
assign w23884 = b[61] & w11196;
assign w23885 = b[60] & w11194;
assign w23886 = w11189 & w11400;
assign w23887 = ~w23884 & ~w23885;
assign w23888 = ~w23883 & w23887;
assign w23889 = ~w23886 & w23888;
assign w23890 = a[62] & ~w23889;
assign w23891 = ~a[62] & w23889;
assign w23892 = ~w23890 & ~w23891;
assign w23893 = w23882 & w23892;
assign w23894 = ~w23882 & ~w23892;
assign w23895 = ~w23893 & ~w23894;
assign w23896 = w23875 & ~w23895;
assign w23897 = ~w23875 & w23895;
assign w23898 = ~w23896 & ~w23897;
assign w23899 = b[62] & w10496;
assign w23900 = b[63] & w10146;
assign w23901 = w10141 & w12156;
assign w23902 = ~w23899 & ~w23900;
assign w23903 = ~w23901 & w23902;
assign w23904 = a[59] & w23903;
assign w23905 = ~a[59] & ~w23903;
assign w23906 = ~w23904 & ~w23905;
assign w23907 = w23898 & ~w23906;
assign w23908 = ~w23898 & w23906;
assign w23909 = ~w23907 & ~w23908;
assign w23910 = ~w23862 & ~w23866;
assign w23911 = ~w23909 & w23910;
assign w23912 = w23909 & ~w23910;
assign w23913 = ~w23911 & ~w23912;
assign w23914 = (~w22175 & w25409) | (~w22175 & w25410) | (w25409 & w25410);
assign w23915 = (w22175 & w25662) | (w22175 & w25663) | (w25662 & w25663);
assign w23916 = ~w23914 & ~w23915;
assign w23917 = ~w23897 & ~w23907;
assign w23918 = b[60] & w11561;
assign w23919 = b[61] & w11194;
assign w23920 = b[62] & w11196;
assign w23921 = w11189 & w11763;
assign w23922 = ~w23919 & ~w23920;
assign w23923 = ~w23918 & w23922;
assign w23924 = ~w23921 & w23923;
assign w23925 = a[62] & ~w23924;
assign w23926 = ~a[62] & w23924;
assign w23927 = ~w23925 & ~w23926;
assign w23928 = w10141 & ~w12154;
assign w23929 = ~w10496 & ~w23928;
assign w23930 = b[63] & ~w23929;
assign w23931 = ~a[59] & ~w23930;
assign w23932 = a[59] & w23930;
assign w23933 = ~w23931 & ~w23932;
assign w23934 = w23927 & w23933;
assign w23935 = ~w23927 & ~w23933;
assign w23936 = ~w23934 & ~w23935;
assign w23937 = ~w23880 & ~w23893;
assign w23938 = b[58] & w11921;
assign w23939 = b[59] & w11923;
assign w23940 = ~w23938 & ~w23939;
assign w23941 = w23878 & ~w23940;
assign w23942 = ~w23878 & w23940;
assign w23943 = ~w23941 & ~w23942;
assign w23944 = w23937 & w23943;
assign w23945 = ~w23937 & ~w23943;
assign w23946 = ~w23944 & ~w23945;
assign w23947 = w23936 & ~w23946;
assign w23948 = ~w23936 & w23946;
assign w23949 = ~w23947 & ~w23948;
assign w23950 = ~w23917 & w23949;
assign w23951 = w23917 & ~w23949;
assign w23952 = ~w23950 & ~w23951;
assign w23953 = (~w22175 & w25411) | (~w22175 & w25412) | (w25411 & w25412);
assign w23954 = (w22175 & w25664) | (w22175 & w25665) | (w25664 & w25665);
assign w23955 = ~w23953 & ~w23954;
assign w23956 = ~w23934 & ~w23947;
assign w23957 = b[59] & w11921;
assign w23958 = b[60] & w11923;
assign w23959 = ~w23957 & ~w23958;
assign w23960 = ~a[59] & ~w23940;
assign w23961 = a[59] & w23940;
assign w23962 = ~w23960 & ~w23961;
assign w23963 = w23959 & ~w23962;
assign w23964 = ~w23959 & w23962;
assign w23965 = ~w23963 & ~w23964;
assign w23966 = b[61] & w11561;
assign w23967 = b[63] & w11196;
assign w23968 = b[62] & w11194;
assign w23969 = w11189 & w12132;
assign w23970 = ~w23967 & ~w23968;
assign w23971 = ~w23966 & w23970;
assign w23972 = ~w23969 & w23971;
assign w23973 = a[62] & ~w23972;
assign w23974 = ~a[62] & w23972;
assign w23975 = ~w23973 & ~w23974;
assign w23976 = w23965 & w23975;
assign w23977 = ~w23965 & ~w23975;
assign w23978 = ~w23976 & ~w23977;
assign w23979 = ~w23941 & ~w23944;
assign w23980 = w23978 & w23979;
assign w23981 = ~w23978 & ~w23979;
assign w23982 = ~w23980 & ~w23981;
assign w23983 = w23956 & ~w23982;
assign w23984 = ~w23956 & w23982;
assign w23985 = ~w23983 & ~w23984;
assign w23986 = (w23335 & w25081) | (w23335 & w25082) | (w25081 & w25082);
assign w23987 = (~w23335 & w25083) | (~w23335 & w25084) | (w25083 & w25084);
assign w23988 = ~w23986 & ~w23987;
assign w23989 = ~w23976 & ~w23980;
assign w23990 = b[60] & w11921;
assign w23991 = b[61] & w11923;
assign w23992 = ~w23990 & ~w23991;
assign w23993 = ~w23960 & ~w23964;
assign w23994 = w23992 & ~w23993;
assign w23995 = ~w23992 & w23993;
assign w23996 = ~w23994 & ~w23995;
assign w23997 = b[62] & w11561;
assign w23998 = b[63] & w11194;
assign w23999 = w11189 & w12156;
assign w24000 = ~w23997 & ~w23998;
assign w24001 = ~w23999 & w24000;
assign w24002 = a[62] & ~w24001;
assign w24003 = ~a[62] & w24001;
assign w24004 = ~w24002 & ~w24003;
assign w24005 = w23996 & w24004;
assign w24006 = ~w23996 & ~w24004;
assign w24007 = ~w24005 & ~w24006;
assign w24008 = w23989 & ~w24007;
assign w24009 = ~w23989 & w24007;
assign w24010 = ~w24008 & ~w24009;
assign w24011 = (~w23335 & w25085) | (~w23335 & w25086) | (w25085 & w25086);
assign w24012 = (w23335 & w25087) | (w23335 & w25088) | (w25087 & w25088);
assign w24013 = ~w24011 & ~w24012;
assign w24014 = ~w23994 & ~w24005;
assign w24015 = b[61] & w11921;
assign w24016 = b[62] & w11923;
assign w24017 = ~w24015 & ~w24016;
assign w24018 = w23992 & ~w24017;
assign w24019 = ~w23992 & w24017;
assign w24020 = ~w24018 & ~w24019;
assign w24021 = w11189 & ~w12154;
assign w24022 = ~w11561 & ~w24021;
assign w24023 = b[63] & ~w24022;
assign w24024 = a[62] & ~w24023;
assign w24025 = ~a[62] & w24023;
assign w24026 = ~w24024 & ~w24025;
assign w24027 = w24020 & ~w24026;
assign w24028 = ~w24020 & w24026;
assign w24029 = ~w24027 & ~w24028;
assign w24030 = w24014 & ~w24029;
assign w24031 = ~w24014 & w24029;
assign w24032 = ~w24030 & ~w24031;
assign w24033 = (~w23335 & w25089) | (~w23335 & w25090) | (w25089 & w25090);
assign w24034 = (w23335 & w25241) | (w23335 & w25242) | (w25241 & w25242);
assign w24035 = ~w24033 & ~w24034;
assign w24036 = ~w24018 & ~w24027;
assign w24037 = b[62] & w11921;
assign w24038 = a[63] & b[63];
assign w24039 = a[62] & ~b[63];
assign w24040 = ~w24038 & ~w24039;
assign w24041 = ~w24037 & ~w24040;
assign w24042 = w23992 & w24041;
assign w24043 = ~w23992 & ~w24041;
assign w24044 = ~w24042 & ~w24043;
assign w24045 = ~w24036 & w24044;
assign w24046 = w24036 & ~w24044;
assign w24047 = ~w24045 & ~w24046;
assign w24048 = (~w20820 & w25709) | (~w20820 & w25710) | (w25709 & w25710);
assign w24049 = (w20820 & w25711) | (w20820 & w25712) | (w25711 & w25712);
assign w24050 = ~w24048 & ~w24049;
assign w24051 = ~w24038 & ~w24043;
assign w24052 = w12128 & w23990;
assign w24053 = ~w24051 & ~w24052;
assign w24054 = (~w20820 & w25713) | (~w20820 & w25714) | (w25713 & w25714);
assign w24055 = (w20820 & w25715) | (w20820 & w25716) | (w25715 & w25716);
assign w24056 = ~w24054 & ~w24055;
assign w24057 = a[0] & b[1];
assign w24058 = w8 & ~w10;
assign w24059 = ~w12 & ~w1;
assign w24060 = w12 & w1;
assign w24061 = ~w12 & w17;
assign w24062 = a[2] & b[0];
assign w24063 = a[0] & b[2];
assign w24064 = w29 & ~w28;
assign w24065 = a[0] & b[3];
assign w24066 = ~b[1] & a[2];
assign w24067 = (a[2] & w39) | (a[2] & w24585) | (w39 & w24585);
assign w24068 = (w47 & w24586) | (w47 & w24587) | (w24586 & w24587);
assign w24069 = w38 & w25757;
assign w24070 = b[0] & a[5];
assign w24071 = ~w69 & ~w57;
assign w24072 = w69 & w57;
assign w24073 = a[0] & b[4];
assign w24074 = ~w5 & w85;
assign w24075 = ~b[2] & a[2];
assign w24076 = ~w34 & ~w52;
assign w24077 = w65 & b[0];
assign w24078 = ~w101 & ~w104;
assign w24079 = ~w78 & ~w77;
assign w24080 = a[0] & b[5];
assign w24081 = ~w119 & ~w120;
assign w24082 = ~w119 & ~a[2];
assign w24083 = ~w117 & ~w122;
assign w24084 = ~w129 & ~w127;
assign w24085 = w65 & b[1];
assign w24086 = (w137 & ~w46) | (w137 & w24588) | (~w46 & w24588);
assign w24087 = w46 & w24589;
assign w24088 = w106 & a[5];
assign w24089 = a[0] & b[6];
assign w24090 = ~w112 & ~w111;
assign w24091 = ~w154 & ~w111;
assign w24092 = ~w154 & w24090;
assign w24093 = ~w5 & w158;
assign w24094 = ~b[4] & a[2];
assign w24095 = a[2] & ~w158;
assign w24096 = a[2] & ~w24093;
assign w24097 = ~w166 & ~w164;
assign w24098 = b[0] & a[8];
assign w24099 = ~w186 & ~w175;
assign w24100 = w186 & w175;
assign w24101 = w65 & b[2];
assign w24102 = a[0] & b[7];
assign w24103 = ~w153 & ~w213;
assign w24104 = w153 & w213;
assign w24105 = ~w5 & w217;
assign w24106 = ~b[5] & a[2];
assign w24107 = a[2] & ~w217;
assign w24108 = a[2] & ~w24105;
assign w24109 = ~b[0] & a[8];
assign w24110 = ~w186 & w229;
assign w24111 = w37 & ~a[5];
assign w24112 = w65 & b[3];
assign w24113 = w251 & a[5];
assign w24114 = ~w253 & ~w254;
assign w24115 = ~w205 & ~w201;
assign w24116 = a[0] & b[8];
assign w24117 = ~w212 & ~w213;
assign w24118 = (~w212 & ~w213) | (~w212 & w24590) | (~w213 & w24590);
assign w24119 = w267 & ~w24117;
assign w24120 = w267 & ~w24118;
assign w24121 = ~w5 & w271;
assign w24122 = ~b[6] & a[2];
assign w24123 = a[2] & ~w271;
assign w24124 = a[2] & ~w24121;
assign w24125 = w170 & ~w223;
assign w24126 = (w287 & ~w46) | (w287 & w24591) | (~w46 & w24591);
assign w24127 = w46 & w24592;
assign w24128 = w65 & b[4];
assign w24129 = ~w304 & a[5];
assign w24130 = w304 & ~a[5];
assign w24131 = ~w258 & ~w256;
assign w24132 = a[0] & b[9];
assign w24133 = ~w266 & ~w319;
assign w24134 = w266 & w319;
assign w24135 = ~w5 & w323;
assign w24136 = ~b[7] & a[2];
assign w24137 = a[2] & ~w323;
assign w24138 = a[2] & ~w24135;
assign w24139 = b[0] & a[11];
assign w24140 = ~w361 & ~w350;
assign w24141 = w361 & w350;
assign w24142 = w65 & b[5];
assign w24143 = ~w66 & w378;
assign w24144 = ~w310 & ~w308;
assign w24145 = a[0] & b[10];
assign w24146 = ~w318 & ~w319;
assign w24147 = (~w318 & ~w319) | (~w318 & w24593) | (~w319 & w24593);
assign w24148 = w394 & ~w24146;
assign w24149 = w394 & ~w24147;
assign w24150 = ~w5 & w398;
assign w24151 = ~b[8] & a[2];
assign w24152 = a[2] & ~w398;
assign w24153 = a[2] & ~w24150;
assign w24154 = ~w331 & ~w330;
assign w24155 = ~w370 & ~w367;
assign w24156 = ~b[0] & a[11];
assign w24157 = ~w361 & w413;
assign w24158 = ~w173 & ~a[8];
assign w24159 = w173 & ~a[7];
assign w24160 = w431 & a[8];
assign w24161 = ~w433 & ~w437;
assign w24162 = w65 & b[6];
assign w24163 = ~w66 & w449;
assign w24164 = ~w386 & ~w384;
assign w24165 = a[0] & b[11];
assign w24166 = ~w393 & ~w24148;
assign w24167 = ~w393 & ~w24149;
assign w24168 = ~w5 & w470;
assign w24169 = ~b[9] & a[2];
assign w24170 = a[2] & ~w470;
assign w24171 = a[2] & ~w24168;
assign w24172 = (w485 & ~w46) | (w485 & w24594) | (~w46 & w24594);
assign w24173 = w46 & w24595;
assign w24174 = ~w502 & a[8];
assign w24175 = w502 & ~a[8];
assign w24176 = ~w441 & ~w440;
assign w24177 = w65 & b[7];
assign w24178 = ~w66 & w517;
assign w24179 = a[0] & b[12];
assign w24180 = ~w465 & ~w464;
assign w24181 = ~w533 & ~w464;
assign w24182 = ~w533 & w24180;
assign w24183 = w533 & w464;
assign w24184 = ~w5 & w537;
assign w24185 = ~b[10] & a[2];
assign w24186 = a[2] & ~w537;
assign w24187 = a[2] & ~w24184;
assign w24188 = ~w478 & ~w476;
assign w24189 = b[0] & a[14];
assign w24190 = ~w576 & ~w565;
assign w24191 = w576 & w565;
assign w24192 = ~w179 & w593;
assign w24193 = ~w508 & ~w506;
assign w24194 = w65 & b[8];
assign w24195 = ~w66 & w609;
assign w24196 = ~w524 & ~w523;
assign w24197 = a[0] & b[13];
assign w24198 = ~w532 & ~w24183;
assign w24199 = (~w532 & w24180) | (~w532 & w24596) | (w24180 & w24596);
assign w24200 = w625 & ~w24198;
assign w24201 = w625 & ~w24199;
assign w24202 = ~w625 & w24198;
assign w24203 = ~w625 & w24199;
assign w24204 = ~w5 & w629;
assign w24205 = ~b[11] & a[2];
assign w24206 = a[2] & ~w629;
assign w24207 = a[2] & ~w24204;
assign w24208 = ~b[0] & a[14];
assign w24209 = ~w576 & w642;
assign w24210 = ~w348 & ~a[11];
assign w24211 = w348 & ~a[10];
assign w24212 = w660 & a[11];
assign w24213 = ~w662 & ~w666;
assign w24214 = ~w585 & ~w582;
assign w24215 = ~w179 & w679;
assign w24216 = w601 & ~w598;
assign w24217 = w65 & b[9];
assign w24218 = ~w66 & w695;
assign w24219 = a[0] & b[14];
assign w24220 = ~w624 & ~w24200;
assign w24221 = ~w624 & ~w24201;
assign w24222 = ~w5 & w715;
assign w24223 = ~b[12] & a[2];
assign w24224 = a[2] & ~w715;
assign w24225 = a[2] & ~w24222;
assign w24226 = ~w637 & ~w636;
assign w24227 = w65 & b[10];
assign w24228 = ~w66 & w733;
assign w24229 = (w742 & ~w46) | (w742 & w24597) | (~w46 & w24597);
assign w24230 = w46 & w24598;
assign w24231 = ~w759 & a[11];
assign w24232 = w759 & ~a[11];
assign w24233 = ~w670 & ~w668;
assign w24234 = ~w179 & w774;
assign w24235 = ~w702 & ~w701;
assign w24236 = a[0] & b[15];
assign w24237 = ~w710 & ~w709;
assign w24238 = w796 & ~w709;
assign w24239 = w796 & w24237;
assign w24240 = ~w5 & w800;
assign w24241 = ~b[13] & a[2];
assign w24242 = ~w765 & ~w763;
assign w24243 = b[0] & a[17];
assign w24244 = ~w839 & ~w828;
assign w24245 = w839 & w828;
assign w24246 = ~w354 & w856;
assign w24247 = ~w179 & w871;
assign w24248 = ~w781 & ~w780;
assign w24249 = w65 & b[11];
assign w24250 = ~w66 & w887;
assign w24251 = a[0] & b[16];
assign w24252 = ~w794 & ~w24238;
assign w24253 = ~w794 & ~w24239;
assign w24254 = ~w902 & ~w24252;
assign w24255 = ~w902 & ~w24253;
assign w24256 = ~w5 & w906;
assign w24257 = ~b[14] & a[2];
assign w24258 = a[2] & ~w906;
assign w24259 = a[2] & ~w24256;
assign w24260 = ~w808 & ~w806;
assign w24261 = w65 & b[12];
assign w24262 = ~w66 & w923;
assign w24263 = ~b[0] & a[17];
assign w24264 = ~w839 & w929;
assign w24265 = ~w563 & ~a[14];
assign w24266 = w563 & ~a[13];
assign w24267 = w947 & a[14];
assign w24268 = ~w949 & ~w953;
assign w24269 = ~w848 & ~w845;
assign w24270 = ~w354 & w966;
assign w24271 = ~w813 & ~w861;
assign w24272 = ~w179 & w982;
assign w24273 = ~w894 & ~w892;
assign w24274 = a[0] & b[17];
assign w24275 = ~w901 & ~w24252;
assign w24276 = ~w901 & ~w24253;
assign w24277 = w900 & ~w1004;
assign w24278 = ~w900 & w1004;
assign w24279 = ~w5 & w1009;
assign w24280 = ~b[15] & a[2];
assign w24281 = a[2] & ~w1009;
assign w24282 = a[2] & ~w24279;
assign w24283 = ~w179 & w1027;
assign w24284 = (w1036 & ~w46) | (w1036 & w24599) | (~w46 & w24599);
assign w24285 = w46 & w24600;
assign w24286 = ~w1053 & a[14];
assign w24287 = w1053 & ~a[14];
assign w24288 = ~w957 & ~w955;
assign w24289 = ~w354 & w1068;
assign w24290 = ~w989 & ~w987;
assign w24291 = w65 & b[13];
assign w24292 = ~w66 & w1090;
assign w24293 = ~a[5] & w1090;
assign w24294 = ~a[5] & w24292;
assign w24295 = a[0] & b[18];
assign w24296 = (~w1003 & ~w1004) | (~w1003 & w24601) | (~w1004 & w24601);
assign w24297 = w1105 & ~w1003;
assign w24298 = w1105 & w24296;
assign w24299 = ~w5 & w1109;
assign w24300 = ~b[16] & a[2];
assign w24301 = ~w1017 & ~w1016;
assign w24302 = w65 & b[14];
assign w24303 = ~w66 & w1126;
assign w24304 = ~w1059 & ~w1057;
assign w24305 = b[0] & a[20];
assign w24306 = ~w1157 & ~w1146;
assign w24307 = w1157 & w1146;
assign w24308 = ~w569 & w1174;
assign w24309 = ~w354 & w1189;
assign w24310 = ~w1075 & ~w1073;
assign w24311 = ~w179 & w1205;
assign w24312 = ~w1097 & ~w1096;
assign w24313 = a[0] & b[19];
assign w24314 = ~w1103 & ~w24297;
assign w24315 = ~w1103 & ~w24298;
assign w24316 = w1228 & ~w24314;
assign w24317 = w1228 & ~w24315;
assign w24318 = ~w5 & w1232;
assign w24319 = ~b[17] & a[2];
assign w24320 = ~w179 & w1250;
assign w24321 = (a[17] & ~w1260) | (a[17] & w24602) | (~w1260 & w24602);
assign w24322 = w1260 & w24603;
assign w24323 = ~b[0] & a[20];
assign w24324 = ~w1157 & w1264;
assign w24325 = ~w1166 & ~w1163;
assign w24326 = ~w569 & w1291;
assign w24327 = ~w1131 & ~w1180;
assign w24328 = ~w354 & w1307;
assign w24329 = ~w1212 & ~w1210;
assign w24330 = w65 & b[15];
assign w24331 = ~w66 & w1329;
assign w24332 = a[0] & b[20];
assign w24333 = ~w1226 & ~w24316;
assign w24334 = ~w1226 & ~w24317;
assign w24335 = ~w1344 & ~w24333;
assign w24336 = ~w1344 & ~w24334;
assign w24337 = w1344 & w24333;
assign w24338 = w1344 & w24334;
assign w24339 = ~w5 & w1348;
assign w24340 = ~b[18] & a[2];
assign w24341 = a[2] & ~w1348;
assign w24342 = a[2] & ~w24339;
assign w24343 = ~w1240 & ~w1239;
assign w24344 = w65 & b[16];
assign w24345 = ~w66 & w1365;
assign w24346 = ~a[5] & w1365;
assign w24347 = ~a[5] & w24345;
assign w24348 = (w1375 & ~w46) | (w1375 & w24742) | (~w46 & w24742);
assign w24349 = w46 & w24743;
assign w24350 = ~w1392 & a[17];
assign w24351 = w1392 & ~a[17];
assign w24352 = ~w1282 & ~w1280;
assign w24353 = w48 & ~w49;
assign w24354 = ~w5 & w123;
assign w24355 = ~w1336 & ~w1334;
assign w24356 = ~w1478 & ~w1477;
assign w24357 = ~w1579 & ~w1577;
assign w24358 = ~w1736 & ~w1734;
assign w24359 = ~w1883 & ~w1881;
assign w24360 = ~w2072 & ~w2070;
assign w24361 = ~w2177 & ~w2175;
assign w24362 = ~w2341 & ~w2339;
assign w24363 = ~w2529 & ~w2528;
assign w24364 = ~w2721 & ~w2720;
assign w24365 = ~w2919 & ~w2917;
assign w24366 = ~w3044 & ~w3043;
assign w24367 = ~w3255 & ~w3254;
assign w24368 = ~w3456 & ~w3455;
assign w24369 = ~w3675 & ~w3674;
assign w24370 = ~w3898 & ~w3897;
assign w24371 = ~w4117 & ~w4116;
assign w24372 = ~w4368 & ~w4367;
assign w24373 = ~w4525 & ~w4523;
assign w24374 = ~w4754 & ~w4753;
assign w24375 = ~w5017 & ~w5016;
assign w24376 = ~w5266 & ~w5265;
assign w24377 = ~w5529 & ~w5528;
assign w24378 = ~w5798 & ~w5796;
assign w24379 = ~w6080 & ~w6078;
assign w24380 = ~w6008 & ~w6006;
assign w24381 = ~w6278 & ~w6276;
assign w24382 = ~w6565 & ~w6564;
assign w24383 = ~w6847 & ~w6845;
assign w24384 = ~w7144 & ~w7143;
assign w24385 = ~w7448 & ~w7447;
assign w24386 = ~w7746 & ~w7745;
assign w24387 = ~w8069 & ~w8067;
assign w24388 = ~w8290 & ~w8288;
assign w24389 = ~w8638 & ~w8637;
assign w24390 = ~w8951 & ~w8949;
assign w24391 = ~w9298 & ~w9297;
assign w24392 = ~w9632 & ~w9631;
assign w24393 = ~w9973 & ~w9971;
assign w24394 = ~w10348 & w10698;
assign w24395 = ~w10640 & ~w10639;
assign w24396 = ~w10977 & ~w10976;
assign w24397 = ~w11349 & ~w11347;
assign w24398 = ~w11412 & w11778;
assign w24399 = ~w11731 & ~w11730;
assign w24400 = ~w11783 & ~w12146;
assign w24401 = ~w12508 & ~w12507;
assign w24402 = ~w12862 & w13209;
assign w24403 = ~w13207 & w13557;
assign w24404 = (~w13556 & ~w13557) | (~w13556 & w24604) | (~w13557 & w24604);
assign w24405 = ~w13903 & ~w13902;
assign w24406 = ~w14244 & ~w14243;
assign w24407 = w14575 & ~w14243;
assign w24408 = ~w14244 & w24407;
assign w24409 = w14573 & w14904;
assign w24410 = ~w14903 & ~w14904;
assign w24411 = (~w14903 & ~w14904) | (~w14903 & w24605) | (~w14904 & w24605);
assign w24412 = (~w15226 & ~w24410) | (~w15226 & w25634) | (~w24410 & w25634);
assign w24413 = (~w15226 & ~w24411) | (~w15226 & w25634) | (~w24411 & w25634);
assign w24414 = w15540 & w15847;
assign w24415 = ~w15844 & ~w15847;
assign w24416 = (~w15844 & ~w15847) | (~w15844 & w24606) | (~w15847 & w24606);
assign w24417 = ~w16150 & w24415;
assign w24418 = ~w16150 & w24416;
assign w24419 = ~w16151 & ~w24417;
assign w24420 = ~w16151 & ~w24418;
assign w24421 = ~w16444 & ~w24419;
assign w24422 = ~w16444 & ~w24420;
assign w24423 = ~w16737 & ~w16734;
assign w24424 = w17026 & w16734;
assign w24425 = (w17026 & w16737) | (w17026 & w24424) | (w16737 & w24424);
assign w24426 = ~w17025 & ~w24424;
assign w24427 = ~w17025 & ~w24425;
assign w24428 = w17305 & ~w24426;
assign w24429 = w17305 & ~w24427;
assign w24430 = ~w17304 & ~w24428;
assign w24431 = ~w17304 & ~w24429;
assign w24432 = w17576 & ~w24430;
assign w24433 = w17576 & ~w24431;
assign w24434 = ~w17575 & ~w24432;
assign w24435 = ~w17575 & ~w24433;
assign w24436 = ~w17844 & w24434;
assign w24437 = ~w17844 & w24435;
assign w24438 = ~w17845 & ~w24436;
assign w24439 = ~w17845 & ~w24437;
assign w24440 = ~w18103 & ~w24438;
assign w24441 = ~w18103 & ~w24439;
assign w24442 = (~w18359 & ~w18361) | (~w18359 & w25413) | (~w18361 & w25413);
assign w24443 = (~w18613 & ~w18614) | (~w18613 & w24744) | (~w18614 & w24744);
assign w24444 = (~w18613 & w24442) | (~w18613 & w24607) | (w24442 & w24607);
assign w24445 = (~w18857 & w24443) | (~w18857 & w24745) | (w24443 & w24745);
assign w24446 = (~w18857 & w24444) | (~w18857 & w24745) | (w24444 & w24745);
assign w24447 = (~w19100 & w24445) | (~w19100 & w25534) | (w24445 & w25534);
assign w24448 = (~w19100 & w24446) | (~w19100 & w25534) | (w24446 & w25534);
assign w24449 = w19341 & w24447;
assign w24450 = w19341 & w24448;
assign w24451 = ~w19340 & ~w24449;
assign w24452 = (~w19340 & ~w24448) | (~w19340 & w25635) | (~w24448 & w25635);
assign w24453 = w19570 & w24451;
assign w24454 = w19570 & w24452;
assign w24455 = ~w19569 & ~w24453;
assign w24456 = ~w19569 & ~w24454;
assign w24457 = w19797 & ~w24455;
assign w24458 = w19797 & ~w24456;
assign w24459 = ~w19795 & ~w24457;
assign w24460 = ~w19795 & ~w24458;
assign w24461 = w20018 & ~w24459;
assign w24462 = w20018 & ~w24460;
assign w24463 = w20017 & w20231;
assign w24464 = ~w20230 & ~w20231;
assign w24465 = ~w20230 & ~w24463;
assign w24466 = w20436 & ~w24464;
assign w24467 = w20436 & ~w24465;
assign w24468 = ~w20435 & ~w24466;
assign w24469 = ~w20435 & ~w24467;
assign w24470 = ~w20630 & w24468;
assign w24471 = ~w20630 & w24469;
assign w24472 = ~w20631 & ~w24470;
assign w24473 = ~w20631 & ~w24471;
assign w24474 = ~w20819 & ~w20817;
assign w24475 = w21007 & w20817;
assign w24476 = (w21007 & w20819) | (w21007 & w24475) | (w20819 & w24475);
assign w24477 = ~w21005 & ~w24475;
assign w24478 = ~w21005 & ~w24476;
assign w24479 = w21191 & w24477;
assign w24480 = ~w24476 & w24746;
assign w24481 = (~w21190 & ~w24477) | (~w21190 & w25636) | (~w24477 & w25636);
assign w24482 = ~w21190 & ~w24480;
assign w24483 = w21369 & w24481;
assign w24484 = w21369 & w24482;
assign w24485 = ~w21367 & ~w24483;
assign w24486 = (~w21367 & ~w24482) | (~w21367 & w25637) | (~w24482 & w25637);
assign w24487 = (w21545 & w24483) | (w21545 & w25666) | (w24483 & w25666);
assign w24488 = w21545 & ~w24486;
assign w24489 = ~w21543 & ~w24487;
assign w24490 = (~w21543 & w24486) | (~w21543 & w25667) | (w24486 & w25667);
assign w24491 = w21715 & w24489;
assign w24492 = w21715 & w24490;
assign w24493 = ~w21714 & ~w24491;
assign w24494 = ~w21714 & ~w24492;
assign w24495 = w21873 & w24493;
assign w24496 = w21873 & w24494;
assign w24497 = ~w21872 & ~w24495;
assign w24498 = ~w21872 & ~w24496;
assign w24499 = w22028 & ~w24497;
assign w24500 = w22028 & ~w24498;
assign w24501 = ~w22026 & ~w24499;
assign w24502 = ~w22026 & ~w24500;
assign w24503 = w22173 & w24501;
assign w24504 = w22173 & w24502;
assign w24505 = ~w22172 & w22309;
assign w24506 = (~w22308 & ~w22309) | (~w22308 & w24608) | (~w22309 & w24608);
assign w24507 = w22445 & w22308;
assign w24508 = w22445 & ~w24506;
assign w24509 = (~w22443 & ~w22445) | (~w22443 & w25243) | (~w22445 & w25243);
assign w24510 = (w24608 & w25535) | (w24608 & w25536) | (w25535 & w25536);
assign w24511 = w22576 & w24509;
assign w24512 = w22576 & w24510;
assign w24513 = (~w22575 & ~w22576) | (~w22575 & w25244) | (~w22576 & w25244);
assign w24514 = ~w22575 & ~w24512;
assign w24515 = (w25244 & w25245) | (w25244 & w25537) | (w25245 & w25537);
assign w24516 = ~w24512 & w25245;
assign w24517 = ~w22701 & ~w24515;
assign w24518 = (~w22701 & w24512) | (~w22701 & w25414) | (w24512 & w25414);
assign w24519 = (w22826 & w24515) | (w22826 & w25638) | (w24515 & w25638);
assign w24520 = (~w24512 & w25638) | (~w24512 & w25639) | (w25638 & w25639);
assign w24521 = ~w22824 & ~w24519;
assign w24522 = ~w22824 & ~w24520;
assign w24523 = ~w24519 & w25668;
assign w24524 = ~w24520 & w25668;
assign w24525 = ~w22943 & ~w24523;
assign w24526 = ~w22943 & ~w24524;
assign w24527 = w23053 & w24525;
assign w24528 = w23053 & w24526;
assign w24529 = ~w23052 & ~w24527;
assign w24530 = ~w23052 & ~w24528;
assign w24531 = w23156 & ~w24529;
assign w24532 = w23156 & ~w24530;
assign w24533 = ~w23155 & ~w24531;
assign w24534 = ~w23155 & ~w24532;
assign w24535 = w23248 & ~w24533;
assign w24536 = w23248 & ~w24534;
assign w24537 = ~w23247 & ~w24535;
assign w24538 = ~w23247 & ~w24536;
assign w24539 = ~w23334 & ~w23333;
assign w24540 = w23418 & w23333;
assign w24541 = (w23418 & w23334) | (w23418 & w24540) | (w23334 & w24540);
assign w24542 = ~w23417 & ~w24540;
assign w24543 = ~w23417 & ~w24541;
assign w24544 = w23497 & w24542;
assign w24545 = ~w23495 & ~w24544;
assign w24546 = (~w23495 & ~w24543) | (~w23495 & w24748) | (~w24543 & w24748);
assign w24547 = ~w24544 & w24909;
assign w24548 = w23569 & w24546;
assign w24549 = ~w23568 & ~w24547;
assign w24550 = (~w23568 & ~w24546) | (~w23568 & w24910) | (~w24546 & w24910);
assign w24551 = (w23639 & w24547) | (w23639 & w25246) | (w24547 & w25246);
assign w24552 = (w24546 & w25246) | (w24546 & w25247) | (w25246 & w25247);
assign w24553 = (~w24546 & w25417) | (~w24546 & w25416) | (w25417 & w25416);
assign w24554 = (w24547 & w25640) | (w24547 & w25641) | (w25640 & w25641);
assign w24555 = (~w23705 & ~w24553) | (~w23705 & w25540) | (~w24553 & w25540);
assign w24556 = w23765 & w24554;
assign w24557 = (~w24553 & w25642) | (~w24553 & w25643) | (w25642 & w25643);
assign w24558 = (~w23763 & ~w24554) | (~w23763 & w25669) | (~w24554 & w25669);
assign w24559 = ~w23763 & ~w24557;
assign w24560 = w23821 & ~w24558;
assign w24561 = (w23821 & w24557) | (w23821 & w25670) | (w24557 & w25670);
assign w24562 = ~w23820 & ~w24560;
assign w24563 = ~w23820 & ~w24561;
assign w24564 = w23871 & ~w24562;
assign w24565 = w23871 & ~w24563;
assign w24566 = ~w23870 & ~w24564;
assign w24567 = ~w23870 & ~w24565;
assign w24568 = w23913 & ~w24566;
assign w24569 = w23913 & ~w24567;
assign w24570 = ~w23912 & ~w24568;
assign w24571 = ~w23912 & ~w24569;
assign w24572 = w23952 & ~w24570;
assign w24573 = w23952 & ~w24571;
assign w24574 = ~w23950 & ~w23984;
assign w24575 = ~w24574 & ~w23983;
assign w24576 = ~w24010 & ~w24009;
assign w24577 = w24032 & w24009;
assign w24578 = w24032 & ~w24576;
assign w24579 = ~w24031 & ~w24577;
assign w24580 = ~w24031 & ~w24578;
assign w24581 = w24047 & w24579;
assign w24582 = w24047 & w24580;
assign w24583 = ~w24046 & ~w24581;
assign w24584 = ~w24046 & ~w24582;
assign w24585 = w40 & a[2];
assign w24586 = ~w38 & a[2];
assign w24587 = ~w38 & w24067;
assign w24588 = ~w66 & w137;
assign w24589 = w66 & ~w137;
assign w24590 = ~w153 & ~w212;
assign w24591 = ~w179 & w287;
assign w24592 = w179 & ~w287;
assign w24593 = ~w266 & ~w318;
assign w24594 = ~w354 & w485;
assign w24595 = w354 & ~w485;
assign w24596 = ~w533 & ~w532;
assign w24597 = ~w569 & w742;
assign w24598 = w569 & ~w742;
assign w24599 = ~w832 & w1036;
assign w24600 = w832 & ~w1036;
assign w24601 = w900 & ~w1003;
assign w24602 = w1258 & a[17];
assign w24603 = ~w1258 & ~a[17];
assign w24604 = w13207 & ~w13556;
assign w24605 = ~w14573 & ~w14903;
assign w24606 = ~w15540 & ~w15844;
assign w24607 = ~w18614 & ~w18613;
assign w24608 = w22172 & ~w22308;
assign w24609 = w94 & ~w91;
assign w24610 = ~w1314 & ~w1312;
assign w24611 = ~w1398 & ~w1396;
assign w24612 = ~w1415 & ~w1413;
assign w24613 = ~w1448 & ~w1447;
assign w24614 = ~w1530 & ~w1527;
assign w24615 = ~w1494 & ~w1545;
assign w24616 = ~w1602 & ~w1601;
assign w24617 = (w1806 & ~w46) | (w1806 & w24749) | (~w46 & w24749);
assign w24618 = w46 & w24750;
assign w24619 = ~w1766 & ~w1765;
assign w24620 = ~w1507 & ~a[23];
assign w24621 = w1507 & ~a[22];
assign w24622 = ~w1968 & ~w1965;
assign w24623 = (w2260 & ~w46) | (w2260 & w24751) | (~w46 & w24751);
assign w24624 = w46 & w24752;
assign w24625 = ~w1945 & ~a[26];
assign w24626 = w1945 & ~a[25];
assign w24627 = ~w2449 & ~w2446;
assign w24628 = ~w2465 & ~w2464;
assign w24629 = w2479 & w2679;
assign w24630 = ~w2555 & ~w2554;
assign w24631 = (w2783 & ~w46) | (w2783 & w24753) | (~w46 & w24753);
assign w24632 = ~w2684 & ~w2682;
assign w24633 = ~w2798 & ~w2796;
assign w24634 = w46 & w24754;
assign w24635 = ~w2855 & ~w2853;
assign w24636 = ~w3075 & ~w3073;
assign w24637 = ~w2426 & ~a[29];
assign w24638 = w2426 & ~a[28];
assign w24639 = w2995 & ~w2988;
assign w24640 = ~w3275 & ~w3273;
assign w24641 = ~w3486 & ~w3484;
assign w24642 = ~w3721 & ~w3719;
assign w24643 = ~w3581 & w3778;
assign w24644 = w3779 & w3990;
assign w24645 = ~w3779 & ~w3990;
assign w24646 = w4240 & b[1];
assign w24647 = w46 & w25091;
assign w24648 = (~a[38] & ~w46) | (~a[38] & w25092) | (~w46 & w25092);
assign w24649 = ~w4463 & ~w4461;
assign w24650 = ~w4479 & ~w4477;
assign w24651 = ~w4519 & ~w4518;
assign w24652 = ~w4578 & ~w4577;
assign w24653 = ~w4708 & ~w4707;
assign w24654 = ~w4646 & ~w4656;
assign w24655 = ~w4725 & ~w4724;
assign w24656 = ~w4748 & ~w4747;
assign w24657 = ~w5011 & ~w5010;
assign w24658 = ~w5260 & ~w5258;
assign w24659 = ~w5523 & ~w5522;
assign w24660 = ~w5791 & ~w5790;
assign w24661 = ~w6057 & ~w6055;
assign w24662 = ~w6345 & ~w6344;
assign w24663 = ~w6545 & ~w6544;
assign w24664 = ~w6522 & ~w6520;
assign w24665 = ~w6502 & ~w6500;
assign w24666 = ~w6516 & ~w6515;
assign w24667 = ~w6552 & ~w6550;
assign w24668 = ~w6609 & ~w6607;
assign w24669 = ~w6804 & ~w6802;
assign w24670 = ~w6775 & ~w6773;
assign w24671 = ~w6834 & ~w6832;
assign w24672 = ~w7122 & ~w7120;
assign w24673 = ~w7425 & ~w7423;
assign w24674 = ~w7732 & ~w7731;
assign w24675 = ~w8039 & ~w8038;
assign w24676 = ~w8359 & ~w8358;
assign w24677 = ~w8694 & ~w8692;
assign w24678 = ~w8921 & ~w8919;
assign w24679 = ~w8909 & ~w8907;
assign w24680 = ~w8880 & ~w8879;
assign w24681 = ~w8903 & ~w8902;
assign w24682 = ~w8995 & ~w8993;
assign w24683 = ~w9259 & ~w9258;
assign w24684 = ~w9236 & ~w9234;
assign w24685 = ~w9217 & ~w9215;
assign w24686 = ~w9602 & ~w9600;
assign w24687 = ~w9953 & ~w9952;
assign w24688 = ~w10308 & ~w10307;
assign w24689 = ~w10327 & ~w10325;
assign w24690 = ~w24394 & ~w10696;
assign w24691 = ~w10680 & ~w10679;
assign w24692 = ~w11019 & ~w11017;
assign w24693 = w10703 & ~w11048;
assign w24694 = ~w11295 & ~w11294;
assign w24695 = ~w11276 & ~w11275;
assign w24696 = ~w11302 & ~w11300;
assign w24697 = ~w11397 & ~w11396;
assign w24698 = ~w11408 & ~w11389;
assign w24699 = ~w11659 & ~w11657;
assign w24700 = ~w11695 & ~w11694;
assign w24701 = ~w12140 & ~w12121;
assign w24702 = ~w11793 & ~w12115;
assign w24703 = ~w12018 & ~w12016;
assign w24704 = ~w12102 & ~w12100;
assign w24705 = ~w12492 & ~w12490;
assign w24706 = (~w13556 & w24604) | (~w13556 & w25248) | (w24604 & w25248);
assign w24707 = (~w13556 & w24404) | (~w13556 & w24402) | (w24404 & w24402);
assign w24708 = ~w13762 & ~w13774;
assign w24709 = ~w13779 & ~w13791;
assign w24710 = ~w13796 & ~w13808;
assign w24711 = ~w13813 & ~w13588;
assign w24712 = ~w13816 & ~w13828;
assign w24713 = ~w13833 & ~w13845;
assign w24714 = ~w13850 & ~w13862;
assign w24715 = ~w13867 & ~w13574;
assign w24716 = ~w13870 & ~w13882;
assign w24717 = ~w1513 & w17535;
assign w24718 = ~w1150 & w17550;
assign w24719 = ~w1513 & w18077;
assign w24720 = ~w12155 & w1150;
assign w24721 = ~w1513 & w18345;
assign w24722 = ~w2980 & w20410;
assign w24723 = ~w12155 & w2980;
assign w24724 = (w24472 & w24473) | (w24472 & w24462) | (w24473 & w24462);
assign w24725 = (w24472 & w24473) | (w24472 & w24461) | (w24473 & w24461);
assign w24726 = ~w12155 & w4923;
assign w24727 = ~w8195 & w23165;
assign w24728 = ~w7312 & w23234;
assign w24729 = ~w8195 & w23257;
assign w24730 = ~w12155 & w7312;
assign w24731 = b[62] & w7312;
assign w24732 = (~w24009 & w24576) | (~w24009 & w23983) | (w24576 & w23983);
assign w24733 = (~w24009 & w24576) | (~w24009 & ~w24575) | (w24576 & ~w24575);
assign w24734 = w24047 & w25761;
assign w24735 = w24047 & w25762;
assign w24736 = ~w24047 & ~w25762;
assign w24737 = ~w24047 & ~w25761;
assign w24738 = w24053 & w25763;
assign w24739 = w24053 & w25764;
assign w24740 = ~w24053 & ~w25763;
assign w24741 = ~w24053 & ~w25764;
assign w24742 = ~w1150 & w1375;
assign w24743 = w1150 & ~w1375;
assign w24744 = ~w18359 & ~w18613;
assign w24745 = ~w18858 & ~w18857;
assign w24746 = ~w21005 & w21191;
assign w24747 = ~w22445 & ~w22443;
assign w24748 = ~w23497 & ~w23495;
assign w24749 = ~w1513 & w1806;
assign w24750 = w1513 & ~w1806;
assign w24751 = ~w1951 & w2260;
assign w24752 = w1951 & ~w2260;
assign w24753 = ~w2432 & w2783;
assign w24754 = w2432 & ~w2966;
assign w24755 = w12187 & w12177;
assign w24756 = (a[20] & ~w1667) | (a[20] & w24911) | (~w1667 & w24911);
assign w24757 = w1667 & w24912;
assign w24758 = ~w1520 & w1671;
assign w24759 = ~w1689 & ~w1687;
assign w24760 = ~w1723 & ~w1721;
assign w24761 = ~w1846 & ~w1844;
assign w24762 = ~w1869 & ~w1868;
assign w24763 = ~w1958 & w2109;
assign w24764 = ~w2129 & ~w2133;
assign w24765 = ~w2041 & ~w2040;
assign w24766 = ~w2137 & ~w2135;
assign w24767 = ~w2207 & ~w2206;
assign w24768 = ~w2389 & ~w2388;
assign w24769 = ~w2439 & w2617;
assign w24770 = ~w2637 & ~w2641;
assign w24771 = ~w2662 & ~w2661;
assign w24772 = w46 & w24913;
assign w24773 = ~w2645 & ~w2643;
assign w24774 = ~w24631 & ~w2968;
assign w24775 = ~w2787 & ~w2965;
assign w24776 = ~w2981 & w3170;
assign w24777 = ~w3189 & ~w3193;
assign w24778 = w2954 & ~w3009;
assign w24779 = w3171 & w3364;
assign w24780 = ~w3171 & ~w3364;
assign w24781 = ~w3197 & ~w3195;
assign w24782 = ~w3231 & ~w3230;
assign w24783 = w3237 & w3433;
assign w24784 = ~w3237 & ~w3433;
assign w24785 = ~w3300 & ~w3299;
assign w24786 = ~w2977 & b[2];
assign w24787 = ~w3400 & ~w3399;
assign w24788 = ~w3439 & ~w3437;
assign w24789 = ~w3658 & ~w3656;
assign w24790 = ~b[0] & a[35];
assign w24791 = ~w3881 & ~w3880;
assign w24792 = w3577 & b[1];
assign w24793 = w46 & w25093;
assign w24794 = (~a[35] & ~w46) | (~a[35] & w25094) | (~w46 & w25094);
assign w24795 = ~w3795 & ~w3793;
assign w24796 = ~w4110 & ~w4109;
assign w24797 = ~w3986 & ~w3991;
assign w24798 = w3577 & b[2];
assign w24799 = ~w4026 & ~w4024;
assign w24800 = ~w4344 & ~w4342;
assign w24801 = w4221 & ~w4251;
assign w24802 = (a[35] & ~w4442) | (a[35] & w25095) | (~w4442 & w25095);
assign w24803 = w4442 & w25096;
assign w24804 = ~w4244 & w4446;
assign w24805 = ~w4593 & ~w4591;
assign w24806 = w4240 & b[2];
assign w24807 = w4675 & ~w4672;
assign w24808 = ~w4922 & b[1];
assign w24809 = w46 & w25097;
assign w24810 = (~a[41] & ~w46) | (~a[41] & w25098) | (~w46 & w25098);
assign w24811 = ~w5177 & ~w5175;
assign w24812 = w6168 & a[44];
assign w24813 = ~w6168 & ~a[44];
assign w24814 = ~w5949 & ~w5948;
assign w24815 = ~w5972 & ~w5971;
assign w24816 = w5977 & ~w6232;
assign w24817 = ~w5977 & w6232;
assign w24818 = ~w6065 & ~w6064;
assign w24819 = ~w6261 & ~w6259;
assign w24820 = ~w6238 & ~w6236;
assign w24821 = ~w6163 & ~w6174;
assign w24822 = ~w6209 & ~w6208;
assign w24823 = ~w6255 & ~w6254;
assign w24824 = ~w6558 & ~w6557;
assign w24825 = ~w6840 & ~w6839;
assign w24826 = w6473 & b[1];
assign w24827 = w46 & w25249;
assign w24828 = (~a[47] & ~w46) | (~a[47] & w25250) | (~w46 & w25250);
assign w24829 = ~w7128 & ~w7127;
assign w24830 = ~w7431 & ~w7429;
assign w24831 = ~w7739 & ~w7737;
assign w24832 = ~w8045 & ~w8044;
assign w24833 = ~w8382 & ~w8380;
assign w24834 = ~w8283 & ~w8282;
assign w24835 = ~w8261 & ~w8259;
assign w24836 = ~w8255 & ~w8253;
assign w24837 = ~w8235 & ~w8233;
assign w24838 = ~w8228 & ~w8227;
assign w24839 = ~w8242 & ~w8240;
assign w24840 = ~w8367 & ~w8365;
assign w24841 = ~w8622 & ~w8620;
assign w24842 = ~w8599 & ~w8598;
assign w24843 = ~w8571 & ~w8569;
assign w24844 = ~w8934 & ~w8932;
assign w24845 = ~w9281 & ~w9280;
assign w24846 = ~w9625 & ~w9624;
assign w24847 = ~w9966 & ~w9965;
assign w24848 = ~w10320 & ~w10319;
assign w24849 = (~w11776 & ~w11778) | (~w11776 & w24914) | (~w11778 & w24914);
assign w24850 = ~w11619 & ~w11617;
assign w24851 = ~w11760 & ~w11759;
assign w24852 = ~w11760 & ~b[62];
assign w24853 = ~w11989 & ~w11987;
assign w24854 = ~w12066 & ~w12065;
assign w24855 = ~w12429 & ~w12428;
assign w24856 = ~w12408 & ~w12406;
assign w24857 = ~w12467 & ~w12466;
assign w24858 = ~w12853 & w25765;
assign w24859 = ~w12496 & w25541;
assign w24860 = (w12496 & w25542) | (w12496 & w25543) | (w25542 & w25543);
assign w24861 = w12853 & ~w12498;
assign w24862 = ~w12522 & ~w12842;
assign w24863 = w12809 & w12892;
assign w24864 = ~w12809 & ~w12892;
assign w24865 = ~w12702 & ~w12700;
assign w24866 = ~w12838 & ~w12837;
assign w24867 = ~w13064 & ~w13052;
assign w24868 = a[23] & ~w17535;
assign w24869 = a[23] & ~w24717;
assign w24870 = ~a[23] & w17535;
assign w24871 = ~a[23] & w24717;
assign w24872 = a[20] & ~w17550;
assign w24873 = a[20] & ~w24718;
assign w24874 = a[23] & ~w18077;
assign w24875 = a[23] & ~w24719;
assign w24876 = ~a[23] & w18077;
assign w24877 = ~a[23] & w24719;
assign w24878 = a[23] & ~w18345;
assign w24879 = a[23] & ~w24721;
assign w24880 = ~a[23] & w18345;
assign w24881 = ~a[23] & w24721;
assign w24882 = a[32] & ~w20410;
assign w24883 = a[32] & ~w24722;
assign w24884 = ~a[32] & w20410;
assign w24885 = ~a[32] & w24722;
assign w24886 = a[53] & ~w23165;
assign w24887 = a[53] & ~w24727;
assign w24888 = ~a[53] & w23165;
assign w24889 = ~a[53] & w24727;
assign w24890 = a[53] & ~w23257;
assign w24891 = a[53] & ~w24729;
assign w24892 = ~a[53] & w23257;
assign w24893 = ~a[53] & w24729;
assign w24894 = ~w8195 & w23343;
assign w24895 = ~w23950 & ~w24573;
assign w24896 = ~w23950 & ~w24572;
assign w24897 = (~w23983 & w24575) | (~w23983 & w24573) | (w24575 & w24573);
assign w24898 = (~w23983 & w24575) | (~w23983 & w24572) | (w24575 & w24572);
assign w24899 = (w24733 & w24732) | (w24733 & ~w24573) | (w24732 & ~w24573);
assign w24900 = (w24733 & w24732) | (w24733 & ~w24572) | (w24732 & ~w24572);
assign w24901 = (w24735 & w24734) | (w24735 & ~w24573) | (w24734 & ~w24573);
assign w24902 = (w24735 & w24734) | (w24735 & ~w24572) | (w24734 & ~w24572);
assign w24903 = (w24737 & w24736) | (w24737 & w24573) | (w24736 & w24573);
assign w24904 = (w24737 & w24736) | (w24737 & w24572) | (w24736 & w24572);
assign w24905 = (w24739 & w24738) | (w24739 & ~w24573) | (w24738 & ~w24573);
assign w24906 = (w24739 & w24738) | (w24739 & ~w24572) | (w24738 & ~w24572);
assign w24907 = (w24741 & w24740) | (w24741 & w24573) | (w24740 & w24573);
assign w24908 = (w24741 & w24740) | (w24741 & w24572) | (w24740 & w24572);
assign w24909 = ~w23495 & w23569;
assign w24910 = ~w23569 & ~w23568;
assign w24911 = w1665 & a[20];
assign w24912 = ~w1665 & ~a[20];
assign w24913 = w2432 & ~w2783;
assign w24914 = w11412 & ~w11776;
assign w24915 = ~b[0] & a[23];
assign w24916 = ~w1829 & ~w1827;
assign w24917 = w1932 & ~w1982;
assign w24918 = ~w2017 & ~w2015;
assign w24919 = ~w2171 & ~w2170;
assign w24920 = ~w2184 & ~w2183;
assign w24921 = ~w2334 & ~w2333;
assign w24922 = ~w2358 & ~w2356;
assign w24923 = ~b[0] & a[29];
assign w24924 = w2635 & a[26];
assign w24925 = ~w2522 & ~w2521;
assign w24926 = ~w2546 & ~w2545;
assign w24927 = ~w2776 & a[26];
assign w24928 = w2776 & ~a[26];
assign w24929 = ~w2715 & ~w2714;
assign w24930 = ~w2745 & ~w2743;
assign w24931 = b[0] & w2966;
assign w24932 = b[0] & ~w24634;
assign w24933 = ~w2815 & ~w2813;
assign w24934 = ~w2848 & ~w2847;
assign w24935 = ~w2895 & ~w2894;
assign w24936 = ~b[0] & a[32];
assign w24937 = w3187 & a[29];
assign w24938 = ~w3068 & ~w3067;
assign w24939 = ~w3123 & ~w3122;
assign w24940 = ~w2977 & b[1];
assign w24941 = w46 & w25099;
assign w24942 = (~a[32] & ~w46) | (~a[32] & w25100) | (~w46 & w25100);
assign w24943 = ~w3269 & ~w3267;
assign w24944 = ~w3360 & ~w3365;
assign w24945 = ~w3479 & ~w3478;
assign w24946 = (a[32] & ~w3774) | (a[32] & w25251) | (~w3774 & w25251);
assign w24947 = w3774 & w25252;
assign w24948 = w3558 & ~w3588;
assign w24949 = ~w3698 & ~w3696;
assign w24950 = ~w3812 & ~w3810;
assign w24951 = ~w3929 & ~w3927;
assign w24952 = ~w4042 & ~w4041;
assign w24953 = ~w4059 & ~w4058;
assign w24954 = w4063 & w4304;
assign w24955 = ~w4126 & ~w4125;
assign w24956 = ~w4309 & ~w4308;
assign w24957 = w3577 & b[3];
assign w24958 = ~b[0] & a[38];
assign w24959 = ~w4281 & ~w4279;
assign w24960 = ~w4550 & ~w4549;
assign w24961 = ~w4776 & ~w4774;
assign w24962 = ~w5029 & ~w5028;
assign w24963 = ~w4980 & ~w4978;
assign w24964 = ~w4958 & ~w4956;
assign w24965 = (a[38] & ~w5156) | (a[38] & w25253) | (~w5156 & w25253);
assign w24966 = w5156 & w25254;
assign w24967 = ~w4926 & w5160;
assign w24968 = ~w4933 & ~w5177;
assign w24969 = w4933 & w5177;
assign w24970 = ~w5289 & ~w5287;
assign w24971 = ~w5216 & ~w5214;
assign w24972 = ~w5193 & ~w5192;
assign w24973 = ~w5398 & ~w5408;
assign w24974 = ~w5559 & ~w5557;
assign w24975 = ~w5671 & w5932;
assign w24976 = ~w5696 & ~w5695;
assign w24977 = w5669 & b[1];
assign w24978 = w5669 & b[2];
assign w24979 = ~w6477 & w6725;
assign w24980 = ~w6742 & ~w6740;
assign w24981 = ~w6996 & ~w7006;
assign w24982 = w7873 & a[50];
assign w24983 = ~w7873 & ~a[50];
assign w24984 = ~w7596 & ~w7594;
assign w24985 = ~w7611 & w7914;
assign w24986 = ~w7629 & ~w7627;
assign w24987 = ~w7755 & ~w7754;
assign w24988 = ~w7987 & ~w7985;
assign w24989 = ~w7958 & ~w7956;
assign w24990 = ~w7942 & ~w7940;
assign w24991 = ~w7868 & ~w7879;
assign w24992 = ~w7936 & ~w7935;
assign w24993 = ~w7981 & ~w7980;
assign w24994 = ~w8296 & ~w8294;
assign w24995 = ~w8277 & ~w8276;
assign w24996 = ~w8644 & ~w8643;
assign w24997 = w8199 & b[1];
assign w24998 = w8836 & a[53];
assign w24999 = ~w8836 & ~a[53];
assign w25000 = ~w8616 & ~w8614;
assign w25001 = ~w8957 & ~w8956;
assign w25002 = ~w8928 & ~w8926;
assign w25003 = ~w9304 & ~w9302;
assign w25004 = ~w9275 & ~w9274;
assign w25005 = ~w9638 & ~w9637;
assign w25006 = ~w9619 & ~w9618;
assign w25007 = ~w9979 & ~w9978;
assign w25008 = ~w9960 & ~w9959;
assign w25009 = ~w10314 & ~w10312;
assign w25010 = w12863 & ~w12507;
assign w25011 = w12863 & w24401;
assign w25012 = ~w12658 & ~w12656;
assign w25013 = ~w12735 & w13077;
assign w25014 = w12735 & ~w13077;
assign w25015 = ~w13047 & ~w13035;
assign w25016 = ~w13023 & ~w13011;
assign w25017 = ~w12915 & ~w13004;
assign w25018 = ~w12905 & ~w13028;
assign w25019 = ~w13414 & ~w13426;
assign w25020 = ~w832 & w16711;
assign w25021 = ~w1951 & w17520;
assign w25022 = ~w1513 & w17817;
assign w25023 = ~w17530 & ~w17540;
assign w25024 = ~w17545 & ~w17555;
assign w25025 = ~w18092 & a[20];
assign w25026 = w18092 & ~a[20];
assign w25027 = ~w18072 & ~w18082;
assign w25028 = ~w1951 & w18125;
assign w25029 = ~w18340 & ~w18350;
assign w25030 = ~w3573 & w20603;
assign w25031 = ~w20405 & ~w20415;
assign w25032 = ~w3573 & w20641;
assign w25033 = w20807 & ~a[32];
assign w25034 = ~w20807 & a[32];
assign w25035 = ~w3573 & w20829;
assign w25036 = ~w4923 & w21724;
assign w25037 = ~w5663 & w22143;
assign w25038 = ~w4923 & w22158;
assign w25039 = ~w5663 & w22182;
assign w25040 = w22297 & ~a[41];
assign w25041 = ~w22297 & a[41];
assign w25042 = ~w7312 & w23061;
assign w25043 = ~w8195 & w23126;
assign w25044 = ~w9158 & w23174;
assign w25045 = a[50] & ~w23234;
assign w25046 = a[50] & ~w24728;
assign w25047 = w23160 & ~w23225;
assign w25048 = ~w9158 & w23266;
assign w25049 = ~w23324 & a[50];
assign w25050 = w23324 & ~a[50];
assign w25051 = a[53] & ~w23343;
assign w25052 = a[53] & ~w24894;
assign w25053 = ~w9158 & w23389;
assign w25054 = ~w23314 & ~w23313;
assign w25055 = ~w7586 & w25766;
assign w25056 = ~w7586 & w25767;
assign w25057 = ~w23327 & ~w23319;
assign w25058 = (~w23333 & w24539) | (~w23333 & w24538) | (w24539 & w24538);
assign w25059 = (~w23333 & w24539) | (~w23333 & w24537) | (w24539 & w24537);
assign w25060 = ~w9158 & w23427;
assign w25061 = ~w8195 & w23482;
assign w25062 = (w24542 & w24543) | (w24542 & w24538) | (w24543 & w24538);
assign w25063 = (w24542 & w24543) | (w24542 & w24537) | (w24543 & w24537);
assign w25064 = ~w9158 & w23506;
assign w25065 = (w24546 & w24545) | (w24546 & ~w24538) | (w24545 & ~w24538);
assign w25066 = (w24546 & w24545) | (w24546 & ~w24537) | (w24545 & ~w24537);
assign w25067 = (w24550 & w24549) | (w24550 & w24538) | (w24549 & w24538);
assign w25068 = (w24550 & w24549) | (w24550 & w24537) | (w24549 & w24537);
assign w25069 = (w24553 & w25758) | (w24553 & w24538) | (w25758 & w24538);
assign w25070 = (w24553 & w25758) | (w24553 & w24537) | (w25758 & w24537);
assign w25071 = (w24555 & w24554) | (w24555 & ~w24538) | (w24554 & ~w24538);
assign w25072 = (w24555 & w24554) | (w24555 & ~w24537) | (w24554 & ~w24537);
assign w25073 = (w24559 & w24558) | (w24559 & w24538) | (w24558 & w24538);
assign w25074 = (w24559 & w24558) | (w24559 & w24537) | (w24558 & w24537);
assign w25075 = (w24563 & w24562) | (w24563 & w24538) | (w24562 & w24538);
assign w25076 = (w24563 & w24562) | (w24563 & w24537) | (w24562 & w24537);
assign w25077 = (w24567 & w24566) | (w24567 & w24538) | (w24566 & w24538);
assign w25078 = (w24567 & w24566) | (w24567 & w24537) | (w24566 & w24537);
assign w25079 = (w24571 & w24570) | (w24571 & w24538) | (w24570 & w24538);
assign w25080 = (w24571 & w24570) | (w24571 & w24537) | (w24570 & w24537);
assign w25081 = ~w23985 & w24896;
assign w25082 = ~w23985 & w24895;
assign w25083 = w23985 & ~w24896;
assign w25084 = w23985 & ~w24895;
assign w25085 = w24010 & w24898;
assign w25086 = w24010 & w24897;
assign w25087 = ~w24010 & ~w24898;
assign w25088 = ~w24010 & ~w24897;
assign w25089 = (w24577 & w24578) | (w24577 & w24898) | (w24578 & w24898);
assign w25090 = (w24577 & w24578) | (w24577 & w24897) | (w24578 & w24897);
assign w25091 = w4236 & a[38];
assign w25092 = ~w4236 & ~a[38];
assign w25093 = w3573 & a[35];
assign w25094 = ~w3573 & ~a[35];
assign w25095 = w4438 & a[35];
assign w25096 = ~w4438 & ~a[35];
assign w25097 = w4923 & a[41];
assign w25098 = ~w4923 & ~a[41];
assign w25099 = w2980 & a[32];
assign w25100 = ~w2980 & ~a[32];
assign w25101 = ~w1823 & a[20];
assign w25102 = w1823 & ~a[20];
assign w25103 = ~w2301 & ~w2300;
assign w25104 = ~w2479 & ~w2484;
assign w25105 = ~w2680 & w2616;
assign w25106 = w2680 & ~w2616;
assign w25107 = ~w2831 & ~w2830;
assign w25108 = ~w3051 & ~w3049;
assign w25109 = ~w3262 & ~w3260;
assign w25110 = ~w3462 & ~w3461;
assign w25111 = ~w2977 & b[3];
assign w25112 = ~w3638 & ~w3637;
assign w25113 = ~w3651 & ~w3650;
assign w25114 = ~w3681 & ~w3679;
assign w25115 = ~w3905 & ~w3903;
assign w25116 = ~w3875 & ~w3874;
assign w25117 = ~w4140 & ~w4138;
assign w25118 = ~w4104 & ~w4103;
assign w25119 = ~w4287 & ~w4285;
assign w25120 = ~w4338 & ~w4336;
assign w25121 = ~w4544 & ~w4542;
assign w25122 = ~w4570 & ~w4568;
assign w25123 = ~w4760 & ~w4758;
assign w25124 = ~w4823 & ~w4822;
assign w25125 = w4240 & b[3];
assign w25126 = ~b[0] & a[41];
assign w25127 = ~w5023 & ~w5021;
assign w25128 = ~w5283 & ~w5282;
assign w25129 = ~w5472 & ~w5471;
assign w25130 = ~w5459 & ~w5458;
assign w25131 = ~w4922 & b[2];
assign w25132 = ~w5536 & ~w5534;
assign w25133 = ~w5716 & ~w5714;
assign w25134 = (a[41] & ~w5928) | (a[41] & w25544) | (~w5928 & w25544);
assign w25135 = w5928 & w25545;
assign w25136 = ~w5678 & w5949;
assign w25137 = w5678 & ~w5949;
assign w25138 = ~w5822 & ~w5821;
assign w25139 = ~w5965 & ~w5964;
assign w25140 = ~w6225 & ~w6224;
assign w25141 = w5980 & ~w6231;
assign w25142 = ~w6539 & ~w6538;
assign w25143 = ~w7041 & ~w7039;
assign w25144 = ~w7064 & ~w7063;
assign w25145 = ~w7353 & ~w7351;
assign w25146 = (a[47] & ~w7575) | (a[47] & w25546) | (~w7575 & w25546);
assign w25147 = w7575 & w25547;
assign w25148 = ~w7315 & w7579;
assign w25149 = ~w7340 & ~w7339;
assign w25150 = ~w7376 & ~w7375;
assign w25151 = ~w7400 & ~w7399;
assign w25152 = ~w7464 & ~w7462;
assign w25153 = ~w7687 & ~w7685;
assign w25154 = ~w7641 & ~w7639;
assign w25155 = ~w7311 & b[1];
assign w25156 = ~w7674 & ~w7672;
assign w25157 = ~w7311 & b[2];
assign w25158 = w7614 & ~w7912;
assign w25159 = ~w8003 & ~w8001;
assign w25160 = ~w8203 & w8508;
assign w25161 = ~w8313 & ~w8312;
assign w25162 = ~w8651 & ~w8649;
assign w25163 = ~w8593 & ~w8591;
assign w25164 = ~w8525 & ~w8524;
assign w25165 = ~w8548 & ~w8546;
assign w25166 = ~w8831 & ~w8842;
assign w25167 = ~w8867 & ~w8865;
assign w25168 = ~w8915 & ~w8914;
assign w25169 = ~w8963 & ~w8961;
assign w25170 = ~w9253 & ~w9251;
assign w25171 = ~w9311 & ~w9309;
assign w25172 = ~w9596 & ~w9594;
assign w25173 = ~w9645 & ~w9643;
assign w25174 = ~w9946 & ~w9945;
assign w25175 = ~w10003 & ~w10001;
assign w25176 = ~w10302 & ~w10300;
assign w25177 = ~w10674 & ~w10673;
assign w25178 = ~w11013 & ~w11011;
assign w25179 = ~w10937 & ~w10935;
assign w25180 = ~w10911 & ~w10910;
assign w25181 = ~w10899 & ~w10898;
assign w25182 = ~w10876 & ~w10874;
assign w25183 = ~w10883 & ~w10881;
assign w25184 = ~w10931 & ~w10929;
assign w25185 = ~w11032 & ~w11031;
assign w25186 = ~w11282 & ~w11280;
assign w25187 = ~w11260 & ~w11258;
assign w25188 = ~w11308 & ~w11306;
assign w25189 = ~w11702 & ~w11700;
assign w25190 = ~w11642 & ~w11640;
assign w25191 = ~w11675 & ~w11674;
assign w25192 = ~w12072 & ~w12071;
assign w25193 = ~w12011 & ~w12009;
assign w25194 = ~w12025 & ~w12024;
assign w25195 = ~w12473 & ~w12471;
assign w25196 = ~w12422 & ~w12420;
assign w25197 = ~w12736 & w25013;
assign w25198 = w25014 & ~w13077;
assign w25199 = (~w13077 & w25014) | (~w13077 & w12736) | (w25014 & w12736);
assign w25200 = ~w12794 & ~w12792;
assign w25201 = w13197 & ~w12837;
assign w25202 = w13197 & w24866;
assign w25203 = ~w13197 & w12837;
assign w25204 = ~w13197 & ~w24866;
assign w25205 = ~w13203 & ~w12880;
assign w25206 = ~w13184 & ~w12893;
assign w25207 = ~w13200 & ~w13198;
assign w25208 = ~w832 & w15561;
assign w25209 = a[23] & ~w17817;
assign w25210 = a[23] & ~w25022;
assign w25211 = ~w17812 & ~w17822;
assign w25212 = a[26] & ~w18125;
assign w25213 = a[26] & ~w25028;
assign w25214 = ~a[26] & w18125;
assign w25215 = ~a[26] & w25028;
assign w25216 = a[35] & ~w20603;
assign w25217 = a[35] & ~w25030;
assign w25218 = ~a[35] & w20603;
assign w25219 = ~a[35] & w25030;
assign w25220 = ~w4236 & w20978;
assign w25221 = a[44] & ~w22143;
assign w25222 = a[44] & ~w25037;
assign w25223 = ~a[44] & w22143;
assign w25224 = ~a[44] & w25037;
assign w25225 = ~a[56] & w23174;
assign w25226 = ~a[56] & w25044;
assign w25227 = ~w10141 & w23183;
assign w25228 = a[56] & ~w23266;
assign w25229 = a[56] & ~w25048;
assign w25230 = ~a[56] & w23266;
assign w25231 = ~a[56] & w25048;
assign w25232 = w23241 & ~w23238;
assign w25233 = a[56] & ~w23389;
assign w25234 = a[56] & ~w25053;
assign w25235 = ~a[56] & w23389;
assign w25236 = ~a[56] & w25053;
assign w25237 = a[56] & ~w23427;
assign w25238 = a[56] & ~w25060;
assign w25239 = ~a[56] & w23427;
assign w25240 = ~a[56] & w25060;
assign w25241 = ~w24032 & w24900;
assign w25242 = ~w24032 & w24899;
assign w25243 = ~w22308 & ~w22443;
assign w25244 = ~w24509 & ~w22575;
assign w25245 = ~w22575 & w22702;
assign w25246 = w23568 & w23639;
assign w25247 = w23639 & ~w24910;
assign w25248 = ~w13557 & ~w13556;
assign w25249 = w6469 & a[47];
assign w25250 = ~w6469 & ~a[47];
assign w25251 = w3770 & a[32];
assign w25252 = ~w3770 & ~a[32];
assign w25253 = w5152 & a[38];
assign w25254 = ~w5152 & ~a[38];
assign w25255 = ~w3851 & ~w3849;
assign w25256 = ~w4063 & ~w4067;
assign w25257 = w4305 & ~w4188;
assign w25258 = ~w4305 & w4188;
assign w25259 = ~w5228 & ~w5226;
assign w25260 = ~w5484 & ~w5483;
assign w25261 = ~w5761 & ~w5760;
assign w25262 = ~w6027 & ~w6026;
assign w25263 = ~w5991 & ~w5990;
assign w25264 = ~w6297 & ~w6295;
assign w25265 = ~w6594 & ~w6592;
assign w25266 = ~w6721 & a[44];
assign w25267 = w6721 & ~a[44];
assign w25268 = w6484 & w6742;
assign w25269 = ~w6484 & ~w6742;
assign w25270 = ~w6876 & ~w6875;
assign w25271 = ~w6821 & ~w6819;
assign w25272 = ~w6758 & ~w6757;
assign w25273 = ~w7181 & ~w7180;
assign w25274 = ~w7099 & ~w7097;
assign w25275 = ~w7057 & ~w7056;
assign w25276 = w6473 & b[2];
assign w25277 = w7322 & w7596;
assign w25278 = ~w7322 & ~w7596;
assign w25279 = ~w7412 & ~w7411;
assign w25280 = ~w7612 & ~w7611;
assign w25281 = ~w7916 & ~w7926;
assign w25282 = w7916 & w7926;
assign w25283 = ~w7710 & ~w7709;
assign w25284 = ~w8016 & ~w8014;
assign w25285 = ~w7929 & ~w7928;
assign w25286 = ~w8248 & ~w8246;
assign w25287 = ~w8335 & ~w8334;
assign w25288 = ~w8577 & ~w8575;
assign w25289 = ~w8664 & ~w8663;
assign w25290 = ~w8986 & ~w8984;
assign w25291 = ~w9341 & ~w9339;
assign w25292 = ~w9589 & ~w9587;
assign w25293 = ~w9929 & ~w9928;
assign w25294 = ~w10285 & ~w10283;
assign w25295 = ~w10668 & ~w10666;
assign w25296 = ~w10996 & ~w10994;
assign w25297 = ~w11368 & ~w11366;
assign w25298 = ~w11237 & ~w11235;
assign w25299 = ~w11221 & ~w11220;
assign w25300 = ~w11254 & ~w11253;
assign w25301 = ~w11384 & ~w11383;
assign w25302 = (~w11396 & w24697) | (~w11396 & ~w11031) | (w24697 & ~w11031);
assign w25303 = (~w11396 & w24697) | (~w11396 & w25185) | (w24697 & w25185);
assign w25304 = ~w11636 & ~w11635;
assign w25305 = ~w11995 & ~w11994;
assign w25306 = ~w12446 & ~w12444;
assign w25307 = ~w12415 & ~w12413;
assign w25308 = ~w12719 & ~w12717;
assign w25309 = ~w12758 & ~w12756;
assign w25310 = ~w12788 & ~w12787;
assign w25311 = ~w13178 & ~w12795;
assign w25312 = ~w13067 & ~w13078;
assign w25313 = a[17] & ~w15561;
assign w25314 = a[17] & ~w25208;
assign w25315 = ~a[17] & w15561;
assign w25316 = ~a[17] & w25208;
assign w25317 = ~w832 & w16161;
assign w25318 = ~w1513 & w17275;
assign w25319 = a[26] & ~w17520;
assign w25320 = a[26] & ~w25021;
assign w25321 = ~w1951 & w17855;
assign w25322 = ~w18087 & ~w18096;
assign w25323 = ~w1951 & w18584;
assign w25324 = ~w18337 & ~w18130;
assign w25325 = ~w3573 & w20399;
assign w25326 = ~w4236 & w20588;
assign w25327 = a[35] & ~w20641;
assign w25328 = a[35] & ~w25032;
assign w25329 = ~a[35] & w20641;
assign w25330 = ~a[35] & w25032;
assign w25331 = ~w4236 & w20789;
assign w25332 = w20610 & ~w20607;
assign w25333 = a[38] & ~w20978;
assign w25334 = a[38] & ~w25220;
assign w25335 = ~a[38] & w20978;
assign w25336 = ~a[38] & w25220;
assign w25337 = ~w5663 & w21666;
assign w25338 = a[41] & ~w21724;
assign w25339 = a[41] & ~w25036;
assign w25340 = ~w5663 & w21732;
assign w25341 = ~w5663 & w21999;
assign w25342 = ~w6469 & w22128;
assign w25343 = w22166 & ~w22163;
assign w25344 = a[44] & ~w22182;
assign w25345 = a[44] & ~w25039;
assign w25346 = ~a[44] & w22182;
assign w25347 = ~a[44] & w25039;
assign w25348 = ~w6469 & w22190;
assign w25349 = w22150 & ~w22147;
assign w25350 = ~w22172 & ~w24504;
assign w25351 = ~w22172 & ~w24503;
assign w25352 = ~w6469 & w22416;
assign w25353 = (~w22308 & w24506) | (~w22308 & w24504) | (w24506 & w24504);
assign w25354 = (~w22308 & w24506) | (~w22308 & w24503) | (w24506 & w24503);
assign w25355 = (w24509 & w24510) | (w24509 & w24504) | (w24510 & w24504);
assign w25356 = (w24509 & w24510) | (w24509 & w24503) | (w24510 & w24503);
assign w25357 = ~w6469 & w22546;
assign w25358 = (w24513 & w24514) | (w24513 & ~w24504) | (w24514 & ~w24504);
assign w25359 = (w24513 & w24514) | (w24513 & ~w24503) | (w24514 & ~w24503);
assign w25360 = (w24517 & w24518) | (w24517 & w24504) | (w24518 & w24504);
assign w25361 = (w24517 & w24518) | (w24517 & w24503) | (w24518 & w24503);
assign w25362 = (w24521 & w24522) | (w24521 & w24504) | (w24522 & w24504);
assign w25363 = (w24521 & w24522) | (w24521 & w24503) | (w24522 & w24503);
assign w25364 = ~w11189 & w22993;
assign w25365 = (w24525 & w24526) | (w24525 & ~w24504) | (w24526 & ~w24504);
assign w25366 = (w24525 & w24526) | (w24525 & ~w24503) | (w24526 & ~w24503);
assign w25367 = ~w9158 & w23071;
assign w25368 = a[53] & ~w23126;
assign w25369 = a[53] & ~w25043;
assign w25370 = (w24529 & w24530) | (w24529 & w24504) | (w24530 & w24504);
assign w25371 = (w24529 & w24530) | (w24529 & w24503) | (w24530 & w24503);
assign w25372 = ~a[59] & w23183;
assign w25373 = ~a[59] & w25227;
assign w25374 = ~w11189 & w23191;
assign w25375 = (w24533 & w24534) | (w24533 & w24504) | (w24534 & w24504);
assign w25376 = (w24533 & w24534) | (w24533 & w24503) | (w24534 & w24503);
assign w25377 = w23169 & ~w23219;
assign w25378 = ~w10141 & w23275;
assign w25379 = ~w11189 & w23292;
assign w25380 = ~w23334 & w24537;
assign w25381 = ~w23334 & w24538;
assign w25382 = w23334 & ~w24537;
assign w25383 = w23334 & ~w24538;
assign w25384 = ~w10141 & w23352;
assign w25385 = (w24540 & w24541) | (w24540 & ~w24537) | (w24541 & ~w24537);
assign w25386 = (w24540 & w24541) | (w24540 & ~w24538) | (w24541 & ~w24538);
assign w25387 = ~w10141 & w23436;
assign w25388 = w23497 & w25063;
assign w25389 = w23497 & w25062;
assign w25390 = w23422 & ~w23473;
assign w25391 = a[56] & ~w23506;
assign w25392 = a[56] & ~w25064;
assign w25393 = ~a[56] & w23506;
assign w25394 = ~a[56] & w25064;
assign w25395 = ~w10141 & w23515;
assign w25396 = w23490 & ~w23487;
assign w25397 = (w24547 & w24548) | (w24547 & ~w24537) | (w24548 & ~w24537);
assign w25398 = (w24547 & w24548) | (w24547 & ~w24538) | (w24548 & ~w24538);
assign w25399 = (w24552 & w24551) | (w24552 & ~w24537) | (w24551 & ~w24537);
assign w25400 = (w24552 & w24551) | (w24552 & ~w24538) | (w24551 & ~w24538);
assign w25401 = w23706 & w25768;
assign w25402 = w23706 & w25769;
assign w25403 = (w24557 & w24556) | (w24557 & ~w24537) | (w24556 & ~w24537);
assign w25404 = (w24557 & w24556) | (w24557 & ~w24538) | (w24556 & ~w24538);
assign w25405 = (w24561 & w24560) | (w24561 & ~w24537) | (w24560 & ~w24537);
assign w25406 = (w24561 & w24560) | (w24561 & ~w24538) | (w24560 & ~w24538);
assign w25407 = w23871 & ~w25076;
assign w25408 = w23871 & ~w25075;
assign w25409 = w23913 & ~w25078;
assign w25410 = w23913 & ~w25077;
assign w25411 = w23952 & ~w25080;
assign w25412 = w23952 & ~w25079;
assign w25413 = w18102 & ~w18359;
assign w25414 = ~w25245 & ~w22701;
assign w25415 = ~w23638 & ~w23639;
assign w25416 = ~w23638 & ~w25246;
assign w25417 = ~w23638 & ~w25247;
assign w25418 = ~w4922 & b[3];
assign w25419 = ~b[0] & a[44];
assign w25420 = ~w7093 & ~w7091;
assign w25421 = ~w7406 & ~w7404;
assign w25422 = ~w7369 & ~w7367;
assign w25423 = w6473 & b[3];
assign w25424 = ~b[0] & a[50];
assign w25425 = ~w7693 & ~w7692;
assign w25426 = ~w7657 & ~w7656;
assign w25427 = ~w8009 & ~w8007;
assign w25428 = ~w7964 & ~w7963;
assign w25429 = ~w8319 & ~w8318;
assign w25430 = ~w8657 & ~w8655;
assign w25431 = ~w8969 & ~w8967;
assign w25432 = ~w9317 & ~w9315;
assign w25433 = ~w9668 & ~w9666;
assign w25434 = ~w9561 & ~w9559;
assign w25435 = ~w9890 & ~w9888;
assign w25436 = ~w10266 & ~w10265;
assign w25437 = (~w13902 & w24405) | (~w13902 & w24706) | (w24405 & w24706);
assign w25438 = (~w13902 & w24405) | (~w13902 & w24707) | (w24405 & w24707);
assign w25439 = ~w14190 & ~w14202;
assign w25440 = ~w14139 & ~w14151;
assign w25441 = ~w14088 & ~w14100;
assign w25442 = ~w14105 & ~w14117;
assign w25443 = ~w14122 & ~w14134;
assign w25444 = ~w14156 & ~w14168;
assign w25445 = ~w14173 & ~w14185;
assign w25446 = ~w14207 & ~w14219;
assign w25447 = ~w1150 & w15573;
assign w25448 = ~w569 & w15831;
assign w25449 = ~w15822 & ~w15566;
assign w25450 = ~w832 & w16123;
assign w25451 = a[17] & ~w16161;
assign w25452 = a[17] & ~w25317;
assign w25453 = ~a[17] & w16161;
assign w25454 = ~a[17] & w25317;
assign w25455 = ~w1150 & w16415;
assign w25456 = ~w1951 & w16662;
assign w25457 = ~w1150 & w16695;
assign w25458 = a[17] & ~w16711;
assign w25459 = a[17] & ~w25020;
assign w25460 = ~a[17] & w16711;
assign w25461 = ~a[17] & w25020;
assign w25462 = ~a[23] & w17275;
assign w25463 = ~a[23] & w25318;
assign w25464 = ~w2432 & w17504;
assign w25465 = ~w1150 & w17833;
assign w25466 = ~w17827 & ~w17838;
assign w25467 = ~a[26] & w17855;
assign w25468 = ~a[26] & w25321;
assign w25469 = a[26] & ~w18584;
assign w25470 = a[26] & ~w25323;
assign w25471 = ~w1513 & w18600;
assign w25472 = ~w18355 & ~w18118;
assign w25473 = ~w1951 & w18624;
assign w25474 = ~w18579 & ~w18589;
assign w25475 = ~w12155 & w1513;
assign w25476 = a[35] & ~w20399;
assign w25477 = a[35] & ~w25325;
assign w25478 = ~w4923 & w20448;
assign w25479 = ~a[38] & w20588;
assign w25480 = ~a[38] & w25326;
assign w25481 = ~w2980 & w20619;
assign w25482 = ~w20613 & ~w20624;
assign w25483 = a[38] & ~w20789;
assign w25484 = a[38] & ~w25331;
assign w25485 = ~a[38] & w20789;
assign w25486 = ~a[38] & w25331;
assign w25487 = ~w20802 & ~w20811;
assign w25488 = a[35] & ~w20829;
assign w25489 = a[35] & ~w25035;
assign w25490 = ~a[35] & w20829;
assign w25491 = ~a[35] & w25035;
assign w25492 = ~w4923 & w20838;
assign w25493 = ~w20799 & ~w20797;
assign w25494 = w2980 & b[62];
assign w25495 = w2980 & ~w24852;
assign w25496 = ~w4236 & w21163;
assign w25497 = ~w20832 & ~w20986;
assign w25498 = ~w3573 & w21179;
assign w25499 = ~w4923 & w21883;
assign w25500 = a[44] & ~w21999;
assign w25501 = a[44] & ~w25341;
assign w25502 = ~w7312 & w22039;
assign w25503 = ~a[47] & w22128;
assign w25504 = ~a[47] & w25342;
assign w25505 = a[47] & ~w22190;
assign w25506 = a[47] & ~w25348;
assign w25507 = ~a[47] & w22190;
assign w25508 = ~a[47] & w25348;
assign w25509 = ~w22292 & ~w22301;
assign w25510 = ~w5663 & w22318;
assign w25511 = a[47] & ~w22416;
assign w25512 = a[47] & ~w25352;
assign w25513 = ~a[47] & w22416;
assign w25514 = ~a[47] & w25352;
assign w25515 = ~w22289 & ~w22287;
assign w25516 = w4923 & b[62];
assign w25517 = w4923 & ~w24852;
assign w25518 = a[47] & ~w22546;
assign w25519 = a[47] & ~w25357;
assign w25520 = ~a[47] & w22546;
assign w25521 = ~a[47] & w25357;
assign w25522 = ~w12155 & w5663;
assign w25523 = ~w11189 & w23362;
assign w25524 = a[59] & ~w23436;
assign w25525 = a[59] & ~w25387;
assign w25526 = ~a[59] & w23436;
assign w25527 = ~a[59] & w25387;
assign w25528 = a[59] & ~w23515;
assign w25529 = a[59] & ~w25395;
assign w25530 = ~a[59] & w23515;
assign w25531 = ~a[59] & w25395;
assign w25532 = ~w12155 & w8195;
assign w25533 = ~w10141 & w23578;
assign w25534 = ~w19102 & ~w19100;
assign w25535 = (~w22443 & w24747) | (~w22443 & ~w22308) | (w24747 & ~w22308);
assign w25536 = (~w22443 & w24747) | (~w22443 & ~w22309) | (w24747 & ~w22309);
assign w25537 = w22702 & ~w22576;
assign w25538 = w23706 & w25415;
assign w25539 = w23706 & w25416;
assign w25540 = ~w23706 & ~w23705;
assign w25541 = ~w12187 & ~w12853;
assign w25542 = w12853 & w12177;
assign w25543 = w12853 & w24755;
assign w25544 = w5924 & a[41];
assign w25545 = ~w5924 & ~a[41];
assign w25546 = w7571 & a[47];
assign w25547 = ~w7571 & ~a[47];
assign w25548 = ~w9204 & ~w9202;
assign w25549 = ~w9538 & ~w9536;
assign w25550 = ~w9877 & ~w9876;
assign w25551 = ~w10254 & ~w10252;
assign w25552 = ~w10617 & ~w10616;
assign w25553 = ~w10954 & ~w10952;
assign w25554 = ~w11325 & ~w11323;
assign w25555 = ~w11708 & ~w11706;
assign w25556 = ~w12079 & ~w12078;
assign w25557 = ~w12479 & ~w12478;
assign w25558 = ~w12847 & ~w12855;
assign w25559 = ~w12811 & w24864;
assign w25560 = (w24413 & w24412) | (w24413 & w24407) | (w24412 & w24407);
assign w25561 = (w24413 & w24412) | (w24413 & w24408) | (w24412 & w24408);
assign w25562 = ~w15523 & ~w15533;
assign w25563 = ~w15520 & ~w15243;
assign w25564 = a[20] & ~w15573;
assign w25565 = a[20] & ~w25447;
assign w25566 = ~w15483 & ~w15257;
assign w25567 = ~w15480 & ~w15271;
assign w25568 = ~w1513 & w15809;
assign w25569 = ~w15503 & ~w15515;
assign w25570 = a[14] & ~w15831;
assign w25571 = a[14] & ~w25448;
assign w25572 = ~a[14] & w15831;
assign w25573 = ~a[14] & w25448;
assign w25574 = a[17] & ~w16123;
assign w25575 = a[17] & ~w25450;
assign w25576 = ~a[20] & w16415;
assign w25577 = ~a[20] & w25455;
assign w25578 = ~w16117 & ~w16127;
assign w25579 = ~w12155 & w569;
assign w25580 = a[20] & ~w16695;
assign w25581 = a[20] & ~w25457;
assign w25582 = ~a[20] & w16695;
assign w25583 = ~a[20] & w25457;
assign w25584 = ~w16424 & ~w16166;
assign w25585 = ~w16705 & ~w16715;
assign w25586 = ~w2432 & w18137;
assign w25587 = ~w18594 & ~w18605;
assign w25588 = a[26] & ~w18624;
assign w25589 = a[26] & ~w25473;
assign w25590 = ~a[26] & w18624;
assign w25591 = ~a[26] & w25473;
assign w25592 = ~w18846 & a[23];
assign w25593 = w18846 & ~a[23];
assign w25594 = ~w4236 & w20242;
assign w25595 = ~a[41] & w20448;
assign w25596 = ~a[41] & w25478;
assign w25597 = ~w6469 & w20551;
assign w25598 = ~w5663 & w20567;
assign w25599 = ~w4923 & w20650;
assign w25600 = ~w5663 & w20659;
assign w25601 = ~w6469 & w20668;
assign w25602 = w20595 & ~w20592;
assign w25603 = a[38] & ~w21163;
assign w25604 = a[38] & ~w25496;
assign w25605 = a[35] & ~w21179;
assign w25606 = a[35] & ~w25498;
assign w25607 = ~w6469 & w21893;
assign w25608 = ~a[50] & w22039;
assign w25609 = ~a[50] & w25502;
assign w25610 = ~w9158 & w22049;
assign w25611 = ~w8195 & w22107;
assign w25612 = ~w7312 & w22199;
assign w25613 = ~w8195 & w22208;
assign w25614 = ~w9158 & w22217;
assign w25615 = w22135 & ~w22132;
assign w25616 = a[44] & ~w22318;
assign w25617 = a[44] & ~w25510;
assign w25618 = ~w7312 & w22327;
assign w25619 = ~w7312 & w22454;
assign w25620 = ~w5663 & w22561;
assign w25621 = w22553 & ~w22550;
assign w25622 = w22689 & ~a[44];
assign w25623 = ~w22689 & a[44];
assign w25624 = w22569 & ~w22566;
assign w25625 = a[59] & ~w23578;
assign w25626 = a[59] & ~w25533;
assign w25627 = ~a[59] & w23578;
assign w25628 = ~a[59] & w25533;
assign w25629 = ~w9158 & w23615;
assign w25630 = ~w23548 & ~w23547;
assign w25631 = w8195 & b[62];
assign w25632 = w8195 & ~w24852;
assign w25633 = ~w23562 & ~w23553;
assign w25634 = ~w15227 & ~w15226;
assign w25635 = ~w19341 & ~w19340;
assign w25636 = ~w21191 & ~w21190;
assign w25637 = ~w21369 & ~w21367;
assign w25638 = w22701 & w22826;
assign w25639 = w22826 & ~w25414;
assign w25640 = ~w23705 & ~w25539;
assign w25641 = ~w23705 & ~w25538;
assign w25642 = w23765 & ~w23705;
assign w25643 = w23765 & w25540;
assign w25644 = (w24538 & w24537) | (w24538 & w24504) | (w24537 & w24504);
assign w25645 = (w24538 & w24537) | (w24538 & w24503) | (w24537 & w24503);
assign w25646 = ~w23418 & w25059;
assign w25647 = ~w23418 & w25058;
assign w25648 = ~w23497 & ~w25063;
assign w25649 = ~w23497 & ~w25062;
assign w25650 = ~w23569 & ~w25066;
assign w25651 = ~w23569 & ~w25065;
assign w25652 = ~w23639 & w25068;
assign w25653 = ~w23639 & w25067;
assign w25654 = ~w23706 & ~w25070;
assign w25655 = ~w23706 & ~w25069;
assign w25656 = ~w23765 & ~w25072;
assign w25657 = ~w23765 & ~w25071;
assign w25658 = ~w23821 & w25074;
assign w25659 = ~w23821 & w25073;
assign w25660 = ~w23871 & w25076;
assign w25661 = ~w23871 & w25075;
assign w25662 = ~w23913 & w25078;
assign w25663 = ~w23913 & w25077;
assign w25664 = ~w23952 & w25080;
assign w25665 = ~w23952 & w25079;
assign w25666 = w21367 & w21545;
assign w25667 = ~w21545 & ~w21543;
assign w25668 = ~w22824 & w22944;
assign w25669 = ~w23765 & ~w23763;
assign w25670 = w23763 & w23821;
assign w25671 = (w24462 & w24461) | (w24462 & ~w24440) | (w24461 & ~w24440);
assign w25672 = (w24462 & w24461) | (w24462 & ~w24441) | (w24461 & ~w24441);
assign w25673 = (~w20817 & w24474) | (~w20817 & ~w24725) | (w24474 & ~w24725);
assign w25674 = (~w20817 & w24474) | (~w20817 & ~w24724) | (w24474 & ~w24724);
assign w25675 = (w24477 & w24478) | (w24477 & ~w24725) | (w24478 & ~w24725);
assign w25676 = (w24477 & w24478) | (w24477 & ~w24724) | (w24478 & ~w24724);
assign w25677 = (w24481 & w24482) | (w24481 & w24725) | (w24482 & w24725);
assign w25678 = (w24481 & w24482) | (w24481 & w24724) | (w24482 & w24724);
assign w25679 = (w24486 & w24485) | (w24486 & ~w24725) | (w24485 & ~w24725);
assign w25680 = (w24486 & w24485) | (w24486 & ~w24724) | (w24485 & ~w24724);
assign w25681 = (w24490 & w24489) | (w24490 & ~w24725) | (w24489 & ~w24725);
assign w25682 = (w24490 & w24489) | (w24490 & ~w24724) | (w24489 & ~w24724);
assign w25683 = (w24494 & w24493) | (w24494 & w24725) | (w24493 & w24725);
assign w25684 = (w24494 & w24493) | (w24494 & w24724) | (w24493 & w24724);
assign w25685 = (w24498 & w24497) | (w24498 & ~w24725) | (w24497 & ~w24725);
assign w25686 = (w24498 & w24497) | (w24498 & ~w24724) | (w24497 & ~w24724);
assign w25687 = (w24502 & w24501) | (w24502 & ~w24725) | (w24501 & ~w24725);
assign w25688 = (w24502 & w24501) | (w24502 & ~w24724) | (w24501 & ~w24724);
assign w25689 = (w24504 & w24503) | (w24504 & ~w24725) | (w24503 & ~w24725);
assign w25690 = (w24504 & w24503) | (w24504 & ~w24724) | (w24503 & ~w24724);
assign w25691 = ~w22309 & ~w25351;
assign w25692 = ~w22309 & ~w25350;
assign w25693 = ~w22445 & w25354;
assign w25694 = ~w22445 & w25353;
assign w25695 = ~w22576 & ~w25356;
assign w25696 = ~w22576 & ~w25355;
assign w25697 = ~w22702 & ~w25359;
assign w25698 = ~w22702 & ~w25358;
assign w25699 = ~w22826 & w25361;
assign w25700 = ~w22826 & w25360;
assign w25701 = ~w22944 & ~w25363;
assign w25702 = ~w22944 & ~w25362;
assign w25703 = ~w23053 & ~w25366;
assign w25704 = ~w23053 & ~w25365;
assign w25705 = ~w23156 & w25371;
assign w25706 = ~w23156 & w25370;
assign w25707 = ~w23248 & w25376;
assign w25708 = ~w23248 & w25375;
assign w25709 = (w24902 & w24901) | (w24902 & w25645) | (w24901 & w25645);
assign w25710 = (w24902 & w24901) | (w24902 & w25644) | (w24901 & w25644);
assign w25711 = (w24904 & w24903) | (w24904 & ~w25645) | (w24903 & ~w25645);
assign w25712 = (w24904 & w24903) | (w24904 & ~w25644) | (w24903 & ~w25644);
assign w25713 = (w24906 & w24905) | (w24906 & w25645) | (w24905 & w25645);
assign w25714 = (w24906 & w24905) | (w24906 & w25644) | (w24905 & w25644);
assign w25715 = (w24908 & w24907) | (w24908 & ~w25645) | (w24907 & ~w25645);
assign w25716 = (w24908 & w24907) | (w24908 & ~w25644) | (w24907 & ~w25644);
assign w25717 = (w111 & ~w24090) | (w111 & ~w113) | (~w24090 & ~w113);
assign w25718 = (~w212 & ~w213) | (~w212 & w25770) | (~w213 & w25770);
assign w25719 = (~w318 & ~w319) | (~w318 & w25771) | (~w319 & w25771);
assign w25720 = (w464 & ~w24180) | (w464 & ~w466) | (~w24180 & ~w466);
assign w25721 = (~w24198 & ~w24199) | (~w24198 & ~w466) | (~w24199 & ~w466);
assign w25722 = (w709 & ~w24237) | (w709 & ~w711) | (~w24237 & ~w711);
assign w25723 = ~w794 & ~w798;
assign w25724 = (w1003 & ~w24296) | (w1003 & ~w1005) | (~w24296 & ~w1005);
assign w25725 = ~w1103 & ~w1107;
assign w25726 = (w12792 & w12795) | (w12792 & ~w25200) | (w12795 & ~w25200);
assign w25727 = (~w12794 & ~w13178) | (~w12794 & w25311) | (~w13178 & w25311);
assign w25728 = w24605 & ~w14577;
assign w25729 = (~w14903 & ~w14904) | (~w14903 & w25728) | (~w14904 & w25728);
assign w25730 = (w15573 & w25447) | (w15573 & ~w9657) | (w25447 & ~w9657);
assign w25731 = w24606 & ~w15542;
assign w25732 = (w16123 & w25450) | (w16123 & ~w11035) | (w25450 & ~w11035);
assign w25733 = (~w16415 & ~w25455) | (~w16415 & ~w10339) | (~w25455 & ~w10339);
assign w25734 = (~w17275 & ~w25318) | (~w17275 & ~w10339) | (~w25318 & ~w10339);
assign w25735 = (w17520 & w25021) | (w17520 & ~w9657) | (w25021 & ~w9657);
assign w25736 = (w17550 & w24718) | (w17550 & ~w11763) | (w24718 & ~w11763);
assign w25737 = (w17817 & w25022) | (w17817 & ~w11035) | (w25022 & ~w11035);
assign w25738 = (~w17855 & ~w25321) | (~w17855 & ~w10339) | (~w25321 & ~w10339);
assign w25739 = (~w24436 & ~w24437) | (~w24436 & ~w16450) | (~w24437 & ~w16450);
assign w25740 = (w18584 & w25323) | (w18584 & ~w11035) | (w25323 & ~w11035);
assign w25741 = (w20399 & w25325) | (w20399 & ~w10371) | (w25325 & ~w10371);
assign w25742 = (~w20448 & ~w25478) | (~w20448 & ~w8998) | (~w25478 & ~w8998);
assign w25743 = (~w20588 & ~w25326) | (~w20588 & ~w9992) | (~w25326 & ~w9992);
assign w25744 = (w21163 & w25496) | (w21163 & ~w11035) | (w25496 & ~w11035);
assign w25745 = (w21179 & w25498) | (w21179 & ~w12132) | (w25498 & ~w12132);
assign w25746 = (w24489 & w24490) | (w24489 & ~w20820) | (w24490 & ~w20820);
assign w25747 = (w21724 & w25036) | (w21724 & ~w11400) | (w25036 & ~w11400);
assign w25748 = (w21999 & w25341) | (w21999 & ~w10371) | (w25341 & ~w10371);
assign w25749 = (~w22039 & ~w25502) | (~w22039 & ~w8998) | (~w25502 & ~w8998);
assign w25750 = (~w22128 & ~w25342) | (~w22128 & ~w9992) | (~w25342 & ~w9992);
assign w25751 = (w22318 & w25510) | (w22318 & ~w11763) | (w25510 & ~w11763);
assign w25752 = (w23126 & w25043) | (w23126 & ~w10371) | (w25043 & ~w10371);
assign w25753 = (~w23174 & ~w25044) | (~w23174 & ~w9992) | (~w25044 & ~w9992);
assign w25754 = (~w23183 & ~w25227) | (~w23183 & ~w8998) | (~w25227 & ~w8998);
assign w25755 = (w23234 & w24728) | (w23234 & ~w12132) | (w24728 & ~w12132);
assign w25756 = (w23343 & w24894) | (w23343 & ~w11763) | (w24894 & ~w11763);
assign w25757 = (~a[2] & ~w24067) | (~a[2] & ~w47) | (~w24067 & ~w47);
assign w25758 = ~w23638 & ~w24551;
assign w25759 = (~w24577 & ~w24578) | (~w24577 & w23983) | (~w24578 & w23983);
assign w25760 = (~w24577 & ~w24578) | (~w24577 & ~w24575) | (~w24578 & ~w24575);
assign w25761 = ~w24031 & w25759;
assign w25762 = ~w24031 & w25760;
assign w25763 = (~w24583 & ~w24584) | (~w24583 & w23983) | (~w24584 & w23983);
assign w25764 = (~w24583 & ~w24584) | (~w24583 & ~w24575) | (~w24584 & ~w24575);
assign w25765 = (~w12177 & ~w24755) | (~w12177 & ~w12496) | (~w24755 & ~w12496);
assign w25766 = ~w7312 | ~w24731;
assign w25767 = (~w24731 & ~w7312) | (~w24731 & ~w11760) | (~w7312 & ~w11760);
assign w25768 = (w24553 & w25758) | (w24553 & w24537) | (w25758 & w24537);
assign w25769 = (w24553 & w25758) | (w24553 & w24538) | (w25758 & w24538);
assign w25770 = w24590 & ~w156;
assign w25771 = w24593 & ~w268;
assign one = 1;
assign f[0] = w0;// level 1
assign f[1] = w16;// level 6
assign f[2] = w33;// level 8
assign f[3] = w56;// level 11
assign f[4] = w97;// level 12
assign f[5] = w133;// level 14
assign f[6] = w169;// level 15
assign f[7] = w228;// level 17
assign f[8] = w283;// level 18
assign f[9] = ~w335;// level 20
assign f[10] = w410;// level 21
assign f[11] = w481;// level 23
assign f[12] = w549;// level 24
assign f[13] = ~w640;// level 26
assign f[14] = w727;// level 27
assign f[15] = ~w811;// level 29
assign f[16] = w918;// level 30
assign f[17] = ~w1021;// level 32
assign f[18] = w1121;// level 33
assign f[19] = ~w1244;// level 35
assign f[20] = w1360;// level 36
assign f[21] = ~w1482;// level 38
assign f[22] = w1630;// level 39
assign f[23] = ~w1770;// level 41
assign f[24] = w1910;// level 42
assign f[25] = w2075;// level 44
assign f[26] = w2234;// level 45
assign f[27] = w2392;// level 47
assign f[28] = w2574;// level 48
assign f[29] = w2748;// level 50
assign f[30] = w2923;// level 51
assign f[31] = ~w3127;// level 53
assign f[32] = w3319;// level 54
assign f[33] = w3513;// level 56
assign f[34] = w3725;// level 58
assign f[35] = w3932;// level 60
assign f[36] = w4144;// level 62
assign f[37] = w4371;// level 63
assign f[38] = w4597;// level 64
assign f[39] = ~w4827;// level 65
assign f[40] = w5073;// level 67
assign f[41] = w5316;// level 69
assign f[42] = w5563;// level 71
assign f[43] = ~w5826;// level 72
assign f[44] = w6084;// level 74
assign f[45] = w6348;// level 75
assign f[46] = w6628;// level 76
assign f[47] = ~w6904;// level 78
assign f[48] = w7185;// level 80
assign f[49] = w7482;// level 81
assign f[50] = w7774;// level 83
assign f[51] = w8072;// level 85
assign f[52] = w8386;// level 86
assign f[53] = w8697;// level 87
assign f[54] = w9013;// level 88
assign f[55] = w9344;// level 90
assign f[56] = w9672;// level 91
assign f[57] = w10006;// level 92
assign f[58] = ~w10354;// level 94
assign f[59] = w10702;// level 96
assign f[60] = w11053;// level 96
assign f[61] = ~w11418;// level 98
assign f[62] = w11782;// level 100
assign f[63] = ~w12150;// level 100
assign f[64] = ~w12512;// level 102
assign f[65] = w12867;// level 103
assign f[66] = ~w13213;// level 104
assign f[67] = w13561;// level 105
assign f[68] = w13907;// level 104
assign f[69] = ~w14247;// level 104
assign f[70] = w14579;// level 105
assign f[71] = w14908;// level 106
assign f[72] = ~w15230;// level 107
assign f[73] = w15545;// level 105
assign f[74] = w15851;// level 106
assign f[75] = w16155;// level 107
assign f[76] = w16449;// level 106
assign f[77] = w16741;// level 107
assign f[78] = w17030;// level 107
assign f[79] = w17309;// level 107
assign f[80] = w17580;// level 107
assign f[81] = w17849;// level 107
assign f[82] = w18108;// level 108
assign f[83] = w18366;// level 109
assign f[84] = w18618;// level 108
assign f[85] = w18862;// level 108
assign f[86] = w19106;// level 108
assign f[87] = ~w19344;// level 108
assign f[88] = w19574;// level 108
assign f[89] = w19801;// level 108
assign f[90] = w20022;// level 108
assign f[91] = w20235;// level 109
assign f[92] = w20440;// level 109
assign f[93] = w20635;// level 109
assign f[94] = w20823;// level 108
assign f[95] = w21011;// level 109
assign f[96] = ~w21194;// level 109
assign f[97] = w21373;// level 109
assign f[98] = w21549;// level 109
assign f[99] = ~w21718;// level 109
assign f[100] = w21877;// level 109
assign f[101] = w22032;// level 109
assign f[102] = ~w22176;// level 109
assign f[103] = w22312;// level 109
assign f[104] = w22448;// level 109
assign f[105] = ~w22579;// level 109
assign f[106] = w22705;// level 109
assign f[107] = w22829;// level 109
assign f[108] = ~w22947;// level 109
assign f[109] = w23056;// level 109
assign f[110] = w23159;// level 109
assign f[111] = w23251;// level 109
assign f[112] = w23338;// level 109
assign f[113] = w23421;// level 109
assign f[114] = ~w23500;// level 109
assign f[115] = w23572;// level 109
assign f[116] = w23642;// level 109
assign f[117] = ~w23709;// level 109
assign f[118] = w23768;// level 109
assign f[119] = w23824;// level 109
assign f[120] = w23874;// level 109
assign f[121] = w23916;// level 109
assign f[122] = w23955;// level 109
assign f[123] = w23988;// level 109
assign f[124] = w24013;// level 109
assign f[125] = w24035;// level 109
assign f[126] = ~w24050;// level 109
assign f[127] = w24056;// level 109
endmodule
