module des_area ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71;
  wire n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
    n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
    n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
    n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
    n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
    n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
    n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
    n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
    n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
    n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
    n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
    n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
    n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
    n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
    n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
    n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
    n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
    n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
    n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
    n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3530, n3531, n3532,
    n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
    n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
    n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
    n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
    n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
    n3828, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
    n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
    n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
    n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
    n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
    n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
    n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
    n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
    n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
    n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
    n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
    n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
    n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
    n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
    n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5081,
    n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
    n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
    n5214, n5215, n5216, n5217, n5218, n5219, n5221, n5222, n5223, n5224,
    n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297;
  assign n442 = ~pi364 & ~pi365;
  assign n443 = ~pi366 & n442;
  assign n444 = ~pi362 & ~pi367;
  assign n445 = ~pi363 & n444;
  assign n446 = n443 & n445;
  assign n447 = pi128 & n446;
  assign n448 = pi366 & n442;
  assign n449 = n445 & n448;
  assign n450 = pi000 & n449;
  assign n451 = ~pi366 & pi367;
  assign n452 = ~pi362 & ~pi363;
  assign n453 = n451 & n452;
  assign n454 = n442 & n453;
  assign n455 = pi090 & ~n454;
  assign n456 = pi000 & n454;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~n449 & ~n457;
  assign n459 = ~n450 & ~n458;
  assign n460 = ~n446 & ~n459;
  assign n461 = ~n447 & ~n460;
  assign n462 = pi364 & ~pi365;
  assign n463 = pi362 & ~pi363;
  assign n464 = n462 & n463;
  assign n465 = pi366 & ~pi367;
  assign n466 = pi360 & ~n465;
  assign n467 = ~pi360 & n465;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~pi360 & ~pi366;
  assign n470 = pi367 & n469;
  assign n471 = pi325 & n470;
  assign n472 = ~pi366 & ~pi367;
  assign n473 = ~pi360 & n472;
  assign n474 = pi360 & n451;
  assign n475 = ~n473 & ~n474;
  assign n476 = pi213 & ~n475;
  assign n477 = ~n471 & ~n476;
  assign n478 = pi360 & n465;
  assign n479 = ~pi360 & ~pi367;
  assign n480 = pi366 & n479;
  assign n481 = ~n478 & ~n480;
  assign n482 = pi269 & ~n481;
  assign n483 = pi360 & n472;
  assign n484 = pi325 & n483;
  assign n485 = ~n482 & ~n484;
  assign n486 = n477 & n485;
  assign n487 = ~n468 & ~n486;
  assign n488 = pi236 & ~n475;
  assign n489 = pi348 & n470;
  assign n490 = ~n488 & ~n489;
  assign n491 = pi348 & n483;
  assign n492 = pi292 & n465;
  assign n493 = ~n491 & ~n492;
  assign n494 = n490 & n493;
  assign n495 = n468 & ~n494;
  assign n496 = ~n487 & ~n495;
  assign n497 = n464 & ~n496;
  assign n498 = pi362 & pi363;
  assign n499 = n442 & n498;
  assign n500 = pi208 & ~n475;
  assign n501 = pi320 & n470;
  assign n502 = ~n500 & ~n501;
  assign n503 = pi320 & n483;
  assign n504 = pi264 & ~n481;
  assign n505 = ~n503 & ~n504;
  assign n506 = n502 & n505;
  assign n507 = n468 & ~n506;
  assign n508 = pi353 & n470;
  assign n509 = pi241 & ~n475;
  assign n510 = ~n508 & ~n509;
  assign n511 = pi297 & ~n481;
  assign n512 = pi353 & n483;
  assign n513 = ~n511 & ~n512;
  assign n514 = n510 & n513;
  assign n515 = ~n468 & ~n514;
  assign n516 = ~n507 & ~n515;
  assign n517 = n499 & ~n516;
  assign n518 = ~n497 & ~n517;
  assign n519 = ~pi364 & pi365;
  assign n520 = n452 & n519;
  assign n521 = pi356 & n470;
  assign n522 = pi244 & ~n475;
  assign n523 = ~n521 & ~n522;
  assign n524 = pi356 & n483;
  assign n525 = pi300 & ~n481;
  assign n526 = ~n524 & ~n525;
  assign n527 = n523 & n526;
  assign n528 = n468 & ~n527;
  assign n529 = pi349 & n470;
  assign n530 = pi237 & ~n475;
  assign n531 = ~n529 & ~n530;
  assign n532 = pi349 & n483;
  assign n533 = pi293 & ~n481;
  assign n534 = ~n532 & ~n533;
  assign n535 = n531 & n534;
  assign n536 = ~n468 & ~n535;
  assign n537 = ~n528 & ~n536;
  assign n538 = n520 & ~n537;
  assign n539 = ~pi362 & pi363;
  assign n540 = n442 & n539;
  assign n541 = pi200 & ~n475;
  assign n542 = pi312 & n483;
  assign n543 = pi256 & ~n481;
  assign n544 = ~n542 & ~n543;
  assign n545 = pi312 & n470;
  assign n546 = n544 & ~n545;
  assign n547 = ~n541 & n546;
  assign n548 = ~n468 & ~n547;
  assign n549 = pi306 & n483;
  assign n550 = pi250 & ~n481;
  assign n551 = ~n549 & ~n550;
  assign n552 = pi306 & n470;
  assign n553 = pi194 & ~n475;
  assign n554 = ~n552 & ~n553;
  assign n555 = n551 & n554;
  assign n556 = n468 & ~n555;
  assign n557 = ~n548 & ~n556;
  assign n558 = n540 & ~n557;
  assign n559 = ~n538 & ~n558;
  assign n560 = n442 & n463;
  assign n561 = pi347 & n470;
  assign n562 = pi235 & ~n475;
  assign n563 = ~n561 & ~n562;
  assign n564 = pi291 & ~n481;
  assign n565 = pi347 & n483;
  assign n566 = ~n564 & ~n565;
  assign n567 = n563 & n566;
  assign n568 = n468 & ~n567;
  assign n569 = pi270 & ~n481;
  assign n570 = pi326 & n483;
  assign n571 = ~n569 & ~n570;
  assign n572 = pi214 & ~n475;
  assign n573 = pi326 & n470;
  assign n574 = ~n572 & ~n573;
  assign n575 = n571 & n574;
  assign n576 = ~n468 & ~n575;
  assign n577 = ~n568 & ~n576;
  assign n578 = n560 & ~n577;
  assign n579 = n498 & n519;
  assign n580 = pi222 & ~n475;
  assign n581 = pi334 & n470;
  assign n582 = ~n580 & ~n581;
  assign n583 = pi334 & n483;
  assign n584 = pi278 & ~n481;
  assign n585 = ~n583 & ~n584;
  assign n586 = n582 & n585;
  assign n587 = ~n468 & ~n586;
  assign n588 = pi339 & n483;
  assign n589 = pi283 & ~n481;
  assign n590 = ~n588 & ~n589;
  assign n591 = pi227 & ~n475;
  assign n592 = pi339 & n470;
  assign n593 = ~n591 & ~n592;
  assign n594 = n590 & n593;
  assign n595 = n468 & ~n594;
  assign n596 = ~n587 & ~n595;
  assign n597 = n579 & ~n596;
  assign n598 = ~n578 & ~n597;
  assign n599 = n559 & n598;
  assign n600 = pi364 & pi365;
  assign n601 = n539 & n600;
  assign n602 = ~n468 & ~n567;
  assign n603 = n468 & ~n575;
  assign n604 = ~n602 & ~n603;
  assign n605 = n601 & ~n604;
  assign n606 = n452 & n600;
  assign n607 = n468 & ~n514;
  assign n608 = ~n468 & ~n506;
  assign n609 = ~n607 & ~n608;
  assign n610 = n606 & ~n609;
  assign n611 = ~n605 & ~n610;
  assign n612 = n599 & n611;
  assign n613 = n462 & n539;
  assign n614 = pi311 & n470;
  assign n615 = pi255 & ~n481;
  assign n616 = ~n614 & ~n615;
  assign n617 = pi311 & n483;
  assign n618 = pi199 & ~n475;
  assign n619 = ~n617 & ~n618;
  assign n620 = n616 & n619;
  assign n621 = ~n468 & ~n620;
  assign n622 = pi223 & ~n475;
  assign n623 = pi335 & n470;
  assign n624 = ~n622 & ~n623;
  assign n625 = pi279 & ~n481;
  assign n626 = pi335 & n483;
  assign n627 = ~n625 & ~n626;
  assign n628 = n624 & n627;
  assign n629 = n468 & ~n628;
  assign n630 = ~n621 & ~n629;
  assign n631 = n613 & ~n630;
  assign n632 = n462 & n498;
  assign n633 = ~n468 & ~n527;
  assign n634 = n468 & ~n535;
  assign n635 = ~n633 & ~n634;
  assign n636 = n632 & ~n635;
  assign n637 = ~n631 & ~n636;
  assign n638 = n519 & n539;
  assign n639 = ~n468 & ~n494;
  assign n640 = n468 & ~n486;
  assign n641 = ~n639 & ~n640;
  assign n642 = n638 & ~n641;
  assign n643 = n463 & n519;
  assign n644 = n468 & ~n620;
  assign n645 = ~n468 & ~n628;
  assign n646 = ~n644 & ~n645;
  assign n647 = n643 & ~n646;
  assign n648 = ~n642 & ~n647;
  assign n649 = n637 & n648;
  assign n650 = n498 & n600;
  assign n651 = pi333 & n470;
  assign n652 = pi221 & ~n475;
  assign n653 = ~n651 & ~n652;
  assign n654 = pi277 & ~n481;
  assign n655 = pi333 & n483;
  assign n656 = ~n654 & ~n655;
  assign n657 = n653 & n656;
  assign n658 = n468 & ~n657;
  assign n659 = pi228 & pi360;
  assign n660 = ~pi366 & n659;
  assign n661 = pi367 & n660;
  assign n662 = pi284 & ~n481;
  assign n663 = pi340 & n470;
  assign n664 = pi228 & n473;
  assign n665 = ~n663 & ~n664;
  assign n666 = pi340 & n483;
  assign n667 = n665 & ~n666;
  assign n668 = ~n662 & n667;
  assign n669 = ~n661 & n668;
  assign n670 = ~n468 & ~n669;
  assign n671 = ~n658 & ~n670;
  assign n672 = n650 & ~n671;
  assign n673 = n463 & n600;
  assign n674 = ~n468 & ~n555;
  assign n675 = n468 & ~n547;
  assign n676 = ~n674 & ~n675;
  assign n677 = n673 & ~n676;
  assign n678 = n452 & n462;
  assign n679 = n468 & ~n586;
  assign n680 = ~n468 & ~n594;
  assign n681 = ~n679 & ~n680;
  assign n682 = n678 & ~n681;
  assign n683 = ~n677 & ~n682;
  assign n684 = n442 & n452;
  assign n685 = ~n468 & ~n657;
  assign n686 = n468 & ~n669;
  assign n687 = ~n685 & ~n686;
  assign n688 = n684 & ~n687;
  assign n689 = n683 & ~n688;
  assign n690 = ~n672 & n689;
  assign n691 = n649 & n690;
  assign n692 = n612 & n691;
  assign n693 = n518 & n692;
  assign n694 = ~n449 & ~n454;
  assign n695 = pi063 & n694;
  assign n696 = pi107 & ~n694;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n446 & ~n697;
  assign n699 = pi189 & n446;
  assign po61 = n698 | n699;
  assign n701 = ~n693 & ~po61;
  assign n702 = n693 & po61;
  assign n703 = ~n701 & ~n702;
  assign n704 = ~pi043 & ~n454;
  assign n705 = ~pi101 & n454;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n449 & n706;
  assign n708 = pi101 & n449;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~n446 & ~n709;
  assign n711 = pi163 & n446;
  assign po35 = n710 | n711;
  assign n713 = ~n537 & n684;
  assign n714 = pi230 & ~n475;
  assign n715 = pi342 & n470;
  assign n716 = ~n714 & ~n715;
  assign n717 = pi286 & ~n481;
  assign n718 = pi342 & n483;
  assign n719 = ~n717 & ~n718;
  assign n720 = n716 & n719;
  assign n721 = n468 & ~n720;
  assign n722 = pi248 & ~n481;
  assign n723 = pi304 & n483;
  assign n724 = ~n722 & ~n723;
  assign n725 = pi192 & ~n475;
  assign n726 = pi304 & n470;
  assign n727 = ~n725 & ~n726;
  assign n728 = n724 & n727;
  assign n729 = ~n468 & ~n728;
  assign n730 = ~n721 & ~n729;
  assign n731 = n601 & ~n730;
  assign n732 = pi299 & ~n481;
  assign n733 = pi355 & n483;
  assign n734 = ~n732 & ~n733;
  assign n735 = pi355 & n470;
  assign n736 = pi243 & ~n475;
  assign n737 = ~n735 & ~n736;
  assign n738 = n734 & n737;
  assign n739 = ~n468 & ~n738;
  assign n740 = pi262 & ~n481;
  assign n741 = pi318 & n483;
  assign n742 = ~n740 & ~n741;
  assign n743 = pi206 & ~n475;
  assign n744 = pi318 & n470;
  assign n745 = ~n743 & ~n744;
  assign n746 = n742 & n745;
  assign n747 = n468 & ~n746;
  assign n748 = ~n739 & ~n747;
  assign n749 = n540 & ~n748;
  assign n750 = pi271 & ~n481;
  assign n751 = pi327 & n483;
  assign n752 = ~n750 & ~n751;
  assign n753 = pi327 & n470;
  assign n754 = pi215 & ~n475;
  assign n755 = ~n753 & ~n754;
  assign n756 = n752 & n755;
  assign n757 = n468 & ~n756;
  assign n758 = pi290 & ~n481;
  assign n759 = pi346 & n483;
  assign n760 = ~n758 & ~n759;
  assign n761 = pi234 & ~n475;
  assign n762 = pi346 & n470;
  assign n763 = ~n761 & ~n762;
  assign n764 = n760 & n763;
  assign n765 = ~n468 & ~n764;
  assign n766 = ~n757 & ~n765;
  assign n767 = n579 & ~n766;
  assign n768 = ~n749 & ~n767;
  assign n769 = n520 & ~n687;
  assign n770 = n768 & ~n769;
  assign n771 = ~n731 & n770;
  assign n772 = ~n713 & n771;
  assign n773 = n468 & ~n738;
  assign n774 = ~n468 & ~n746;
  assign n775 = ~n773 & ~n774;
  assign n776 = n673 & ~n775;
  assign n777 = ~n635 & n650;
  assign n778 = pi249 & ~n481;
  assign n779 = pi193 & ~n475;
  assign n780 = ~n778 & ~n779;
  assign n781 = pi305 & n483;
  assign n782 = pi305 & n470;
  assign n783 = ~n781 & ~n782;
  assign n784 = n780 & n783;
  assign n785 = ~n468 & ~n784;
  assign n786 = pi313 & n483;
  assign n787 = pi257 & ~n481;
  assign n788 = ~n786 & ~n787;
  assign n789 = pi201 & ~n475;
  assign n790 = pi313 & n470;
  assign n791 = ~n789 & ~n790;
  assign n792 = n788 & n791;
  assign n793 = n468 & ~n792;
  assign n794 = ~n785 & ~n793;
  assign n795 = n638 & ~n794;
  assign n796 = ~n777 & ~n795;
  assign n797 = ~n468 & ~n756;
  assign n798 = n468 & ~n764;
  assign n799 = ~n797 & ~n798;
  assign n800 = n678 & ~n799;
  assign n801 = n632 & ~n671;
  assign n802 = ~n800 & ~n801;
  assign n803 = n796 & n802;
  assign n804 = pi276 & ~n481;
  assign n805 = pi332 & n483;
  assign n806 = ~n804 & ~n805;
  assign n807 = pi220 & ~n475;
  assign n808 = pi332 & n470;
  assign n809 = ~n807 & ~n808;
  assign n810 = n806 & n809;
  assign n811 = n468 & ~n810;
  assign n812 = pi341 & n483;
  assign n813 = pi285 & ~n481;
  assign n814 = ~n812 & ~n813;
  assign n815 = pi341 & n470;
  assign n816 = pi229 & ~n475;
  assign n817 = ~n815 & ~n816;
  assign n818 = n814 & n817;
  assign n819 = ~n468 & ~n818;
  assign n820 = ~n811 & ~n819;
  assign n821 = n499 & ~n820;
  assign n822 = ~n468 & ~n720;
  assign n823 = n468 & ~n728;
  assign n824 = ~n822 & ~n823;
  assign n825 = n560 & ~n824;
  assign n826 = ~n821 & ~n825;
  assign n827 = ~n468 & ~n810;
  assign n828 = n468 & ~n818;
  assign n829 = ~n827 & ~n828;
  assign n830 = n606 & ~n829;
  assign n831 = n468 & ~n784;
  assign n832 = ~n468 & ~n792;
  assign n833 = ~n831 & ~n832;
  assign n834 = n464 & ~n833;
  assign n835 = ~n830 & ~n834;
  assign n836 = n826 & n835;
  assign n837 = pi319 & n483;
  assign n838 = pi263 & ~n481;
  assign n839 = ~n837 & ~n838;
  assign n840 = pi207 & ~n475;
  assign n841 = pi319 & n470;
  assign n842 = ~n840 & ~n841;
  assign n843 = n839 & n842;
  assign n844 = n468 & ~n843;
  assign n845 = pi298 & ~n481;
  assign n846 = pi354 & n483;
  assign n847 = ~n845 & ~n846;
  assign n848 = pi354 & n470;
  assign n849 = pi242 & ~n475;
  assign n850 = ~n848 & ~n849;
  assign n851 = n847 & n850;
  assign n852 = ~n468 & ~n851;
  assign n853 = ~n844 & ~n852;
  assign n854 = n613 & ~n853;
  assign n855 = ~n468 & ~n843;
  assign n856 = n468 & ~n851;
  assign n857 = ~n855 & ~n856;
  assign n858 = n643 & ~n857;
  assign n859 = ~n854 & ~n858;
  assign n860 = n836 & n859;
  assign n861 = n803 & n860;
  assign n862 = ~n776 & n861;
  assign n863 = n772 & n862;
  assign n864 = po35 & n863;
  assign n865 = ~po35 & ~n863;
  assign n866 = ~n864 & ~n865;
  assign n867 = pi139 & n446;
  assign n868 = pi049 & ~n454;
  assign n869 = pi119 & n454;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n449 & ~n870;
  assign n872 = pi119 & n449;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n446 & ~n873;
  assign po11 = n867 | n874;
  assign n876 = ~n640 & ~n774;
  assign n877 = n684 & ~n876;
  assign n878 = ~n602 & ~n757;
  assign n879 = n643 & ~n878;
  assign n880 = ~n877 & ~n879;
  assign n881 = ~n487 & ~n747;
  assign n882 = n650 & ~n881;
  assign n883 = ~n568 & ~n797;
  assign n884 = n613 & ~n883;
  assign n885 = ~n882 & ~n884;
  assign n886 = n880 & n885;
  assign n887 = ~n556 & ~n832;
  assign n888 = n632 & ~n887;
  assign n889 = ~n528 & ~n765;
  assign n890 = n673 & ~n889;
  assign n891 = ~n888 & ~n890;
  assign n892 = ~n739 & ~n844;
  assign n893 = n678 & ~n892;
  assign n894 = ~n685 & ~n828;
  assign n895 = n638 & ~n894;
  assign n896 = ~n893 & ~n895;
  assign n897 = n891 & n896;
  assign n898 = ~n773 & ~n855;
  assign n899 = n579 & ~n898;
  assign n900 = ~n822 & ~n831;
  assign n901 = n499 & ~n900;
  assign n902 = ~n899 & ~n901;
  assign n903 = ~n633 & ~n798;
  assign n904 = n540 & ~n903;
  assign n905 = ~n621 & ~n811;
  assign n906 = n560 & ~n905;
  assign n907 = ~n904 & ~n906;
  assign n908 = n902 & n907;
  assign n909 = n897 & n908;
  assign n910 = n886 & n909;
  assign n911 = ~n644 & ~n827;
  assign n912 = n601 & ~n911;
  assign n913 = ~n721 & ~n785;
  assign n914 = n606 & ~n913;
  assign n915 = ~n912 & ~n914;
  assign n916 = ~n658 & ~n819;
  assign n917 = n464 & ~n916;
  assign n918 = ~n674 & ~n793;
  assign n919 = n520 & ~n918;
  assign n920 = ~n917 & ~n919;
  assign n921 = n915 & n920;
  assign n922 = n910 & n921;
  assign n923 = ~po11 & ~n922;
  assign n924 = po11 & n922;
  assign n925 = ~n923 & ~n924;
  assign n926 = ~n568 & ~n680;
  assign n927 = n638 & ~n926;
  assign n928 = ~n633 & ~n679;
  assign n929 = n673 & ~n928;
  assign n930 = ~n927 & ~n929;
  assign n931 = ~n507 & ~n621;
  assign n932 = n606 & ~n931;
  assign n933 = ~n487 & ~n556;
  assign n934 = n579 & ~n933;
  assign n935 = ~n932 & ~n934;
  assign n936 = ~n639 & ~n721;
  assign n937 = n560 & ~n936;
  assign n938 = ~n495 & ~n822;
  assign n939 = n601 & ~n938;
  assign n940 = ~n937 & ~n939;
  assign n941 = n935 & n940;
  assign n942 = ~n548 & ~n844;
  assign n943 = n520 & ~n942;
  assign n944 = ~n595 & ~n602;
  assign n945 = n464 & ~n944;
  assign n946 = ~n943 & ~n945;
  assign n947 = ~n528 & ~n587;
  assign n948 = n540 & ~n947;
  assign n949 = ~n608 & ~n644;
  assign n950 = n499 & ~n949;
  assign n951 = ~n948 & ~n950;
  assign n952 = n946 & n951;
  assign n953 = n941 & n952;
  assign n954 = ~n629 & ~n739;
  assign n955 = n684 & ~n954;
  assign n956 = ~n645 & ~n773;
  assign n957 = n650 & ~n956;
  assign n958 = ~n955 & ~n957;
  assign n959 = ~n640 & ~n674;
  assign n960 = n678 & ~n959;
  assign n961 = ~n675 & ~n855;
  assign n962 = n632 & ~n961;
  assign n963 = ~n960 & ~n962;
  assign n964 = ~n607 & ~n685;
  assign n965 = n613 & ~n964;
  assign n966 = ~n515 & ~n658;
  assign n967 = n643 & ~n966;
  assign n968 = ~n965 & ~n967;
  assign n969 = n963 & n968;
  assign n970 = n958 & n969;
  assign n971 = n953 & n970;
  assign n972 = n930 & n971;
  assign n973 = pi075 & n449;
  assign n974 = ~pi059 & ~n454;
  assign n975 = ~pi075 & n454;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n449 & n976;
  assign n978 = ~n973 & ~n977;
  assign n979 = ~n446 & ~n978;
  assign n980 = pi131 & n446;
  assign po03 = n979 | n980;
  assign n982 = n972 & po03;
  assign n983 = ~n972 & ~po03;
  assign n984 = ~n982 & ~n983;
  assign n985 = ~n925 & n984;
  assign n986 = n866 & n985;
  assign n987 = n703 & n986;
  assign n988 = ~n639 & ~n856;
  assign n989 = n673 & ~n988;
  assign n990 = ~n680 & ~n811;
  assign n991 = n632 & ~n990;
  assign n992 = ~n989 & ~n991;
  assign n993 = ~n607 & ~n774;
  assign n994 = n643 & ~n993;
  assign n995 = ~n515 & ~n747;
  assign n996 = n613 & ~n995;
  assign n997 = ~n994 & ~n996;
  assign n998 = n992 & n997;
  assign n999 = ~n608 & ~n757;
  assign n1000 = n684 & ~n999;
  assign n1001 = ~n507 & ~n797;
  assign n1002 = n650 & ~n1001;
  assign n1003 = ~n1000 & ~n1002;
  assign n1004 = ~n587 & ~n793;
  assign n1005 = n601 & ~n1004;
  assign n1006 = ~n595 & ~n827;
  assign n1007 = n520 & ~n1006;
  assign n1008 = ~n1005 & ~n1007;
  assign n1009 = ~n495 & ~n852;
  assign n1010 = n540 & ~n1009;
  assign n1011 = ~n548 & ~n823;
  assign n1012 = n464 & ~n1011;
  assign n1013 = ~n1010 & ~n1012;
  assign n1014 = n1008 & n1013;
  assign n1015 = ~n645 & ~n686;
  assign n1016 = n606 & ~n1015;
  assign n1017 = ~n679 & ~n832;
  assign n1018 = n560 & ~n1017;
  assign n1019 = ~n1016 & ~n1018;
  assign n1020 = ~n629 & ~n670;
  assign n1021 = n499 & ~n1020;
  assign n1022 = ~n536 & ~n603;
  assign n1023 = n579 & ~n1022;
  assign n1024 = ~n1021 & ~n1023;
  assign n1025 = n1019 & n1024;
  assign n1026 = n1014 & n1025;
  assign n1027 = ~n576 & ~n634;
  assign n1028 = n678 & ~n1027;
  assign n1029 = ~n675 & ~n729;
  assign n1030 = n638 & ~n1029;
  assign n1031 = ~n1028 & ~n1030;
  assign n1032 = n1026 & n1031;
  assign n1033 = n1003 & n1032;
  assign n1034 = n998 & n1033;
  assign n1035 = pi155 & n446;
  assign n1036 = pi111 & n449;
  assign n1037 = pi031 & ~n454;
  assign n1038 = pi111 & n454;
  assign n1039 = ~n1037 & ~n1038;
  assign n1040 = ~n449 & ~n1039;
  assign n1041 = ~n1036 & ~n1040;
  assign n1042 = ~n446 & ~n1041;
  assign po27 = n1035 | n1042;
  assign n1044 = n1034 & po27;
  assign n1045 = ~n1034 & ~po27;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = ~n925 & ~n1046;
  assign n1048 = pi042 & ~n454;
  assign n1049 = pi084 & n454;
  assign n1050 = ~n1048 & ~n1049;
  assign n1051 = ~n449 & ~n1050;
  assign n1052 = pi084 & n449;
  assign n1053 = ~n1051 & ~n1052;
  assign n1054 = ~n446 & n1053;
  assign n1055 = ~pi147 & n446;
  assign po19 = ~n1054 & ~n1055;
  assign n1057 = ~n679 & ~n822;
  assign n1058 = n613 & ~n1057;
  assign n1059 = ~n548 & ~n831;
  assign n1060 = n650 & ~n1059;
  assign n1061 = ~n1058 & ~n1060;
  assign n1062 = ~n587 & ~n721;
  assign n1063 = n643 & ~n1062;
  assign n1064 = ~n556 & ~n621;
  assign n1065 = n678 & ~n1064;
  assign n1066 = ~n1063 & ~n1065;
  assign n1067 = n1061 & n1066;
  assign n1068 = ~n602 & ~n640;
  assign n1069 = n606 & ~n1068;
  assign n1070 = ~n495 & ~n739;
  assign n1071 = n632 & ~n1070;
  assign n1072 = ~n1069 & ~n1071;
  assign n1073 = ~n487 & ~n568;
  assign n1074 = n499 & ~n1073;
  assign n1075 = n1072 & ~n1074;
  assign n1076 = ~n675 & ~n785;
  assign n1077 = n684 & ~n1076;
  assign n1078 = ~n639 & ~n773;
  assign n1079 = n520 & ~n1078;
  assign n1080 = ~n1077 & ~n1079;
  assign n1081 = ~n595 & ~n685;
  assign n1082 = n673 & ~n1081;
  assign n1083 = n1080 & ~n1082;
  assign n1084 = ~n607 & ~n855;
  assign n1085 = n601 & ~n1084;
  assign n1086 = ~n507 & ~n633;
  assign n1087 = n464 & ~n1086;
  assign n1088 = ~n1085 & ~n1087;
  assign n1089 = ~n658 & ~n680;
  assign n1090 = n540 & ~n1089;
  assign n1091 = ~n515 & ~n844;
  assign n1092 = n560 & ~n1091;
  assign n1093 = ~n1090 & ~n1092;
  assign n1094 = n1088 & n1093;
  assign n1095 = ~n644 & ~n674;
  assign n1096 = n579 & ~n1095;
  assign n1097 = ~n528 & ~n608;
  assign n1098 = n638 & ~n1097;
  assign n1099 = ~n1096 & ~n1098;
  assign n1100 = n1094 & n1099;
  assign n1101 = n1083 & n1100;
  assign n1102 = n1075 & n1101;
  assign n1103 = n1067 & n1102;
  assign n1104 = ~po19 & ~n1103;
  assign n1105 = po19 & n1103;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~n866 & n984;
  assign n1108 = n1106 & n1107;
  assign n1109 = n1047 & n1108;
  assign n1110 = ~n703 & n866;
  assign n1111 = n984 & n1110;
  assign n1112 = n925 & ~n1046;
  assign n1113 = n1111 & n1112;
  assign n1114 = ~n1046 & ~n1106;
  assign n1115 = n925 & n984;
  assign n1116 = ~n703 & n1115;
  assign n1117 = ~n866 & ~n984;
  assign n1118 = n703 & n1117;
  assign n1119 = ~n1116 & ~n1118;
  assign n1120 = n1114 & ~n1119;
  assign n1121 = ~n703 & ~n984;
  assign n1122 = n1047 & ~n1106;
  assign n1123 = n1121 & n1122;
  assign n1124 = ~n1120 & ~n1123;
  assign n1125 = ~n1113 & n1124;
  assign n1126 = ~n1109 & n1125;
  assign n1127 = n703 & ~n1106;
  assign n1128 = n925 & ~n984;
  assign n1129 = n1127 & n1128;
  assign n1130 = n1126 & ~n1129;
  assign n1131 = ~n987 & n1130;
  assign n1132 = n703 & n984;
  assign n1133 = n866 & n1132;
  assign n1134 = ~n925 & ~n984;
  assign n1135 = ~n866 & n1134;
  assign n1136 = ~n703 & ~n866;
  assign n1137 = n925 & n1136;
  assign n1138 = ~n1135 & ~n1137;
  assign n1139 = ~n1121 & n1138;
  assign n1140 = ~n1133 & n1139;
  assign n1141 = n1106 & ~n1140;
  assign n1142 = ~n703 & n985;
  assign n1143 = n703 & n866;
  assign n1144 = ~n984 & n1143;
  assign n1145 = ~n1142 & ~n1144;
  assign n1146 = ~n1106 & ~n1145;
  assign n1147 = ~n1141 & ~n1146;
  assign n1148 = ~n986 & n1147;
  assign n1149 = n703 & n1107;
  assign n1150 = n925 & n1149;
  assign n1151 = n1148 & ~n1150;
  assign n1152 = n1046 & ~n1151;
  assign n1153 = ~n984 & n1110;
  assign n1154 = ~n925 & n1153;
  assign n1155 = ~n984 & n1136;
  assign n1156 = n925 & n1155;
  assign n1157 = ~n1150 & ~n1156;
  assign n1158 = ~n1154 & n1157;
  assign n1159 = n1106 & ~n1158;
  assign n1160 = ~n1152 & ~n1159;
  assign n1161 = n1131 & n1160;
  assign n1162 = n461 & ~n1161;
  assign n1163 = ~n461 & n1161;
  assign po00 = n1162 | n1163;
  assign n1165 = pi129 & n446;
  assign n1166 = ~pi001 & ~n454;
  assign n1167 = ~pi106 & n454;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~n449 & n1168;
  assign n1170 = pi106 & n449;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = ~n446 & ~n1171;
  assign po01 = n1165 | n1172;
  assign n1174 = pi071 & ~n454;
  assign n1175 = ~pi058 & n454;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = ~n449 & ~n1176;
  assign n1178 = ~pi058 & n449;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = ~n446 & ~n1179;
  assign n1181 = pi130 & n446;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = pi011 & ~n449;
  assign n1184 = ~n454 & n1183;
  assign n1185 = pi112 & ~n449;
  assign n1186 = n454 & n1185;
  assign n1187 = pi112 & n449;
  assign n1188 = ~n1186 & ~n1187;
  assign n1189 = ~n1184 & n1188;
  assign n1190 = ~n446 & ~n1189;
  assign n1191 = pi159 & n446;
  assign po31 = n1190 | n1191;
  assign n1193 = pi258 & ~n481;
  assign n1194 = pi314 & n483;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = pi314 & n470;
  assign n1197 = pi202 & ~n475;
  assign n1198 = ~n1196 & ~n1197;
  assign n1199 = n1195 & n1198;
  assign n1200 = n468 & ~n1199;
  assign n1201 = pi338 & n483;
  assign n1202 = pi282 & ~n481;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = pi338 & n470;
  assign n1205 = pi226 & ~n475;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = n1203 & n1206;
  assign n1208 = ~n468 & ~n1207;
  assign n1209 = ~n1200 & ~n1208;
  assign n1210 = n673 & ~n1209;
  assign n1211 = pi205 & ~n475;
  assign n1212 = pi317 & n470;
  assign n1213 = pi317 & n483;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = pi261 & ~n481;
  assign n1216 = n1214 & ~n1215;
  assign n1217 = ~n1211 & n1216;
  assign n1218 = ~n468 & ~n1217;
  assign n1219 = pi310 & n470;
  assign n1220 = pi254 & ~n481;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = pi310 & n483;
  assign n1223 = pi198 & ~n475;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = n1221 & n1224;
  assign n1226 = n468 & ~n1225;
  assign n1227 = ~n1218 & ~n1226;
  assign n1228 = n650 & ~n1227;
  assign n1229 = ~n1210 & ~n1228;
  assign n1230 = pi287 & ~n481;
  assign n1231 = pi343 & n483;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = pi343 & n470;
  assign n1234 = pi231 & ~n475;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = n1232 & n1235;
  assign n1237 = ~n468 & ~n1236;
  assign n1238 = pi309 & n483;
  assign n1239 = pi253 & ~n481;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = pi197 & ~n475;
  assign n1242 = pi309 & n470;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = n1240 & n1243;
  assign n1245 = n468 & ~n1244;
  assign n1246 = ~n1237 & ~n1245;
  assign n1247 = n678 & ~n1246;
  assign n1248 = pi337 & n470;
  assign n1249 = pi225 & ~n475;
  assign n1250 = ~n1248 & ~n1249;
  assign n1251 = pi281 & ~n481;
  assign n1252 = pi337 & n483;
  assign n1253 = ~n1251 & ~n1252;
  assign n1254 = n1250 & n1253;
  assign n1255 = n468 & ~n1254;
  assign n1256 = pi259 & ~n481;
  assign n1257 = pi315 & n483;
  assign n1258 = ~n1256 & ~n1257;
  assign n1259 = pi315 & n470;
  assign n1260 = pi203 & ~n475;
  assign n1261 = ~n1259 & ~n1260;
  assign n1262 = n1258 & n1261;
  assign n1263 = ~n468 & ~n1262;
  assign n1264 = ~n1255 & ~n1263;
  assign n1265 = n613 & ~n1264;
  assign n1266 = ~n1247 & ~n1265;
  assign n1267 = n1229 & n1266;
  assign n1268 = n468 & ~n1217;
  assign n1269 = ~n468 & ~n1225;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = n684 & ~n1270;
  assign n1272 = pi351 & n483;
  assign n1273 = pi351 & n470;
  assign n1274 = pi295 & ~n481;
  assign n1275 = pi239 & ~n475;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = ~n1273 & n1276;
  assign n1278 = ~n1272 & n1277;
  assign n1279 = n468 & ~n1278;
  assign n1280 = pi302 & ~n481;
  assign n1281 = pi358 & n483;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = pi358 & n470;
  assign n1284 = pi246 & ~n475;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = n1282 & n1285;
  assign n1287 = ~n468 & ~n1286;
  assign n1288 = ~n1279 & ~n1287;
  assign n1289 = n632 & ~n1288;
  assign n1290 = ~n1271 & ~n1289;
  assign n1291 = ~n468 & ~n1278;
  assign n1292 = n468 & ~n1286;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n520 & ~n1293;
  assign n1295 = pi352 & n483;
  assign n1296 = pi296 & ~n481;
  assign n1297 = pi352 & n470;
  assign n1298 = pi240 & ~n475;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = ~n1296 & n1299;
  assign n1301 = ~n1295 & n1300;
  assign n1302 = ~n468 & ~n1301;
  assign n1303 = pi245 & ~n475;
  assign n1304 = pi357 & n470;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = pi301 & ~n481;
  assign n1307 = pi357 & n483;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = n1305 & n1308;
  assign n1310 = n468 & ~n1309;
  assign n1311 = ~n1302 & ~n1310;
  assign n1312 = n606 & ~n1311;
  assign n1313 = pi328 & n470;
  assign n1314 = pi216 & ~n475;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = pi272 & ~n481;
  assign n1317 = pi328 & n483;
  assign n1318 = ~n1316 & ~n1317;
  assign n1319 = n1315 & n1318;
  assign n1320 = n468 & ~n1319;
  assign n1321 = pi324 & n470;
  assign n1322 = pi212 & ~n475;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = pi268 & ~n481;
  assign n1325 = pi324 & n483;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = n1323 & n1326;
  assign n1328 = ~n468 & ~n1327;
  assign n1329 = ~n1320 & ~n1328;
  assign n1330 = n601 & ~n1329;
  assign n1331 = n468 & ~n1301;
  assign n1332 = ~n468 & ~n1309;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = n499 & ~n1333;
  assign n1335 = ~n1330 & ~n1334;
  assign n1336 = ~n1312 & n1335;
  assign n1337 = ~n1294 & n1336;
  assign n1338 = n468 & ~n1207;
  assign n1339 = ~n468 & ~n1199;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = n540 & ~n1340;
  assign n1342 = pi211 & ~n475;
  assign n1343 = pi323 & n470;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = pi267 & ~n481;
  assign n1346 = pi323 & n483;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = n1344 & n1347;
  assign n1349 = n468 & ~n1348;
  assign n1350 = pi329 & n483;
  assign n1351 = pi273 & ~n481;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = pi217 & ~n475;
  assign n1354 = pi329 & n470;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = n1352 & n1355;
  assign n1357 = ~n468 & ~n1356;
  assign n1358 = ~n1349 & ~n1357;
  assign n1359 = n464 & ~n1358;
  assign n1360 = ~n1341 & ~n1359;
  assign n1361 = n468 & ~n1327;
  assign n1362 = ~n468 & ~n1319;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n560 & ~n1363;
  assign n1365 = n468 & ~n1236;
  assign n1366 = ~n468 & ~n1244;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = n579 & ~n1367;
  assign n1369 = ~n1364 & ~n1368;
  assign n1370 = n1360 & n1369;
  assign n1371 = n1337 & n1370;
  assign n1372 = ~n468 & ~n1254;
  assign n1373 = n468 & ~n1262;
  assign n1374 = ~n1372 & ~n1373;
  assign n1375 = n643 & ~n1374;
  assign n1376 = ~n468 & ~n1348;
  assign n1377 = n468 & ~n1356;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = n638 & ~n1378;
  assign n1380 = ~n1375 & ~n1379;
  assign n1381 = n1371 & n1380;
  assign n1382 = n1290 & n1381;
  assign n1383 = n1267 & n1382;
  assign n1384 = po31 & ~n1383;
  assign n1385 = ~po31 & n1383;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = pi196 & ~n475;
  assign n1388 = pi308 & n470;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = pi308 & n483;
  assign n1391 = pi252 & ~n481;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = n1389 & n1392;
  assign n1394 = ~n468 & ~n1393;
  assign n1395 = pi331 & n470;
  assign n1396 = pi219 & ~n475;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = pi275 & ~n481;
  assign n1399 = pi331 & n483;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = n1397 & n1400;
  assign n1402 = n468 & ~n1401;
  assign n1403 = ~n1394 & ~n1402;
  assign n1404 = n678 & ~n1403;
  assign n1405 = pi204 & ~n475;
  assign n1406 = pi316 & n470;
  assign n1407 = ~n1405 & ~n1406;
  assign n1408 = pi260 & ~n481;
  assign n1409 = pi316 & n483;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = n1407 & n1410;
  assign n1412 = n468 & ~n1411;
  assign n1413 = ~n1376 & ~n1412;
  assign n1414 = n632 & ~n1413;
  assign n1415 = ~n1404 & ~n1414;
  assign n1416 = pi303 & ~n481;
  assign n1417 = pi359 & n483;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = pi359 & n470;
  assign n1420 = pi247 & ~n475;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = n1418 & n1421;
  assign n1423 = n468 & ~n1422;
  assign n1424 = ~n1372 & ~n1423;
  assign n1425 = n613 & ~n1424;
  assign n1426 = ~n468 & ~n1422;
  assign n1427 = ~n1255 & ~n1426;
  assign n1428 = n643 & ~n1427;
  assign n1429 = ~n1425 & ~n1428;
  assign n1430 = n1415 & n1429;
  assign n1431 = pi251 & ~n481;
  assign n1432 = pi307 & n483;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = pi195 & ~n475;
  assign n1435 = pi307 & n470;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = n1433 & n1436;
  assign n1438 = n468 & ~n1437;
  assign n1439 = ~n1332 & ~n1438;
  assign n1440 = n684 & ~n1439;
  assign n1441 = ~n468 & ~n1437;
  assign n1442 = ~n1310 & ~n1441;
  assign n1443 = n650 & ~n1442;
  assign n1444 = ~n1440 & ~n1443;
  assign n1445 = pi210 & ~n475;
  assign n1446 = pi322 & n470;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = pi322 & n483;
  assign n1449 = pi266 & ~n481;
  assign n1450 = ~n1448 & ~n1449;
  assign n1451 = n1447 & n1450;
  assign n1452 = ~n468 & ~n1451;
  assign n1453 = ~n1268 & ~n1452;
  assign n1454 = n499 & ~n1453;
  assign n1455 = n1444 & ~n1454;
  assign n1456 = pi350 & n470;
  assign n1457 = pi238 & ~n475;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = pi294 & ~n481;
  assign n1460 = pi350 & n483;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = n1458 & n1461;
  assign n1463 = n468 & ~n1462;
  assign n1464 = ~n1339 & ~n1463;
  assign n1465 = n601 & ~n1464;
  assign n1466 = pi345 & n470;
  assign n1467 = pi233 & ~n475;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = pi345 & n483;
  assign n1470 = pi289 & ~n481;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = n1468 & n1471;
  assign n1473 = n468 & ~n1472;
  assign n1474 = ~n1291 & ~n1473;
  assign n1475 = n464 & ~n1474;
  assign n1476 = ~n1465 & ~n1475;
  assign n1477 = ~n468 & ~n1472;
  assign n1478 = ~n1279 & ~n1477;
  assign n1479 = n638 & ~n1478;
  assign n1480 = n1476 & ~n1479;
  assign n1481 = pi336 & n470;
  assign n1482 = pi224 & ~n475;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = pi280 & ~n481;
  assign n1485 = pi336 & n483;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = n1483 & n1486;
  assign n1488 = n468 & ~n1487;
  assign n1489 = ~n1362 & ~n1488;
  assign n1490 = n673 & ~n1489;
  assign n1491 = ~n468 & ~n1487;
  assign n1492 = ~n1320 & ~n1491;
  assign n1493 = n540 & ~n1492;
  assign n1494 = ~n468 & ~n1462;
  assign n1495 = ~n1200 & ~n1494;
  assign n1496 = n560 & ~n1495;
  assign n1497 = ~n1493 & ~n1496;
  assign n1498 = ~n1490 & n1497;
  assign n1499 = ~n468 & ~n1411;
  assign n1500 = ~n1349 & ~n1499;
  assign n1501 = n520 & ~n1500;
  assign n1502 = n468 & ~n1393;
  assign n1503 = ~n468 & ~n1401;
  assign n1504 = ~n1502 & ~n1503;
  assign n1505 = n579 & ~n1504;
  assign n1506 = ~n1501 & ~n1505;
  assign n1507 = n468 & ~n1451;
  assign n1508 = ~n1218 & ~n1507;
  assign n1509 = n606 & ~n1508;
  assign n1510 = n1506 & ~n1509;
  assign n1511 = n1498 & n1510;
  assign n1512 = n1480 & n1511;
  assign n1513 = n1455 & n1512;
  assign n1514 = n1430 & n1513;
  assign n1515 = pi151 & n446;
  assign n1516 = pi007 & ~n454;
  assign n1517 = pi076 & n454;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n449 & ~n1518;
  assign n1520 = pi076 & n449;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n446 & ~n1521;
  assign po23 = n1515 | n1522;
  assign n1524 = ~n1514 & ~po23;
  assign n1525 = n1514 & po23;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = pi135 & n446;
  assign n1528 = pi108 & ~n446;
  assign n1529 = n449 & n1528;
  assign n1530 = ~n1527 & ~n1529;
  assign n1531 = pi056 & ~n454;
  assign n1532 = pi108 & n454;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n446 & ~n449;
  assign n1535 = ~n1533 & n1534;
  assign po07 = ~n1530 | n1535;
  assign n1537 = ~n1269 & ~n1473;
  assign n1538 = n643 & ~n1537;
  assign n1539 = ~n1438 & ~n1499;
  assign n1540 = n678 & ~n1539;
  assign n1541 = ~n1263 & ~n1502;
  assign n1542 = n650 & ~n1541;
  assign n1543 = ~n1540 & ~n1542;
  assign n1544 = ~n1287 & ~n1507;
  assign n1545 = n560 & ~n1544;
  assign n1546 = ~n1328 & ~n1402;
  assign n1547 = n520 & ~n1546;
  assign n1548 = ~n1545 & ~n1547;
  assign n1549 = pi218 & ~n475;
  assign n1550 = pi330 & n470;
  assign n1551 = pi330 & n483;
  assign n1552 = ~n1550 & ~n1551;
  assign n1553 = pi274 & ~n481;
  assign n1554 = n1552 & ~n1553;
  assign n1555 = ~n1549 & n1554;
  assign n1556 = n468 & ~n1555;
  assign n1557 = ~n1494 & ~n1556;
  assign n1558 = n606 & ~n1557;
  assign n1559 = pi265 & ~n481;
  assign n1560 = pi321 & n483;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = pi321 & n470;
  assign n1563 = pi209 & ~n475;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = n1561 & n1564;
  assign n1566 = n468 & ~n1565;
  assign n1567 = ~n1426 & ~n1566;
  assign n1568 = n464 & ~n1567;
  assign n1569 = ~n1558 & ~n1568;
  assign n1570 = n1548 & n1569;
  assign n1571 = n1543 & n1570;
  assign n1572 = pi344 & n470;
  assign n1573 = pi232 & ~n475;
  assign n1574 = ~n1572 & ~n1573;
  assign n1575 = pi344 & n483;
  assign n1576 = pi288 & ~n481;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = n1574 & n1577;
  assign n1579 = n468 & ~n1578;
  assign n1580 = ~n1491 & ~n1579;
  assign n1581 = n673 & ~n1580;
  assign n1582 = ~n1361 & ~n1503;
  assign n1583 = n632 & ~n1582;
  assign n1584 = ~n1581 & ~n1583;
  assign n1585 = ~n1226 & ~n1477;
  assign n1586 = n613 & ~n1585;
  assign n1587 = n1584 & ~n1586;
  assign n1588 = ~n468 & ~n1565;
  assign n1589 = ~n1423 & ~n1588;
  assign n1590 = n638 & ~n1589;
  assign n1591 = ~n1373 & ~n1394;
  assign n1592 = n684 & ~n1591;
  assign n1593 = ~n1590 & ~n1592;
  assign n1594 = ~n468 & ~n1555;
  assign n1595 = ~n1463 & ~n1594;
  assign n1596 = n499 & ~n1595;
  assign n1597 = ~n1292 & ~n1452;
  assign n1598 = n601 & ~n1597;
  assign n1599 = ~n1596 & ~n1598;
  assign n1600 = ~n1412 & ~n1441;
  assign n1601 = n579 & ~n1600;
  assign n1602 = ~n468 & ~n1578;
  assign n1603 = ~n1488 & ~n1602;
  assign n1604 = n540 & ~n1603;
  assign n1605 = ~n1601 & ~n1604;
  assign n1606 = n1599 & n1605;
  assign n1607 = n1593 & n1606;
  assign n1608 = n1587 & n1607;
  assign n1609 = n1571 & n1608;
  assign n1610 = ~n1538 & n1609;
  assign n1611 = ~po07 & ~n1610;
  assign n1612 = ~n1538 & n1607;
  assign n1613 = n1587 & n1612;
  assign n1614 = n1571 & n1613;
  assign n1615 = po07 & n1614;
  assign n1616 = ~n1611 & ~n1615;
  assign n1617 = pi167 & n446;
  assign n1618 = ~pi019 & ~n454;
  assign n1619 = ~pi104 & n454;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = ~n449 & n1620;
  assign n1622 = pi104 & n449;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = ~n446 & ~n1623;
  assign po39 = n1617 | n1624;
  assign n1626 = ~n1320 & ~n1376;
  assign n1627 = n606 & ~n1626;
  assign n1628 = ~n1279 & ~n1332;
  assign n1629 = n464 & ~n1628;
  assign n1630 = ~n1627 & ~n1629;
  assign n1631 = ~n1349 & ~n1362;
  assign n1632 = n499 & ~n1631;
  assign n1633 = ~n1218 & ~n1245;
  assign n1634 = n540 & ~n1633;
  assign n1635 = ~n1632 & ~n1634;
  assign n1636 = ~n1365 & ~n1394;
  assign n1637 = n643 & ~n1636;
  assign n1638 = ~n1357 & ~n1507;
  assign n1639 = n632 & ~n1638;
  assign n1640 = ~n1637 & ~n1639;
  assign n1641 = ~n1237 & ~n1502;
  assign n1642 = n613 & ~n1641;
  assign n1643 = ~n1255 & ~n1339;
  assign n1644 = n678 & ~n1643;
  assign n1645 = ~n1642 & ~n1644;
  assign n1646 = n1640 & n1645;
  assign n1647 = ~n1208 & ~n1473;
  assign n1648 = n684 & ~n1647;
  assign n1649 = ~n1338 & ~n1477;
  assign n1650 = n650 & ~n1649;
  assign n1651 = ~n1268 & ~n1366;
  assign n1652 = n673 & ~n1651;
  assign n1653 = ~n1291 & ~n1310;
  assign n1654 = n638 & ~n1653;
  assign n1655 = ~n1652 & ~n1654;
  assign n1656 = ~n1650 & n1655;
  assign n1657 = ~n1648 & n1656;
  assign n1658 = n1646 & n1657;
  assign n1659 = ~n1377 & ~n1452;
  assign n1660 = n520 & ~n1659;
  assign n1661 = ~n1302 & ~n1402;
  assign n1662 = n601 & ~n1661;
  assign n1663 = ~n1660 & ~n1662;
  assign n1664 = ~n1331 & ~n1503;
  assign n1665 = n560 & ~n1664;
  assign n1666 = ~n1200 & ~n1372;
  assign n1667 = n579 & ~n1666;
  assign n1668 = ~n1665 & ~n1667;
  assign n1669 = n1663 & n1668;
  assign n1670 = n1658 & n1669;
  assign n1671 = n1635 & n1670;
  assign n1672 = n1630 & n1671;
  assign n1673 = ~po39 & ~n1672;
  assign n1674 = po39 & n1672;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~n1263 & ~n1349;
  assign n1677 = n673 & ~n1676;
  assign n1678 = ~n1269 & ~n1320;
  assign n1679 = n632 & ~n1678;
  assign n1680 = ~n1677 & ~n1679;
  assign n1681 = ~n1332 & ~n1338;
  assign n1682 = n638 & ~n1681;
  assign n1683 = ~n1302 & ~n1365;
  assign n1684 = n678 & ~n1683;
  assign n1685 = ~n1682 & ~n1684;
  assign n1686 = n1680 & n1685;
  assign n1687 = ~n1291 & ~n1579;
  assign n1688 = n650 & ~n1687;
  assign n1689 = ~n1200 & ~n1328;
  assign n1690 = n613 & ~n1689;
  assign n1691 = ~n1339 & ~n1361;
  assign n1692 = n643 & ~n1691;
  assign n1693 = ~n1690 & ~n1692;
  assign n1694 = ~n1279 & ~n1602;
  assign n1695 = n684 & ~n1694;
  assign n1696 = n1693 & ~n1695;
  assign n1697 = ~n1688 & n1696;
  assign n1698 = n1686 & n1697;
  assign n1699 = ~n1208 & ~n1310;
  assign n1700 = n464 & ~n1699;
  assign n1701 = ~n1237 & ~n1331;
  assign n1702 = n579 & ~n1701;
  assign n1703 = ~n1700 & ~n1702;
  assign n1704 = ~n1255 & ~n1287;
  assign n1705 = n601 & ~n1704;
  assign n1706 = ~n1245 & ~n1357;
  assign n1707 = n606 & ~n1706;
  assign n1708 = ~n1705 & ~n1707;
  assign n1709 = n1703 & n1708;
  assign n1710 = ~n1226 & ~n1362;
  assign n1711 = n520 & ~n1710;
  assign n1712 = ~n1373 & ~n1376;
  assign n1713 = n540 & ~n1712;
  assign n1714 = ~n1711 & ~n1713;
  assign n1715 = ~n1292 & ~n1372;
  assign n1716 = n560 & ~n1715;
  assign n1717 = ~n1366 & ~n1377;
  assign n1718 = n499 & ~n1717;
  assign n1719 = ~n1716 & ~n1718;
  assign n1720 = n1714 & n1719;
  assign n1721 = n1709 & n1720;
  assign n1722 = n1698 & n1721;
  assign n1723 = pi052 & ~n454;
  assign n1724 = pi086 & n454;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = ~n449 & ~n1725;
  assign n1727 = pi086 & n449;
  assign n1728 = ~n1726 & ~n1727;
  assign n1729 = ~n446 & ~n1728;
  assign n1730 = pi185 & n446;
  assign po57 = n1729 | n1730;
  assign n1732 = ~n1722 & ~po57;
  assign n1733 = n1722 & po57;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = n1675 & n1734;
  assign n1736 = ~n1675 & ~n1734;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1616 & ~n1737;
  assign n1739 = pi017 & ~n454;
  assign n1740 = pi114 & n454;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = n1534 & ~n1741;
  assign n1743 = pi143 & n446;
  assign n1744 = pi114 & ~n446;
  assign n1745 = n449 & n1744;
  assign n1746 = ~n1743 & ~n1745;
  assign po15 = n1742 | ~n1746;
  assign n1748 = ~n1503 & ~n1507;
  assign n1749 = n678 & ~n1748;
  assign n1750 = ~n1291 & ~n1423;
  assign n1751 = n673 & ~n1750;
  assign n1752 = ~n1749 & ~n1751;
  assign n1753 = ~n1372 & ~n1412;
  assign n1754 = n601 & ~n1753;
  assign n1755 = ~n1394 & ~n1473;
  assign n1756 = n606 & ~n1755;
  assign n1757 = ~n1754 & ~n1756;
  assign n1758 = ~n1200 & ~n1441;
  assign n1759 = n520 & ~n1758;
  assign n1760 = ~n1218 & ~n1488;
  assign n1761 = n464 & ~n1760;
  assign n1762 = ~n1759 & ~n1761;
  assign n1763 = n1757 & n1762;
  assign n1764 = n1752 & n1763;
  assign n1765 = ~n1376 & ~n1556;
  assign n1766 = n684 & ~n1765;
  assign n1767 = ~n1268 & ~n1491;
  assign n1768 = n638 & ~n1767;
  assign n1769 = ~n1766 & ~n1768;
  assign n1770 = ~n1320 & ~n1494;
  assign n1771 = n643 & ~n1770;
  assign n1772 = ~n1339 & ~n1438;
  assign n1773 = n632 & ~n1772;
  assign n1774 = ~n1771 & ~n1773;
  assign n1775 = n1769 & n1774;
  assign n1776 = n1764 & n1775;
  assign n1777 = ~n1255 & ~n1499;
  assign n1778 = n560 & ~n1777;
  assign n1779 = ~n1402 & ~n1452;
  assign n1780 = n579 & ~n1779;
  assign n1781 = ~n1778 & ~n1780;
  assign n1782 = ~n1279 & ~n1426;
  assign n1783 = n540 & ~n1782;
  assign n1784 = ~n1477 & ~n1502;
  assign n1785 = n499 & ~n1784;
  assign n1786 = ~n1783 & ~n1785;
  assign n1787 = n1781 & n1786;
  assign n1788 = ~n1362 & ~n1463;
  assign n1789 = n613 & ~n1788;
  assign n1790 = ~n1349 & ~n1594;
  assign n1791 = n650 & ~n1790;
  assign n1792 = ~n1789 & ~n1791;
  assign n1793 = n1787 & n1792;
  assign n1794 = n1776 & n1793;
  assign n1795 = po15 & ~n1794;
  assign n1796 = n1775 & n1793;
  assign n1797 = n1764 & n1796;
  assign n1798 = ~po15 & n1797;
  assign n1799 = ~n1795 & ~n1798;
  assign n1800 = n1736 & n1799;
  assign n1801 = ~n1738 & ~n1800;
  assign n1802 = ~n1526 & ~n1801;
  assign n1803 = n1386 & n1802;
  assign n1804 = ~n1616 & n1799;
  assign n1805 = n1735 & n1804;
  assign n1806 = ~n1734 & ~n1799;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = n1616 & ~n1734;
  assign n1809 = n1807 & ~n1808;
  assign n1810 = n1526 & ~n1809;
  assign n1811 = n1616 & ~n1799;
  assign n1812 = n1675 & n1811;
  assign n1813 = n1616 & ~n1675;
  assign n1814 = n1734 & n1813;
  assign n1815 = n1799 & n1814;
  assign n1816 = ~n1812 & ~n1815;
  assign n1817 = ~n1526 & n1734;
  assign n1818 = ~n1799 & n1817;
  assign n1819 = ~n1526 & n1804;
  assign n1820 = ~n1734 & n1819;
  assign n1821 = ~n1818 & ~n1820;
  assign n1822 = n1816 & n1821;
  assign n1823 = ~n1810 & n1822;
  assign n1824 = ~n1386 & ~n1823;
  assign n1825 = n1675 & ~n1734;
  assign n1826 = ~n1616 & n1825;
  assign n1827 = ~n1799 & n1826;
  assign n1828 = ~n1616 & ~n1675;
  assign n1829 = n1734 & n1828;
  assign n1830 = n1616 & n1735;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = n1526 & ~n1831;
  assign n1833 = ~n1827 & ~n1832;
  assign n1834 = ~n1799 & n1814;
  assign n1835 = n1833 & ~n1834;
  assign n1836 = n1386 & ~n1835;
  assign n1837 = n1616 & n1736;
  assign n1838 = ~n1799 & n1837;
  assign n1839 = n1616 & n1825;
  assign n1840 = n1799 & n1839;
  assign n1841 = ~n1838 & ~n1840;
  assign n1842 = n1526 & ~n1841;
  assign n1843 = ~n1836 & ~n1842;
  assign n1844 = ~n1824 & n1843;
  assign n1845 = ~n1803 & n1844;
  assign n1846 = ~n1182 & n1845;
  assign n1847 = n1182 & ~n1845;
  assign po02 = n1846 | n1847;
  assign n1849 = pi132 & n446;
  assign n1850 = pi127 & ~n454;
  assign n1851 = pi046 & n454;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~n449 & ~n1852;
  assign n1854 = pi046 & n449;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = ~n446 & ~n1855;
  assign n1857 = ~n1849 & ~n1856;
  assign n1858 = n1799 & n1830;
  assign n1859 = ~n1799 & n1839;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1526 & ~n1860;
  assign n1862 = ~n1616 & n1675;
  assign n1863 = ~n1675 & n1811;
  assign n1864 = ~n1862 & ~n1863;
  assign n1865 = ~n1837 & n1864;
  assign n1866 = n1526 & ~n1865;
  assign n1867 = ~n1828 & ~n1839;
  assign n1868 = ~n1526 & ~n1867;
  assign n1869 = ~n1866 & ~n1868;
  assign n1870 = n1738 & ~n1799;
  assign n1871 = ~n1858 & ~n1870;
  assign n1872 = n1869 & n1871;
  assign n1873 = n1386 & ~n1872;
  assign n1874 = ~n1826 & ~n1829;
  assign n1875 = ~n1830 & ~n1837;
  assign n1876 = n1874 & n1875;
  assign n1877 = ~n1799 & ~n1876;
  assign n1878 = ~n1815 & ~n1877;
  assign n1879 = n1526 & n1799;
  assign n1880 = ~n1867 & n1879;
  assign n1881 = n1878 & ~n1880;
  assign n1882 = ~n1386 & ~n1881;
  assign n1883 = ~n1873 & ~n1882;
  assign n1884 = ~n1861 & n1883;
  assign n1885 = ~n1857 & n1884;
  assign n1886 = n1857 & ~n1884;
  assign po04 = n1885 | n1886;
  assign n1888 = pi047 & ~n454;
  assign n1889 = pi125 & n454;
  assign n1890 = ~n1888 & ~n1889;
  assign n1891 = ~n449 & ~n1890;
  assign n1892 = pi125 & n449;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = ~n446 & ~n1893;
  assign n1895 = pi133 & n446;
  assign po05 = n1894 | n1895;
  assign n1897 = pi134 & n446;
  assign n1898 = pi055 & n449;
  assign n1899 = pi097 & ~n454;
  assign n1900 = pi055 & n454;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = ~n449 & ~n1901;
  assign n1903 = ~n1898 & ~n1902;
  assign n1904 = ~n446 & ~n1903;
  assign n1905 = ~n1897 & ~n1904;
  assign n1906 = ~n1291 & ~n1556;
  assign n1907 = n601 & ~n1906;
  assign n1908 = ~n1320 & ~n1588;
  assign n1909 = n520 & ~n1908;
  assign n1910 = ~n1907 & ~n1909;
  assign n1911 = ~n1463 & ~n1503;
  assign n1912 = n464 & ~n1911;
  assign n1913 = ~n1473 & ~n1491;
  assign n1914 = n579 & ~n1913;
  assign n1915 = ~n1912 & ~n1914;
  assign n1916 = n1910 & n1915;
  assign n1917 = ~n1362 & ~n1566;
  assign n1918 = n632 & ~n1917;
  assign n1919 = ~n1255 & ~n1602;
  assign n1920 = n650 & ~n1919;
  assign n1921 = ~n1918 & ~n1920;
  assign n1922 = ~n1372 & ~n1579;
  assign n1923 = n684 & ~n1922;
  assign n1924 = ~n1402 & ~n1494;
  assign n1925 = n638 & ~n1924;
  assign n1926 = ~n1923 & ~n1925;
  assign n1927 = ~n1394 & ~n1412;
  assign n1928 = n673 & ~n1927;
  assign n1929 = ~n1268 & ~n1441;
  assign n1930 = n643 & ~n1929;
  assign n1931 = ~n1928 & ~n1930;
  assign n1932 = n1926 & n1931;
  assign n1933 = ~n1218 & ~n1438;
  assign n1934 = n613 & ~n1933;
  assign n1935 = ~n1477 & ~n1488;
  assign n1936 = n678 & ~n1935;
  assign n1937 = ~n1934 & ~n1936;
  assign n1938 = n1932 & n1937;
  assign n1939 = n1921 & n1938;
  assign n1940 = ~n1279 & ~n1594;
  assign n1941 = n560 & ~n1940;
  assign n1942 = ~n1423 & ~n1452;
  assign n1943 = n606 & ~n1942;
  assign n1944 = ~n1941 & ~n1943;
  assign n1945 = ~n1499 & ~n1502;
  assign n1946 = n540 & ~n1945;
  assign n1947 = ~n1426 & ~n1507;
  assign n1948 = n499 & ~n1947;
  assign n1949 = ~n1946 & ~n1948;
  assign n1950 = n1944 & n1949;
  assign n1951 = n1939 & n1950;
  assign n1952 = n1916 & n1951;
  assign n1953 = po61 & n1952;
  assign n1954 = ~po61 & ~n1952;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = ~n1310 & ~n1366;
  assign n1957 = n678 & ~n1956;
  assign n1958 = ~n1208 & ~n1320;
  assign n1959 = n613 & ~n1958;
  assign n1960 = ~n1338 & ~n1362;
  assign n1961 = n643 & ~n1960;
  assign n1962 = ~n1959 & ~n1961;
  assign n1963 = ~n1292 & ~n1394;
  assign n1964 = n650 & ~n1963;
  assign n1965 = n1962 & ~n1964;
  assign n1966 = ~n1957 & n1965;
  assign n1967 = ~n1372 & ~n1377;
  assign n1968 = n540 & ~n1967;
  assign n1969 = ~n1200 & ~n1302;
  assign n1970 = n464 & ~n1969;
  assign n1971 = ~n1968 & ~n1970;
  assign n1972 = ~n1291 & ~n1373;
  assign n1973 = n560 & ~n1972;
  assign n1974 = ~n1365 & ~n1376;
  assign n1975 = n499 & ~n1974;
  assign n1976 = ~n1973 & ~n1975;
  assign n1977 = n1971 & n1976;
  assign n1978 = ~n1263 & ~n1279;
  assign n1979 = n601 & ~n1978;
  assign n1980 = ~n1245 & ~n1332;
  assign n1981 = n579 & ~n1980;
  assign n1982 = ~n1979 & ~n1981;
  assign n1983 = ~n1237 & ~n1349;
  assign n1984 = n606 & ~n1983;
  assign n1985 = n1982 & ~n1984;
  assign n1986 = ~n1218 & ~n1361;
  assign n1987 = n520 & ~n1986;
  assign n1988 = ~n1287 & ~n1502;
  assign n1989 = n684 & ~n1988;
  assign n1990 = ~n1268 & ~n1328;
  assign n1991 = n632 & ~n1990;
  assign n1992 = ~n1989 & ~n1991;
  assign n1993 = ~n1987 & n1992;
  assign n1994 = ~n1255 & ~n1357;
  assign n1995 = n673 & ~n1994;
  assign n1996 = ~n1331 & ~n1339;
  assign n1997 = n638 & ~n1996;
  assign n1998 = ~n1995 & ~n1997;
  assign n1999 = n1993 & n1998;
  assign n2000 = n1985 & n1999;
  assign n2001 = n1977 & n2000;
  assign n2002 = n1966 & n2001;
  assign n2003 = pi157 & n446;
  assign n2004 = pi121 & ~n446;
  assign n2005 = n449 & n2004;
  assign n2006 = ~n2003 & ~n2005;
  assign n2007 = pi034 & ~n454;
  assign n2008 = pi121 & n454;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = n1534 & ~n2009;
  assign po29 = ~n2006 | n2010;
  assign n2012 = ~n2002 & ~po29;
  assign n2013 = n2002 & po29;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = pi173 & n446;
  assign n2016 = pi123 & n454;
  assign n2017 = pi016 & ~n454;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = ~n449 & ~n2018;
  assign n2020 = pi123 & n449;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = ~n446 & ~n2021;
  assign po45 = n2015 | n2022;
  assign n2024 = ~n1287 & ~n1349;
  assign n2025 = n613 & ~n2024;
  assign n2026 = ~n1331 & ~n1357;
  assign n2027 = n678 & ~n2026;
  assign n2028 = ~n1292 & ~n1376;
  assign n2029 = n643 & ~n2028;
  assign n2030 = ~n2027 & ~n2029;
  assign n2031 = n632 & ~n1919;
  assign n2032 = n2030 & ~n2031;
  assign n2033 = ~n2025 & n2032;
  assign n2034 = ~n1208 & ~n1365;
  assign n2035 = n606 & ~n2034;
  assign n2036 = ~n1302 & ~n1377;
  assign n2037 = n579 & ~n2036;
  assign n2038 = ~n2035 & ~n2037;
  assign n2039 = ~n1366 & ~n1373;
  assign n2040 = n638 & ~n2039;
  assign n2041 = n2038 & ~n2040;
  assign n2042 = n520 & ~n1922;
  assign n2043 = n684 & ~n1908;
  assign n2044 = n650 & ~n1917;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = ~n2042 & n2045;
  assign n2047 = ~n1200 & ~n1269;
  assign n2048 = n601 & ~n2047;
  assign n2049 = ~n1237 & ~n1338;
  assign n2050 = n499 & ~n2049;
  assign n2051 = ~n1226 & ~n1339;
  assign n2052 = n560 & ~n2051;
  assign n2053 = ~n2050 & ~n2052;
  assign n2054 = ~n2048 & n2053;
  assign n2055 = n2046 & n2054;
  assign n2056 = ~n1332 & ~n1361;
  assign n2057 = n540 & ~n2056;
  assign n2058 = ~n1245 & ~n1263;
  assign n2059 = n464 & ~n2058;
  assign n2060 = ~n2057 & ~n2059;
  assign n2061 = ~n1310 & ~n1328;
  assign n2062 = n673 & ~n2061;
  assign n2063 = n2060 & ~n2062;
  assign n2064 = n2055 & n2063;
  assign n2065 = n2041 & n2064;
  assign n2066 = n2033 & n2065;
  assign n2067 = po45 & ~n2066;
  assign n2068 = ~po45 & n2066;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = pi165 & n446;
  assign n2071 = ~pi023 & ~n454;
  assign n2072 = ~pi105 & n454;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n449 & n2073;
  assign n2075 = pi105 & n449;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = ~n446 & ~n2076;
  assign po37 = n2070 | n2077;
  assign n2079 = ~n1349 & ~n1503;
  assign n2080 = n540 & ~n2079;
  assign n2081 = ~n1218 & ~n1255;
  assign n2082 = n499 & ~n2081;
  assign n2083 = ~n2080 & ~n2082;
  assign n2084 = ~n1339 & ~n1502;
  assign n2085 = n464 & ~n2084;
  assign n2086 = ~n1291 & ~n1320;
  assign n2087 = n579 & ~n2086;
  assign n2088 = ~n2085 & ~n2087;
  assign n2089 = ~n1310 & ~n1452;
  assign n2090 = n643 & ~n2089;
  assign n2091 = ~n1237 & ~n1488;
  assign n2092 = n632 & ~n2091;
  assign n2093 = ~n2090 & ~n2092;
  assign n2094 = ~n1376 & ~n1402;
  assign n2095 = n673 & ~n2094;
  assign n2096 = ~n1332 & ~n1507;
  assign n2097 = n613 & ~n2096;
  assign n2098 = ~n2095 & ~n2097;
  assign n2099 = n2093 & n2098;
  assign n2100 = ~n1331 & ~n1426;
  assign n2101 = n650 & ~n2100;
  assign n2102 = ~n1279 & ~n1362;
  assign n2103 = n678 & ~n2102;
  assign n2104 = ~n1200 & ~n1394;
  assign n2105 = n638 & ~n2104;
  assign n2106 = ~n2103 & ~n2105;
  assign n2107 = ~n1302 & ~n1423;
  assign n2108 = n684 & ~n2107;
  assign n2109 = n2106 & ~n2108;
  assign n2110 = ~n2101 & n2109;
  assign n2111 = n2099 & n2110;
  assign n2112 = ~n1365 & ~n1491;
  assign n2113 = n520 & ~n2112;
  assign n2114 = ~n1366 & ~n1473;
  assign n2115 = n601 & ~n2114;
  assign n2116 = ~n2113 & ~n2115;
  assign n2117 = ~n1268 & ~n1372;
  assign n2118 = n606 & ~n2117;
  assign n2119 = ~n1245 & ~n1477;
  assign n2120 = n560 & ~n2119;
  assign n2121 = ~n2118 & ~n2120;
  assign n2122 = n2116 & n2121;
  assign n2123 = n2111 & n2122;
  assign n2124 = n2088 & n2123;
  assign n2125 = n2083 & n2124;
  assign n2126 = po37 & n2125;
  assign n2127 = ~po37 & ~n2125;
  assign n2128 = ~n2126 & ~n2127;
  assign n2129 = ~n2069 & ~n2128;
  assign n2130 = ~n2014 & n2129;
  assign n2131 = ~n1423 & ~n1441;
  assign n2132 = n499 & ~n2131;
  assign n2133 = ~n1412 & ~n1494;
  assign n2134 = n678 & ~n2133;
  assign n2135 = n650 & ~n1990;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = ~n1488 & ~n1594;
  assign n2138 = n638 & ~n2137;
  assign n2139 = ~n1477 & ~n1566;
  assign n2140 = n673 & ~n2139;
  assign n2141 = ~n2138 & ~n2140;
  assign n2142 = n2136 & n2141;
  assign n2143 = ~n2132 & n2142;
  assign n2144 = ~n1473 & ~n1588;
  assign n2145 = n540 & ~n2144;
  assign n2146 = ~n1269 & ~n1402;
  assign n2147 = n560 & ~n2146;
  assign n2148 = ~n2145 & ~n2147;
  assign n2149 = ~n1226 & ~n1503;
  assign n2150 = n601 & ~n2149;
  assign n2151 = n2148 & ~n2150;
  assign n2152 = ~n1426 & ~n1438;
  assign n2153 = n606 & ~n2152;
  assign n2154 = n520 & ~n1988;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = ~n1491 & ~n1556;
  assign n2157 = n464 & ~n2156;
  assign n2158 = n2155 & ~n2157;
  assign n2159 = n632 & ~n1963;
  assign n2160 = ~n1452 & ~n1579;
  assign n2161 = n613 & ~n2160;
  assign n2162 = ~n1507 & ~n1602;
  assign n2163 = n643 & ~n2162;
  assign n2164 = ~n2161 & ~n2163;
  assign n2165 = n684 & ~n1986;
  assign n2166 = n2164 & ~n2165;
  assign n2167 = ~n2159 & n2166;
  assign n2168 = ~n1463 & ~n1499;
  assign n2169 = n579 & ~n2168;
  assign n2170 = n2167 & ~n2169;
  assign n2171 = n2158 & n2170;
  assign n2172 = n2151 & n2171;
  assign n2173 = n2143 & n2172;
  assign n2174 = po03 & n2173;
  assign n2175 = ~po03 & ~n2173;
  assign n2176 = ~n2174 & ~n2175;
  assign n2177 = n2014 & ~n2176;
  assign n2178 = n2128 & n2177;
  assign n2179 = ~n2069 & n2178;
  assign n2180 = ~n2130 & ~n2179;
  assign n2181 = ~n1218 & ~n1349;
  assign n2182 = n638 & ~n2181;
  assign n2183 = ~n1332 & ~n1502;
  assign n2184 = n673 & ~n2183;
  assign n2185 = ~n2182 & ~n2184;
  assign n2186 = ~n1357 & ~n1488;
  assign n2187 = n684 & ~n2186;
  assign n2188 = n2185 & ~n2187;
  assign n2189 = ~n1268 & ~n1376;
  assign n2190 = n464 & ~n2189;
  assign n2191 = n2188 & ~n2190;
  assign n2192 = ~n1200 & ~n1291;
  assign n2193 = n499 & ~n2192;
  assign n2194 = ~n1320 & ~n1372;
  assign n2195 = n678 & ~n2194;
  assign n2196 = ~n1377 & ~n1491;
  assign n2197 = n650 & ~n2196;
  assign n2198 = ~n2195 & ~n2197;
  assign n2199 = ~n1302 & ~n1473;
  assign n2200 = n632 & ~n2199;
  assign n2201 = ~n1366 & ~n1402;
  assign n2202 = n613 & ~n2201;
  assign n2203 = ~n1245 & ~n1503;
  assign n2204 = n643 & ~n2203;
  assign n2205 = ~n2202 & ~n2204;
  assign n2206 = ~n2200 & n2205;
  assign n2207 = n2198 & n2206;
  assign n2208 = ~n2193 & n2207;
  assign n2209 = ~n1331 & ~n1477;
  assign n2210 = n520 & ~n2209;
  assign n2211 = ~n1237 & ~n1507;
  assign n2212 = n601 & ~n2211;
  assign n2213 = ~n2210 & ~n2212;
  assign n2214 = n2208 & n2213;
  assign n2215 = ~n1365 & ~n1452;
  assign n2216 = n560 & ~n2215;
  assign n2217 = ~n1255 & ~n1362;
  assign n2218 = n579 & ~n2217;
  assign n2219 = ~n2216 & ~n2218;
  assign n2220 = ~n1279 & ~n1339;
  assign n2221 = n606 & ~n2220;
  assign n2222 = ~n1310 & ~n1394;
  assign n2223 = n540 & ~n2222;
  assign n2224 = ~n2221 & ~n2223;
  assign n2225 = n2219 & n2224;
  assign n2226 = n2214 & n2225;
  assign n2227 = n2191 & n2226;
  assign n2228 = pi009 & ~n449;
  assign n2229 = ~n454 & n2228;
  assign n2230 = pi080 & ~n449;
  assign n2231 = n454 & n2230;
  assign n2232 = pi080 & n449;
  assign n2233 = ~n2231 & ~n2232;
  assign n2234 = ~n2229 & n2233;
  assign n2235 = ~n446 & ~n2234;
  assign n2236 = pi181 & n446;
  assign po53 = n2235 | n2236;
  assign n2238 = ~n2227 & ~po53;
  assign n2239 = n2227 & po53;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = ~po03 & n2173;
  assign n2242 = po03 & ~n2173;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = ~n2014 & ~n2243;
  assign n2245 = n2128 & n2244;
  assign n2246 = n2069 & n2128;
  assign n2247 = ~n2243 & n2246;
  assign n2248 = ~n2014 & n2246;
  assign n2249 = ~n2247 & ~n2248;
  assign n2250 = ~n2245 & n2249;
  assign n2251 = ~n2240 & ~n2250;
  assign n2252 = n2180 & ~n2251;
  assign n2253 = n1955 & ~n2252;
  assign n2254 = n2069 & n2178;
  assign n2255 = ~n2128 & n2177;
  assign n2256 = ~n2069 & n2255;
  assign n2257 = ~n2014 & ~n2176;
  assign n2258 = n2069 & n2257;
  assign n2259 = ~n2256 & ~n2258;
  assign n2260 = n2240 & ~n2259;
  assign n2261 = ~n2069 & n2128;
  assign n2262 = ~n2243 & n2261;
  assign n2263 = n2014 & n2262;
  assign n2264 = n2069 & n2245;
  assign n2265 = ~n2263 & ~n2264;
  assign n2266 = n2069 & n2177;
  assign n2267 = n2014 & ~n2243;
  assign n2268 = ~n2128 & n2267;
  assign n2269 = ~n2266 & ~n2268;
  assign n2270 = ~n2240 & ~n2269;
  assign n2271 = n2265 & ~n2270;
  assign n2272 = ~n2260 & n2271;
  assign n2273 = ~n2254 & n2272;
  assign n2274 = ~n1955 & ~n2273;
  assign n2275 = ~n2069 & ~n2240;
  assign n2276 = n2178 & n2275;
  assign n2277 = n2257 & n2275;
  assign n2278 = ~n2128 & n2277;
  assign n2279 = ~n2276 & ~n2278;
  assign n2280 = n2129 & ~n2243;
  assign n2281 = ~n2014 & n2280;
  assign n2282 = ~n2263 & ~n2281;
  assign n2283 = n2128 & n2257;
  assign n2284 = ~n2069 & n2283;
  assign n2285 = n2282 & ~n2284;
  assign n2286 = n2240 & ~n2285;
  assign n2287 = n2014 & n2069;
  assign n2288 = ~n2128 & n2287;
  assign n2289 = ~n2128 & ~n2243;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = n1955 & ~n2290;
  assign n2292 = n2240 & n2291;
  assign n2293 = ~n2286 & ~n2292;
  assign n2294 = n2279 & n2293;
  assign n2295 = ~n2274 & n2294;
  assign n2296 = ~n2253 & n2295;
  assign n2297 = ~n1905 & n2296;
  assign n2298 = n1905 & ~n2296;
  assign po06 = n2297 | n2298;
  assign n2300 = pi136 & n446;
  assign n2301 = pi035 & n449;
  assign n2302 = pi088 & ~n454;
  assign n2303 = pi035 & n454;
  assign n2304 = ~n2302 & ~n2303;
  assign n2305 = ~n449 & ~n2304;
  assign n2306 = ~n2301 & ~n2305;
  assign n2307 = ~n446 & ~n2306;
  assign n2308 = ~n2300 & ~n2307;
  assign n2309 = ~n1955 & ~n2240;
  assign n2310 = ~n2128 & n2243;
  assign n2311 = ~n2130 & ~n2310;
  assign n2312 = n2309 & ~n2311;
  assign n2313 = ~n2240 & n2255;
  assign n2314 = n2069 & n2313;
  assign n2315 = n2069 & n2283;
  assign n2316 = n2246 & n2267;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = ~n2240 & ~n2317;
  assign n2319 = ~n2314 & ~n2318;
  assign n2320 = ~n2264 & ~n2288;
  assign n2321 = ~n2069 & n2240;
  assign n2322 = n2128 & n2321;
  assign n2323 = ~n2244 & n2322;
  assign n2324 = n2128 & n2240;
  assign n2325 = n2243 & n2324;
  assign n2326 = n2014 & n2325;
  assign n2327 = ~n2323 & ~n2326;
  assign n2328 = n2320 & n2327;
  assign n2329 = ~n1955 & ~n2328;
  assign n2330 = n2240 & n2264;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = n2319 & n2331;
  assign n2333 = ~n2312 & n2332;
  assign n2334 = n2240 & n2244;
  assign n2335 = ~n2069 & n2334;
  assign n2336 = ~n2069 & n2245;
  assign n2337 = ~n2128 & n2244;
  assign n2338 = n2069 & n2337;
  assign n2339 = ~n2069 & n2267;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = ~n2240 & ~n2340;
  assign n2342 = ~n2336 & ~n2341;
  assign n2343 = ~n2179 & ~n2315;
  assign n2344 = ~n2128 & n2257;
  assign n2345 = n2240 & n2344;
  assign n2346 = n2343 & ~n2345;
  assign n2347 = n2342 & n2346;
  assign n2348 = ~n2335 & n2347;
  assign n2349 = n1955 & ~n2348;
  assign n2350 = n2333 & ~n2349;
  assign n2351 = n2069 & n2240;
  assign n2352 = n2268 & n2351;
  assign n2353 = n2350 & ~n2352;
  assign n2354 = ~n2308 & n2353;
  assign n2355 = n2308 & ~n2353;
  assign po08 = n2354 | n2355;
  assign n2357 = pi137 & n446;
  assign n2358 = pi027 & ~n454;
  assign n2359 = pi099 & n454;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~n449 & ~n2360;
  assign n2362 = pi099 & n449;
  assign n2363 = ~n2361 & ~n2362;
  assign n2364 = ~n446 & ~n2363;
  assign po09 = n2357 | n2364;
  assign n2366 = pi138 & n446;
  assign n2367 = ~pi118 & ~n454;
  assign n2368 = ~pi048 & n454;
  assign n2369 = ~n2367 & ~n2368;
  assign n2370 = ~n449 & ~n2369;
  assign n2371 = ~pi048 & n449;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~n446 & ~n2372;
  assign n2374 = ~n2366 & ~n2373;
  assign n2375 = pi183 & n446;
  assign n2376 = pi109 & ~n446;
  assign n2377 = n449 & n2376;
  assign n2378 = ~n2375 & ~n2377;
  assign n2379 = pi005 & ~n454;
  assign n2380 = pi109 & n454;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = n1534 & ~n2381;
  assign po55 = ~n2378 | n2382;
  assign n2384 = ~n1579 & ~n1588;
  assign n2385 = n678 & ~n2384;
  assign n2386 = n632 & ~n2196;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = ~n1287 & ~n1438;
  assign n2389 = n638 & ~n2388;
  assign n2390 = ~n1361 & ~n1499;
  assign n2391 = n673 & ~n2390;
  assign n2392 = ~n2389 & ~n2391;
  assign n2393 = n2387 & n2392;
  assign n2394 = n520 & ~n2186;
  assign n2395 = ~n1269 & ~n1556;
  assign n2396 = n499 & ~n2395;
  assign n2397 = ~n2394 & ~n2396;
  assign n2398 = ~n1338 & ~n1426;
  assign n2399 = n601 & ~n2398;
  assign n2400 = ~n1292 & ~n1441;
  assign n2401 = n464 & ~n2400;
  assign n2402 = ~n2399 & ~n2401;
  assign n2403 = n2397 & n2402;
  assign n2404 = ~n1328 & ~n1412;
  assign n2405 = n540 & ~n2404;
  assign n2406 = ~n1208 & ~n1423;
  assign n2407 = n560 & ~n2406;
  assign n2408 = ~n2405 & ~n2407;
  assign n2409 = ~n1226 & ~n1594;
  assign n2410 = n606 & ~n2409;
  assign n2411 = ~n1566 & ~n1602;
  assign n2412 = n579 & ~n2411;
  assign n2413 = ~n2410 & ~n2412;
  assign n2414 = n2408 & n2413;
  assign n2415 = ~n1263 & ~n1463;
  assign n2416 = n643 & ~n2415;
  assign n2417 = ~n1373 & ~n1494;
  assign n2418 = n613 & ~n2417;
  assign n2419 = ~n2416 & ~n2418;
  assign n2420 = n684 & ~n2209;
  assign n2421 = n650 & ~n2199;
  assign n2422 = ~n2420 & ~n2421;
  assign n2423 = n2419 & n2422;
  assign n2424 = n2414 & n2423;
  assign n2425 = n2403 & n2424;
  assign n2426 = n2393 & n2425;
  assign n2427 = ~po55 & ~n2426;
  assign n2428 = po55 & n2426;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = n520 & ~n1694;
  assign n2431 = ~n1463 & ~n1477;
  assign n2432 = n606 & ~n2431;
  assign n2433 = ~n2430 & ~n2432;
  assign n2434 = ~n1218 & ~n1566;
  assign n2435 = n601 & ~n2434;
  assign n2436 = n2433 & ~n2435;
  assign n2437 = ~n1402 & ~n1441;
  assign n2438 = n540 & ~n2437;
  assign n2439 = ~n1499 & ~n1507;
  assign n2440 = n638 & ~n2439;
  assign n2441 = ~n1423 & ~n1491;
  assign n2442 = n678 & ~n2441;
  assign n2443 = ~n2440 & ~n2442;
  assign n2444 = ~n2438 & n2443;
  assign n2445 = ~n1473 & ~n1494;
  assign n2446 = n499 & ~n2445;
  assign n2447 = n684 & ~n1710;
  assign n2448 = n632 & ~n1687;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = ~n1268 & ~n1588;
  assign n2451 = n560 & ~n2450;
  assign n2452 = n2449 & ~n2451;
  assign n2453 = ~n2446 & n2452;
  assign n2454 = ~n1394 & ~n1556;
  assign n2455 = n613 & ~n2454;
  assign n2456 = ~n1502 & ~n1594;
  assign n2457 = n643 & ~n2456;
  assign n2458 = ~n2455 & ~n2457;
  assign n2459 = ~n1438 & ~n1503;
  assign n2460 = n673 & ~n2459;
  assign n2461 = n650 & ~n1678;
  assign n2462 = ~n2460 & ~n2461;
  assign n2463 = n2458 & n2462;
  assign n2464 = ~n1426 & ~n1488;
  assign n2465 = n579 & ~n2464;
  assign n2466 = ~n1412 & ~n1452;
  assign n2467 = n464 & ~n2466;
  assign n2468 = ~n2465 & ~n2467;
  assign n2469 = n2463 & n2468;
  assign n2470 = n2453 & n2469;
  assign n2471 = n2444 & n2470;
  assign n2472 = n2436 & n2471;
  assign n2473 = ~po39 & n2472;
  assign n2474 = po39 & ~n2472;
  assign n2475 = ~n2473 & ~n2474;
  assign n2476 = ~n1310 & ~n1376;
  assign n2477 = n579 & ~n2476;
  assign n2478 = ~n1218 & ~n1338;
  assign n2479 = n560 & ~n2478;
  assign n2480 = ~n2477 & ~n2479;
  assign n2481 = n520 & ~n1591;
  assign n2482 = ~n1331 & ~n1362;
  assign n2483 = n540 & ~n2482;
  assign n2484 = ~n2481 & ~n2483;
  assign n2485 = ~n1208 & ~n1268;
  assign n2486 = n601 & ~n2485;
  assign n2487 = ~n1237 & ~n1255;
  assign n2488 = n464 & ~n2487;
  assign n2489 = ~n2486 & ~n2488;
  assign n2490 = ~n1200 & ~n1366;
  assign n2491 = n606 & ~n2490;
  assign n2492 = ~n1245 & ~n1339;
  assign n2493 = n499 & ~n2492;
  assign n2494 = ~n2491 & ~n2493;
  assign n2495 = n2489 & n2494;
  assign n2496 = n684 & ~n1546;
  assign n2497 = n632 & ~n1541;
  assign n2498 = ~n2496 & ~n2497;
  assign n2499 = n2495 & n2498;
  assign n2500 = n2484 & n2499;
  assign n2501 = n2480 & n2500;
  assign n2502 = ~n1302 & ~n1320;
  assign n2503 = n673 & ~n2502;
  assign n2504 = ~n1365 & ~n1372;
  assign n2505 = n638 & ~n2504;
  assign n2506 = ~n2503 & ~n2505;
  assign n2507 = ~n1332 & ~n1349;
  assign n2508 = n678 & ~n2507;
  assign n2509 = ~n1279 & ~n1357;
  assign n2510 = n613 & ~n2509;
  assign n2511 = ~n1291 & ~n1377;
  assign n2512 = n643 & ~n2511;
  assign n2513 = ~n2510 & ~n2512;
  assign n2514 = n650 & ~n1582;
  assign n2515 = n2513 & ~n2514;
  assign n2516 = ~n2508 & n2515;
  assign n2517 = n2506 & n2516;
  assign n2518 = n2501 & n2517;
  assign n2519 = ~po31 & ~n2518;
  assign n2520 = po31 & n2516;
  assign n2521 = n2506 & n2520;
  assign n2522 = n2501 & n2521;
  assign n2523 = ~n2519 & ~n2522;
  assign n2524 = n632 & ~n1442;
  assign n2525 = n684 & ~n1500;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = ~n1302 & ~n1579;
  assign n2528 = n540 & ~n2527;
  assign n2529 = n2526 & ~n2528;
  assign n2530 = ~n1328 & ~n1373;
  assign n2531 = n678 & ~n2530;
  assign n2532 = n650 & ~n1413;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = ~n1365 & ~n1588;
  assign n2535 = n613 & ~n2534;
  assign n2536 = ~n1237 & ~n1566;
  assign n2537 = n643 & ~n2536;
  assign n2538 = ~n2535 & ~n2537;
  assign n2539 = n2533 & n2538;
  assign n2540 = ~n1269 & ~n1377;
  assign n2541 = n464 & ~n2540;
  assign n2542 = n2539 & ~n2541;
  assign n2543 = ~n1208 & ~n1292;
  assign n2544 = n499 & ~n2543;
  assign n2545 = ~n1287 & ~n1338;
  assign n2546 = n606 & ~n2545;
  assign n2547 = ~n1226 & ~n1357;
  assign n2548 = n638 & ~n2547;
  assign n2549 = ~n1331 & ~n1602;
  assign n2550 = n673 & ~n2549;
  assign n2551 = ~n2548 & ~n2550;
  assign n2552 = ~n2546 & n2551;
  assign n2553 = ~n2544 & n2552;
  assign n2554 = n520 & ~n1439;
  assign n2555 = ~n1263 & ~n1361;
  assign n2556 = n579 & ~n2555;
  assign n2557 = ~n2554 & ~n2556;
  assign n2558 = ~n1245 & ~n1594;
  assign n2559 = n601 & ~n2558;
  assign n2560 = ~n1366 & ~n1556;
  assign n2561 = n560 & ~n2560;
  assign n2562 = ~n2559 & ~n2561;
  assign n2563 = n2557 & n2562;
  assign n2564 = n2553 & n2563;
  assign n2565 = n2542 & n2564;
  assign n2566 = n2529 & n2565;
  assign n2567 = ~po05 & n2566;
  assign n2568 = po05 & ~n2566;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = ~n2523 & ~n2569;
  assign n2571 = ~n2475 & n2570;
  assign n2572 = ~n2429 & n2571;
  assign n2573 = ~n449 & n454;
  assign n2574 = pi102 & n2573;
  assign n2575 = pi102 & n449;
  assign n2576 = pi032 & ~n454;
  assign n2577 = ~n449 & n2576;
  assign n2578 = ~n2575 & ~n2577;
  assign n2579 = ~n2574 & n2578;
  assign n2580 = ~n446 & ~n2579;
  assign n2581 = pi191 & n446;
  assign po63 = n2580 | n2581;
  assign n2583 = ~n1338 & ~n1499;
  assign n2584 = n613 & ~n2583;
  assign n2585 = ~n1208 & ~n1412;
  assign n2586 = n643 & ~n2585;
  assign n2587 = ~n2584 & ~n2586;
  assign n2588 = n520 & ~n2107;
  assign n2589 = ~n1287 & ~n1566;
  assign n2590 = n499 & ~n2589;
  assign n2591 = ~n2588 & ~n2590;
  assign n2592 = ~n1377 & ~n1494;
  assign n2593 = n601 & ~n2592;
  assign n2594 = ~n1269 & ~n1579;
  assign n2595 = n579 & ~n2594;
  assign n2596 = ~n2593 & ~n2595;
  assign n2597 = n2591 & n2596;
  assign n2598 = ~n1292 & ~n1588;
  assign n2599 = n606 & ~n2598;
  assign n2600 = ~n1361 & ~n1594;
  assign n2601 = n464 & ~n2600;
  assign n2602 = ~n2599 & ~n2601;
  assign n2603 = ~n1263 & ~n1438;
  assign n2604 = n540 & ~n2603;
  assign n2605 = ~n1357 & ~n1463;
  assign n2606 = n560 & ~n2605;
  assign n2607 = ~n2604 & ~n2606;
  assign n2608 = n2602 & n2607;
  assign n2609 = n2597 & n2608;
  assign n2610 = n2587 & n2609;
  assign n2611 = ~n1373 & ~n1441;
  assign n2612 = n673 & ~n2611;
  assign n2613 = n650 & ~n2091;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = ~n1226 & ~n1602;
  assign n2616 = n678 & ~n2615;
  assign n2617 = n632 & ~n2100;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n1328 & ~n1556;
  assign n2620 = n638 & ~n2619;
  assign n2621 = n684 & ~n2112;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = n2618 & n2622;
  assign n2624 = n2614 & n2623;
  assign n2625 = n2610 & n2624;
  assign n2626 = ~po63 & n2625;
  assign n2627 = po63 & ~n2625;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~n2475 & n2569;
  assign n2630 = n2475 & n2570;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = n2429 & ~n2631;
  assign n2633 = ~n1394 & ~n1579;
  assign n2634 = n601 & ~n2633;
  assign n2635 = ~n1412 & ~n1491;
  assign n2636 = n606 & ~n2635;
  assign n2637 = ~n2634 & ~n2636;
  assign n2638 = ~n1507 & ~n1594;
  assign n2639 = n540 & ~n2638;
  assign n2640 = n520 & ~n1270;
  assign n2641 = ~n2639 & ~n2640;
  assign n2642 = ~n1502 & ~n1602;
  assign n2643 = n560 & ~n2642;
  assign n2644 = ~n1488 & ~n1499;
  assign n2645 = n499 & ~n2644;
  assign n2646 = ~n2643 & ~n2645;
  assign n2647 = n2641 & n2646;
  assign n2648 = ~n1452 & ~n1556;
  assign n2649 = n673 & ~n2648;
  assign n2650 = n684 & ~n1293;
  assign n2651 = ~n2649 & ~n2650;
  assign n2652 = ~n1426 & ~n1463;
  assign n2653 = n678 & ~n2652;
  assign n2654 = ~n1441 & ~n1473;
  assign n2655 = n638 & ~n2654;
  assign n2656 = ~n2653 & ~n2655;
  assign n2657 = n2651 & n2656;
  assign n2658 = n632 & ~n1227;
  assign n2659 = ~n1503 & ~n1566;
  assign n2660 = n613 & ~n2659;
  assign n2661 = ~n1402 & ~n1588;
  assign n2662 = n643 & ~n2661;
  assign n2663 = ~n2660 & ~n2662;
  assign n2664 = n650 & ~n1288;
  assign n2665 = n2663 & ~n2664;
  assign n2666 = ~n2658 & n2665;
  assign n2667 = n2657 & n2666;
  assign n2668 = ~n1438 & ~n1477;
  assign n2669 = n464 & ~n2668;
  assign n2670 = ~n1423 & ~n1494;
  assign n2671 = n579 & ~n2670;
  assign n2672 = ~n2669 & ~n2671;
  assign n2673 = n2667 & n2672;
  assign n2674 = n2647 & n2673;
  assign n2675 = n2637 & n2674;
  assign n2676 = pi103 & n449;
  assign n2677 = pi045 & ~n454;
  assign n2678 = pi103 & n454;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n449 & ~n2679;
  assign n2681 = ~n2676 & ~n2680;
  assign n2682 = ~n446 & ~n2681;
  assign n2683 = pi175 & n446;
  assign po47 = n2682 | n2683;
  assign n2685 = n2675 & po47;
  assign n2686 = ~n2675 & ~po47;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = n2523 & ~n2569;
  assign n2689 = ~n2687 & n2688;
  assign n2690 = n2523 & n2569;
  assign n2691 = n2475 & n2690;
  assign n2692 = ~n2689 & ~n2691;
  assign n2693 = ~n2429 & ~n2692;
  assign n2694 = ~n2632 & ~n2693;
  assign n2695 = n2475 & ~n2523;
  assign n2696 = n2687 & n2695;
  assign n2697 = n2569 & n2696;
  assign n2698 = n2694 & ~n2697;
  assign n2699 = ~n2628 & ~n2698;
  assign n2700 = ~n2475 & n2687;
  assign n2701 = n2523 & n2700;
  assign n2702 = n2569 & n2701;
  assign n2703 = n2475 & ~n2687;
  assign n2704 = ~n2523 & n2703;
  assign n2705 = ~n2429 & n2687;
  assign n2706 = ~n2475 & n2705;
  assign n2707 = ~n2523 & n2706;
  assign n2708 = ~n2704 & ~n2707;
  assign n2709 = n2569 & n2703;
  assign n2710 = n2708 & ~n2709;
  assign n2711 = ~n2475 & n2688;
  assign n2712 = n2429 & n2711;
  assign n2713 = n2475 & n2688;
  assign n2714 = n2687 & n2713;
  assign n2715 = ~n2712 & ~n2714;
  assign n2716 = n2710 & n2715;
  assign n2717 = ~n2702 & n2716;
  assign n2718 = n2628 & ~n2717;
  assign n2719 = ~n2523 & n2569;
  assign n2720 = ~n2475 & n2719;
  assign n2721 = ~n2687 & n2720;
  assign n2722 = n2687 & n2688;
  assign n2723 = ~n2721 & ~n2722;
  assign n2724 = n2429 & ~n2723;
  assign n2725 = ~n2718 & ~n2724;
  assign n2726 = ~n2699 & n2725;
  assign n2727 = ~n2572 & n2726;
  assign n2728 = n2374 & ~n2727;
  assign n2729 = ~n2374 & n2727;
  assign po10 = n2728 | n2729;
  assign n2731 = n2014 & n2246;
  assign n2732 = ~n2284 & ~n2731;
  assign n2733 = n2069 & n2344;
  assign n2734 = n2069 & n2334;
  assign n2735 = n2014 & n2129;
  assign n2736 = ~n2255 & ~n2735;
  assign n2737 = n2240 & ~n2736;
  assign n2738 = ~n2734 & ~n2737;
  assign n2739 = n2069 & ~n2240;
  assign n2740 = n2267 & n2739;
  assign n2741 = ~n2240 & n2344;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = n2738 & n2742;
  assign n2744 = ~n2733 & n2743;
  assign n2745 = n2732 & n2744;
  assign n2746 = ~n1955 & ~n2745;
  assign n2747 = ~n2255 & ~n2264;
  assign n2748 = ~n2069 & n2177;
  assign n2749 = n2747 & ~n2748;
  assign n2750 = ~n2240 & ~n2749;
  assign n2751 = n2282 & ~n2352;
  assign n2752 = n2240 & n2283;
  assign n2753 = n2751 & ~n2752;
  assign n2754 = ~n2750 & n2753;
  assign n2755 = n1955 & ~n2754;
  assign n2756 = n2282 & ~n2733;
  assign n2757 = ~n2240 & ~n2756;
  assign n2758 = ~n2014 & n2128;
  assign n2759 = n2321 & n2758;
  assign n2760 = n2069 & n2326;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = ~n2757 & n2761;
  assign n2763 = ~n2755 & n2762;
  assign n2764 = ~n2746 & n2763;
  assign n2765 = pi115 & ~n454;
  assign n2766 = pi038 & n454;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = ~n449 & ~n2767;
  assign n2769 = pi038 & n449;
  assign n2770 = ~n2768 & ~n2769;
  assign n2771 = ~n446 & ~n2770;
  assign n2772 = pi140 & n446;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = ~n2764 & n2773;
  assign n2775 = n2764 & ~n2773;
  assign po12 = n2774 | n2775;
  assign n2777 = pi141 & n446;
  assign n2778 = pi041 & ~n454;
  assign n2779 = pi113 & n454;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = ~n449 & ~n2780;
  assign n2782 = pi113 & n449;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = ~n446 & ~n2783;
  assign po13 = n2777 | n2784;
  assign n2786 = pi142 & n446;
  assign n2787 = pi120 & ~n454;
  assign n2788 = pi022 & n454;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = ~n449 & ~n2789;
  assign n2791 = pi022 & n449;
  assign n2792 = ~n2790 & ~n2791;
  assign n2793 = ~n446 & ~n2792;
  assign n2794 = ~n2786 & ~n2793;
  assign n2795 = ~n2631 & ~n2687;
  assign n2796 = ~n2429 & n2475;
  assign n2797 = ~n2687 & n2796;
  assign n2798 = ~n2569 & n2797;
  assign n2799 = n2687 & n2690;
  assign n2800 = ~n2475 & n2523;
  assign n2801 = n2687 & n2800;
  assign n2802 = ~n2630 & ~n2801;
  assign n2803 = ~n2799 & n2802;
  assign n2804 = ~n2429 & ~n2803;
  assign n2805 = n2429 & n2687;
  assign n2806 = n2713 & n2805;
  assign n2807 = ~n2804 & ~n2806;
  assign n2808 = ~n2798 & n2807;
  assign n2809 = ~n2795 & n2808;
  assign n2810 = n2571 & n2687;
  assign n2811 = n2809 & ~n2810;
  assign n2812 = n2628 & ~n2811;
  assign n2813 = ~n2687 & n2691;
  assign n2814 = ~n2475 & ~n2687;
  assign n2815 = n2688 & n2814;
  assign n2816 = ~n2800 & ~n2814;
  assign n2817 = n2429 & ~n2816;
  assign n2818 = ~n2815 & ~n2817;
  assign n2819 = ~n2813 & n2818;
  assign n2820 = ~n2628 & ~n2819;
  assign n2821 = n2630 & ~n2687;
  assign n2822 = ~n2810 & ~n2821;
  assign n2823 = ~n2429 & ~n2822;
  assign n2824 = n2569 & n2695;
  assign n2825 = ~n2713 & ~n2719;
  assign n2826 = n2687 & ~n2825;
  assign n2827 = ~n2824 & ~n2826;
  assign n2828 = ~n2429 & ~n2827;
  assign n2829 = ~n2628 & n2828;
  assign n2830 = ~n2687 & n2800;
  assign n2831 = ~n2697 & ~n2830;
  assign n2832 = n2429 & ~n2831;
  assign n2833 = ~n2829 & ~n2832;
  assign n2834 = ~n2823 & n2833;
  assign n2835 = ~n2820 & n2834;
  assign n2836 = ~n2812 & n2835;
  assign n2837 = n2794 & ~n2836;
  assign n2838 = ~n2794 & n2836;
  assign po14 = n2837 | n2838;
  assign n2840 = pi144 & n446;
  assign n2841 = pi036 & n449;
  assign n2842 = pi069 & ~n454;
  assign n2843 = pi036 & n454;
  assign n2844 = ~n2842 & ~n2843;
  assign n2845 = ~n449 & ~n2844;
  assign n2846 = ~n2841 & ~n2845;
  assign n2847 = ~n446 & ~n2846;
  assign n2848 = ~n2840 & ~n2847;
  assign n2849 = ~n757 & ~n855;
  assign n2850 = n638 & ~n2849;
  assign n2851 = ~n644 & ~n729;
  assign n2852 = n684 & ~n2851;
  assign n2853 = ~n2850 & ~n2852;
  assign n2854 = ~n633 & ~n747;
  assign n2855 = n560 & ~n2854;
  assign n2856 = ~n528 & ~n774;
  assign n2857 = n601 & ~n2856;
  assign n2858 = ~n2855 & ~n2857;
  assign n2859 = ~n602 & ~n856;
  assign n2860 = n520 & ~n2859;
  assign n2861 = ~n811 & ~n822;
  assign n2862 = n540 & ~n2861;
  assign n2863 = ~n2860 & ~n2862;
  assign n2864 = n2858 & n2863;
  assign n2865 = ~n785 & ~n828;
  assign n2866 = n579 & ~n2865;
  assign n2867 = ~n739 & ~n798;
  assign n2868 = n499 & ~n2867;
  assign n2869 = ~n2866 & ~n2868;
  assign n2870 = ~n765 & ~n773;
  assign n2871 = n606 & ~n2870;
  assign n2872 = ~n797 & ~n844;
  assign n2873 = n464 & ~n2872;
  assign n2874 = ~n2871 & ~n2873;
  assign n2875 = n2869 & n2874;
  assign n2876 = n2864 & n2875;
  assign n2877 = ~n568 & ~n852;
  assign n2878 = n632 & ~n2877;
  assign n2879 = ~n721 & ~n827;
  assign n2880 = n673 & ~n2879;
  assign n2881 = ~n2878 & ~n2880;
  assign n2882 = ~n685 & ~n793;
  assign n2883 = n643 & ~n2882;
  assign n2884 = ~n621 & ~n823;
  assign n2885 = n650 & ~n2884;
  assign n2886 = ~n2883 & ~n2885;
  assign n2887 = n2881 & n2886;
  assign n2888 = ~n658 & ~n832;
  assign n2889 = n613 & ~n2888;
  assign n2890 = ~n819 & ~n831;
  assign n2891 = n678 & ~n2890;
  assign n2892 = ~n2889 & ~n2891;
  assign n2893 = n2887 & n2892;
  assign n2894 = n2876 & n2893;
  assign n2895 = n2853 & n2894;
  assign n2896 = po57 & n2895;
  assign n2897 = ~po57 & ~n2895;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = ~n670 & ~n747;
  assign n2900 = n606 & ~n2899;
  assign n2901 = ~n686 & ~n774;
  assign n2902 = n499 & ~n2901;
  assign n2903 = ~n2900 & ~n2902;
  assign n2904 = ~n823 & ~n852;
  assign n2905 = n579 & ~n2904;
  assign n2906 = ~n495 & ~n819;
  assign n2907 = n520 & ~n2906;
  assign n2908 = ~n2905 & ~n2907;
  assign n2909 = n2903 & n2908;
  assign n2910 = ~n536 & ~n793;
  assign n2911 = n464 & ~n2910;
  assign n2912 = ~n675 & ~n765;
  assign n2913 = n560 & ~n2912;
  assign n2914 = ~n2911 & ~n2913;
  assign n2915 = ~n548 & ~n798;
  assign n2916 = n601 & ~n2915;
  assign n2917 = ~n603 & ~n827;
  assign n2918 = n540 & ~n2917;
  assign n2919 = ~n2916 & ~n2918;
  assign n2920 = n2914 & n2919;
  assign n2921 = n2909 & n2920;
  assign n2922 = ~n639 & ~n828;
  assign n2923 = n632 & ~n2922;
  assign n2924 = ~n607 & ~n785;
  assign n2925 = n650 & ~n2924;
  assign n2926 = ~n2923 & ~n2925;
  assign n2927 = ~n515 & ~n831;
  assign n2928 = n684 & ~n2927;
  assign n2929 = ~n729 & ~n856;
  assign n2930 = n678 & ~n2929;
  assign n2931 = ~n2928 & ~n2930;
  assign n2932 = ~n645 & ~n757;
  assign n2933 = n613 & ~n2932;
  assign n2934 = ~n629 & ~n797;
  assign n2935 = n643 & ~n2934;
  assign n2936 = ~n2933 & ~n2935;
  assign n2937 = n2931 & n2936;
  assign n2938 = ~n576 & ~n811;
  assign n2939 = n673 & ~n2938;
  assign n2940 = ~n634 & ~n832;
  assign n2941 = n638 & ~n2940;
  assign n2942 = ~n2939 & ~n2941;
  assign n2943 = n2937 & n2942;
  assign n2944 = n2926 & n2943;
  assign n2945 = n2921 & n2944;
  assign n2946 = pi085 & ~n694;
  assign n2947 = pi030 & n694;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = ~n446 & ~n2948;
  assign n2950 = pi177 & n446;
  assign po49 = n2949 | n2950;
  assign n2952 = n2945 & po49;
  assign n2953 = ~n2945 & ~po49;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = ~n773 & ~n827;
  assign n2956 = n464 & ~n2955;
  assign n2957 = ~n658 & ~n852;
  assign n2958 = n601 & ~n2957;
  assign n2959 = ~n798 & ~n819;
  assign n2960 = n579 & ~n2959;
  assign n2961 = ~n2958 & ~n2960;
  assign n2962 = ~n633 & ~n823;
  assign n2963 = n520 & ~n2962;
  assign n2964 = n2961 & ~n2963;
  assign n2965 = ~n2956 & n2964;
  assign n2966 = ~n528 & ~n729;
  assign n2967 = n632 & ~n2966;
  assign n2968 = ~n765 & ~n828;
  assign n2969 = n678 & ~n2968;
  assign n2970 = ~n2967 & ~n2969;
  assign n2971 = ~n797 & ~n831;
  assign n2972 = n606 & ~n2971;
  assign n2973 = n2970 & ~n2972;
  assign n2974 = ~n602 & ~n686;
  assign n2975 = n650 & ~n2974;
  assign n2976 = ~n739 & ~n811;
  assign n2977 = n638 & ~n2976;
  assign n2978 = ~n2975 & ~n2977;
  assign n2979 = ~n721 & ~n774;
  assign n2980 = n613 & ~n2979;
  assign n2981 = ~n747 & ~n822;
  assign n2982 = n643 & ~n2981;
  assign n2983 = ~n2980 & ~n2982;
  assign n2984 = n2978 & n2983;
  assign n2985 = ~n568 & ~n670;
  assign n2986 = n684 & ~n2985;
  assign n2987 = ~n832 & ~n844;
  assign n2988 = n673 & ~n2987;
  assign n2989 = ~n2986 & ~n2988;
  assign n2990 = ~n685 & ~n856;
  assign n2991 = n560 & ~n2990;
  assign n2992 = n2989 & ~n2991;
  assign n2993 = ~n793 & ~n855;
  assign n2994 = n540 & ~n2993;
  assign n2995 = ~n757 & ~n785;
  assign n2996 = n499 & ~n2995;
  assign n2997 = ~n2994 & ~n2996;
  assign n2998 = n2992 & n2997;
  assign n2999 = n2984 & n2998;
  assign n3000 = n2973 & n2999;
  assign n3001 = n2965 & n3000;
  assign n3002 = pi124 & n449;
  assign n3003 = pi013 & ~n454;
  assign n3004 = pi124 & n454;
  assign n3005 = ~n3003 & ~n3004;
  assign n3006 = ~n449 & ~n3005;
  assign n3007 = ~n3002 & ~n3006;
  assign n3008 = ~n446 & ~n3007;
  assign n3009 = pi161 & n446;
  assign po33 = n3008 | n3009;
  assign n3011 = n3001 & po33;
  assign n3012 = n2961 & n2992;
  assign n3013 = n2984 & n3012;
  assign n3014 = n2973 & n3013;
  assign n3015 = ~n2956 & ~n2963;
  assign n3016 = n2997 & n3015;
  assign n3017 = n3014 & n3016;
  assign n3018 = ~po33 & ~n3017;
  assign n3019 = ~n3011 & ~n3018;
  assign n3020 = ~n640 & ~n827;
  assign n3021 = n650 & ~n3020;
  assign n3022 = ~n507 & ~n832;
  assign n3023 = n520 & ~n3022;
  assign n3024 = ~n576 & ~n629;
  assign n3025 = n579 & ~n3024;
  assign n3026 = ~n3023 & ~n3025;
  assign n3027 = ~n3021 & n3026;
  assign n3028 = ~n680 & ~n747;
  assign n3029 = n601 & ~n3028;
  assign n3030 = ~n595 & ~n774;
  assign n3031 = n560 & ~n3030;
  assign n3032 = ~n3029 & ~n3031;
  assign n3033 = ~n487 & ~n811;
  assign n3034 = n684 & ~n3033;
  assign n3035 = n3032 & ~n3034;
  assign n3036 = ~n495 & ~n670;
  assign n3037 = n638 & ~n3036;
  assign n3038 = n3035 & ~n3037;
  assign n3039 = n3027 & n3038;
  assign n3040 = ~n603 & ~n645;
  assign n3041 = n678 & ~n3040;
  assign n3042 = ~n608 & ~n793;
  assign n3043 = n632 & ~n3042;
  assign n3044 = ~n607 & ~n729;
  assign n3045 = n540 & ~n3044;
  assign n3046 = ~n639 & ~n686;
  assign n3047 = n464 & ~n3046;
  assign n3048 = ~n3045 & ~n3047;
  assign n3049 = ~n3043 & n3048;
  assign n3050 = ~n587 & ~n856;
  assign n3051 = n613 & ~n3050;
  assign n3052 = ~n548 & ~n634;
  assign n3053 = n606 & ~n3052;
  assign n3054 = ~n536 & ~n675;
  assign n3055 = n499 & ~n3054;
  assign n3056 = ~n3053 & ~n3055;
  assign n3057 = ~n3051 & n3056;
  assign n3058 = ~n515 & ~n823;
  assign n3059 = n673 & ~n3058;
  assign n3060 = ~n679 & ~n852;
  assign n3061 = n643 & ~n3060;
  assign n3062 = ~n3059 & ~n3061;
  assign n3063 = n3057 & n3062;
  assign n3064 = n3049 & n3063;
  assign n3065 = ~n3041 & n3064;
  assign n3066 = n3039 & n3065;
  assign n3067 = po07 & ~n3066;
  assign n3068 = ~po07 & n3066;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = ~n3019 & n3069;
  assign n3071 = pi081 & n454;
  assign n3072 = pi024 & ~n454;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = ~n449 & ~n3073;
  assign n3075 = pi081 & n449;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = ~n446 & ~n3076;
  assign n3078 = pi153 & n446;
  assign po25 = n3077 | n3078;
  assign n3080 = ~n658 & ~n739;
  assign n3081 = n606 & ~n3080;
  assign n3082 = ~n602 & ~n828;
  assign n3083 = n540 & ~n3082;
  assign n3084 = ~n3081 & ~n3083;
  assign n3085 = ~n721 & ~n855;
  assign n3086 = n678 & ~n3085;
  assign n3087 = n650 & ~n3042;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = ~n621 & ~n798;
  assign n3090 = n643 & ~n3089;
  assign n3091 = ~n568 & ~n819;
  assign n3092 = n673 & ~n3091;
  assign n3093 = ~n3090 & ~n3092;
  assign n3094 = n3088 & n3093;
  assign n3095 = n632 & ~n3020;
  assign n3096 = ~n644 & ~n765;
  assign n3097 = n613 & ~n3096;
  assign n3098 = ~n633 & ~n831;
  assign n3099 = n638 & ~n3098;
  assign n3100 = ~n3097 & ~n3099;
  assign n3101 = n684 & ~n3022;
  assign n3102 = n3100 & ~n3101;
  assign n3103 = ~n3095 & n3102;
  assign n3104 = n3094 & n3103;
  assign n3105 = ~n556 & ~n797;
  assign n3106 = n601 & ~n3105;
  assign n3107 = ~n674 & ~n757;
  assign n3108 = n560 & ~n3107;
  assign n3109 = ~n3106 & ~n3108;
  assign n3110 = n520 & ~n3033;
  assign n3111 = ~n822 & ~n844;
  assign n3112 = n579 & ~n3111;
  assign n3113 = ~n3110 & ~n3112;
  assign n3114 = n3109 & n3113;
  assign n3115 = ~n685 & ~n773;
  assign n3116 = n499 & ~n3115;
  assign n3117 = ~n528 & ~n785;
  assign n3118 = n464 & ~n3117;
  assign n3119 = ~n3116 & ~n3118;
  assign n3120 = n3114 & n3119;
  assign n3121 = n3104 & n3120;
  assign n3122 = n3084 & n3121;
  assign n3123 = po25 & n3122;
  assign n3124 = ~po25 & ~n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = n3069 & n3125;
  assign n3127 = ~n608 & ~n721;
  assign n3128 = n540 & ~n3127;
  assign n3129 = ~n640 & ~n685;
  assign n3130 = n464 & ~n3129;
  assign n3131 = ~n3128 & ~n3130;
  assign n3132 = ~n587 & ~n773;
  assign n3133 = n560 & ~n3132;
  assign n3134 = ~n528 & ~n674;
  assign n3135 = n499 & ~n3134;
  assign n3136 = ~n3133 & ~n3135;
  assign n3137 = ~n568 & ~n621;
  assign n3138 = n579 & ~n3137;
  assign n3139 = n3136 & ~n3138;
  assign n3140 = ~n487 & ~n658;
  assign n3141 = n638 & ~n3140;
  assign n3142 = ~n595 & ~n855;
  assign n3143 = n613 & ~n3142;
  assign n3144 = ~n602 & ~n644;
  assign n3145 = n678 & ~n3144;
  assign n3146 = ~n3143 & ~n3145;
  assign n3147 = n632 & ~n2924;
  assign n3148 = n3146 & ~n3147;
  assign n3149 = ~n3141 & n3148;
  assign n3150 = n650 & ~n2922;
  assign n3151 = ~n507 & ~n822;
  assign n3152 = n673 & ~n3151;
  assign n3153 = ~n680 & ~n844;
  assign n3154 = n643 & ~n3153;
  assign n3155 = ~n3152 & ~n3154;
  assign n3156 = n684 & ~n2906;
  assign n3157 = n3155 & ~n3156;
  assign n3158 = ~n3150 & n3157;
  assign n3159 = n3149 & n3158;
  assign n3160 = n520 & ~n2927;
  assign n3161 = ~n679 & ~n739;
  assign n3162 = n601 & ~n3161;
  assign n3163 = ~n3160 & ~n3162;
  assign n3164 = ~n556 & ~n633;
  assign n3165 = n606 & ~n3164;
  assign n3166 = n3163 & ~n3165;
  assign n3167 = n3159 & n3166;
  assign n3168 = n3139 & n3167;
  assign n3169 = n3131 & n3168;
  assign n3170 = pi057 & ~n449;
  assign n3171 = ~n454 & n3170;
  assign n3172 = pi079 & ~n449;
  assign n3173 = n454 & n3172;
  assign n3174 = pi079 & n449;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = ~n3171 & n3175;
  assign n3177 = ~n446 & ~n3176;
  assign n3178 = pi169 & n446;
  assign po41 = n3177 | n3178;
  assign n3180 = n3169 & po41;
  assign n3181 = ~n3169 & ~po41;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = n3126 & n3182;
  assign n3184 = ~n3070 & ~n3183;
  assign n3185 = n3019 & ~n3069;
  assign n3186 = ~n3182 & n3185;
  assign n3187 = n3184 & ~n3186;
  assign n3188 = n2954 & ~n3187;
  assign n3189 = ~n3069 & ~n3125;
  assign n3190 = ~n3019 & n3189;
  assign n3191 = n3182 & n3190;
  assign n3192 = ~n3188 & ~n3191;
  assign n3193 = ~n2898 & ~n3192;
  assign n3194 = ~po25 & n3122;
  assign n3195 = po25 & ~n3122;
  assign n3196 = ~n3194 & ~n3195;
  assign n3197 = ~n3069 & ~n3196;
  assign n3198 = ~n3019 & ~n3182;
  assign n3199 = n3197 & n3198;
  assign n3200 = n3069 & ~n3125;
  assign n3201 = n3019 & n3200;
  assign n3202 = n3182 & n3201;
  assign n3203 = ~n3199 & ~n3202;
  assign n3204 = ~n2954 & ~n3203;
  assign n3205 = ~n3019 & ~n3069;
  assign n3206 = ~n3182 & n3205;
  assign n3207 = ~n3019 & n3182;
  assign n3208 = ~n3196 & n3207;
  assign n3209 = n3069 & n3208;
  assign n3210 = n3185 & n3196;
  assign n3211 = n3182 & n3210;
  assign n3212 = ~n3209 & ~n3211;
  assign n3213 = n3019 & n3126;
  assign n3214 = ~n3210 & ~n3213;
  assign n3215 = ~n3019 & n3196;
  assign n3216 = ~n3182 & n3215;
  assign n3217 = n3214 & ~n3216;
  assign n3218 = ~n2954 & ~n3217;
  assign n3219 = ~n3182 & n3201;
  assign n3220 = n3019 & n3197;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = n2954 & ~n3221;
  assign n3223 = ~n3218 & ~n3222;
  assign n3224 = n3212 & n3223;
  assign n3225 = ~n3206 & n3224;
  assign n3226 = n2898 & ~n3225;
  assign n3227 = n2954 & n3182;
  assign n3228 = n3070 & n3227;
  assign n3229 = ~n2954 & n3182;
  assign n3230 = n3197 & n3229;
  assign n3231 = ~n2954 & n3201;
  assign n3232 = ~n3230 & ~n3231;
  assign n3233 = ~n2898 & ~n3232;
  assign n3234 = ~n3228 & ~n3233;
  assign n3235 = n3019 & ~n3182;
  assign n3236 = n3126 & n3235;
  assign n3237 = ~n2954 & n3236;
  assign n3238 = n3234 & ~n3237;
  assign n3239 = ~n3226 & n3238;
  assign n3240 = ~n3204 & n3239;
  assign n3241 = ~n3193 & n3240;
  assign n3242 = ~n2848 & n3241;
  assign n3243 = n2848 & ~n3241;
  assign po16 = n3242 | n3243;
  assign n3245 = pi082 & n449;
  assign n3246 = pi044 & ~n454;
  assign n3247 = pi082 & n454;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = ~n449 & ~n3248;
  assign n3250 = ~n3245 & ~n3249;
  assign n3251 = ~n446 & ~n3250;
  assign n3252 = pi145 & n446;
  assign po17 = n3251 | n3252;
  assign n3254 = pi146 & n446;
  assign n3255 = pi037 & n449;
  assign n3256 = pi067 & ~n454;
  assign n3257 = pi037 & n454;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = ~n449 & ~n3258;
  assign n3260 = ~n3255 & ~n3259;
  assign n3261 = ~n446 & ~n3260;
  assign n3262 = ~n3254 & ~n3261;
  assign n3263 = ~n621 & ~n831;
  assign n3264 = n540 & ~n3263;
  assign n3265 = ~n528 & ~n855;
  assign n3266 = n606 & ~n3265;
  assign n3267 = ~n3264 & ~n3266;
  assign n3268 = ~n633 & ~n844;
  assign n3269 = n499 & ~n3268;
  assign n3270 = ~n685 & ~n721;
  assign n3271 = n579 & ~n3270;
  assign n3272 = ~n3269 & ~n3271;
  assign n3273 = ~n640 & ~n765;
  assign n3274 = n601 & ~n3273;
  assign n3275 = n520 & ~n999;
  assign n3276 = ~n3274 & ~n3275;
  assign n3277 = ~n487 & ~n798;
  assign n3278 = n560 & ~n3277;
  assign n3279 = ~n568 & ~n739;
  assign n3280 = n464 & ~n3279;
  assign n3281 = ~n3278 & ~n3280;
  assign n3282 = n3276 & n3281;
  assign n3283 = n3272 & n3282;
  assign n3284 = n3267 & n3283;
  assign n3285 = n650 & ~n990;
  assign n3286 = n632 & ~n1001;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n556 & ~n819;
  assign n3289 = n613 & ~n3288;
  assign n3290 = n684 & ~n1006;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = ~n674 & ~n828;
  assign n3293 = n643 & ~n3292;
  assign n3294 = ~n644 & ~n785;
  assign n3295 = n673 & ~n3294;
  assign n3296 = ~n3293 & ~n3295;
  assign n3297 = n3291 & n3296;
  assign n3298 = ~n658 & ~n822;
  assign n3299 = n678 & ~n3298;
  assign n3300 = ~n602 & ~n773;
  assign n3301 = n638 & ~n3300;
  assign n3302 = ~n3299 & ~n3301;
  assign n3303 = n3297 & n3302;
  assign n3304 = n3287 & n3303;
  assign n3305 = n3284 & n3304;
  assign n3306 = pi187 & n446;
  assign n3307 = pi077 & ~n694;
  assign n3308 = pi061 & n694;
  assign n3309 = ~n3307 & ~n3308;
  assign n3310 = ~n446 & ~n3309;
  assign po59 = n3306 | n3310;
  assign n3312 = n3305 & po59;
  assign n3313 = ~n3305 & ~po59;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n629 & ~n819;
  assign n3316 = n560 & ~n3315;
  assign n3317 = ~n823 & ~n832;
  assign n3318 = n499 & ~n3317;
  assign n3319 = ~n3316 & ~n3318;
  assign n3320 = ~n686 & ~n827;
  assign n3321 = n638 & ~n3320;
  assign n3322 = n650 & ~n1070;
  assign n3323 = ~n3321 & ~n3322;
  assign n3324 = ~n576 & ~n798;
  assign n3325 = n613 & ~n3324;
  assign n3326 = n684 & ~n1078;
  assign n3327 = ~n3325 & ~n3326;
  assign n3328 = n3323 & n3327;
  assign n3329 = ~n603 & ~n765;
  assign n3330 = n643 & ~n3329;
  assign n3331 = n632 & ~n1059;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = ~n747 & ~n852;
  assign n3334 = n678 & ~n3333;
  assign n3335 = ~n536 & ~n757;
  assign n3336 = n673 & ~n3335;
  assign n3337 = ~n3334 & ~n3336;
  assign n3338 = n3332 & n3337;
  assign n3339 = n3328 & n3338;
  assign n3340 = n520 & ~n1076;
  assign n3341 = ~n670 & ~n811;
  assign n3342 = n464 & ~n3341;
  assign n3343 = ~n3340 & ~n3342;
  assign n3344 = ~n634 & ~n797;
  assign n3345 = n540 & ~n3344;
  assign n3346 = ~n774 & ~n856;
  assign n3347 = n579 & ~n3346;
  assign n3348 = ~n3345 & ~n3347;
  assign n3349 = n3343 & n3348;
  assign n3350 = ~n645 & ~n828;
  assign n3351 = n601 & ~n3350;
  assign n3352 = ~n729 & ~n793;
  assign n3353 = n606 & ~n3352;
  assign n3354 = ~n3351 & ~n3353;
  assign n3355 = n3349 & n3354;
  assign n3356 = n3339 & n3355;
  assign n3357 = n3319 & n3356;
  assign n3358 = pi100 & ~n694;
  assign n3359 = pi015 & n694;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = ~n446 & ~n3360;
  assign n3362 = pi171 & n446;
  assign po43 = n3361 | n3362;
  assign n3364 = ~n3357 & ~po43;
  assign n3365 = n3357 & po43;
  assign n3366 = ~n3364 & ~n3365;
  assign n3367 = ~n729 & ~n773;
  assign n3368 = n613 & ~n3367;
  assign n3369 = ~n739 & ~n823;
  assign n3370 = n643 & ~n3369;
  assign n3371 = ~n3368 & ~n3370;
  assign n3372 = ~n774 & ~n828;
  assign n3373 = n464 & ~n3372;
  assign n3374 = ~n797 & ~n811;
  assign n3375 = n579 & ~n3374;
  assign n3376 = ~n3373 & ~n3375;
  assign n3377 = ~n765 & ~n793;
  assign n3378 = n499 & ~n3377;
  assign n3379 = ~n785 & ~n856;
  assign n3380 = n540 & ~n3379;
  assign n3381 = ~n3378 & ~n3380;
  assign n3382 = n3376 & n3381;
  assign n3383 = ~n686 & ~n855;
  assign n3384 = n560 & ~n3383;
  assign n3385 = ~n798 & ~n832;
  assign n3386 = n606 & ~n3385;
  assign n3387 = ~n3384 & ~n3386;
  assign n3388 = ~n634 & ~n822;
  assign n3389 = n520 & ~n3388;
  assign n3390 = ~n670 & ~n844;
  assign n3391 = n601 & ~n3390;
  assign n3392 = ~n3389 & ~n3391;
  assign n3393 = n3387 & n3392;
  assign n3394 = n3382 & n3393;
  assign n3395 = ~n757 & ~n827;
  assign n3396 = n678 & ~n3395;
  assign n3397 = ~n747 & ~n819;
  assign n3398 = n638 & ~n3397;
  assign n3399 = ~n3396 & ~n3398;
  assign n3400 = ~n831 & ~n852;
  assign n3401 = n673 & ~n3400;
  assign n3402 = ~n576 & ~n658;
  assign n3403 = n684 & ~n3402;
  assign n3404 = ~n3401 & ~n3403;
  assign n3405 = n3399 & n3404;
  assign n3406 = ~n603 & ~n685;
  assign n3407 = n650 & ~n3406;
  assign n3408 = ~n536 & ~n721;
  assign n3409 = n632 & ~n3408;
  assign n3410 = ~n3407 & ~n3409;
  assign n3411 = n3405 & n3410;
  assign n3412 = n3394 & n3411;
  assign n3413 = n3371 & n3412;
  assign n3414 = ~po35 & ~n3413;
  assign n3415 = po35 & n3413;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = ~n587 & ~n757;
  assign n3418 = n650 & ~n3417;
  assign n3419 = ~n679 & ~n797;
  assign n3420 = n684 & ~n3419;
  assign n3421 = ~n3418 & ~n3420;
  assign n3422 = ~n568 & ~n822;
  assign n3423 = n606 & ~n3422;
  assign n3424 = n3421 & ~n3423;
  assign n3425 = ~n640 & ~n785;
  assign n3426 = n613 & ~n3425;
  assign n3427 = ~n595 & ~n765;
  assign n3428 = n632 & ~n3427;
  assign n3429 = ~n3426 & ~n3428;
  assign n3430 = ~n487 & ~n831;
  assign n3431 = n643 & ~n3430;
  assign n3432 = ~n556 & ~n739;
  assign n3433 = n673 & ~n3432;
  assign n3434 = ~n3431 & ~n3433;
  assign n3435 = n3429 & n3434;
  assign n3436 = ~n644 & ~n855;
  assign n3437 = n464 & ~n3436;
  assign n3438 = n3435 & ~n3437;
  assign n3439 = ~n621 & ~n844;
  assign n3440 = n638 & ~n3439;
  assign n3441 = ~n528 & ~n685;
  assign n3442 = n678 & ~n3441;
  assign n3443 = ~n3440 & ~n3442;
  assign n3444 = ~n602 & ~n721;
  assign n3445 = n499 & ~n3444;
  assign n3446 = n3443 & ~n3445;
  assign n3447 = ~n633 & ~n658;
  assign n3448 = n579 & ~n3447;
  assign n3449 = n3446 & ~n3448;
  assign n3450 = ~n680 & ~n798;
  assign n3451 = n520 & ~n3450;
  assign n3452 = ~n608 & ~n828;
  assign n3453 = n560 & ~n3452;
  assign n3454 = ~n3451 & ~n3453;
  assign n3455 = ~n674 & ~n773;
  assign n3456 = n540 & ~n3455;
  assign n3457 = ~n507 & ~n819;
  assign n3458 = n601 & ~n3457;
  assign n3459 = ~n3456 & ~n3458;
  assign n3460 = n3454 & n3459;
  assign n3461 = n3449 & n3460;
  assign n3462 = n3438 & n3461;
  assign n3463 = n3424 & n3462;
  assign n3464 = ~po01 & ~n3463;
  assign n3465 = po01 & n3463;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = ~n536 & ~n595;
  assign n3468 = n540 & ~n3467;
  assign n3469 = ~n607 & ~n645;
  assign n3470 = n499 & ~n3469;
  assign n3471 = ~n3468 & ~n3470;
  assign n3472 = ~n556 & ~n852;
  assign n3473 = n520 & ~n3472;
  assign n3474 = ~n487 & ~n823;
  assign n3475 = n601 & ~n3474;
  assign n3476 = ~n3473 & ~n3475;
  assign n3477 = ~n640 & ~n729;
  assign n3478 = n560 & ~n3477;
  assign n3479 = ~n495 & ~n548;
  assign n3480 = n579 & ~n3479;
  assign n3481 = ~n3478 & ~n3480;
  assign n3482 = n3476 & n3481;
  assign n3483 = ~n621 & ~n747;
  assign n3484 = n684 & ~n3483;
  assign n3485 = ~n639 & ~n675;
  assign n3486 = n678 & ~n3485;
  assign n3487 = ~n674 & ~n856;
  assign n3488 = n632 & ~n3487;
  assign n3489 = ~n3486 & ~n3488;
  assign n3490 = ~n644 & ~n774;
  assign n3491 = n650 & ~n3490;
  assign n3492 = n3489 & ~n3491;
  assign n3493 = ~n3484 & n3492;
  assign n3494 = ~n576 & ~n679;
  assign n3495 = n638 & ~n3494;
  assign n3496 = ~n634 & ~n680;
  assign n3497 = n673 & ~n3496;
  assign n3498 = ~n608 & ~n686;
  assign n3499 = n613 & ~n3498;
  assign n3500 = ~n3497 & ~n3499;
  assign n3501 = ~n507 & ~n670;
  assign n3502 = n643 & ~n3501;
  assign n3503 = n3500 & ~n3502;
  assign n3504 = ~n3495 & n3503;
  assign n3505 = n3493 & n3504;
  assign n3506 = ~n587 & ~n603;
  assign n3507 = n464 & ~n3506;
  assign n3508 = ~n515 & ~n629;
  assign n3509 = n606 & ~n3508;
  assign n3510 = ~n3507 & ~n3509;
  assign n3511 = n3505 & n3510;
  assign n3512 = n3482 & n3511;
  assign n3513 = n3471 & n3512;
  assign n3514 = ~po27 & ~n3513;
  assign n3515 = po27 & n3513;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = n3466 & n3516;
  assign n3518 = n3416 & n3517;
  assign n3519 = n3366 & n3518;
  assign n3520 = pi054 & ~n449;
  assign n3521 = ~n454 & n3520;
  assign n3522 = pi078 & ~n449;
  assign n3523 = n454 & n3522;
  assign n3524 = pi078 & n449;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = ~n3521 & n3525;
  assign n3527 = ~n446 & ~n3526;
  assign n3528 = pi179 & n446;
  assign po51 = n3527 | n3528;
  assign n3530 = ~n670 & ~n679;
  assign n3531 = n540 & ~n3530;
  assign n3532 = ~n645 & ~n675;
  assign n3533 = n579 & ~n3532;
  assign n3534 = ~n3531 & ~n3533;
  assign n3535 = n520 & ~n876;
  assign n3536 = ~n608 & ~n856;
  assign n3537 = n601 & ~n3536;
  assign n3538 = ~n3535 & ~n3537;
  assign n3539 = ~n507 & ~n852;
  assign n3540 = n560 & ~n3539;
  assign n3541 = ~n515 & ~n634;
  assign n3542 = n464 & ~n3541;
  assign n3543 = ~n3540 & ~n3542;
  assign n3544 = n3538 & n3543;
  assign n3545 = ~n587 & ~n686;
  assign n3546 = n673 & ~n3545;
  assign n3547 = n684 & ~n918;
  assign n3548 = ~n3546 & ~n3547;
  assign n3549 = ~n680 & ~n823;
  assign n3550 = n613 & ~n3549;
  assign n3551 = ~n595 & ~n729;
  assign n3552 = n643 & ~n3551;
  assign n3553 = ~n3550 & ~n3552;
  assign n3554 = n3548 & n3553;
  assign n3555 = n650 & ~n887;
  assign n3556 = ~n536 & ~n607;
  assign n3557 = n638 & ~n3556;
  assign n3558 = ~n548 & ~n629;
  assign n3559 = n678 & ~n3558;
  assign n3560 = ~n3557 & ~n3559;
  assign n3561 = n632 & ~n881;
  assign n3562 = n3560 & ~n3561;
  assign n3563 = ~n3555 & n3562;
  assign n3564 = n3554 & n3563;
  assign n3565 = ~n603 & ~n639;
  assign n3566 = n606 & ~n3565;
  assign n3567 = ~n495 & ~n576;
  assign n3568 = n499 & ~n3567;
  assign n3569 = ~n3566 & ~n3568;
  assign n3570 = n3564 & n3569;
  assign n3571 = n3544 & n3570;
  assign n3572 = n3534 & n3571;
  assign n3573 = po51 & n3572;
  assign n3574 = ~po51 & ~n3572;
  assign n3575 = ~n3573 & ~n3574;
  assign n3576 = ~n3416 & n3516;
  assign n3577 = n3366 & n3516;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = ~n3466 & ~n3516;
  assign n3580 = n3416 & n3579;
  assign n3581 = n3578 & ~n3580;
  assign n3582 = n3575 & ~n3581;
  assign n3583 = ~n3416 & n3579;
  assign n3584 = n3466 & ~n3516;
  assign n3585 = n3416 & n3584;
  assign n3586 = ~n3583 & ~n3585;
  assign n3587 = ~n3575 & ~n3586;
  assign n3588 = ~n3582 & ~n3587;
  assign n3589 = ~n3519 & n3588;
  assign n3590 = ~n3314 & ~n3589;
  assign n3591 = ~n3416 & n3584;
  assign n3592 = n3575 & n3591;
  assign n3593 = ~n3366 & ~n3466;
  assign n3594 = n3416 & n3593;
  assign n3595 = ~n3366 & n3591;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = ~n3366 & n3516;
  assign n3598 = n3416 & n3597;
  assign n3599 = n3575 & n3598;
  assign n3600 = n3366 & n3585;
  assign n3601 = n3366 & n3583;
  assign n3602 = ~n3575 & n3576;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = ~n3600 & n3603;
  assign n3605 = ~n3599 & n3604;
  assign n3606 = n3596 & n3605;
  assign n3607 = ~n3592 & n3606;
  assign n3608 = n3314 & ~n3607;
  assign n3609 = n3575 & n3595;
  assign n3610 = ~n3366 & ~n3575;
  assign n3611 = n3466 & n3576;
  assign n3612 = n3610 & n3611;
  assign n3613 = ~n3466 & n3516;
  assign n3614 = n3610 & n3613;
  assign n3615 = n3416 & n3614;
  assign n3616 = ~n3612 & ~n3615;
  assign n3617 = ~n3609 & n3616;
  assign n3618 = ~n3608 & n3617;
  assign n3619 = ~n3590 & n3618;
  assign n3620 = ~n3262 & n3619;
  assign n3621 = n3262 & ~n3619;
  assign po18 = n3620 | n3621;
  assign n3623 = pi148 & n446;
  assign n3624 = pi068 & ~n454;
  assign n3625 = pi002 & n454;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = ~n449 & ~n3626;
  assign n3628 = pi002 & n449;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = ~n446 & ~n3629;
  assign n3631 = ~n3623 & ~n3630;
  assign n3632 = n3366 & n3517;
  assign n3633 = ~n3366 & n3416;
  assign n3634 = ~n3466 & n3633;
  assign n3635 = ~n3516 & n3634;
  assign n3636 = ~n3632 & ~n3635;
  assign n3637 = n3575 & ~n3636;
  assign n3638 = n3583 & n3610;
  assign n3639 = ~n3615 & ~n3638;
  assign n3640 = ~n3609 & n3639;
  assign n3641 = n3416 & ~n3516;
  assign n3642 = n3366 & n3641;
  assign n3643 = ~n3518 & ~n3642;
  assign n3644 = ~n3416 & n3613;
  assign n3645 = ~n3366 & n3644;
  assign n3646 = n3643 & ~n3645;
  assign n3647 = n3575 & ~n3646;
  assign n3648 = ~n3366 & n3611;
  assign n3649 = ~n3366 & n3585;
  assign n3650 = ~n3416 & ~n3516;
  assign n3651 = ~n3613 & ~n3650;
  assign n3652 = n3366 & ~n3651;
  assign n3653 = ~n3649 & ~n3652;
  assign n3654 = ~n3648 & n3653;
  assign n3655 = ~n3575 & ~n3654;
  assign n3656 = ~n3647 & ~n3655;
  assign n3657 = n3314 & ~n3656;
  assign n3658 = n3575 & n3576;
  assign n3659 = n3366 & n3658;
  assign n3660 = ~n3592 & ~n3659;
  assign n3661 = ~n3366 & n3575;
  assign n3662 = ~n3516 & n3661;
  assign n3663 = ~n3598 & ~n3642;
  assign n3664 = ~n3575 & ~n3663;
  assign n3665 = ~n3614 & ~n3664;
  assign n3666 = ~n3662 & n3665;
  assign n3667 = n3416 & n3613;
  assign n3668 = ~n3366 & n3667;
  assign n3669 = n3366 & n3466;
  assign n3670 = ~n3416 & n3669;
  assign n3671 = n3516 & n3670;
  assign n3672 = ~n3668 & ~n3671;
  assign n3673 = n3666 & n3672;
  assign n3674 = n3660 & n3673;
  assign n3675 = ~n3314 & ~n3674;
  assign n3676 = ~n3657 & ~n3675;
  assign n3677 = n3640 & n3676;
  assign n3678 = ~n3637 & n3677;
  assign n3679 = n3631 & n3678;
  assign n3680 = ~n3631 & ~n3678;
  assign po20 = n3679 | n3680;
  assign n3682 = pi083 & n449;
  assign n3683 = pi003 & ~n454;
  assign n3684 = pi083 & n454;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = ~n449 & ~n3685;
  assign n3687 = ~n3682 & ~n3686;
  assign n3688 = ~n446 & ~n3687;
  assign n3689 = pi149 & n446;
  assign po21 = n3688 | n3689;
  assign n3691 = n866 & ~n984;
  assign n3692 = ~n1121 & ~n3691;
  assign n3693 = n925 & ~n3692;
  assign n3694 = ~n925 & n1110;
  assign n3695 = ~n1149 & ~n3694;
  assign n3696 = n1106 & ~n3695;
  assign n3697 = n866 & n925;
  assign n3698 = ~n1144 & ~n3697;
  assign n3699 = ~n1136 & n3698;
  assign n3700 = ~n1106 & ~n3699;
  assign n3701 = ~n3696 & ~n3700;
  assign n3702 = ~n3693 & n3701;
  assign n3703 = ~n1046 & ~n3702;
  assign n3704 = ~n1106 & n1111;
  assign n3705 = n925 & n1118;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = ~n925 & n1143;
  assign n3708 = n984 & n1136;
  assign n3709 = ~n3707 & ~n3708;
  assign n3710 = n1106 & ~n3709;
  assign n3711 = ~n987 & ~n3710;
  assign n3712 = n3706 & n3711;
  assign n3713 = n1046 & ~n3712;
  assign n3714 = ~n3703 & ~n3713;
  assign n3715 = ~n925 & n1106;
  assign n3716 = n1118 & n3715;
  assign n3717 = n1106 & n1110;
  assign n3718 = n925 & n3717;
  assign n3719 = ~n984 & n3718;
  assign n3720 = ~n3716 & ~n3719;
  assign n3721 = ~n925 & n1155;
  assign n3722 = n925 & n1144;
  assign n3723 = ~n925 & n1149;
  assign n3724 = ~n3722 & ~n3723;
  assign n3725 = ~n3721 & n3724;
  assign n3726 = ~n1106 & ~n3725;
  assign n3727 = n3720 & ~n3726;
  assign n3728 = n3714 & n3727;
  assign n3729 = pi004 & n449;
  assign n3730 = pi072 & ~n454;
  assign n3731 = pi004 & n454;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = ~n449 & ~n3732;
  assign n3734 = ~n3729 & ~n3733;
  assign n3735 = ~n446 & ~n3734;
  assign n3736 = pi150 & n446;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = ~n3728 & n3737;
  assign n3739 = n3720 & ~n3737;
  assign n3740 = ~n3726 & n3739;
  assign n3741 = n3714 & n3740;
  assign po22 = n3738 | n3741;
  assign n3743 = n2475 & n2687;
  assign n3744 = n2570 & n3743;
  assign n3745 = ~n2687 & n2713;
  assign n3746 = ~n2687 & n2719;
  assign n3747 = ~n2571 & ~n3746;
  assign n3748 = ~n2429 & ~n3747;
  assign n3749 = ~n3745 & ~n3748;
  assign n3750 = ~n3744 & n3749;
  assign n3751 = n2429 & ~n2687;
  assign n3752 = n2523 & n3751;
  assign n3753 = n2687 & n2720;
  assign n3754 = ~n2711 & ~n3753;
  assign n3755 = ~n2691 & n3754;
  assign n3756 = n2429 & ~n3755;
  assign n3757 = ~n3752 & ~n3756;
  assign n3758 = n3750 & n3757;
  assign n3759 = ~n2628 & ~n3758;
  assign n3760 = ~n2713 & ~n2824;
  assign n3761 = n2687 & ~n3760;
  assign n3762 = ~n2702 & ~n3761;
  assign n3763 = n2628 & ~n3762;
  assign n3764 = ~n2687 & n2690;
  assign n3765 = ~n2800 & ~n3764;
  assign n3766 = ~n2630 & n3765;
  assign n3767 = ~n2429 & n2628;
  assign n3768 = ~n3766 & n3767;
  assign n3769 = ~n3763 & ~n3768;
  assign n3770 = n2429 & n2628;
  assign n3771 = ~n3747 & n3770;
  assign n3772 = ~n2523 & n3743;
  assign n3773 = ~n2702 & ~n3772;
  assign n3774 = ~n2429 & ~n3773;
  assign n3775 = ~n3771 & ~n3774;
  assign n3776 = n3769 & n3775;
  assign n3777 = ~n3759 & n3776;
  assign n3778 = pi070 & ~n454;
  assign n3779 = pi020 & n454;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = ~n449 & ~n3780;
  assign n3782 = pi020 & n449;
  assign n3783 = ~n3781 & ~n3782;
  assign n3784 = ~n446 & ~n3783;
  assign n3785 = pi152 & n446;
  assign n3786 = ~n3784 & ~n3785;
  assign n3787 = ~n3777 & n3786;
  assign n3788 = n3777 & ~n3786;
  assign po24 = n3787 | n3788;
  assign n3790 = pi154 & n446;
  assign n3791 = pi116 & ~n454;
  assign n3792 = pi029 & n454;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = ~n449 & ~n3793;
  assign n3795 = pi029 & n449;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = ~n446 & ~n3796;
  assign n3798 = ~n3790 & ~n3797;
  assign n3799 = ~n2289 & ~n2748;
  assign n3800 = ~n2240 & ~n3799;
  assign n3801 = n2069 & n2268;
  assign n3802 = n2128 & n2267;
  assign n3803 = n2240 & n3802;
  assign n3804 = ~n2345 & ~n3803;
  assign n3805 = ~n3801 & n3804;
  assign n3806 = ~n2759 & n3805;
  assign n3807 = ~n3800 & n3806;
  assign n3808 = ~n2284 & ~n2733;
  assign n3809 = n3807 & n3808;
  assign n3810 = ~n1955 & ~n3809;
  assign n3811 = ~n2264 & ~n2326;
  assign n3812 = ~n2248 & ~n2288;
  assign n3813 = ~n2240 & ~n3812;
  assign n3814 = n2240 & n2337;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = ~n2278 & n3815;
  assign n3817 = ~n2263 & n3816;
  assign n3818 = n3811 & n3817;
  assign n3819 = n1955 & ~n3818;
  assign n3820 = ~n3810 & ~n3819;
  assign n3821 = ~n2240 & n2264;
  assign n3822 = ~n2256 & ~n2733;
  assign n3823 = n2240 & ~n3822;
  assign n3824 = ~n2760 & ~n3823;
  assign n3825 = ~n3821 & n3824;
  assign n3826 = n3820 & n3825;
  assign n3827 = ~n3798 & n3826;
  assign n3828 = n3798 & ~n3826;
  assign po26 = n3827 | n3828;
  assign n3830 = pi033 & n449;
  assign n3831 = pi110 & ~n454;
  assign n3832 = pi033 & n454;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = ~n449 & ~n3833;
  assign n3835 = ~n3830 & ~n3834;
  assign n3836 = ~n446 & ~n3835;
  assign n3837 = pi156 & n446;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = ~n515 & ~n811;
  assign n3840 = n601 & ~n3839;
  assign n3841 = ~n576 & ~n823;
  assign n3842 = n606 & ~n3841;
  assign n3843 = ~n3840 & ~n3842;
  assign n3844 = ~n607 & ~n827;
  assign n3845 = n560 & ~n3844;
  assign n3846 = ~n634 & ~n670;
  assign n3847 = n579 & ~n3846;
  assign n3848 = ~n3845 & ~n3847;
  assign n3849 = n520 & ~n3419;
  assign n3850 = ~n675 & ~n774;
  assign n3851 = n540 & ~n3850;
  assign n3852 = ~n3849 & ~n3851;
  assign n3853 = ~n603 & ~n729;
  assign n3854 = n499 & ~n3853;
  assign n3855 = ~n645 & ~n856;
  assign n3856 = n464 & ~n3855;
  assign n3857 = ~n3854 & ~n3856;
  assign n3858 = n3852 & n3857;
  assign n3859 = n3848 & n3858;
  assign n3860 = n3843 & n3859;
  assign n3861 = n650 & ~n3427;
  assign n3862 = n684 & ~n3450;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~n548 & ~n747;
  assign n3865 = n673 & ~n3864;
  assign n3866 = n632 & ~n3417;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = ~n629 & ~n852;
  assign n3869 = n638 & ~n3868;
  assign n3870 = ~n495 & ~n832;
  assign n3871 = n643 & ~n3870;
  assign n3872 = ~n3869 & ~n3871;
  assign n3873 = n3867 & n3872;
  assign n3874 = ~n536 & ~n686;
  assign n3875 = n678 & ~n3874;
  assign n3876 = ~n639 & ~n793;
  assign n3877 = n613 & ~n3876;
  assign n3878 = ~n3875 & ~n3877;
  assign n3879 = n3873 & n3878;
  assign n3880 = n3863 & n3879;
  assign n3881 = n3860 & n3880;
  assign n3882 = po25 & n3881;
  assign n3883 = ~po25 & ~n3881;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = ~n621 & ~n679;
  assign n3886 = n464 & ~n3885;
  assign n3887 = ~n556 & ~n680;
  assign n3888 = n499 & ~n3887;
  assign n3889 = ~n3886 & ~n3888;
  assign n3890 = ~n675 & ~n685;
  assign n3891 = n601 & ~n3890;
  assign n3892 = ~n595 & ~n674;
  assign n3893 = n606 & ~n3892;
  assign n3894 = ~n3891 & ~n3893;
  assign n3895 = ~n645 & ~n721;
  assign n3896 = n520 & ~n3895;
  assign n3897 = ~n608 & ~n640;
  assign n3898 = n579 & ~n3897;
  assign n3899 = ~n3896 & ~n3898;
  assign n3900 = ~n515 & ~n568;
  assign n3901 = n540 & ~n3900;
  assign n3902 = ~n548 & ~n658;
  assign n3903 = n560 & ~n3902;
  assign n3904 = ~n3901 & ~n3903;
  assign n3905 = n3899 & n3904;
  assign n3906 = ~n487 & ~n507;
  assign n3907 = n678 & ~n3906;
  assign n3908 = ~n576 & ~n844;
  assign n3909 = n650 & ~n3908;
  assign n3910 = ~n3907 & ~n3909;
  assign n3911 = ~n587 & ~n644;
  assign n3912 = n638 & ~n3911;
  assign n3913 = ~n602 & ~n607;
  assign n3914 = n673 & ~n3913;
  assign n3915 = ~n3912 & ~n3914;
  assign n3916 = n3910 & n3915;
  assign n3917 = ~n603 & ~n855;
  assign n3918 = n684 & ~n3917;
  assign n3919 = ~n495 & ~n633;
  assign n3920 = n613 & ~n3919;
  assign n3921 = ~n528 & ~n639;
  assign n3922 = n643 & ~n3921;
  assign n3923 = ~n3920 & ~n3922;
  assign n3924 = ~n629 & ~n822;
  assign n3925 = n632 & ~n3924;
  assign n3926 = n3923 & ~n3925;
  assign n3927 = ~n3918 & n3926;
  assign n3928 = n3916 & n3927;
  assign n3929 = n3905 & n3928;
  assign n3930 = n3894 & n3929;
  assign n3931 = n3889 & n3930;
  assign n3932 = ~po09 & n3931;
  assign n3933 = po09 & ~n3931;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = ~n607 & ~n765;
  assign n3936 = n520 & ~n3935;
  assign n3937 = ~n634 & ~n852;
  assign n3938 = n499 & ~n3937;
  assign n3939 = ~n3936 & ~n3938;
  assign n3940 = ~n536 & ~n856;
  assign n3941 = n606 & ~n3940;
  assign n3942 = ~n495 & ~n797;
  assign n3943 = n560 & ~n3942;
  assign n3944 = ~n3941 & ~n3943;
  assign n3945 = ~n639 & ~n757;
  assign n3946 = n601 & ~n3945;
  assign n3947 = ~n576 & ~n747;
  assign n3948 = n464 & ~n3947;
  assign n3949 = ~n3946 & ~n3948;
  assign n3950 = n3944 & n3949;
  assign n3951 = ~n679 & ~n819;
  assign n3952 = n650 & ~n3951;
  assign n3953 = ~n603 & ~n774;
  assign n3954 = n638 & ~n3953;
  assign n3955 = ~n3952 & ~n3954;
  assign n3956 = ~n645 & ~n793;
  assign n3957 = n673 & ~n3956;
  assign n3958 = ~n675 & ~n827;
  assign n3959 = n643 & ~n3958;
  assign n3960 = ~n3957 & ~n3959;
  assign n3961 = n3955 & n3960;
  assign n3962 = ~n548 & ~n811;
  assign n3963 = n613 & ~n3962;
  assign n3964 = ~n515 & ~n798;
  assign n3965 = n632 & ~n3964;
  assign n3966 = ~n3963 & ~n3965;
  assign n3967 = ~n587 & ~n828;
  assign n3968 = n684 & ~n3967;
  assign n3969 = ~n670 & ~n823;
  assign n3970 = n678 & ~n3969;
  assign n3971 = ~n3968 & ~n3970;
  assign n3972 = n3966 & n3971;
  assign n3973 = n3961 & n3972;
  assign n3974 = ~n686 & ~n729;
  assign n3975 = n579 & ~n3974;
  assign n3976 = ~n629 & ~n832;
  assign n3977 = n540 & ~n3976;
  assign n3978 = ~n3975 & ~n3977;
  assign n3979 = n3973 & n3978;
  assign n3980 = n3950 & n3979;
  assign n3981 = n3939 & n3980;
  assign n3982 = ~po01 & ~n3981;
  assign n3983 = po01 & n3981;
  assign n3984 = ~n3982 & ~n3983;
  assign n3985 = ~n602 & ~n793;
  assign n3986 = n560 & ~n3985;
  assign n3987 = ~n568 & ~n832;
  assign n3988 = n601 & ~n3987;
  assign n3989 = ~n739 & ~n831;
  assign n3990 = n579 & ~n3989;
  assign n3991 = ~n3988 & ~n3990;
  assign n3992 = ~n819 & ~n844;
  assign n3993 = n606 & ~n3992;
  assign n3994 = n520 & ~n3483;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = n3991 & n3995;
  assign n3997 = ~n3986 & n3996;
  assign n3998 = n684 & ~n3472;
  assign n3999 = ~n658 & ~n797;
  assign n4000 = n673 & ~n3999;
  assign n4001 = ~n3998 & ~n4000;
  assign n4002 = ~n721 & ~n765;
  assign n4003 = n464 & ~n4002;
  assign n4004 = n4001 & ~n4003;
  assign n4005 = ~n528 & ~n827;
  assign n4006 = n613 & ~n4005;
  assign n4007 = ~n773 & ~n785;
  assign n4008 = n678 & ~n4007;
  assign n4009 = ~n4006 & ~n4008;
  assign n4010 = ~n828 & ~n855;
  assign n4011 = n499 & ~n4010;
  assign n4012 = n4009 & ~n4011;
  assign n4013 = n650 & ~n3487;
  assign n4014 = n632 & ~n3490;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = ~n633 & ~n811;
  assign n4017 = n643 & ~n4016;
  assign n4018 = ~n798 & ~n822;
  assign n4019 = n638 & ~n4018;
  assign n4020 = ~n4017 & ~n4019;
  assign n4021 = n4015 & n4020;
  assign n4022 = ~n685 & ~n757;
  assign n4023 = n540 & ~n4022;
  assign n4024 = n4021 & ~n4023;
  assign n4025 = n4012 & n4024;
  assign n4026 = n4004 & n4025;
  assign n4027 = n3997 & n4026;
  assign n4028 = po59 & ~n4027;
  assign n4029 = ~po59 & n4027;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = ~n729 & ~n828;
  assign n4032 = n673 & ~n4031;
  assign n4033 = ~n686 & ~n785;
  assign n4034 = n643 & ~n4033;
  assign n4035 = ~n765 & ~n856;
  assign n4036 = n638 & ~n4035;
  assign n4037 = ~n4034 & ~n4036;
  assign n4038 = n632 & ~n3908;
  assign n4039 = n4037 & ~n4038;
  assign n4040 = ~n4032 & n4039;
  assign n4041 = n520 & ~n3917;
  assign n4042 = ~n536 & ~n773;
  assign n4043 = n601 & ~n4042;
  assign n4044 = ~n4041 & ~n4043;
  assign n4045 = ~n757 & ~n774;
  assign n4046 = n606 & ~n4045;
  assign n4047 = ~n747 & ~n797;
  assign n4048 = n499 & ~n4047;
  assign n4049 = ~n4046 & ~n4048;
  assign n4050 = n4044 & n4049;
  assign n4051 = ~n670 & ~n831;
  assign n4052 = n613 & ~n4051;
  assign n4053 = ~n811 & ~n832;
  assign n4054 = n678 & ~n4053;
  assign n4055 = ~n4052 & ~n4054;
  assign n4056 = n650 & ~n3924;
  assign n4057 = n684 & ~n3895;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = ~n793 & ~n827;
  assign n4060 = n579 & ~n4059;
  assign n4061 = ~n798 & ~n852;
  assign n4062 = n464 & ~n4061;
  assign n4063 = ~n4060 & ~n4062;
  assign n4064 = ~n819 & ~n823;
  assign n4065 = n540 & ~n4064;
  assign n4066 = ~n634 & ~n739;
  assign n4067 = n560 & ~n4066;
  assign n4068 = ~n4065 & ~n4067;
  assign n4069 = n4063 & n4068;
  assign n4070 = n4058 & n4069;
  assign n4071 = n4055 & n4070;
  assign n4072 = n4050 & n4071;
  assign n4073 = n4040 & n4072;
  assign n4074 = po33 & ~n4073;
  assign n4075 = ~po33 & n4073;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~n4030 & n4076;
  assign n4078 = ~n3984 & n4077;
  assign n4079 = ~n3934 & n4078;
  assign n4080 = n632 & ~n2974;
  assign n4081 = ~n487 & ~n629;
  assign n4082 = n673 & ~n4081;
  assign n4083 = ~n556 & ~n576;
  assign n4084 = n643 & ~n4083;
  assign n4085 = ~n507 & ~n548;
  assign n4086 = n638 & ~n4085;
  assign n4087 = ~n4084 & ~n4086;
  assign n4088 = ~n595 & ~n639;
  assign n4089 = n499 & ~n4088;
  assign n4090 = n4087 & ~n4089;
  assign n4091 = ~n4082 & n4090;
  assign n4092 = ~n4080 & n4091;
  assign n4093 = ~n515 & ~n679;
  assign n4094 = n579 & ~n4093;
  assign n4095 = ~n536 & ~n644;
  assign n4096 = n560 & ~n4095;
  assign n4097 = ~n4094 & ~n4096;
  assign n4098 = n684 & ~n2962;
  assign n4099 = ~n603 & ~n674;
  assign n4100 = n613 & ~n4099;
  assign n4101 = ~n587 & ~n607;
  assign n4102 = n678 & ~n4101;
  assign n4103 = ~n4100 & ~n4102;
  assign n4104 = n650 & ~n2966;
  assign n4105 = n4103 & ~n4104;
  assign n4106 = ~n4098 & n4105;
  assign n4107 = n4097 & n4106;
  assign n4108 = ~n608 & ~n675;
  assign n4109 = n464 & ~n4108;
  assign n4110 = ~n621 & ~n634;
  assign n4111 = n601 & ~n4110;
  assign n4112 = n520 & ~n2985;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = ~n4109 & n4113;
  assign n4115 = ~n640 & ~n645;
  assign n4116 = n540 & ~n4115;
  assign n4117 = ~n495 & ~n680;
  assign n4118 = n606 & ~n4117;
  assign n4119 = ~n4116 & ~n4118;
  assign n4120 = n4114 & n4119;
  assign n4121 = n4107 & n4120;
  assign n4122 = n4092 & n4121;
  assign n4123 = po17 & n4122;
  assign n4124 = ~po17 & ~n4122;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = ~n3934 & ~n3984;
  assign n4127 = ~n4076 & n4126;
  assign n4128 = n4030 & n4127;
  assign n4129 = ~n4125 & n4128;
  assign n4130 = ~n4030 & ~n4076;
  assign n4131 = ~n3984 & n4130;
  assign n4132 = n3934 & n4131;
  assign n4133 = n3984 & ~n4030;
  assign n4134 = n4030 & n4076;
  assign n4135 = ~n3984 & n4134;
  assign n4136 = n3934 & n4135;
  assign n4137 = ~n4133 & ~n4136;
  assign n4138 = n4125 & ~n4137;
  assign n4139 = ~n4132 & ~n4138;
  assign n4140 = ~n3934 & n3984;
  assign n4141 = n4076 & n4140;
  assign n4142 = n4030 & n4141;
  assign n4143 = n4139 & ~n4142;
  assign n4144 = ~n4129 & n4143;
  assign n4145 = ~n4079 & n4144;
  assign n4146 = n4030 & ~n4076;
  assign n4147 = n3984 & n4146;
  assign n4148 = n3934 & n4147;
  assign n4149 = n4145 & ~n4148;
  assign n4150 = n3884 & ~n4149;
  assign n4151 = ~n3984 & n4146;
  assign n4152 = n4125 & n4151;
  assign n4153 = ~n3984 & n4076;
  assign n4154 = ~n3934 & ~n4030;
  assign n4155 = n3984 & ~n4076;
  assign n4156 = ~n4154 & ~n4155;
  assign n4157 = ~n4153 & n4156;
  assign n4158 = ~n4125 & ~n4157;
  assign n4159 = n3984 & n4134;
  assign n4160 = n3934 & n4159;
  assign n4161 = ~n4030 & n4127;
  assign n4162 = ~n3984 & n4030;
  assign n4163 = n4076 & n4162;
  assign n4164 = ~n3934 & n4163;
  assign n4165 = ~n4161 & ~n4164;
  assign n4166 = ~n3934 & n4147;
  assign n4167 = n4165 & ~n4166;
  assign n4168 = n3934 & n4078;
  assign n4169 = n4167 & ~n4168;
  assign n4170 = ~n4160 & n4169;
  assign n4171 = ~n4158 & n4170;
  assign n4172 = ~n4152 & n4171;
  assign n4173 = ~n3884 & ~n4172;
  assign n4174 = ~n4150 & ~n4173;
  assign n4175 = ~n3838 & n4174;
  assign n4176 = n3838 & ~n4174;
  assign po28 = n4175 | n4176;
  assign n4178 = pi158 & n446;
  assign n4179 = pi010 & n449;
  assign n4180 = pi122 & ~n454;
  assign n4181 = pi010 & n454;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n449 & ~n4182;
  assign n4184 = ~n4179 & ~n4183;
  assign n4185 = ~n446 & ~n4184;
  assign n4186 = ~n4178 & ~n4185;
  assign n4187 = n3517 & n3661;
  assign n4188 = ~n3635 & ~n4187;
  assign n4189 = n3416 & n3669;
  assign n4190 = ~n3366 & ~n3516;
  assign n4191 = ~n3594 & ~n4190;
  assign n4192 = ~n3575 & ~n4191;
  assign n4193 = ~n4189 & ~n4192;
  assign n4194 = n4188 & n4193;
  assign n4195 = n3314 & ~n4194;
  assign n4196 = n3517 & n3610;
  assign n4197 = n3366 & n3591;
  assign n4198 = ~n3580 & ~n4197;
  assign n4199 = ~n3575 & ~n4198;
  assign n4200 = ~n3667 & ~n3671;
  assign n4201 = ~n3366 & n3584;
  assign n4202 = n4200 & ~n4201;
  assign n4203 = n3575 & ~n4202;
  assign n4204 = ~n3645 & ~n4203;
  assign n4205 = ~n4199 & n4204;
  assign n4206 = ~n4196 & n4205;
  assign n4207 = ~n3314 & ~n4206;
  assign n4208 = ~n3518 & ~n3644;
  assign n4209 = n3366 & ~n4208;
  assign n4210 = ~n3366 & n3579;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = ~n3575 & ~n4211;
  assign n4213 = n3586 & ~n3667;
  assign n4214 = n3366 & ~n4213;
  assign n4215 = n3575 & n4214;
  assign n4216 = ~n4212 & ~n4215;
  assign n4217 = ~n4207 & n4216;
  assign n4218 = ~n4195 & n4217;
  assign n4219 = ~n4186 & n4218;
  assign n4220 = n4186 & ~n4218;
  assign po30 = n4219 | n4220;
  assign n4222 = pi160 & n446;
  assign n4223 = pi126 & ~n454;
  assign n4224 = pi012 & n454;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = ~n449 & ~n4225;
  assign n4227 = pi012 & n449;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = ~n446 & ~n4228;
  assign n4230 = ~n4222 & ~n4229;
  assign n4231 = n3416 & n3661;
  assign n4232 = n3466 & n4231;
  assign n4233 = ~n3645 & ~n4232;
  assign n4234 = ~n3517 & ~n3579;
  assign n4235 = n3366 & ~n4234;
  assign n4236 = ~n3583 & ~n4235;
  assign n4237 = ~n3575 & ~n4236;
  assign n4238 = ~n3366 & n3641;
  assign n4239 = ~n3585 & ~n4238;
  assign n4240 = n3366 & n3667;
  assign n4241 = n4239 & ~n4240;
  assign n4242 = n3575 & ~n4241;
  assign n4243 = ~n3614 & ~n4242;
  assign n4244 = ~n3595 & n4243;
  assign n4245 = ~n4237 & n4244;
  assign n4246 = ~n3601 & ~n3671;
  assign n4247 = n4245 & n4246;
  assign n4248 = n3314 & ~n4247;
  assign n4249 = ~n3416 & n3593;
  assign n4250 = n3366 & n3580;
  assign n4251 = ~n4249 & ~n4250;
  assign n4252 = n4208 & n4251;
  assign n4253 = n3575 & ~n4252;
  assign n4254 = ~n4197 & ~n4253;
  assign n4255 = ~n3314 & ~n4254;
  assign n4256 = ~n3314 & ~n3575;
  assign n4257 = ~n3366 & n3517;
  assign n4258 = ~n4238 & ~n4257;
  assign n4259 = ~n4240 & n4258;
  assign n4260 = n4256 & ~n4259;
  assign n4261 = ~n4255 & ~n4260;
  assign n4262 = ~n4248 & n4261;
  assign n4263 = n4233 & n4262;
  assign n4264 = n4230 & n4263;
  assign n4265 = ~n4230 & ~n4263;
  assign po32 = n4264 | n4265;
  assign n4267 = pi039 & n449;
  assign n4268 = pi094 & ~n454;
  assign n4269 = pi039 & n454;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = ~n449 & ~n4270;
  assign n4272 = ~n4267 & ~n4271;
  assign n4273 = ~n446 & ~n4272;
  assign n4274 = pi162 & n446;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = ~n2954 & n3220;
  assign n4277 = ~n3182 & n4276;
  assign n4278 = n2954 & n3216;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = ~n2954 & ~n3182;
  assign n4281 = n3197 & n4280;
  assign n4282 = n3189 & n3229;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = ~n3231 & n4283;
  assign n4285 = n3019 & n3196;
  assign n4286 = n3182 & n4285;
  assign n4287 = ~n3209 & ~n4286;
  assign n4288 = ~n3019 & n3200;
  assign n4289 = ~n3182 & n4288;
  assign n4290 = n4287 & ~n4289;
  assign n4291 = ~n3182 & n3220;
  assign n4292 = ~n3019 & ~n3196;
  assign n4293 = n3182 & n4292;
  assign n4294 = ~n3213 & ~n4293;
  assign n4295 = n2954 & ~n4294;
  assign n4296 = ~n4291 & ~n4295;
  assign n4297 = n4290 & n4296;
  assign n4298 = n4284 & n4297;
  assign n4299 = ~n2898 & ~n4298;
  assign n4300 = ~n3182 & n3190;
  assign n4301 = ~n3213 & ~n4288;
  assign n4302 = n3182 & ~n4301;
  assign n4303 = ~n4300 & ~n4302;
  assign n4304 = n3019 & ~n3196;
  assign n4305 = n3182 & n4304;
  assign n4306 = ~n3206 & ~n3210;
  assign n4307 = ~n4305 & n4306;
  assign n4308 = n2954 & ~n4307;
  assign n4309 = n3126 & ~n3182;
  assign n4310 = n3197 & n3207;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = ~n2954 & ~n4311;
  assign n4313 = ~n4308 & ~n4312;
  assign n4314 = n4303 & n4313;
  assign n4315 = n2898 & ~n4314;
  assign n4316 = ~n4299 & ~n4315;
  assign n4317 = n4279 & n4316;
  assign n4318 = ~n4275 & n4317;
  assign n4319 = n4275 & ~n4317;
  assign po34 = n4318 | n4319;
  assign n4321 = ~n2720 & ~n2813;
  assign n4322 = ~n3744 & n4321;
  assign n4323 = n3767 & ~n4322;
  assign n4324 = ~n2702 & ~n2815;
  assign n4325 = ~n2429 & ~n4324;
  assign n4326 = ~n4323 & ~n4325;
  assign n4327 = ~n2721 & ~n2798;
  assign n4328 = n2569 & n3743;
  assign n4329 = ~n2713 & ~n4328;
  assign n4330 = ~n2429 & ~n4329;
  assign n4331 = n4327 & ~n4330;
  assign n4332 = ~n2702 & n4331;
  assign n4333 = ~n2815 & n4332;
  assign n4334 = n2570 & n2687;
  assign n4335 = ~n2709 & ~n4334;
  assign n4336 = n2429 & ~n4335;
  assign n4337 = ~n2810 & ~n4336;
  assign n4338 = n4333 & n4337;
  assign n4339 = ~n2628 & ~n4338;
  assign n4340 = ~n2475 & n3751;
  assign n4341 = n2690 & n4340;
  assign n4342 = n2571 & ~n2687;
  assign n4343 = n2523 & n3743;
  assign n4344 = ~n2722 & ~n4343;
  assign n4345 = n2429 & ~n4344;
  assign n4346 = n2429 & n2570;
  assign n4347 = ~n2687 & n4346;
  assign n4348 = n2429 & ~n3760;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = ~n4345 & n4349;
  assign n4351 = ~n4342 & n4350;
  assign n4352 = ~n4341 & n4351;
  assign n4353 = n2628 & ~n4352;
  assign n4354 = ~n4339 & ~n4353;
  assign n4355 = n4326 & n4354;
  assign n4356 = pi091 & ~n454;
  assign n4357 = pi025 & n454;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = ~n449 & ~n4358;
  assign n4360 = pi025 & n449;
  assign n4361 = ~n4359 & ~n4360;
  assign n4362 = ~n446 & ~n4361;
  assign n4363 = pi164 & n446;
  assign n4364 = ~n4362 & ~n4363;
  assign n4365 = ~n4355 & ~n4364;
  assign n4366 = n4355 & n4364;
  assign po36 = n4365 | n4366;
  assign n4368 = pi166 & n446;
  assign n4369 = pi093 & ~n454;
  assign n4370 = pi018 & n454;
  assign n4371 = ~n4369 & ~n4370;
  assign n4372 = ~n449 & ~n4371;
  assign n4373 = pi018 & n449;
  assign n4374 = ~n4372 & ~n4373;
  assign n4375 = ~n446 & ~n4374;
  assign n4376 = ~n4368 & ~n4375;
  assign n4377 = ~n3202 & ~n4289;
  assign n4378 = ~n3191 & n4377;
  assign n4379 = ~n3199 & n4378;
  assign n4380 = n2954 & ~n4379;
  assign n4381 = n3182 & n3220;
  assign n4382 = n3182 & n3200;
  assign n4383 = ~n3185 & ~n4382;
  assign n4384 = ~n2954 & ~n4383;
  assign n4385 = ~n3196 & n4280;
  assign n4386 = ~n4384 & ~n4385;
  assign n4387 = ~n3190 & ~n3209;
  assign n4388 = n2954 & ~n4387;
  assign n4389 = n4386 & ~n4388;
  assign n4390 = ~n3236 & n4389;
  assign n4391 = ~n4381 & n4390;
  assign n4392 = ~n2898 & ~n4391;
  assign n4393 = ~n4380 & ~n4392;
  assign n4394 = n2898 & n3229;
  assign n4395 = n4292 & n4394;
  assign n4396 = ~n2954 & n3216;
  assign n4397 = ~n3197 & ~n4292;
  assign n4398 = ~n3182 & ~n4397;
  assign n4399 = n3019 & n3069;
  assign n4400 = n3182 & n4399;
  assign n4401 = ~n4398 & ~n4400;
  assign n4402 = ~n3201 & n4401;
  assign n4403 = n2954 & ~n4402;
  assign n4404 = ~n3211 & ~n4403;
  assign n4405 = ~n4396 & n4404;
  assign n4406 = n2898 & ~n4405;
  assign n4407 = ~n4395 & ~n4406;
  assign n4408 = n4393 & n4407;
  assign n4409 = ~n3237 & n4408;
  assign n4410 = n4376 & n4409;
  assign n4411 = ~n4376 & ~n4409;
  assign po38 = n4410 | n4411;
  assign n4413 = pi168 & n446;
  assign n4414 = pi066 & ~n454;
  assign n4415 = ~pi050 & n454;
  assign n4416 = ~n4414 & ~n4415;
  assign n4417 = ~n449 & ~n4416;
  assign n4418 = ~pi050 & n449;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = ~n446 & ~n4419;
  assign n4421 = ~n4413 & ~n4420;
  assign n4422 = ~n1269 & ~n1423;
  assign n4423 = n540 & ~n4422;
  assign n4424 = ~n1338 & ~n1503;
  assign n4425 = n684 & ~n4424;
  assign n4426 = ~n4423 & ~n4425;
  assign n4427 = ~n1463 & ~n1602;
  assign n4428 = n638 & ~n4427;
  assign n4429 = ~n1292 & ~n1491;
  assign n4430 = n613 & ~n4429;
  assign n4431 = ~n1287 & ~n1488;
  assign n4432 = n643 & ~n4431;
  assign n4433 = ~n4430 & ~n4432;
  assign n4434 = ~n1263 & ~n1507;
  assign n4435 = n520 & ~n4434;
  assign n4436 = n4433 & ~n4435;
  assign n4437 = ~n4428 & n4436;
  assign n4438 = n4426 & n4437;
  assign n4439 = ~n1373 & ~n1452;
  assign n4440 = n632 & ~n4439;
  assign n4441 = ~n1438 & ~n1594;
  assign n4442 = n579 & ~n4441;
  assign n4443 = ~n4440 & ~n4442;
  assign n4444 = ~n1328 & ~n1473;
  assign n4445 = n560 & ~n4444;
  assign n4446 = n4443 & ~n4445;
  assign n4447 = ~n1494 & ~n1579;
  assign n4448 = n464 & ~n4447;
  assign n4449 = ~n1412 & ~n1588;
  assign n4450 = n499 & ~n4449;
  assign n4451 = ~n1208 & ~n1402;
  assign n4452 = n650 & ~n4451;
  assign n4453 = ~n4450 & ~n4452;
  assign n4454 = ~n4448 & n4453;
  assign n4455 = n4446 & n4454;
  assign n4456 = ~n1361 & ~n1477;
  assign n4457 = n601 & ~n4456;
  assign n4458 = ~n1226 & ~n1426;
  assign n4459 = n673 & ~n4458;
  assign n4460 = ~n1499 & ~n1566;
  assign n4461 = n606 & ~n4460;
  assign n4462 = ~n1441 & ~n1556;
  assign n4463 = n678 & ~n4462;
  assign n4464 = ~n4461 & ~n4463;
  assign n4465 = ~n4459 & n4464;
  assign n4466 = ~n4457 & n4465;
  assign n4467 = n4455 & n4466;
  assign n4468 = n4438 & n4467;
  assign n4469 = po21 & n4468;
  assign n4470 = ~po21 & ~n4468;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = ~n1302 & ~n1412;
  assign n4473 = n560 & ~n4472;
  assign n4474 = ~n1226 & ~n1287;
  assign n4475 = n579 & ~n4474;
  assign n4476 = ~n4473 & ~n4475;
  assign n4477 = ~n1208 & ~n1556;
  assign n4478 = n540 & ~n4477;
  assign n4479 = ~n1373 & ~n1588;
  assign n4480 = n464 & ~n4479;
  assign n4481 = ~n4478 & ~n4480;
  assign n4482 = ~n1331 & ~n1499;
  assign n4483 = n601 & ~n4482;
  assign n4484 = ~n1361 & ~n1602;
  assign n4485 = n606 & ~n4484;
  assign n4486 = ~n4483 & ~n4485;
  assign n4487 = n4481 & n4486;
  assign n4488 = ~n1269 & ~n1292;
  assign n4489 = n678 & ~n4488;
  assign n4490 = ~n1245 & ~n1426;
  assign n4491 = n684 & ~n4490;
  assign n4492 = ~n4489 & ~n4491;
  assign n4493 = ~n1357 & ~n1438;
  assign n4494 = n643 & ~n4493;
  assign n4495 = ~n1366 & ~n1423;
  assign n4496 = n650 & ~n4495;
  assign n4497 = ~n4494 & ~n4496;
  assign n4498 = n4492 & n4497;
  assign n4499 = ~n1377 & ~n1441;
  assign n4500 = n613 & ~n4499;
  assign n4501 = ~n1365 & ~n1494;
  assign n4502 = n632 & ~n4501;
  assign n4503 = ~n4500 & ~n4502;
  assign n4504 = ~n1263 & ~n1566;
  assign n4505 = n638 & ~n4504;
  assign n4506 = ~n1338 & ~n1594;
  assign n4507 = n673 & ~n4506;
  assign n4508 = ~n4505 & ~n4507;
  assign n4509 = n4503 & n4508;
  assign n4510 = n4498 & n4509;
  assign n4511 = ~n1237 & ~n1463;
  assign n4512 = n520 & ~n4511;
  assign n4513 = ~n1328 & ~n1579;
  assign n4514 = n499 & ~n4513;
  assign n4515 = ~n4512 & ~n4514;
  assign n4516 = n4510 & n4515;
  assign n4517 = n4487 & n4516;
  assign n4518 = n4476 & n4517;
  assign n4519 = ~po37 & n4518;
  assign n4520 = po37 & ~n4518;
  assign n4521 = ~n4519 & ~n4520;
  assign n4522 = ~n1245 & ~n1499;
  assign n4523 = n632 & ~n4522;
  assign n4524 = ~n1208 & ~n1579;
  assign n4525 = n638 & ~n4524;
  assign n4526 = ~n4523 & ~n4525;
  assign n4527 = ~n1302 & ~n1556;
  assign n4528 = n643 & ~n4527;
  assign n4529 = ~n1377 & ~n1588;
  assign n4530 = n673 & ~n4529;
  assign n4531 = ~n4528 & ~n4530;
  assign n4532 = ~n1287 & ~n1361;
  assign n4533 = n678 & ~n4532;
  assign n4534 = ~n1310 & ~n1494;
  assign n4535 = n684 & ~n4534;
  assign n4536 = ~n4533 & ~n4535;
  assign n4537 = ~n1332 & ~n1463;
  assign n4538 = n650 & ~n4537;
  assign n4539 = ~n1331 & ~n1594;
  assign n4540 = n613 & ~n4539;
  assign n4541 = ~n4538 & ~n4540;
  assign n4542 = n4536 & n4541;
  assign n4543 = ~n1366 & ~n1412;
  assign n4544 = n520 & ~n4543;
  assign n4545 = ~n1226 & ~n1263;
  assign n4546 = n499 & ~n4545;
  assign n4547 = ~n4544 & ~n4546;
  assign n4548 = ~n1357 & ~n1566;
  assign n4549 = n540 & ~n4548;
  assign n4550 = ~n1269 & ~n1373;
  assign n4551 = n606 & ~n4550;
  assign n4552 = ~n4549 & ~n4551;
  assign n4553 = n4547 & n4552;
  assign n4554 = ~n1237 & ~n1438;
  assign n4555 = n560 & ~n4554;
  assign n4556 = ~n1292 & ~n1328;
  assign n4557 = n579 & ~n4556;
  assign n4558 = ~n4555 & ~n4557;
  assign n4559 = ~n1365 & ~n1441;
  assign n4560 = n601 & ~n4559;
  assign n4561 = ~n1338 & ~n1602;
  assign n4562 = n464 & ~n4561;
  assign n4563 = ~n4560 & ~n4562;
  assign n4564 = n4558 & n4563;
  assign n4565 = n4553 & n4564;
  assign n4566 = n4542 & n4565;
  assign n4567 = n4531 & n4566;
  assign n4568 = n4526 & n4567;
  assign n4569 = ~po63 & n4568;
  assign n4570 = po63 & ~n4568;
  assign n4571 = ~n4569 & ~n4570;
  assign n4572 = ~n4521 & ~n4571;
  assign n4573 = ~n1292 & ~n1366;
  assign n4574 = n540 & ~n4573;
  assign n4575 = ~n1349 & ~n1602;
  assign n4576 = n601 & ~n4575;
  assign n4577 = ~n4574 & ~n4576;
  assign n4578 = ~n1245 & ~n1287;
  assign n4579 = n673 & ~n4578;
  assign n4580 = ~n1226 & ~n1332;
  assign n4581 = n643 & ~n4580;
  assign n4582 = ~n1208 & ~n1377;
  assign n4583 = n678 & ~n4582;
  assign n4584 = ~n4581 & ~n4583;
  assign n4585 = ~n1372 & ~n1556;
  assign n4586 = n650 & ~n4585;
  assign n4587 = n4584 & ~n4586;
  assign n4588 = ~n4579 & n4587;
  assign n4589 = ~n1255 & ~n1594;
  assign n4590 = n684 & ~n4589;
  assign n4591 = ~n1269 & ~n1310;
  assign n4592 = n613 & ~n4591;
  assign n4593 = ~n1237 & ~n1361;
  assign n4594 = n638 & ~n4593;
  assign n4595 = ~n4592 & ~n4594;
  assign n4596 = ~n1200 & ~n1588;
  assign n4597 = n632 & ~n4596;
  assign n4598 = n4595 & ~n4597;
  assign n4599 = ~n4590 & n4598;
  assign n4600 = n4588 & n4599;
  assign n4601 = ~n1339 & ~n1566;
  assign n4602 = n520 & ~n4601;
  assign n4603 = ~n1338 & ~n1357;
  assign n4604 = n579 & ~n4603;
  assign n4605 = ~n4602 & ~n4604;
  assign n4606 = ~n1376 & ~n1579;
  assign n4607 = n560 & ~n4606;
  assign n4608 = ~n1302 & ~n1373;
  assign n4609 = n499 & ~n4608;
  assign n4610 = ~n4607 & ~n4609;
  assign n4611 = n4605 & n4610;
  assign n4612 = ~n1263 & ~n1331;
  assign n4613 = n606 & ~n4612;
  assign n4614 = ~n1328 & ~n1365;
  assign n4615 = n464 & ~n4614;
  assign n4616 = ~n4613 & ~n4615;
  assign n4617 = n4611 & n4616;
  assign n4618 = n4600 & n4617;
  assign n4619 = n4577 & n4618;
  assign n4620 = po13 & n4619;
  assign n4621 = ~po13 & ~n4619;
  assign n4622 = ~n4620 & ~n4621;
  assign n4623 = ~n1566 & ~n1594;
  assign n4624 = n678 & ~n4623;
  assign n4625 = ~n1269 & ~n1412;
  assign n4626 = n638 & ~n4625;
  assign n4627 = ~n4624 & ~n4626;
  assign n4628 = ~n1373 & ~n1491;
  assign n4629 = n601 & ~n4628;
  assign n4630 = n520 & ~n1647;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = ~n1441 & ~n1579;
  assign n4633 = n606 & ~n4632;
  assign n4634 = ~n1556 & ~n1588;
  assign n4635 = n579 & ~n4634;
  assign n4636 = ~n4633 & ~n4635;
  assign n4637 = n4631 & n4636;
  assign n4638 = ~n1438 & ~n1602;
  assign n4639 = n499 & ~n4638;
  assign n4640 = ~n1226 & ~n1499;
  assign n4641 = n464 & ~n4640;
  assign n4642 = ~n4639 & ~n4641;
  assign n4643 = ~n1287 & ~n1463;
  assign n4644 = n540 & ~n4643;
  assign n4645 = ~n1263 & ~n1488;
  assign n4646 = n560 & ~n4645;
  assign n4647 = ~n4644 & ~n4646;
  assign n4648 = n4642 & n4647;
  assign n4649 = n4637 & n4648;
  assign n4650 = n632 & ~n1649;
  assign n4651 = ~n1292 & ~n1494;
  assign n4652 = n673 & ~n4651;
  assign n4653 = ~n4650 & ~n4652;
  assign n4654 = n684 & ~n1659;
  assign n4655 = ~n1328 & ~n1423;
  assign n4656 = n643 & ~n4655;
  assign n4657 = ~n4654 & ~n4656;
  assign n4658 = n4653 & n4657;
  assign n4659 = ~n1361 & ~n1426;
  assign n4660 = n613 & ~n4659;
  assign n4661 = n650 & ~n1638;
  assign n4662 = ~n4660 & ~n4661;
  assign n4663 = n4658 & n4662;
  assign n4664 = n4649 & n4663;
  assign n4665 = n4627 & n4664;
  assign n4666 = ~po05 & n4665;
  assign n4667 = po05 & ~n4665;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = n4622 & n4668;
  assign n4670 = n4572 & n4669;
  assign n4671 = n4471 & n4670;
  assign n4672 = n4622 & ~n4668;
  assign n4673 = n4521 & n4672;
  assign n4674 = ~n4471 & n4673;
  assign n4675 = ~n1488 & ~n1503;
  assign n4676 = n606 & ~n4675;
  assign n4677 = ~n1477 & ~n1507;
  assign n4678 = n579 & ~n4677;
  assign n4679 = ~n4676 & ~n4678;
  assign n4680 = n684 & ~n4601;
  assign n4681 = ~n1218 & ~n1463;
  assign n4682 = n673 & ~n4681;
  assign n4683 = ~n4680 & ~n4682;
  assign n4684 = ~n1291 & ~n1412;
  assign n4685 = n613 & ~n4684;
  assign n4686 = ~n1279 & ~n1499;
  assign n4687 = n643 & ~n4686;
  assign n4688 = ~n4685 & ~n4687;
  assign n4689 = n4683 & n4688;
  assign n4690 = ~n1452 & ~n1473;
  assign n4691 = n678 & ~n4690;
  assign n4692 = ~n1426 & ~n1502;
  assign n4693 = n638 & ~n4692;
  assign n4694 = ~n4691 & ~n4693;
  assign n4695 = n650 & ~n4596;
  assign n4696 = n632 & ~n4585;
  assign n4697 = ~n4695 & ~n4696;
  assign n4698 = n4694 & n4697;
  assign n4699 = n4689 & n4698;
  assign n4700 = n4679 & n4699;
  assign n4701 = ~n1402 & ~n1491;
  assign n4702 = n499 & ~n4701;
  assign n4703 = ~n1394 & ~n1423;
  assign n4704 = n464 & ~n4703;
  assign n4705 = ~n4702 & ~n4704;
  assign n4706 = ~n1362 & ~n1438;
  assign n4707 = n601 & ~n4706;
  assign n4708 = n520 & ~n4589;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = ~n1268 & ~n1494;
  assign n4711 = n540 & ~n4710;
  assign n4712 = ~n1320 & ~n1441;
  assign n4713 = n560 & ~n4712;
  assign n4714 = ~n4711 & ~n4713;
  assign n4715 = n4709 & n4714;
  assign n4716 = n4705 & n4715;
  assign n4717 = n4700 & n4716;
  assign n4718 = po29 & n4717;
  assign n4719 = ~po29 & ~n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~n4622 & n4668;
  assign n4722 = n4521 & n4571;
  assign n4723 = ~n4572 & ~n4722;
  assign n4724 = n4721 & ~n4723;
  assign n4725 = ~n4571 & n4668;
  assign n4726 = ~n4572 & ~n4725;
  assign n4727 = ~n4622 & ~n4726;
  assign n4728 = ~n4521 & n4571;
  assign n4729 = ~n4668 & n4728;
  assign n4730 = ~n4727 & ~n4729;
  assign n4731 = ~n4471 & ~n4730;
  assign n4732 = ~n4724 & ~n4731;
  assign n4733 = ~n4622 & ~n4668;
  assign n4734 = n4521 & n4733;
  assign n4735 = n4622 & ~n4726;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = n4471 & ~n4736;
  assign n4738 = n4668 & n4728;
  assign n4739 = n4622 & n4738;
  assign n4740 = ~n4737 & ~n4739;
  assign n4741 = n4732 & n4740;
  assign n4742 = ~n4720 & ~n4741;
  assign n4743 = ~n4674 & ~n4742;
  assign n4744 = n4521 & ~n4571;
  assign n4745 = n4721 & n4744;
  assign n4746 = n4471 & n4745;
  assign n4747 = ~n4622 & n4728;
  assign n4748 = n4622 & n4722;
  assign n4749 = ~n4747 & ~n4748;
  assign n4750 = n4471 & ~n4749;
  assign n4751 = ~n4746 & ~n4750;
  assign n4752 = n4571 & n4672;
  assign n4753 = ~n4673 & ~n4752;
  assign n4754 = n4751 & n4753;
  assign n4755 = n4720 & ~n4754;
  assign n4756 = ~n4571 & n4622;
  assign n4757 = ~n4668 & n4722;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n4471 & n4720;
  assign n4760 = ~n4758 & n4759;
  assign n4761 = ~n4755 & ~n4760;
  assign n4762 = n4743 & n4761;
  assign n4763 = ~n4671 & n4762;
  assign n4764 = n4421 & n4763;
  assign n4765 = ~n4421 & ~n4763;
  assign po40 = n4764 | n4765;
  assign n4767 = n3934 & n4125;
  assign n4768 = n4153 & n4767;
  assign n4769 = ~n4128 & ~n4142;
  assign n4770 = ~n4078 & n4769;
  assign n4771 = n4125 & ~n4770;
  assign n4772 = ~n4768 & ~n4771;
  assign n4773 = ~n3934 & ~n4125;
  assign n4774 = n4133 & n4773;
  assign n4775 = n4772 & ~n4774;
  assign n4776 = n3984 & n4030;
  assign n4777 = ~n4125 & n4776;
  assign n4778 = n3934 & n4777;
  assign n4779 = ~n4132 & ~n4147;
  assign n4780 = ~n4125 & ~n4779;
  assign n4781 = ~n3984 & ~n4030;
  assign n4782 = ~n3934 & n4781;
  assign n4783 = n3984 & n4130;
  assign n4784 = n3934 & n4783;
  assign n4785 = ~n4782 & ~n4784;
  assign n4786 = n4125 & ~n4785;
  assign n4787 = ~n4128 & ~n4136;
  assign n4788 = ~n4786 & n4787;
  assign n4789 = ~n4780 & n4788;
  assign n4790 = n3884 & ~n4789;
  assign n4791 = n3934 & ~n4125;
  assign n4792 = n4146 & n4791;
  assign n4793 = ~n4148 & ~n4168;
  assign n4794 = n3934 & ~n3984;
  assign n4795 = ~n4030 & n4794;
  assign n4796 = n4125 & n4795;
  assign n4797 = ~n4076 & n4140;
  assign n4798 = ~n4030 & n4797;
  assign n4799 = ~n4796 & ~n4798;
  assign n4800 = n3984 & n4077;
  assign n4801 = ~n4164 & ~n4800;
  assign n4802 = ~n3934 & n4130;
  assign n4803 = n4801 & ~n4802;
  assign n4804 = ~n4125 & ~n4803;
  assign n4805 = n4799 & ~n4804;
  assign n4806 = n4793 & n4805;
  assign n4807 = ~n4792 & n4806;
  assign n4808 = ~n3884 & ~n4807;
  assign n4809 = ~n4790 & ~n4808;
  assign n4810 = ~n4778 & n4809;
  assign n4811 = n4775 & n4810;
  assign n4812 = pi096 & ~n454;
  assign n4813 = pi014 & n454;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = ~n449 & ~n4814;
  assign n4816 = pi014 & n449;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = ~n446 & ~n4817;
  assign n4819 = pi170 & n446;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~n4811 & n4820;
  assign n4822 = n4811 & ~n4820;
  assign po42 = n4821 | n4822;
  assign n4824 = pi172 & n446;
  assign n4825 = pi021 & n449;
  assign n4826 = pi117 & ~n454;
  assign n4827 = pi021 & n454;
  assign n4828 = ~n4826 & ~n4827;
  assign n4829 = ~n449 & ~n4828;
  assign n4830 = ~n4825 & ~n4829;
  assign n4831 = ~n446 & ~n4830;
  assign n4832 = ~n4824 & ~n4831;
  assign n4833 = ~n925 & n1144;
  assign n4834 = ~n1149 & ~n1153;
  assign n4835 = n925 & n1110;
  assign n4836 = ~n3707 & ~n4835;
  assign n4837 = n4834 & n4836;
  assign n4838 = n1106 & ~n4837;
  assign n4839 = ~n1106 & n1133;
  assign n4840 = n925 & n4839;
  assign n4841 = ~n1106 & n1155;
  assign n4842 = ~n3704 & ~n4841;
  assign n4843 = ~n925 & ~n4842;
  assign n4844 = ~n4840 & ~n4843;
  assign n4845 = ~n3705 & ~n3723;
  assign n4846 = n4844 & n4845;
  assign n4847 = ~n4838 & n4846;
  assign n4848 = ~n4833 & n4847;
  assign n4849 = n1046 & ~n4848;
  assign n4850 = n925 & n1153;
  assign n4851 = n925 & n3708;
  assign n4852 = ~n4850 & ~n4851;
  assign n4853 = ~n1106 & ~n4852;
  assign n4854 = ~n4849 & ~n4853;
  assign n4855 = ~n866 & n985;
  assign n4856 = ~n703 & n4855;
  assign n4857 = ~n987 & ~n1153;
  assign n4858 = n925 & n1107;
  assign n4859 = ~n925 & n1118;
  assign n4860 = ~n4858 & ~n4859;
  assign n4861 = n4857 & n4860;
  assign n4862 = ~n1106 & ~n4861;
  assign n4863 = n925 & n1143;
  assign n4864 = ~n1142 & ~n4863;
  assign n4865 = ~n1155 & n4864;
  assign n4866 = n1106 & ~n4865;
  assign n4867 = ~n3722 & ~n4866;
  assign n4868 = ~n4862 & n4867;
  assign n4869 = ~n4856 & n4868;
  assign n4870 = ~n1046 & ~n4869;
  assign n4871 = ~n1156 & ~n3723;
  assign n4872 = n1106 & ~n4871;
  assign n4873 = ~n4870 & ~n4872;
  assign n4874 = n4854 & n4873;
  assign n4875 = ~n4832 & n4874;
  assign n4876 = n4832 & ~n4874;
  assign po44 = n4875 | n4876;
  assign n4878 = pi040 & n449;
  assign n4879 = pi092 & ~n454;
  assign n4880 = pi040 & n454;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = ~n449 & ~n4881;
  assign n4883 = ~n4878 & ~n4882;
  assign n4884 = ~n446 & ~n4883;
  assign n4885 = pi174 & n446;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = n4720 & n4757;
  assign n4888 = n4622 & n4887;
  assign n4889 = ~n4668 & n4744;
  assign n4890 = n4471 & n4889;
  assign n4891 = ~n4521 & n4668;
  assign n4892 = n4622 & n4728;
  assign n4893 = ~n4891 & ~n4892;
  assign n4894 = n4471 & ~n4893;
  assign n4895 = ~n4890 & ~n4894;
  assign n4896 = n4720 & ~n4895;
  assign n4897 = ~n4888 & ~n4896;
  assign n4898 = ~n4668 & ~n4723;
  assign n4899 = ~n4622 & n4898;
  assign n4900 = ~n4471 & n4672;
  assign n4901 = n4728 & n4900;
  assign n4902 = ~n4471 & ~n4622;
  assign n4903 = n4738 & n4902;
  assign n4904 = ~n4901 & ~n4903;
  assign n4905 = n4669 & ~n4723;
  assign n4906 = ~n4571 & n4673;
  assign n4907 = ~n4745 & ~n4906;
  assign n4908 = ~n4905 & n4907;
  assign n4909 = n4904 & n4908;
  assign n4910 = n4471 & ~n4622;
  assign n4911 = ~n4668 & n4910;
  assign n4912 = n4571 & n4911;
  assign n4913 = n4909 & ~n4912;
  assign n4914 = ~n4899 & n4913;
  assign n4915 = ~n4720 & ~n4914;
  assign n4916 = ~n4622 & n4722;
  assign n4917 = n4668 & n4916;
  assign n4918 = ~n4521 & n4669;
  assign n4919 = ~n4917 & ~n4918;
  assign n4920 = n4471 & ~n4919;
  assign n4921 = ~n4521 & n4733;
  assign n4922 = ~n4571 & ~n4668;
  assign n4923 = ~n4521 & n4922;
  assign n4924 = n4668 & n4744;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = ~n4921 & n4925;
  assign n4927 = n4759 & ~n4926;
  assign n4928 = ~n4920 & ~n4927;
  assign n4929 = ~n4915 & n4928;
  assign n4930 = n4897 & n4929;
  assign n4931 = ~n4886 & n4930;
  assign n4932 = n4886 & ~n4930;
  assign po46 = n4931 | n4932;
  assign n4934 = pi176 & n446;
  assign n4935 = pi026 & n449;
  assign n4936 = pi074 & ~n454;
  assign n4937 = pi026 & n454;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = ~n449 & ~n4938;
  assign n4940 = ~n4935 & ~n4939;
  assign n4941 = ~n446 & ~n4940;
  assign n4942 = ~n4934 & ~n4941;
  assign n4943 = n1735 & n1879;
  assign n4944 = n1526 & ~n1799;
  assign n4945 = n1734 & n4944;
  assign n4946 = n1813 & n4945;
  assign n4947 = n1825 & n4944;
  assign n4948 = n1616 & n4947;
  assign n4949 = ~n4946 & ~n4948;
  assign n4950 = ~n4943 & n4949;
  assign n4951 = n1386 & ~n4950;
  assign n4952 = ~n1799 & n1829;
  assign n4953 = n1616 & n1799;
  assign n4954 = ~n1734 & n4953;
  assign n4955 = ~n4952 & ~n4954;
  assign n4956 = ~n1800 & n4955;
  assign n4957 = n1386 & ~n4956;
  assign n4958 = ~n1526 & n4957;
  assign n4959 = ~n1799 & n1830;
  assign n4960 = ~n1675 & n4953;
  assign n4961 = ~n4959 & ~n4960;
  assign n4962 = ~n1827 & n4961;
  assign n4963 = ~n1526 & ~n4962;
  assign n4964 = n1799 & n1837;
  assign n4965 = ~n1805 & ~n4964;
  assign n4966 = n1386 & ~n4965;
  assign n4967 = ~n4963 & ~n4966;
  assign n4968 = ~n4958 & n4967;
  assign n4969 = ~n4951 & n4968;
  assign n4970 = n1526 & n1825;
  assign n4971 = n1799 & n4970;
  assign n4972 = n1736 & ~n1799;
  assign n4973 = ~n1862 & ~n4972;
  assign n4974 = n1526 & ~n4973;
  assign n4975 = n1799 & n1829;
  assign n4976 = ~n1826 & ~n4975;
  assign n4977 = ~n4974 & n4976;
  assign n4978 = ~n4971 & n4977;
  assign n4979 = ~n1616 & n1806;
  assign n4980 = n1616 & n1817;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = n4978 & n4981;
  assign n4983 = ~n1386 & ~n4982;
  assign n4984 = n1526 & n1734;
  assign n4985 = n1804 & n4984;
  assign n4986 = ~n1616 & ~n1799;
  assign n4987 = n1526 & n4986;
  assign n4988 = n1736 & n4987;
  assign n4989 = ~n4985 & ~n4988;
  assign n4990 = ~n4983 & n4989;
  assign n4991 = n4969 & n4990;
  assign n4992 = ~n4942 & n4991;
  assign n4993 = n4942 & ~n4991;
  assign po48 = n4992 | n4993;
  assign n4995 = pi178 & n446;
  assign n4996 = pi065 & ~n454;
  assign n4997 = pi053 & n454;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = ~n449 & ~n4998;
  assign n5000 = pi053 & n449;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = ~n446 & ~n5001;
  assign n5003 = ~n4995 & ~n5002;
  assign n5004 = n1799 & n1826;
  assign n5005 = ~n1815 & ~n5004;
  assign n5006 = ~n1526 & ~n5005;
  assign n5007 = ~n4985 & ~n5006;
  assign n5008 = ~n1526 & ~n1799;
  assign n5009 = n1830 & n5008;
  assign n5010 = ~n1386 & ~n1526;
  assign n5011 = ~n1837 & ~n4952;
  assign n5012 = ~n1826 & n5011;
  assign n5013 = n5010 & ~n5012;
  assign n5014 = ~n5009 & ~n5013;
  assign n5015 = n1526 & n1837;
  assign n5016 = n1799 & n5015;
  assign n5017 = ~n1805 & ~n4988;
  assign n5018 = n1526 & n1839;
  assign n5019 = n5017 & ~n5018;
  assign n5020 = ~n4946 & n5019;
  assign n5021 = ~n1386 & ~n5020;
  assign n5022 = ~n5016 & ~n5021;
  assign n5023 = ~n1799 & n4970;
  assign n5024 = ~n1812 & ~n5023;
  assign n5025 = ~n5015 & n5024;
  assign n5026 = ~n1675 & n1804;
  assign n5027 = n1616 & n1734;
  assign n5028 = n1735 & ~n1799;
  assign n5029 = ~n5027 & ~n5028;
  assign n5030 = ~n1526 & ~n5029;
  assign n5031 = ~n5026 & ~n5030;
  assign n5032 = n5025 & n5031;
  assign n5033 = n1386 & ~n5032;
  assign n5034 = n5022 & ~n5033;
  assign n5035 = n5014 & n5034;
  assign n5036 = n5007 & n5035;
  assign n5037 = n5003 & n5036;
  assign n5038 = ~n5003 & ~n5036;
  assign po50 = n5037 | n5038;
  assign n5040 = ~n3211 & ~n4300;
  assign n5041 = n2954 & ~n5040;
  assign n5042 = ~n2898 & ~n2954;
  assign n5043 = n4292 & n5042;
  assign n5044 = ~n3019 & n3126;
  assign n5045 = ~n3182 & n5044;
  assign n5046 = n3069 & n3235;
  assign n5047 = ~n4304 & ~n5046;
  assign n5048 = ~n3190 & n5047;
  assign n5049 = n2954 & ~n5048;
  assign n5050 = ~n5045 & ~n5049;
  assign n5051 = ~n2898 & ~n5050;
  assign n5052 = ~n5043 & ~n5051;
  assign n5053 = n2954 & n4288;
  assign n5054 = n3205 & n3229;
  assign n5055 = ~n4310 & ~n5054;
  assign n5056 = ~n3182 & n4304;
  assign n5057 = n5055 & ~n5056;
  assign n5058 = ~n3202 & n5057;
  assign n5059 = ~n5053 & n5058;
  assign n5060 = n2898 & ~n5059;
  assign n5061 = ~n3182 & n3210;
  assign n5062 = ~n3202 & ~n5061;
  assign n5063 = ~n4289 & n5062;
  assign n5064 = ~n4293 & n5063;
  assign n5065 = ~n2954 & ~n5064;
  assign n5066 = ~n5060 & ~n5065;
  assign n5067 = n5052 & n5066;
  assign n5068 = ~n5041 & n5067;
  assign n5069 = pi064 & ~n454;
  assign n5070 = pi008 & n454;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = ~n449 & ~n5071;
  assign n5073 = pi008 & n449;
  assign n5074 = ~n5072 & ~n5073;
  assign n5075 = ~n446 & ~n5074;
  assign n5076 = pi180 & n446;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n5068 & n5077;
  assign n5079 = n5068 & ~n5077;
  assign po52 = n5078 | n5079;
  assign n5081 = ~n4077 & ~n4146;
  assign n5082 = n3984 & ~n5081;
  assign n5083 = ~n3934 & n5082;
  assign n5084 = ~n4161 & ~n5083;
  assign n5085 = n4030 & n4794;
  assign n5086 = ~n5082 & ~n5085;
  assign n5087 = ~n3934 & n4077;
  assign n5088 = ~n3934 & n4776;
  assign n5089 = ~n5087 & ~n5088;
  assign n5090 = n5086 & n5089;
  assign n5091 = ~n4125 & ~n5090;
  assign n5092 = n3934 & n4130;
  assign n5093 = ~n4160 & ~n5092;
  assign n5094 = n4125 & ~n5093;
  assign n5095 = ~n5091 & ~n5094;
  assign n5096 = n5084 & n5095;
  assign n5097 = n3884 & ~n5096;
  assign n5098 = ~n3934 & n4134;
  assign n5099 = ~n4798 & ~n5098;
  assign n5100 = n4125 & ~n5099;
  assign n5101 = n3934 & ~n5081;
  assign n5102 = n4125 & n5101;
  assign n5103 = ~n3984 & n4125;
  assign n5104 = ~n5081 & n5103;
  assign n5105 = ~n5102 & ~n5104;
  assign n5106 = ~n5100 & n5105;
  assign n5107 = ~n3884 & ~n5106;
  assign n5108 = ~n5097 & ~n5107;
  assign n5109 = ~n4125 & ~n5093;
  assign n5110 = ~n4164 & ~n5109;
  assign n5111 = ~n3884 & ~n5110;
  assign n5112 = pi006 & n449;
  assign n5113 = pi098 & ~n454;
  assign n5114 = pi006 & n454;
  assign n5115 = ~n5113 & ~n5114;
  assign n5116 = ~n449 & ~n5115;
  assign n5117 = ~n5112 & ~n5116;
  assign n5118 = ~n446 & ~n5117;
  assign n5119 = pi182 & n446;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = n4125 & n4164;
  assign n5122 = ~n4125 & ~n5084;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = ~n5120 & n5123;
  assign n5125 = ~n5111 & n5124;
  assign n5126 = n5108 & n5125;
  assign n5127 = ~n5097 & n5123;
  assign n5128 = ~n5111 & n5127;
  assign n5129 = ~n5107 & n5128;
  assign n5130 = n5120 & ~n5129;
  assign po54 = n5126 | n5130;
  assign n5132 = pi051 & n449;
  assign n5133 = pi089 & ~n454;
  assign n5134 = pi051 & n454;
  assign n5135 = ~n5133 & ~n5134;
  assign n5136 = ~n449 & ~n5135;
  assign n5137 = ~n5132 & ~n5136;
  assign n5138 = ~n446 & ~n5137;
  assign n5139 = pi184 & n446;
  assign n5140 = ~n5138 & ~n5139;
  assign n5141 = ~n4784 & ~n5088;
  assign n5142 = ~n4125 & ~n5141;
  assign n5143 = n4125 & n4128;
  assign n5144 = ~n5142 & ~n5143;
  assign n5145 = n3934 & n4155;
  assign n5146 = ~n5087 & ~n5145;
  assign n5147 = ~n4135 & n5146;
  assign n5148 = n4125 & ~n5147;
  assign n5149 = ~n3984 & n5101;
  assign n5150 = ~n4161 & ~n5149;
  assign n5151 = ~n4159 & n5150;
  assign n5152 = ~n4125 & ~n5151;
  assign n5153 = ~n3934 & n4800;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = ~n5148 & n5154;
  assign n5156 = n3884 & ~n5155;
  assign n5157 = n3934 & n4077;
  assign n5158 = ~n4131 & ~n5157;
  assign n5159 = n4125 & ~n5158;
  assign n5160 = ~n4142 & ~n5159;
  assign n5161 = ~n4128 & ~n4798;
  assign n5162 = ~n3934 & n4153;
  assign n5163 = ~n4155 & ~n5162;
  assign n5164 = ~n4135 & n5163;
  assign n5165 = ~n4125 & ~n5164;
  assign n5166 = n3934 & n4800;
  assign n5167 = ~n5165 & ~n5166;
  assign n5168 = n5161 & n5167;
  assign n5169 = n5160 & n5168;
  assign n5170 = ~n3884 & ~n5169;
  assign n5171 = ~n5156 & ~n5170;
  assign n5172 = n5144 & n5171;
  assign n5173 = ~n5140 & n5172;
  assign n5174 = n5140 & ~n5172;
  assign po56 = n5173 | n5174;
  assign n5176 = pi186 & n446;
  assign n5177 = pi073 & ~n454;
  assign n5178 = pi060 & n454;
  assign n5179 = ~n5177 & ~n5178;
  assign n5180 = ~n449 & ~n5179;
  assign n5181 = pi060 & n449;
  assign n5182 = ~n5180 & ~n5181;
  assign n5183 = ~n446 & ~n5182;
  assign n5184 = ~n5176 & ~n5183;
  assign n5185 = ~n4471 & n4622;
  assign n5186 = n4923 & n5185;
  assign n5187 = ~n4668 & n4756;
  assign n5188 = ~n4892 & ~n5187;
  assign n5189 = n4471 & ~n5188;
  assign n5190 = ~n4745 & ~n4903;
  assign n5191 = ~n5189 & n5190;
  assign n5192 = n4668 & n4910;
  assign n5193 = ~n4728 & n5192;
  assign n5194 = ~n4471 & ~n4721;
  assign n5195 = ~n4723 & n5194;
  assign n5196 = ~n5193 & ~n5195;
  assign n5197 = n5191 & n5196;
  assign n5198 = n4720 & ~n5197;
  assign n5199 = ~n4571 & n4669;
  assign n5200 = ~n4747 & ~n5199;
  assign n5201 = ~n4748 & ~n4757;
  assign n5202 = n5200 & n5201;
  assign n5203 = n4471 & ~n5202;
  assign n5204 = n4669 & n4744;
  assign n5205 = ~n5203 & ~n5204;
  assign n5206 = ~n4720 & ~n5205;
  assign n5207 = ~n4724 & ~n4892;
  assign n5208 = ~n4889 & n5207;
  assign n5209 = ~n4471 & ~n4720;
  assign n5210 = ~n5208 & n5209;
  assign n5211 = ~n4746 & ~n5210;
  assign n5212 = n4471 & n4729;
  assign n5213 = ~n4622 & n5212;
  assign n5214 = n5211 & ~n5213;
  assign n5215 = ~n5206 & n5214;
  assign n5216 = ~n5198 & n5215;
  assign n5217 = ~n5186 & n5216;
  assign n5218 = ~n5184 & n5217;
  assign n5219 = n5184 & ~n5217;
  assign po58 = n5218 | n5219;
  assign n5221 = n4572 & n4668;
  assign n5222 = ~n4729 & ~n5221;
  assign n5223 = n4471 & ~n5222;
  assign n5224 = ~n4890 & ~n4917;
  assign n5225 = ~n4738 & ~n4923;
  assign n5226 = ~n4916 & n5225;
  assign n5227 = ~n4471 & ~n5226;
  assign n5228 = n5224 & ~n5227;
  assign n5229 = ~n5223 & n5228;
  assign n5230 = ~n4720 & ~n5229;
  assign n5231 = n4622 & n4729;
  assign n5232 = ~n4622 & n4744;
  assign n5233 = ~n4748 & ~n5232;
  assign n5234 = ~n4471 & ~n5233;
  assign n5235 = ~n5231 & ~n5234;
  assign n5236 = n4471 & n4757;
  assign n5237 = ~n4738 & ~n5236;
  assign n5238 = n4925 & n5237;
  assign n5239 = ~n4622 & ~n5238;
  assign n5240 = n5235 & ~n5239;
  assign n5241 = n4720 & ~n5240;
  assign n5242 = n4668 & n4748;
  assign n5243 = ~n4906 & ~n5242;
  assign n5244 = n4471 & ~n5243;
  assign n5245 = ~n4471 & n4725;
  assign n5246 = n4622 & n5245;
  assign n5247 = ~n5244 & ~n5246;
  assign n5248 = ~n5241 & n5247;
  assign n5249 = ~n5230 & n5248;
  assign n5250 = pi095 & ~n454;
  assign n5251 = pi062 & n454;
  assign n5252 = ~n5250 & ~n5251;
  assign n5253 = ~n449 & ~n5252;
  assign n5254 = pi062 & n449;
  assign n5255 = ~n5253 & ~n5254;
  assign n5256 = ~n446 & ~n5255;
  assign n5257 = pi188 & n446;
  assign n5258 = ~n5256 & ~n5257;
  assign n5259 = ~n5249 & n5258;
  assign n5260 = n5247 & ~n5258;
  assign n5261 = ~n5241 & n5260;
  assign n5262 = ~n5230 & n5261;
  assign po60 = n5259 | n5262;
  assign n5264 = pi190 & n446;
  assign n5265 = pi028 & n449;
  assign n5266 = pi087 & ~n454;
  assign n5267 = pi028 & n454;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n449 & ~n5268;
  assign n5270 = ~n5265 & ~n5269;
  assign n5271 = ~n446 & ~n5270;
  assign n5272 = ~n5264 & ~n5271;
  assign n5273 = n1111 & n3715;
  assign n5274 = n925 & n1108;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = ~n1106 & n3705;
  assign n5277 = n5275 & ~n5276;
  assign n5278 = ~n1144 & ~n3721;
  assign n5279 = n1106 & ~n5278;
  assign n5280 = n4852 & ~n5279;
  assign n5281 = ~n925 & n1127;
  assign n5282 = n5280 & ~n5281;
  assign n5283 = n1046 & ~n5282;
  assign n5284 = n1106 & n1133;
  assign n5285 = ~n1111 & ~n1144;
  assign n5286 = ~n3694 & n5285;
  assign n5287 = ~n1106 & ~n5286;
  assign n5288 = ~n1142 & ~n3716;
  assign n5289 = ~n5287 & n5288;
  assign n5290 = n1157 & n5289;
  assign n5291 = ~n5284 & n5290;
  assign n5292 = ~n1046 & ~n5291;
  assign n5293 = ~n5283 & ~n5292;
  assign n5294 = n5277 & n5293;
  assign n5295 = ~n3719 & n5294;
  assign n5296 = ~n5272 & n5295;
  assign n5297 = n5272 & ~n5295;
  assign po62 = n5296 | n5297;
  assign po65 = 1'b1;
  assign po64 = pi361;
  assign po66 = po20;
  assign po67 = po36;
  assign po68 = po62;
  assign po69 = po16;
  assign po70 = po10;
  assign po71 = po58;
endmodule


