module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926, pi927, pi928, pi929, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288, po289, po290, po291, po292, po293, po294, po295, po296, po297, po298, po299, po300, po301, po302, po303, po304, po305, po306, po307, po308, po309, po310, po311, po312, po313, po314, po315, po316, po317, po318, po319, po320, po321, po322, po323, po324, po325, po326, po327, po328, po329, po330, po331, po332, po333, po334, po335, po336, po337, po338, po339, po340, po341, po342, po343, po344, po345, po346, po347, po348, po349, po350, po351, po352, po353, po354, po355, po356, po357, po358, po359, po360, po361, po362, po363, po364, po365, po366, po367, po368, po369, po370, po371, po372, po373, po374, po375, po376, po377, po378, po379, po380, po381, po382, po383, po384, po385, po386, po387, po388, po389, po390, po391, po392, po393, po394, po395, po396, po397, po398, po399, po400, po401, po402, po403, po404, po405, po406, po407, po408, po409, po410, po411, po412, po413, po414, po415, po416, po417, po418, po419, po420, po421, po422, po423, po424, po425, po426, po427, po428, po429, po430, po431, po432, po433, po434, po435, po436, po437, po438, po439, po440, po441, po442, po443, po444, po445, po446, po447, po448, po449, po450, po451, po452, po453, po454, po455, po456, po457, po458, po459, po460, po461, po462, po463, po464, po465, po466, po467, po468, po469, po470, po471, po472, po473, po474, po475, po476, po477, po478, po479, po480, po481, po482, po483, po484, po485, po486, po487, po488, po489, po490, po491, po492, po493, po494, po495, po496, po497, po498, po499, po500, po501, po502, po503, po504, po505, po506, po507, po508, po509, po510, po511, po512, po513, po514, po515, po516, po517, po518, po519, po520, po521, po522, po523, po524, po525, po526, po527, po528, po529, po530, po531, po532, po533, po534, po535, po536, po537, po538, po539, po540, po541, po542, po543, po544, po545, po546, po547, po548, po549, po550, po551, po552, po553, po554, po555, po556, po557, po558, po559, po560, po561, po562, po563, po564, po565, po566, po567, po568, po569, po570, po571, po572, po573, po574, po575, po576, po577, po578, po579, po580, po581, po582, po583, po584, po585, po586, po587, po588, po589, po590, po591, po592, po593, po594, po595, po596, po597, po598, po599, po600, po601, po602, po603, po604, po605, po606, po607, po608, po609, po610, po611, po612, po613, po614, po615, po616, po617, po618, po619, po620, po621, po622, po623, po624, po625, po626, po627, po628, po629, po630, po631, po632, po633, po634, po635, po636, po637, po638, po639, po640, po641, po642, po643, po644, po645, po646, po647, po648, po649, po650, po651, po652, po653, po654, po655, po656, po657, po658, po659, po660, po661, po662, po663, po664, po665, po666, po667, po668, po669, po670, po671, po672, po673, po674, po675, po676, po677, po678, po679, po680, po681, po682, po683, po684, po685, po686, po687, po688, po689, po690, po691, po692, po693, po694, po695, po696, po697, po698, po699, po700, po701, po702, po703, po704, po705, po706, po707, po708, po709, po710, po711, po712, po713, po714, po715, po716, po717, po718, po719, po720, po721, po722, po723, po724, po725, po726, po727, po728, po729, po730, po731, po732, po733, po734, po735, po736, po737, po738, po739, po740, po741, po742, po743, po744, po745, po746, po747, po748, po749, po750, po751, po752, po753, po754, po755, po756, po757, po758, po759, po760, po761, po762, po763, po764, po765, po766, po767, po768, po769, po770, po771, po772, po773, po774, po775, po776, po777, po778, po779, po780, po781, po782, po783, po784, po785, po786, po787, po788, po789, po790, po791, po792, po793, po794, po795, po796, po797, po798, po799, po800, po801, po802, po803, po804, po805, po806, po807, po808, po809, po810, po811, po812, po813, po814, po815, po816, po817, po818);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926, pi927, pi928, pi929;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257, po258, po259, po260, po261, po262, po263, po264, po265, po266, po267, po268, po269, po270, po271, po272, po273, po274, po275, po276, po277, po278, po279, po280, po281, po282, po283, po284, po285, po286, po287, po288, po289, po290, po291, po292, po293, po294, po295, po296, po297, po298, po299, po300, po301, po302, po303, po304, po305, po306, po307, po308, po309, po310, po311, po312, po313, po314, po315, po316, po317, po318, po319, po320, po321, po322, po323, po324, po325, po326, po327, po328, po329, po330, po331, po332, po333, po334, po335, po336, po337, po338, po339, po340, po341, po342, po343, po344, po345, po346, po347, po348, po349, po350, po351, po352, po353, po354, po355, po356, po357, po358, po359, po360, po361, po362, po363, po364, po365, po366, po367, po368, po369, po370, po371, po372, po373, po374, po375, po376, po377, po378, po379, po380, po381, po382, po383, po384, po385, po386, po387, po388, po389, po390, po391, po392, po393, po394, po395, po396, po397, po398, po399, po400, po401, po402, po403, po404, po405, po406, po407, po408, po409, po410, po411, po412, po413, po414, po415, po416, po417, po418, po419, po420, po421, po422, po423, po424, po425, po426, po427, po428, po429, po430, po431, po432, po433, po434, po435, po436, po437, po438, po439, po440, po441, po442, po443, po444, po445, po446, po447, po448, po449, po450, po451, po452, po453, po454, po455, po456, po457, po458, po459, po460, po461, po462, po463, po464, po465, po466, po467, po468, po469, po470, po471, po472, po473, po474, po475, po476, po477, po478, po479, po480, po481, po482, po483, po484, po485, po486, po487, po488, po489, po490, po491, po492, po493, po494, po495, po496, po497, po498, po499, po500, po501, po502, po503, po504, po505, po506, po507, po508, po509, po510, po511, po512, po513, po514, po515, po516, po517, po518, po519, po520, po521, po522, po523, po524, po525, po526, po527, po528, po529, po530, po531, po532, po533, po534, po535, po536, po537, po538, po539, po540, po541, po542, po543, po544, po545, po546, po547, po548, po549, po550, po551, po552, po553, po554, po555, po556, po557, po558, po559, po560, po561, po562, po563, po564, po565, po566, po567, po568, po569, po570, po571, po572, po573, po574, po575, po576, po577, po578, po579, po580, po581, po582, po583, po584, po585, po586, po587, po588, po589, po590, po591, po592, po593, po594, po595, po596, po597, po598, po599, po600, po601, po602, po603, po604, po605, po606, po607, po608, po609, po610, po611, po612, po613, po614, po615, po616, po617, po618, po619, po620, po621, po622, po623, po624, po625, po626, po627, po628, po629, po630, po631, po632, po633, po634, po635, po636, po637, po638, po639, po640, po641, po642, po643, po644, po645, po646, po647, po648, po649, po650, po651, po652, po653, po654, po655, po656, po657, po658, po659, po660, po661, po662, po663, po664, po665, po666, po667, po668, po669, po670, po671, po672, po673, po674, po675, po676, po677, po678, po679, po680, po681, po682, po683, po684, po685, po686, po687, po688, po689, po690, po691, po692, po693, po694, po695, po696, po697, po698, po699, po700, po701, po702, po703, po704, po705, po706, po707, po708, po709, po710, po711, po712, po713, po714, po715, po716, po717, po718, po719, po720, po721, po722, po723, po724, po725, po726, po727, po728, po729, po730, po731, po732, po733, po734, po735, po736, po737, po738, po739, po740, po741, po742, po743, po744, po745, po746, po747, po748, po749, po750, po751, po752, po753, po754, po755, po756, po757, po758, po759, po760, po761, po762, po763, po764, po765, po766, po767, po768, po769, po770, po771, po772, po773, po774, po775, po776, po777, po778, po779, po780, po781, po782, po783, po784, po785, po786, po787, po788, po789, po790, po791, po792, po793, po794, po795, po796, po797, po798, po799, po800, po801, po802, po803, po804, po805, po806, po807, po808, po809, po810, po811, po812, po813, po814, po815, po816, po817, po818;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546;
assign w0 = ~pi553 & pi554;
assign w1 = ~pi668 & w0;
assign w2 = (pi000 & ~w0) | (pi000 & w8690) | (~w0 & w8690);
assign w3 = ~pi559 & pi665;
assign w4 = ~pi550 & pi555;
assign w5 = pi550 & ~pi555;
assign w6 = ~pi551 & ~pi558;
assign w7 = pi551 & pi558;
assign w8 = ~w6 & ~w7;
assign w9 = ~pi390 & ~pi557;
assign w10 = pi390 & pi557;
assign w11 = ~w9 & ~w10;
assign w12 = ~pi552 & ~pi556;
assign w13 = pi552 & pi556;
assign w14 = ~w12 & ~w13;
assign w15 = ~w4 & ~w5;
assign w16 = ~w8 & w15;
assign w17 = ~w11 & ~w14;
assign w18 = w16 & w17;
assign w19 = w3 & ~w18;
assign w20 = ~pi555 & ~pi557;
assign w21 = ~pi556 & ~pi558;
assign w22 = w20 & w21;
assign w23 = pi559 & ~w22;
assign w24 = ~pi550 & ~pi551;
assign w25 = ~pi552 & w24;
assign w26 = ~w23 & ~w25;
assign w27 = ~w19 & ~w26;
assign w28 = ~w19 & w8691;
assign w29 = (pi000 & w19) | (pi000 & w8692) | (w19 & w8692);
assign w30 = w1 & ~w28;
assign w31 = (~w2 & ~w30) | (~w2 & w8693) | (~w30 & w8693);
assign w32 = pi005 & ~pi006;
assign w33 = pi006 & ~pi008;
assign w34 = ~w32 & ~w33;
assign w35 = ~pi005 & pi006;
assign w36 = pi007 & ~w35;
assign w37 = ~w34 & w36;
assign w38 = w34 & ~w36;
assign w39 = ~w37 & ~w38;
assign w40 = pi178 & ~pi195;
assign w41 = ~pi178 & pi195;
assign w42 = ~w40 & ~w41;
assign w43 = w39 & ~w42;
assign w44 = pi007 & pi008;
assign w45 = w35 & w44;
assign w46 = pi006 & pi007;
assign w47 = pi007 & ~pi008;
assign w48 = pi005 & pi008;
assign w49 = ~w33 & ~w47;
assign w50 = (~w46 & ~w49) | (~w46 & w8694) | (~w49 & w8694);
assign w51 = ~w45 & ~w50;
assign w52 = (pi190 & w50) | (pi190 & w8695) | (w50 & w8695);
assign w53 = w43 & ~w52;
assign w54 = ~w43 & w52;
assign w55 = ~w53 & ~w54;
assign w56 = pi006 & w48;
assign w57 = w48 & w8696;
assign w58 = ~pi007 & ~pi008;
assign w59 = w35 & w58;
assign w60 = ~w32 & w58;
assign w61 = ~w35 & ~w48;
assign w62 = ~w60 & w61;
assign w63 = ~w57 & ~w59;
assign w64 = ~w62 & w63;
assign w65 = pi195 & ~w64;
assign w66 = w32 & ~w58;
assign w67 = pi005 & ~w47;
assign w68 = ~w34 & ~w67;
assign w69 = ~w35 & ~w44;
assign w70 = ~w46 & ~w69;
assign w71 = ~w68 & ~w70;
assign w72 = ~w66 & w71;
assign w73 = (pi164 & ~w71) | (pi164 & w8697) | (~w71 & w8697);
assign w74 = w65 & ~w73;
assign w75 = ~w65 & w73;
assign w76 = ~w74 & ~w75;
assign w77 = w55 & ~w76;
assign w78 = ~w55 & w76;
assign w79 = ~w77 & ~w78;
assign w80 = pi164 & ~pi195;
assign w81 = ~pi164 & pi195;
assign w82 = ~w80 & ~w81;
assign w83 = w39 & ~w82;
assign w84 = (~w42 & w50) | (~w42 & w8698) | (w50 & w8698);
assign w85 = (pi190 & ~w71) | (pi190 & w8699) | (~w71 & w8699);
assign w86 = w84 & ~w85;
assign w87 = ~w84 & w85;
assign w88 = ~w86 & ~w87;
assign w89 = pi164 & ~w64;
assign w90 = w88 & ~w89;
assign w91 = ~w88 & w89;
assign w92 = ~w90 & ~w91;
assign w93 = w83 & w92;
assign w94 = ~w83 & ~w92;
assign w95 = ~w93 & ~w94;
assign w96 = ~w79 & ~w95;
assign w97 = w79 & w95;
assign w98 = ~w96 & ~w97;
assign w99 = ~pi553 & ~pi554;
assign w100 = ~pi668 & w99;
assign w101 = pi553 & ~pi554;
assign w102 = pi668 & w99;
assign w103 = ~w1 & ~w101;
assign w104 = ~w102 & w103;
assign w105 = w103 & w8700;
assign w106 = ~w23 & w104;
assign w107 = ~w19 & w106;
assign w108 = ~w105 & ~w107;
assign w109 = (pi673 & w107) | (pi673 & w8701) | (w107 & w8701);
assign w110 = (~w42 & ~w71) | (~w42 & w8702) | (~w71 & w8702);
assign w111 = (~w82 & w50) | (~w82 & w8703) | (w50 & w8703);
assign w112 = w110 & ~w111;
assign w113 = ~w110 & w111;
assign w114 = ~w112 & ~w113;
assign w115 = pi190 & w64;
assign w116 = ~pi164 & w39;
assign w117 = w115 & ~w116;
assign w118 = ~pi190 & ~w39;
assign w119 = ~w116 & ~w118;
assign w120 = ~w115 & ~w119;
assign w121 = ~w117 & ~w120;
assign w122 = w114 & ~w121;
assign w123 = ~w114 & w121;
assign w124 = ~w122 & ~w123;
assign w125 = (pi195 & ~w71) | (pi195 & w8704) | (~w71 & w8704);
assign w126 = pi178 & ~w64;
assign w127 = w125 & ~w126;
assign w128 = ~w125 & w126;
assign w129 = ~w127 & ~w128;
assign w130 = (pi164 & w50) | (pi164 & w8705) | (w50 & w8705);
assign w131 = pi190 & w39;
assign w132 = w130 & ~w131;
assign w133 = ~w130 & w131;
assign w134 = ~w132 & ~w133;
assign w135 = w129 & w134;
assign w136 = ~w129 & ~w134;
assign w137 = ~w135 & ~w136;
assign w138 = w124 & w137;
assign w139 = ~w124 & ~w137;
assign w140 = ~w138 & ~w139;
assign w141 = ~pi008 & w32;
assign w142 = pi007 & ~w69;
assign w143 = ~w56 & ~w141;
assign w144 = ~w142 & w143;
assign w145 = pi110 & ~w144;
assign w146 = pi007 & w68;
assign w147 = ~pi007 & pi008;
assign w148 = ~pi006 & ~w147;
assign w149 = ~w35 & ~w148;
assign w150 = (pi165 & w146) | (pi165 & w8706) | (w146 & w8706);
assign w151 = ~w145 & w150;
assign w152 = w145 & ~w150;
assign w153 = ~w151 & ~w152;
assign w154 = (pi132 & ~w71) | (pi132 & w8707) | (~w71 & w8707);
assign w155 = pi192 & ~w59;
assign w156 = ~w66 & w155;
assign w157 = ~w154 & ~w156;
assign w158 = w51 & w71;
assign w159 = ~w154 & ~w158;
assign w160 = w156 & ~w159;
assign w161 = ~w157 & ~w160;
assign w162 = w153 & ~w161;
assign w163 = ~w153 & w161;
assign w164 = ~w162 & ~w163;
assign w165 = w79 & w164;
assign w166 = ~w79 & ~w164;
assign w167 = ~w165 & ~w166;
assign w168 = ~w140 & ~w167;
assign w169 = w140 & w167;
assign w170 = ~w168 & ~w169;
assign w171 = w109 & w170;
assign w172 = pi165 & w39;
assign w173 = pi132 & ~w64;
assign w174 = w172 & ~w173;
assign w175 = ~w172 & w173;
assign w176 = ~w174 & ~w175;
assign w177 = (pi192 & ~w71) | (pi192 & w8708) | (~w71 & w8708);
assign w178 = (pi110 & w50) | (pi110 & w8709) | (w50 & w8709);
assign w179 = w177 & ~w178;
assign w180 = ~w177 & w178;
assign w181 = ~w179 & ~w180;
assign w182 = w176 & w181;
assign w183 = ~w176 & ~w181;
assign w184 = ~w182 & ~w183;
assign w185 = w137 & w184;
assign w186 = ~w137 & ~w184;
assign w187 = ~w185 & ~w186;
assign w188 = (pi165 & ~w71) | (pi165 & w8710) | (~w71 & w8710);
assign w189 = (pi132 & w50) | (pi132 & w8711) | (w50 & w8711);
assign w190 = w188 & ~w189;
assign w191 = ~w188 & w189;
assign w192 = ~w190 & ~w191;
assign w193 = pi192 & ~w144;
assign w194 = (pi110 & w146) | (pi110 & w8712) | (w146 & w8712);
assign w195 = w193 & ~w194;
assign w196 = ~w193 & w194;
assign w197 = ~w195 & ~w196;
assign w198 = w192 & w197;
assign w199 = ~w192 & ~w197;
assign w200 = ~w198 & ~w199;
assign w201 = ~w187 & w200;
assign w202 = (~w109 & ~w187) | (~w109 & w8713) | (~w187 & w8713);
assign w203 = ~w201 & w202;
assign w204 = (~w203 & ~w170) | (~w203 & w8714) | (~w170 & w8714);
assign w205 = w98 & w204;
assign w206 = ~w98 & ~w204;
assign w207 = ~w205 & ~w206;
assign w208 = (pi133 & w19) | (pi133 & w8715) | (w19 & w8715);
assign w209 = ~w19 & w8716;
assign w210 = ~w208 & ~w209;
assign w211 = w207 & ~w210;
assign w212 = ~w207 & w210;
assign w213 = ~w211 & ~w212;
assign w214 = (pi045 & w19) | (pi045 & w8717) | (w19 & w8717);
assign w215 = ~w19 & w8718;
assign w216 = ~w214 & ~w215;
assign w217 = ~w19 & w8719;
assign w218 = (~pi012 & w19) | (~pi012 & w8720) | (w19 & w8720);
assign w219 = ~w217 & ~w218;
assign w220 = w216 & ~w219;
assign w221 = ~w216 & w219;
assign w222 = ~w220 & ~w221;
assign w223 = w213 & ~w222;
assign w224 = ~w213 & w222;
assign w225 = ~w223 & ~w224;
assign w226 = ~w31 & ~w225;
assign w227 = (~pi000 & ~w0) | (~pi000 & w8721) | (~w0 & w8721);
assign w228 = (~w227 & ~w30) | (~w227 & w8722) | (~w30 & w8722);
assign w229 = w225 & w228;
assign w230 = ~w226 & ~w229;
assign w231 = w124 & w184;
assign w232 = ~w124 & ~w184;
assign w233 = ~w231 & ~w232;
assign w234 = w95 & w233;
assign w235 = (~w109 & w233) | (~w109 & w8723) | (w233 & w8723);
assign w236 = ~w234 & w235;
assign w237 = ~w170 & ~w236;
assign w238 = w170 & w236;
assign w239 = ~w237 & ~w238;
assign w240 = (pi192 & w146) | (pi192 & w8724) | (w146 & w8724);
assign w241 = pi110 & ~w72;
assign w242 = w240 & ~w241;
assign w243 = ~w240 & w241;
assign w244 = ~w242 & ~w243;
assign w245 = pi132 & w39;
assign w246 = (pi165 & w50) | (pi165 & w8725) | (w50 & w8725);
assign w247 = w245 & ~w246;
assign w248 = ~w245 & w246;
assign w249 = ~w247 & ~w248;
assign w250 = w244 & w249;
assign w251 = ~w244 & ~w249;
assign w252 = ~w250 & ~w251;
assign w253 = w239 & w252;
assign w254 = ~w239 & ~w252;
assign w255 = ~w253 & ~w254;
assign w256 = (pi134 & w19) | (pi134 & w8726) | (w19 & w8726);
assign w257 = ~w19 & w8727;
assign w258 = ~w256 & ~w257;
assign w259 = ~w255 & w258;
assign w260 = w255 & ~w258;
assign w261 = ~w259 & ~w260;
assign w262 = ~w19 & w8728;
assign w263 = (~pi044 & w19) | (~pi044 & w8729) | (w19 & w8729);
assign w264 = ~w262 & ~w263;
assign w265 = w261 & ~w264;
assign w266 = ~w261 & w264;
assign w267 = ~w265 & ~w266;
assign w268 = (~pi001 & ~w0) | (~pi001 & w8730) | (~w0 & w8730);
assign w269 = (pi013 & w19) | (pi013 & w8731) | (w19 & w8731);
assign w270 = ~w19 & w8732;
assign w271 = ~w269 & ~w270;
assign w272 = ~w19 & w8733;
assign w273 = (~pi001 & w19) | (~pi001 & w8734) | (w19 & w8734);
assign w274 = ~w272 & ~w273;
assign w275 = w271 & ~w274;
assign w276 = ~w271 & w274;
assign w277 = ~w275 & ~w276;
assign w278 = (~w268 & ~w277) | (~w268 & w8735) | (~w277 & w8735);
assign w279 = ~w267 & ~w278;
assign w280 = (~w268 & w277) | (~w268 & w8735) | (w277 & w8735);
assign w281 = w267 & ~w280;
assign w282 = ~w279 & ~w281;
assign w283 = (pi048 & w19) | (pi048 & w8736) | (w19 & w8736);
assign w284 = ~w19 & w8737;
assign w285 = ~w283 & ~w284;
assign w286 = ~w19 & w8738;
assign w287 = (~pi014 & w19) | (~pi014 & w8739) | (w19 & w8739);
assign w288 = ~w286 & ~w287;
assign w289 = w285 & ~w288;
assign w290 = ~w285 & w288;
assign w291 = ~w289 & ~w290;
assign w292 = w200 & ~w252;
assign w293 = ~w200 & w252;
assign w294 = ~w292 & ~w293;
assign w295 = w167 & w294;
assign w296 = ~w167 & ~w294;
assign w297 = ~w295 & ~w296;
assign w298 = ~w109 & w297;
assign w299 = ~w95 & ~w140;
assign w300 = w95 & w140;
assign w301 = ~w299 & ~w300;
assign w302 = w298 & w301;
assign w303 = ~w109 & ~w297;
assign w304 = ~w301 & w303;
assign w305 = ~w302 & ~w304;
assign w306 = ~w140 & ~w200;
assign w307 = (w109 & ~w140) | (w109 & w8740) | (~w140 & w8740);
assign w308 = ~w306 & w307;
assign w309 = ~w19 & w8741;
assign w310 = (~pi167 & w19) | (~pi167 & w8742) | (w19 & w8742);
assign w311 = ~w309 & ~w310;
assign w312 = w305 & w8743;
assign w313 = (w311 & ~w305) | (w311 & w8744) | (~w305 & w8744);
assign w314 = ~w312 & ~w313;
assign w315 = ~w291 & ~w314;
assign w316 = w291 & w314;
assign w317 = ~w315 & ~w316;
assign w318 = (~pi002 & w19) | (~pi002 & w8745) | (w19 & w8745);
assign w319 = ~w19 & w8746;
assign w320 = w1 & ~w318;
assign w321 = ~w319 & w320;
assign w322 = ~w317 & w321;
assign w323 = ~w314 & w8747;
assign w324 = w1 & w291;
assign w325 = (~pi002 & ~w0) | (~pi002 & w8748) | (~w0 & w8748);
assign w326 = (~w325 & ~w320) | (~w325 & w8749) | (~w320 & w8749);
assign w327 = (w326 & ~w314) | (w326 & w8750) | (~w314 & w8750);
assign w328 = ~w323 & w327;
assign w329 = ~w322 & ~w328;
assign w330 = (pi049 & w19) | (pi049 & w8751) | (w19 & w8751);
assign w331 = ~w19 & w8752;
assign w332 = ~w330 & ~w331;
assign w333 = ~w19 & w8753;
assign w334 = (~pi015 & w19) | (~pi015 & w8754) | (w19 & w8754);
assign w335 = ~w333 & ~w334;
assign w336 = w332 & ~w335;
assign w337 = ~w332 & w335;
assign w338 = ~w336 & ~w337;
assign w339 = w137 & ~w252;
assign w340 = ~w137 & w252;
assign w341 = ~w339 & ~w340;
assign w342 = w167 & w341;
assign w343 = ~w167 & ~w341;
assign w344 = ~w342 & ~w343;
assign w345 = w200 & w344;
assign w346 = ~w200 & ~w344;
assign w347 = ~w345 & ~w346;
assign w348 = w109 & w347;
assign w349 = w98 & w137;
assign w350 = ~w98 & ~w137;
assign w351 = ~w349 & ~w350;
assign w352 = ~w109 & w351;
assign w353 = ~w19 & w8755;
assign w354 = (~pi166 & w19) | (~pi166 & w8756) | (w19 & w8756);
assign w355 = ~w353 & ~w354;
assign w356 = ~w348 & w8757;
assign w357 = (w355 & w348) | (w355 & w8758) | (w348 & w8758);
assign w358 = ~w356 & ~w357;
assign w359 = ~w338 & w358;
assign w360 = w358 & w8759;
assign w361 = w1 & w338;
assign w362 = (pi003 & ~w0) | (pi003 & w8760) | (~w0 & w8760);
assign w363 = (~pi003 & w19) | (~pi003 & w8761) | (w19 & w8761);
assign w364 = ~w19 & w8762;
assign w365 = w1 & ~w363;
assign w366 = ~w364 & w365;
assign w367 = (~w362 & ~w365) | (~w362 & w8763) | (~w365 & w8763);
assign w368 = (w367 & w358) | (w367 & w8764) | (w358 & w8764);
assign w369 = ~w360 & w368;
assign w370 = w338 & ~w358;
assign w371 = ~w359 & ~w370;
assign w372 = w366 & ~w371;
assign w373 = ~w369 & ~w372;
assign w374 = (pi004 & ~w0) | (pi004 & w8765) | (~w0 & w8765);
assign w375 = ~w19 & w8766;
assign w376 = (pi004 & w19) | (pi004 & w8767) | (w19 & w8767);
assign w377 = w1 & ~w375;
assign w378 = (~w374 & ~w377) | (~w374 & w8768) | (~w377 & w8768);
assign w379 = w79 & w140;
assign w380 = ~w79 & ~w140;
assign w381 = ~w379 & ~w380;
assign w382 = w344 & w381;
assign w383 = ~w344 & ~w381;
assign w384 = ~w382 & ~w383;
assign w385 = (pi155 & w19) | (pi155 & w8769) | (w19 & w8769);
assign w386 = ~w19 & w8770;
assign w387 = ~w385 & ~w386;
assign w388 = w384 & ~w387;
assign w389 = ~w384 & w387;
assign w390 = ~w388 & ~w389;
assign w391 = w164 & w301;
assign w392 = ~w164 & ~w301;
assign w393 = ~w391 & ~w392;
assign w394 = ~w303 & w393;
assign w395 = ~w298 & ~w393;
assign w396 = ~w394 & ~w395;
assign w397 = ~w348 & ~w396;
assign w398 = w390 & w397;
assign w399 = ~w390 & ~w397;
assign w400 = ~w398 & ~w399;
assign w401 = (pi057 & w19) | (pi057 & w8771) | (w19 & w8771);
assign w402 = ~w19 & w8772;
assign w403 = ~w401 & ~w402;
assign w404 = ~w19 & w8773;
assign w405 = (~pi016 & w19) | (~pi016 & w8774) | (w19 & w8774);
assign w406 = ~w404 & ~w405;
assign w407 = w403 & ~w406;
assign w408 = ~w403 & w406;
assign w409 = ~w407 & ~w408;
assign w410 = w400 & w409;
assign w411 = ~w400 & ~w409;
assign w412 = ~w410 & ~w411;
assign w413 = ~w378 & ~w412;
assign w414 = (~pi004 & ~w0) | (~pi004 & w8775) | (~w0 & w8775);
assign w415 = (~w414 & ~w377) | (~w414 & w8776) | (~w377 & w8776);
assign w416 = w412 & w415;
assign w417 = ~w413 & ~w416;
assign w418 = (~w23 & w18) | (~w23 & w8777) | (w18 & w8777);
assign w419 = w100 & ~w418;
assign w420 = (pi199 & w19) | (pi199 & w8778) | (w19 & w8778);
assign w421 = ~w19 & w8779;
assign w422 = ~w420 & ~w421;
assign w423 = w419 & ~w422;
assign w424 = ~pi668 & w101;
assign w425 = w101 & w8780;
assign w426 = w99 & w8781;
assign w427 = pi668 & w101;
assign w428 = w101 & w8782;
assign w429 = ~w425 & ~w426;
assign w430 = ~w428 & w429;
assign w431 = ~w19 & w8783;
assign w432 = w101 & w8784;
assign w433 = w101 & w8785;
assign w434 = w99 & w8760;
assign w435 = ~w432 & ~w433;
assign w436 = ~w434 & w435;
assign w437 = (~w436 & w19) | (~w436 & w8786) | (w19 & w8786);
assign w438 = w108 & w8787;
assign w439 = ~w423 & w438;
assign w440 = pi565 & ~pi566;
assign w441 = pi563 & pi567;
assign w442 = w440 & w441;
assign w443 = pi658 & w442;
assign w444 = ~pi563 & ~pi567;
assign w445 = pi565 & pi566;
assign w446 = w444 & w445;
assign w447 = pi534 & w446;
assign w448 = ~pi565 & pi566;
assign w449 = ~pi563 & pi567;
assign w450 = w448 & w449;
assign w451 = pi593 & w450;
assign w452 = w441 & w445;
assign w453 = pi538 & w452;
assign w454 = w445 & w449;
assign w455 = pi539 & w454;
assign w456 = w441 & w448;
assign w457 = pi577 & w456;
assign w458 = ~pi565 & ~pi566;
assign w459 = w441 & w458;
assign w460 = pi570 & w459;
assign w461 = w440 & w444;
assign w462 = pi619 & w461;
assign w463 = pi563 & ~pi567;
assign w464 = w448 & w463;
assign w465 = pi598 & w464;
assign w466 = ~pi556 & pi558;
assign w467 = pi555 & ~pi557;
assign w468 = w466 & w467;
assign w469 = pi673 & ~w468;
assign w470 = w445 & w463;
assign w471 = pi533 & w470;
assign w472 = w444 & w448;
assign w473 = pi639 & w472;
assign w474 = w449 & w458;
assign w475 = pi573 & w474;
assign w476 = w458 & w463;
assign w477 = pi629 & w476;
assign w478 = w440 & w449;
assign w479 = pi622 & w478;
assign w480 = ~w443 & ~w447;
assign w481 = ~w451 & ~w453;
assign w482 = ~w455 & ~w457;
assign w483 = ~w460 & ~w462;
assign w484 = ~w465 & w469;
assign w485 = ~w471 & ~w473;
assign w486 = ~w475 & ~w477;
assign w487 = ~w479 & w486;
assign w488 = w484 & w485;
assign w489 = w482 & w483;
assign w490 = w480 & w481;
assign w491 = w489 & w490;
assign w492 = w487 & w488;
assign w493 = w491 & w492;
assign w494 = pi370 & w464;
assign w495 = pi320 & w472;
assign w496 = pi329 & w454;
assign w497 = pi278 & w478;
assign w498 = pi256 & w452;
assign w499 = pi284 & w474;
assign w500 = pi260 & w450;
assign w501 = pi391 & w476;
assign w502 = pi302 & w461;
assign w503 = pi361 & w456;
assign w504 = pi360 & w470;
assign w505 = pi362 & w459;
assign w506 = pi381 & w442;
assign w507 = pi311 & w446;
assign w508 = ~w469 & ~w494;
assign w509 = ~w495 & ~w496;
assign w510 = ~w497 & ~w498;
assign w511 = ~w499 & ~w500;
assign w512 = ~w501 & ~w502;
assign w513 = ~w503 & ~w504;
assign w514 = ~w505 & ~w506;
assign w515 = ~w507 & w514;
assign w516 = w512 & w513;
assign w517 = w510 & w511;
assign w518 = w508 & w509;
assign w519 = w517 & w518;
assign w520 = w515 & w516;
assign w521 = w519 & w520;
assign w522 = ~w493 & ~w521;
assign w523 = ~pi562 & pi673;
assign w524 = w22 & w523;
assign w525 = ~pi673 & w466;
assign w526 = ~pi562 & w467;
assign w527 = w525 & w526;
assign w528 = ~w524 & ~w527;
assign w529 = pi666 & pi673;
assign w530 = ~pi435 & ~w529;
assign w531 = ~pi666 & pi673;
assign w532 = ~w468 & w531;
assign w533 = ~w530 & ~w532;
assign w534 = w528 & w533;
assign w535 = w444 & w458;
assign w536 = ~pi568 & w535;
assign w537 = w534 & w536;
assign w538 = (~pi280 & w468) | (~pi280 & w8788) | (w468 & w8788);
assign w539 = ~w468 & w8789;
assign w540 = ~w538 & ~w539;
assign w541 = w534 & w8790;
assign w542 = w440 & w463;
assign w543 = (~pi398 & w468) | (~pi398 & w8791) | (w468 & w8791);
assign w544 = ~w468 & w8792;
assign w545 = w542 & ~w543;
assign w546 = ~w544 & w545;
assign w547 = (~w546 & w107) | (~w546 & w8793) | (w107 & w8793);
assign w548 = ~w541 & w547;
assign w549 = ~w522 & w548;
assign w550 = ~w439 & ~w549;
assign w551 = pi355 & w470;
assign w552 = pi316 & w472;
assign w553 = pi401 & w456;
assign w554 = pi342 & w459;
assign w555 = pi257 & w450;
assign w556 = pi276 & w474;
assign w557 = pi327 & w454;
assign w558 = pi378 & w442;
assign w559 = pi365 & w476;
assign w560 = pi371 & w464;
assign w561 = ~w469 & ~w551;
assign w562 = ~w552 & ~w553;
assign w563 = ~w554 & ~w555;
assign w564 = ~w556 & ~w557;
assign w565 = ~w558 & ~w559;
assign w566 = ~w560 & w565;
assign w567 = w563 & w564;
assign w568 = w561 & w562;
assign w569 = w567 & w568;
assign w570 = w566 & w569;
assign w571 = pi608 & w450;
assign w572 = pi466 & w454;
assign w573 = pi610 & w464;
assign w574 = pi572 & w474;
assign w575 = pi627 & w456;
assign w576 = pi467 & w470;
assign w577 = pi616 & w442;
assign w578 = pi654 & w472;
assign w579 = pi664 & w459;
assign w580 = pi597 & w476;
assign w581 = w469 & ~w571;
assign w582 = ~w572 & ~w573;
assign w583 = ~w574 & ~w575;
assign w584 = ~w576 & ~w577;
assign w585 = ~w578 & ~w579;
assign w586 = ~w580 & w585;
assign w587 = w583 & w584;
assign w588 = w581 & w582;
assign w589 = w587 & w588;
assign w590 = w586 & w589;
assign w591 = ~w570 & ~w590;
assign w592 = w535 & w8794;
assign w593 = w534 & w592;
assign w594 = pi637 & w478;
assign w595 = pi630 & w542;
assign w596 = pi468 & w446;
assign w597 = pi656 & w461;
assign w598 = pi469 & w452;
assign w599 = w469 & ~w594;
assign w600 = ~w595 & ~w596;
assign w601 = ~w597 & ~w598;
assign w602 = w600 & w601;
assign w603 = w599 & w602;
assign w604 = ~w593 & w603;
assign w605 = w535 & w8795;
assign w606 = w534 & w605;
assign w607 = pi275 & w478;
assign w608 = pi253 & w461;
assign w609 = pi309 & w446;
assign w610 = pi384 & w542;
assign w611 = pi326 & w452;
assign w612 = ~w469 & ~w607;
assign w613 = ~w608 & ~w609;
assign w614 = ~w610 & ~w611;
assign w615 = w613 & w614;
assign w616 = w612 & w615;
assign w617 = ~w606 & w616;
assign w618 = ~w604 & ~w617;
assign w619 = ~w591 & ~w618;
assign w620 = ~w108 & ~w619;
assign w621 = (pi196 & w19) | (pi196 & w8796) | (w19 & w8796);
assign w622 = ~w19 & w8797;
assign w623 = ~w621 & ~w622;
assign w624 = w419 & ~w623;
assign w625 = w101 & w8798;
assign w626 = w99 & w8799;
assign w627 = w101 & w8800;
assign w628 = ~w625 & ~w626;
assign w629 = ~w627 & w628;
assign w630 = (w629 & w19) | (w629 & w8801) | (w19 & w8801);
assign w631 = w99 & w8802;
assign w632 = w101 & w8803;
assign w633 = w101 & w8804;
assign w634 = ~w631 & ~w632;
assign w635 = ~w633 & w634;
assign w636 = ~w19 & w8805;
assign w637 = ~w630 & ~w636;
assign w638 = ~w624 & ~w637;
assign w639 = ~w620 & w638;
assign w640 = w535 & w8806;
assign w641 = w534 & w640;
assign w642 = pi403 & w476;
assign w643 = pi286 & w461;
assign w644 = pi271 & w478;
assign w645 = pi304 & w450;
assign w646 = pi343 & w442;
assign w647 = pi258 & w446;
assign w648 = pi323 & w454;
assign w649 = ~w469 & ~w642;
assign w650 = ~w643 & ~w644;
assign w651 = ~w645 & ~w646;
assign w652 = ~w647 & ~w648;
assign w653 = w651 & w652;
assign w654 = w649 & w650;
assign w655 = w653 & w654;
assign w656 = ~w641 & w655;
assign w657 = w535 & w8807;
assign w658 = w534 & w657;
assign w659 = pi521 & w446;
assign w660 = pi652 & w478;
assign w661 = pi659 & w450;
assign w662 = pi651 & w476;
assign w663 = pi587 & w442;
assign w664 = pi523 & w454;
assign w665 = pi586 & w461;
assign w666 = w469 & ~w659;
assign w667 = ~w660 & ~w661;
assign w668 = ~w662 & ~w663;
assign w669 = ~w664 & ~w665;
assign w670 = w668 & w669;
assign w671 = w666 & w667;
assign w672 = w670 & w671;
assign w673 = ~w658 & w672;
assign w674 = ~w656 & ~w673;
assign w675 = pi354 & w456;
assign w676 = pi303 & w452;
assign w677 = pi386 & w470;
assign w678 = pi377 & w459;
assign w679 = pi383 & w542;
assign w680 = pi392 & w472;
assign w681 = pi367 & w464;
assign w682 = pi265 & w474;
assign w683 = ~w469 & ~w675;
assign w684 = ~w676 & ~w677;
assign w685 = ~w678 & ~w679;
assign w686 = ~w680 & ~w681;
assign w687 = ~w682 & w686;
assign w688 = w684 & w685;
assign w689 = w683 & w688;
assign w690 = w687 & w689;
assign w691 = pi518 & w470;
assign w692 = pi588 & w456;
assign w693 = pi635 & w464;
assign w694 = pi606 & w459;
assign w695 = pi600 & w472;
assign w696 = pi596 & w542;
assign w697 = pi571 & w474;
assign w698 = pi520 & w452;
assign w699 = w469 & ~w691;
assign w700 = ~w692 & ~w693;
assign w701 = ~w694 & ~w695;
assign w702 = ~w696 & ~w697;
assign w703 = ~w698 & w702;
assign w704 = w700 & w701;
assign w705 = w699 & w704;
assign w706 = w703 & w705;
assign w707 = ~w690 & ~w706;
assign w708 = ~w674 & ~w707;
assign w709 = w109 & w708;
assign w710 = w639 & ~w709;
assign w711 = (pi827 & w23) | (pi827 & w8808) | (w23 & w8808);
assign w712 = ~w19 & w711;
assign w713 = pi202 & w3;
assign w714 = ~w18 & w713;
assign w715 = ~w23 & w8809;
assign w716 = ~w714 & ~w715;
assign w717 = ~w712 & w716;
assign w718 = w419 & ~w717;
assign w719 = w101 & w8810;
assign w720 = w99 & w8811;
assign w721 = w101 & w8812;
assign w722 = ~w719 & ~w720;
assign w723 = ~w721 & w722;
assign w724 = ~w19 & w8813;
assign w725 = w101 & w8814;
assign w726 = w99 & w8815;
assign w727 = w101 & w8816;
assign w728 = ~w725 & ~w726;
assign w729 = ~w727 & w728;
assign w730 = (w729 & w19) | (w729 & w8817) | (w19 & w8817);
assign w731 = ~w724 & ~w730;
assign w732 = ~w718 & ~w731;
assign w733 = w708 & w732;
assign w734 = w109 & ~w733;
assign w735 = ~w639 & ~w734;
assign w736 = ~w710 & ~w735;
assign w737 = ~w550 & w736;
assign w738 = w109 & w550;
assign w739 = w535 & w8818;
assign w740 = w534 & w739;
assign w741 = pi661 & w472;
assign w742 = pi618 & w542;
assign w743 = pi646 & w461;
assign w744 = pi649 & w474;
assign w745 = pi547 & w470;
assign w746 = pi614 & w476;
assign w747 = pi546 & w452;
assign w748 = w469 & ~w741;
assign w749 = ~w742 & ~w743;
assign w750 = ~w744 & ~w745;
assign w751 = ~w746 & ~w747;
assign w752 = w750 & w751;
assign w753 = w748 & w749;
assign w754 = w752 & w753;
assign w755 = ~w740 & w754;
assign w756 = w535 & w8819;
assign w757 = w534 & w756;
assign w758 = pi254 & w474;
assign w759 = pi321 & w472;
assign w760 = pi255 & w461;
assign w761 = pi375 & w476;
assign w762 = pi363 & w470;
assign w763 = pi308 & w452;
assign w764 = pi385 & w542;
assign w765 = ~w469 & ~w758;
assign w766 = ~w759 & ~w760;
assign w767 = ~w761 & ~w762;
assign w768 = ~w763 & ~w764;
assign w769 = w767 & w768;
assign w770 = w765 & w766;
assign w771 = w769 & w770;
assign w772 = ~w757 & w771;
assign w773 = ~w755 & ~w772;
assign w774 = pi632 & w464;
assign w775 = pi548 & w446;
assign w776 = pi589 & w456;
assign w777 = pi611 & w459;
assign w778 = pi662 & w450;
assign w779 = pi605 & w478;
assign w780 = pi549 & w454;
assign w781 = pi617 & w442;
assign w782 = w469 & ~w774;
assign w783 = ~w775 & ~w776;
assign w784 = ~w777 & ~w778;
assign w785 = ~w779 & ~w780;
assign w786 = ~w781 & w785;
assign w787 = w783 & w784;
assign w788 = w782 & w787;
assign w789 = w786 & w788;
assign w790 = pi331 & w454;
assign w791 = pi279 & w478;
assign w792 = pi261 & w450;
assign w793 = pi372 & w464;
assign w794 = pi382 & w442;
assign w795 = pi399 & w456;
assign w796 = pi344 & w459;
assign w797 = pi313 & w446;
assign w798 = ~w469 & ~w790;
assign w799 = ~w791 & ~w792;
assign w800 = ~w793 & ~w794;
assign w801 = ~w795 & ~w796;
assign w802 = ~w797 & w801;
assign w803 = w799 & w800;
assign w804 = w798 & w803;
assign w805 = w802 & w804;
assign w806 = ~w789 & ~w805;
assign w807 = ~w773 & ~w806;
assign w808 = ~w108 & ~w807;
assign w809 = (pi201 & w19) | (pi201 & w8820) | (w19 & w8820);
assign w810 = ~w19 & w8821;
assign w811 = ~w809 & ~w810;
assign w812 = w419 & ~w811;
assign w813 = w99 & w8765;
assign w814 = w101 & w8822;
assign w815 = w101 & w8823;
assign w816 = ~w813 & ~w814;
assign w817 = ~w815 & w816;
assign w818 = (w817 & w19) | (w817 & w8824) | (w19 & w8824);
assign w819 = w99 & w8825;
assign w820 = w101 & w8826;
assign w821 = w101 & w8827;
assign w822 = ~w819 & ~w820;
assign w823 = ~w821 & w822;
assign w824 = ~w19 & w8828;
assign w825 = ~w818 & ~w824;
assign w826 = ~w812 & ~w825;
assign w827 = ~w808 & w826;
assign w828 = ~w808 & w8829;
assign w829 = ~w738 & ~w828;
assign w830 = ~w736 & ~w829;
assign w831 = ~w737 & ~w830;
assign w832 = pi580 & w464;
assign w833 = pi579 & w459;
assign w834 = pi602 & w472;
assign w835 = pi525 & w454;
assign w836 = pi519 & w470;
assign w837 = pi657 & w476;
assign w838 = w469 & ~w832;
assign w839 = ~w833 & ~w834;
assign w840 = ~w835 & ~w836;
assign w841 = ~w837 & w840;
assign w842 = w838 & w839;
assign w843 = w841 & w842;
assign w844 = pi397 & w476;
assign w845 = pi407 & w470;
assign w846 = pi282 & w454;
assign w847 = pi345 & w459;
assign w848 = pi314 & w472;
assign w849 = pi395 & w464;
assign w850 = ~w469 & ~w844;
assign w851 = ~w845 & ~w846;
assign w852 = ~w847 & ~w848;
assign w853 = ~w849 & w852;
assign w854 = w850 & w851;
assign w855 = w853 & w854;
assign w856 = ~w843 & ~w855;
assign w857 = ~w468 & w8830;
assign w858 = (~pi269 & w468) | (~pi269 & w8831) | (w468 & w8831);
assign w859 = ~w857 & ~w858;
assign w860 = w534 & w8832;
assign w861 = pi285 & w461;
assign w862 = pi312 & w452;
assign w863 = pi273 & w478;
assign w864 = pi356 & w456;
assign w865 = pi267 & w474;
assign w866 = pi406 & w542;
assign w867 = pi305 & w450;
assign w868 = pi262 & w446;
assign w869 = pi317 & w442;
assign w870 = ~w469 & ~w861;
assign w871 = ~w862 & ~w863;
assign w872 = ~w864 & ~w865;
assign w873 = ~w866 & ~w867;
assign w874 = ~w868 & ~w869;
assign w875 = w873 & w874;
assign w876 = w871 & w872;
assign w877 = w870 & w876;
assign w878 = w875 & w877;
assign w879 = pi591 & w474;
assign w880 = pi524 & w452;
assign w881 = pi638 & w478;
assign w882 = pi650 & w442;
assign w883 = pi641 & w542;
assign w884 = pi603 & w450;
assign w885 = pi522 & w446;
assign w886 = pi626 & w461;
assign w887 = pi634 & w456;
assign w888 = w469 & ~w879;
assign w889 = ~w880 & ~w881;
assign w890 = ~w882 & ~w883;
assign w891 = ~w884 & ~w885;
assign w892 = ~w886 & ~w887;
assign w893 = w891 & w892;
assign w894 = w889 & w890;
assign w895 = w888 & w894;
assign w896 = w893 & w895;
assign w897 = ~w878 & ~w896;
assign w898 = ~w856 & ~w860;
assign w899 = ~w897 & w898;
assign w900 = ~w108 & ~w899;
assign w901 = (pi010 & w19) | (pi010 & w8833) | (w19 & w8833);
assign w902 = ~w19 & w8834;
assign w903 = ~w901 & ~w902;
assign w904 = w102 & ~w903;
assign w905 = (pi828 & w23) | (pi828 & w8835) | (w23 & w8835);
assign w906 = ~w19 & w905;
assign w907 = pi203 & w3;
assign w908 = ~w18 & w907;
assign w909 = ~w23 & w8836;
assign w910 = ~w908 & ~w909;
assign w911 = ~w906 & w910;
assign w912 = w419 & ~w911;
assign w913 = w101 & w8837;
assign w914 = w101 & w8838;
assign w915 = ~w913 & ~w914;
assign w916 = (w915 & w19) | (w915 & w8839) | (w19 & w8839);
assign w917 = w101 & w8840;
assign w918 = w101 & w8841;
assign w919 = ~w917 & ~w918;
assign w920 = ~w19 & w8842;
assign w921 = ~w916 & ~w920;
assign w922 = ~w912 & ~w921;
assign w923 = ~w904 & w922;
assign w924 = ~w900 & w923;
assign w925 = w827 & ~w924;
assign w926 = ~w827 & w924;
assign w927 = w109 & ~w925;
assign w928 = (w109 & w620) | (w109 & w8843) | (w620 & w8843);
assign w929 = (pi198 & w19) | (pi198 & w8844) | (w19 & w8844);
assign w930 = ~w19 & w8845;
assign w931 = ~w929 & ~w930;
assign w932 = w419 & ~w931;
assign w933 = w101 & w8846;
assign w934 = w99 & w8847;
assign w935 = w101 & w8848;
assign w936 = ~w933 & ~w934;
assign w937 = ~w935 & w936;
assign w938 = ~w19 & w8849;
assign w939 = w101 & w8850;
assign w940 = w99 & w8851;
assign w941 = w101 & w8852;
assign w942 = ~w939 & ~w940;
assign w943 = ~w941 & w942;
assign w944 = (~w943 & w19) | (~w943 & w8853) | (w19 & w8853);
assign w945 = w108 & w8854;
assign w946 = ~w932 & w945;
assign w947 = pi578 & w464;
assign w948 = pi645 & w461;
assign w949 = pi655 & w476;
assign w950 = pi585 & w456;
assign w951 = pi612 & w474;
assign w952 = pi575 & w478;
assign w953 = pi613 & w542;
assign w954 = pi530 & w454;
assign w955 = pi590 & w472;
assign w956 = pi531 & w470;
assign w957 = pi609 & w442;
assign w958 = pi544 & w452;
assign w959 = pi543 & w446;
assign w960 = pi592 & w450;
assign w961 = pi628 & w459;
assign w962 = w469 & ~w947;
assign w963 = ~w948 & ~w949;
assign w964 = ~w950 & ~w951;
assign w965 = ~w952 & ~w953;
assign w966 = ~w954 & ~w955;
assign w967 = ~w956 & ~w957;
assign w968 = ~w958 & ~w959;
assign w969 = ~w960 & ~w961;
assign w970 = w968 & w969;
assign w971 = w966 & w967;
assign w972 = w964 & w965;
assign w973 = w962 & w963;
assign w974 = w972 & w973;
assign w975 = w970 & w971;
assign w976 = w974 & w975;
assign w977 = pi358 & w470;
assign w978 = pi369 & w464;
assign w979 = pi380 & w442;
assign w980 = pi297 & w452;
assign w981 = pi301 & w461;
assign w982 = pi351 & w459;
assign w983 = pi259 & w450;
assign w984 = pi328 & w474;
assign w985 = pi318 & w472;
assign w986 = pi402 & w542;
assign w987 = pi393 & w476;
assign w988 = pi263 & w446;
assign w989 = pi359 & w456;
assign w990 = pi283 & w454;
assign w991 = pi325 & w478;
assign w992 = ~w469 & ~w977;
assign w993 = ~w978 & ~w979;
assign w994 = ~w980 & ~w981;
assign w995 = ~w982 & ~w983;
assign w996 = ~w984 & ~w985;
assign w997 = ~w986 & ~w987;
assign w998 = ~w988 & ~w989;
assign w999 = ~w990 & ~w991;
assign w1000 = w998 & w999;
assign w1001 = w996 & w997;
assign w1002 = w994 & w995;
assign w1003 = w992 & w993;
assign w1004 = w1002 & w1003;
assign w1005 = w1000 & w1001;
assign w1006 = w1004 & w1005;
assign w1007 = ~w976 & ~w1006;
assign w1008 = (~pi277 & w468) | (~pi277 & w8855) | (w468 & w8855);
assign w1009 = ~w468 & w8856;
assign w1010 = ~w1008 & ~w1009;
assign w1011 = w534 & w8857;
assign w1012 = ~w108 & ~w1011;
assign w1013 = ~w1007 & w1012;
assign w1014 = ~w946 & ~w1013;
assign w1015 = ~w109 & ~w1014;
assign w1016 = ~w928 & ~w1015;
assign w1017 = (w1016 & ~w927) | (w1016 & w8858) | (~w927 & w8858);
assign w1018 = w927 & w8859;
assign w1019 = ~w1017 & ~w1018;
assign w1020 = w831 & w1019;
assign w1021 = ~w831 & ~w1019;
assign w1022 = ~w1020 & ~w1021;
assign w1023 = w736 & ~w827;
assign w1024 = w109 & w807;
assign w1025 = (~w1024 & ~w924) | (~w1024 & w8860) | (~w924 & w8860);
assign w1026 = ~w736 & ~w1025;
assign w1027 = ~w1023 & ~w1026;
assign w1028 = w535 & w8861;
assign w1029 = w534 & w1028;
assign w1030 = pi574 & w476;
assign w1031 = pi620 & w459;
assign w1032 = pi535 & w470;
assign w1033 = pi595 & w456;
assign w1034 = pi648 & w478;
assign w1035 = pi527 & w454;
assign w1036 = pi643 & w442;
assign w1037 = w469 & ~w1030;
assign w1038 = ~w1031 & ~w1032;
assign w1039 = ~w1033 & ~w1034;
assign w1040 = ~w1035 & ~w1036;
assign w1041 = w1039 & w1040;
assign w1042 = w1037 & w1038;
assign w1043 = w1041 & w1042;
assign w1044 = ~w1029 & w1043;
assign w1045 = w535 & w8862;
assign w1046 = w534 & w1045;
assign w1047 = pi400 & w470;
assign w1048 = pi374 & w442;
assign w1049 = pi376 & w459;
assign w1050 = pi299 & w478;
assign w1051 = pi353 & w456;
assign w1052 = pi352 & w476;
assign w1053 = pi264 & w454;
assign w1054 = ~w469 & ~w1047;
assign w1055 = ~w1048 & ~w1049;
assign w1056 = ~w1050 & ~w1051;
assign w1057 = ~w1052 & ~w1053;
assign w1058 = w1056 & w1057;
assign w1059 = w1054 & w1055;
assign w1060 = w1058 & w1059;
assign w1061 = ~w1046 & w1060;
assign w1062 = ~w1044 & ~w1061;
assign w1063 = pi623 & w464;
assign w1064 = pi582 & w450;
assign w1065 = pi541 & w446;
assign w1066 = pi540 & w452;
assign w1067 = pi599 & w472;
assign w1068 = pi583 & w542;
assign w1069 = pi569 & w474;
assign w1070 = pi604 & w461;
assign w1071 = w469 & ~w1063;
assign w1072 = ~w1064 & ~w1065;
assign w1073 = ~w1066 & ~w1067;
assign w1074 = ~w1068 & ~w1069;
assign w1075 = ~w1070 & w1074;
assign w1076 = w1072 & w1073;
assign w1077 = w1071 & w1076;
assign w1078 = w1075 & w1077;
assign w1079 = pi266 & w452;
assign w1080 = pi330 & w461;
assign w1081 = pi408 & w542;
assign w1082 = pi366 & w464;
assign w1083 = pi307 & w450;
assign w1084 = pi373 & w472;
assign w1085 = pi310 & w474;
assign w1086 = pi306 & w446;
assign w1087 = ~w469 & ~w1079;
assign w1088 = ~w1080 & ~w1081;
assign w1089 = ~w1082 & ~w1083;
assign w1090 = ~w1084 & ~w1085;
assign w1091 = ~w1086 & w1090;
assign w1092 = w1088 & w1089;
assign w1093 = w1087 & w1092;
assign w1094 = w1091 & w1093;
assign w1095 = ~w1078 & ~w1094;
assign w1096 = ~w1062 & ~w1095;
assign w1097 = ~w108 & ~w1096;
assign w1098 = (pi200 & w19) | (pi200 & w8863) | (w19 & w8863);
assign w1099 = ~w19 & w8864;
assign w1100 = ~w1098 & ~w1099;
assign w1101 = w419 & ~w1100;
assign w1102 = w101 & w8865;
assign w1103 = w99 & w8866;
assign w1104 = w101 & w8867;
assign w1105 = ~w1102 & ~w1103;
assign w1106 = ~w1104 & w1105;
assign w1107 = (w1106 & w19) | (w1106 & w8868) | (w19 & w8868);
assign w1108 = w101 & w8869;
assign w1109 = w99 & w8870;
assign w1110 = w101 & w8871;
assign w1111 = ~w1108 & ~w1109;
assign w1112 = ~w1110 & w1111;
assign w1113 = ~w19 & w8872;
assign w1114 = ~w1107 & ~w1113;
assign w1115 = ~w1101 & ~w1114;
assign w1116 = ~w1097 & w1115;
assign w1117 = ~w1014 & ~w1116;
assign w1118 = w1014 & w1116;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = w109 & w924;
assign w1121 = (pi197 & w19) | (pi197 & w8873) | (w19 & w8873);
assign w1122 = ~w19 & w8874;
assign w1123 = ~w1121 & ~w1122;
assign w1124 = w419 & ~w1123;
assign w1125 = w101 & w8875;
assign w1126 = w99 & w8876;
assign w1127 = w101 & w8877;
assign w1128 = ~w1125 & ~w1126;
assign w1129 = ~w1127 & w1128;
assign w1130 = ~w19 & w8878;
assign w1131 = w101 & w8879;
assign w1132 = w101 & w8880;
assign w1133 = w99 & w8690;
assign w1134 = ~w1131 & ~w1132;
assign w1135 = ~w1133 & w1134;
assign w1136 = (~w1135 & w19) | (~w1135 & w8881) | (w19 & w8881);
assign w1137 = w108 & w8882;
assign w1138 = ~w1124 & w1137;
assign w1139 = pi633 & w542;
assign w1140 = pi631 & w461;
assign w1141 = pi644 & w450;
assign w1142 = pi510 & w454;
assign w1143 = pi621 & w476;
assign w1144 = pi509 & w446;
assign w1145 = pi576 & w456;
assign w1146 = pi581 & w459;
assign w1147 = pi493 & w452;
assign w1148 = pi607 & w478;
assign w1149 = pi625 & w464;
assign w1150 = w469 & ~w1139;
assign w1151 = ~w1140 & ~w1141;
assign w1152 = ~w1142 & ~w1143;
assign w1153 = ~w1144 & ~w1145;
assign w1154 = ~w1146 & ~w1147;
assign w1155 = ~w1148 & ~w1149;
assign w1156 = w1154 & w1155;
assign w1157 = w1152 & w1153;
assign w1158 = w1150 & w1151;
assign w1159 = w1157 & w1158;
assign w1160 = w1156 & w1159;
assign w1161 = pi357 & w456;
assign w1162 = pi340 & w446;
assign w1163 = pi379 & w459;
assign w1164 = pi274 & w478;
assign w1165 = pi319 & w454;
assign w1166 = pi368 & w464;
assign w1167 = pi405 & w542;
assign w1168 = pi364 & w476;
assign w1169 = pi287 & w461;
assign w1170 = pi270 & w452;
assign w1171 = pi341 & w450;
assign w1172 = ~w469 & ~w1161;
assign w1173 = ~w1162 & ~w1163;
assign w1174 = ~w1164 & ~w1165;
assign w1175 = ~w1166 & ~w1167;
assign w1176 = ~w1168 & ~w1169;
assign w1177 = ~w1170 & ~w1171;
assign w1178 = w1176 & w1177;
assign w1179 = w1174 & w1175;
assign w1180 = w1172 & w1173;
assign w1181 = w1179 & w1180;
assign w1182 = w1178 & w1181;
assign w1183 = ~w1160 & ~w1182;
assign w1184 = ~w468 & w8883;
assign w1185 = (~pi272 & w468) | (~pi272 & w8884) | (w468 & w8884);
assign w1186 = ~w1184 & ~w1185;
assign w1187 = w534 & w8885;
assign w1188 = pi584 & w472;
assign w1189 = pi511 & w470;
assign w1190 = pi636 & w474;
assign w1191 = pi663 & w442;
assign w1192 = w469 & ~w1188;
assign w1193 = ~w1189 & ~w1190;
assign w1194 = ~w1191 & w1193;
assign w1195 = w1192 & w1194;
assign w1196 = pi404 & w470;
assign w1197 = pi268 & w474;
assign w1198 = pi315 & w472;
assign w1199 = pi346 & w442;
assign w1200 = ~w469 & ~w1196;
assign w1201 = ~w1197 & ~w1198;
assign w1202 = ~w1199 & w1201;
assign w1203 = w1200 & w1202;
assign w1204 = ~w1195 & ~w1203;
assign w1205 = ~w108 & ~w1187;
assign w1206 = ~w1204 & w1205;
assign w1207 = ~w1183 & w1206;
assign w1208 = ~w1138 & ~w1207;
assign w1209 = ~w1207 & w8886;
assign w1210 = w109 & ~w924;
assign w1211 = w1119 & w1210;
assign w1212 = (~w1209 & w1119) | (~w1209 & w8887) | (w1119 & w8887);
assign w1213 = ~w1211 & w1212;
assign w1214 = ~w1027 & w1213;
assign w1215 = w1027 & ~w1213;
assign w1216 = ~w1214 & ~w1215;
assign w1217 = w1022 & ~w1216;
assign w1218 = ~w1022 & w1216;
assign w1219 = ~w1217 & ~w1218;
assign w1220 = ~w550 & ~w1208;
assign w1221 = w550 & w1208;
assign w1222 = ~w1220 & ~w1221;
assign w1223 = ~w108 & ~w708;
assign w1224 = ~w718 & w8888;
assign w1225 = ~w1223 & w1224;
assign w1226 = (w109 & w1097) | (w109 & w8889) | (w1097 & w8889);
assign w1227 = ~w1225 & ~w1226;
assign w1228 = w1222 & ~w1227;
assign w1229 = ~w1097 & w8890;
assign w1230 = ~w1225 & ~w1229;
assign w1231 = ~w1222 & ~w1230;
assign w1232 = ~w1228 & ~w1231;
assign w1233 = ~w831 & w1232;
assign w1234 = w831 & ~w1232;
assign w1235 = ~w1233 & ~w1234;
assign w1236 = ~w620 & w8891;
assign w1237 = ~w734 & ~w1236;
assign w1238 = w1222 & ~w1237;
assign w1239 = ~w709 & ~w1236;
assign w1240 = ~w1222 & ~w1239;
assign w1241 = ~w1238 & ~w1240;
assign w1242 = w1027 & ~w1241;
assign w1243 = ~w1027 & w1241;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = ~w1235 & w1244;
assign w1246 = w1235 & ~w1244;
assign w1247 = ~w1245 & ~w1246;
assign w1248 = w1219 & ~w1247;
assign w1249 = ~w1027 & ~w1232;
assign w1250 = w1027 & w1232;
assign w1251 = ~w1249 & ~w1250;
assign w1252 = ~w109 & ~w550;
assign w1253 = (w109 & w1207) | (w109 & w8892) | (w1207 & w8892);
assign w1254 = ~w1252 & ~w1253;
assign w1255 = w1119 & ~w1254;
assign w1256 = ~w1207 & w8893;
assign w1257 = ~w1252 & ~w1256;
assign w1258 = ~w1119 & ~w1257;
assign w1259 = ~w1255 & ~w1258;
assign w1260 = w1241 & ~w1259;
assign w1261 = ~w1241 & w1259;
assign w1262 = ~w1260 & ~w1261;
assign w1263 = ~w1019 & w1262;
assign w1264 = w1019 & ~w1262;
assign w1265 = ~w1263 & ~w1264;
assign w1266 = ~w1251 & ~w1265;
assign w1267 = w1248 & ~w1266;
assign w1268 = ~w1248 & w1266;
assign w1269 = ~w1267 & ~w1268;
assign w1270 = (~w109 & w1097) | (~w109 & w8894) | (w1097 & w8894);
assign w1271 = w109 & w1014;
assign w1272 = ~w1270 & ~w1271;
assign w1273 = (w1272 & ~w927) | (w1272 & w8895) | (~w927 & w8895);
assign w1274 = w927 & w8896;
assign w1275 = ~w1273 & ~w1274;
assign w1276 = ~w1019 & w1275;
assign w1277 = w1019 & ~w1275;
assign w1278 = ~w1276 & ~w1277;
assign w1279 = w1027 & ~w1259;
assign w1280 = ~w1027 & w1259;
assign w1281 = ~w1279 & ~w1280;
assign w1282 = ~w1235 & w1281;
assign w1283 = w1244 & ~w1262;
assign w1284 = ~w1282 & ~w1283;
assign w1285 = ~w1278 & ~w1284;
assign w1286 = w1235 & ~w1281;
assign w1287 = w1244 & w1281;
assign w1288 = w1278 & ~w1286;
assign w1289 = ~w1287 & w1288;
assign w1290 = ~w1285 & ~w1289;
assign w1291 = ~w1021 & w1027;
assign w1292 = ~w1020 & ~w1027;
assign w1293 = ~w1291 & ~w1292;
assign w1294 = w1290 & ~w1293;
assign w1295 = ~w1290 & w1293;
assign w1296 = ~w1294 & ~w1295;
assign w1297 = w1269 & w1296;
assign w1298 = ~w1269 & ~w1296;
assign w1299 = ~w1297 & ~w1298;
assign w1300 = w1278 & w1281;
assign w1301 = ~w1278 & ~w1281;
assign w1302 = ~w1300 & ~w1301;
assign w1303 = ~w1022 & w1302;
assign w1304 = w1235 & w1262;
assign w1305 = w1019 & ~w1244;
assign w1306 = w1304 & ~w1305;
assign w1307 = ~w1283 & ~w1305;
assign w1308 = ~w1304 & ~w1307;
assign w1309 = ~w1306 & ~w1308;
assign w1310 = w1303 & ~w1309;
assign w1311 = ~w1303 & w1309;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = w1022 & w1213;
assign w1314 = (~w1250 & w1022) | (~w1250 & w8897) | (w1022 & w8897);
assign w1315 = ~w1313 & w1314;
assign w1316 = ~w1249 & ~w1315;
assign w1317 = w1312 & w1316;
assign w1318 = ~w1312 & ~w1316;
assign w1319 = ~w1317 & ~w1318;
assign w1320 = ~w1235 & ~w1265;
assign w1321 = ~w1022 & w1244;
assign w1322 = ~w1265 & w8898;
assign w1323 = ~w1022 & ~w1247;
assign w1324 = ~w1320 & w1323;
assign w1325 = ~w1322 & ~w1324;
assign w1326 = w1219 & ~w1302;
assign w1327 = w1235 & w1259;
assign w1328 = ~w1235 & ~w1259;
assign w1329 = ~w1327 & ~w1328;
assign w1330 = w1241 & ~w1251;
assign w1331 = (~w1330 & w1329) | (~w1330 & w8899) | (w1329 & w8899);
assign w1332 = w1326 & ~w1331;
assign w1333 = ~w1326 & w1331;
assign w1334 = ~w1332 & ~w1333;
assign w1335 = ~w1325 & w1334;
assign w1336 = w1325 & ~w1334;
assign w1337 = ~w1335 & ~w1336;
assign w1338 = ~w1235 & ~w1262;
assign w1339 = ~w1304 & ~w1338;
assign w1340 = ~w1244 & w1339;
assign w1341 = ~w1022 & w1251;
assign w1342 = (~w1276 & ~w1262) | (~w1276 & w8900) | (~w1262 & w8900);
assign w1343 = w1341 & ~w1342;
assign w1344 = ~w1341 & w1342;
assign w1345 = ~w1343 & ~w1344;
assign w1346 = w1219 & w1235;
assign w1347 = w1345 & ~w1346;
assign w1348 = ~w1345 & w1346;
assign w1349 = ~w1347 & ~w1348;
assign w1350 = w1340 & w1349;
assign w1351 = ~w1340 & ~w1349;
assign w1352 = ~w1350 & ~w1351;
assign w1353 = w187 & ~w384;
assign w1354 = ~w187 & w384;
assign w1355 = ~w1353 & ~w1354;
assign w1356 = (~w303 & w384) | (~w303 & w8901) | (w384 & w8901);
assign w1357 = w1355 & w1356;
assign w1358 = ~w1355 & ~w1356;
assign w1359 = ~w1357 & ~w1358;
assign w1360 = (pi017 & w19) | (pi017 & w8902) | (w19 & w8902);
assign w1361 = ~w19 & w8903;
assign w1362 = ~w1360 & ~w1361;
assign w1363 = (pi056 & w19) | (pi056 & w8904) | (w19 & w8904);
assign w1364 = ~w19 & w8905;
assign w1365 = ~w1363 & ~w1364;
assign w1366 = (pi136 & w19) | (pi136 & w8906) | (w19 & w8906);
assign w1367 = ~w19 & w8907;
assign w1368 = ~w1366 & ~w1367;
assign w1369 = w1365 & ~w1368;
assign w1370 = ~w1365 & w1368;
assign w1371 = ~w1369 & ~w1370;
assign w1372 = w1362 & w1371;
assign w1373 = ~w1362 & ~w1371;
assign w1374 = ~w1372 & ~w1373;
assign w1375 = w1359 & ~w1374;
assign w1376 = ~w1359 & w1374;
assign w1377 = ~w1375 & ~w1376;
assign w1378 = (~pi009 & w19) | (~pi009 & w8908) | (w19 & w8908);
assign w1379 = ~w19 & w8909;
assign w1380 = w1 & ~w1378;
assign w1381 = ~w1379 & w1380;
assign w1382 = ~w1377 & w1381;
assign w1383 = ~w1359 & w8910;
assign w1384 = w1 & ~w1374;
assign w1385 = (pi009 & ~w0) | (pi009 & w8866) | (~w0 & w8866);
assign w1386 = (~w1385 & ~w1380) | (~w1385 & w8911) | (~w1380 & w8911);
assign w1387 = (w1386 & ~w1359) | (w1386 & w8912) | (~w1359 & w8912);
assign w1388 = ~w1383 & w1387;
assign w1389 = ~w1382 & ~w1388;
assign w1390 = ~w109 & ~w164;
assign w1391 = ~w1355 & w1390;
assign w1392 = ~w109 & w164;
assign w1393 = (~w171 & ~w1355) | (~w171 & w8913) | (~w1355 & w8913);
assign w1394 = ~w1391 & w1393;
assign w1395 = (pi188 & w19) | (pi188 & w8914) | (w19 & w8914);
assign w1396 = ~w19 & w8915;
assign w1397 = ~w1395 & ~w1396;
assign w1398 = (pi046 & w19) | (pi046 & w8916) | (w19 & w8916);
assign w1399 = ~w19 & w8917;
assign w1400 = ~w1398 & ~w1399;
assign w1401 = w1397 & ~w1400;
assign w1402 = ~w1397 & w1400;
assign w1403 = ~w1401 & ~w1402;
assign w1404 = ~w19 & w8918;
assign w1405 = (~pi042 & w19) | (~pi042 & w8919) | (w19 & w8919);
assign w1406 = ~w1404 & ~w1405;
assign w1407 = w1403 & ~w1406;
assign w1408 = ~w1403 & w1406;
assign w1409 = ~w1407 & ~w1408;
assign w1410 = w1 & w1409;
assign w1411 = ~w1394 & w1410;
assign w1412 = w1 & ~w1409;
assign w1413 = (w1412 & w1355) | (w1412 & w8920) | (w1355 & w8920);
assign w1414 = w1393 & w1413;
assign w1415 = w1 & w903;
assign w1416 = (~pi010 & ~w0) | (~pi010 & w8921) | (~w0 & w8921);
assign w1417 = (~w1416 & ~w903) | (~w1416 & w8922) | (~w903 & w8922);
assign w1418 = ~w1414 & w1417;
assign w1419 = ~w1411 & w1418;
assign w1420 = w903 & w1414;
assign w1421 = w1409 & w1415;
assign w1422 = ~w1394 & w1421;
assign w1423 = ~w1420 & ~w1422;
assign w1424 = ~w1419 & w1423;
assign w1425 = (~pi011 & ~w0) | (~pi011 & w8923) | (~w0 & w8923);
assign w1426 = ~w19 & w8924;
assign w1427 = (pi011 & w19) | (pi011 & w8925) | (w19 & w8925);
assign w1428 = w1 & ~w1426;
assign w1429 = (~w1425 & ~w1428) | (~w1425 & w8926) | (~w1428 & w8926);
assign w1430 = (pi176 & w19) | (pi176 & w8927) | (w19 & w8927);
assign w1431 = ~w19 & w8928;
assign w1432 = ~w1430 & ~w1431;
assign w1433 = (pi043 & w19) | (pi043 & w8929) | (w19 & w8929);
assign w1434 = ~w19 & w8930;
assign w1435 = ~w1433 & ~w1434;
assign w1436 = (pi047 & w19) | (pi047 & w8931) | (w19 & w8931);
assign w1437 = ~w19 & w8932;
assign w1438 = ~w1436 & ~w1437;
assign w1439 = w1435 & ~w1438;
assign w1440 = ~w1435 & w1438;
assign w1441 = ~w1439 & ~w1440;
assign w1442 = w1432 & w1441;
assign w1443 = ~w1432 & ~w1441;
assign w1444 = ~w1442 & ~w1443;
assign w1445 = w109 & ~w381;
assign w1446 = w233 & w347;
assign w1447 = ~w233 & ~w347;
assign w1448 = ~w1446 & ~w1447;
assign w1449 = (~w1445 & w1448) | (~w1445 & w8933) | (w1448 & w8933);
assign w1450 = w1444 & ~w1449;
assign w1451 = (w1448 & w8934) | (w1448 & w8935) | (w8934 & w8935);
assign w1452 = ~w1450 & ~w1451;
assign w1453 = (~w1429 & w1450) | (~w1429 & w8936) | (w1450 & w8936);
assign w1454 = (pi011 & ~w0) | (pi011 & w8815) | (~w0 & w8815);
assign w1455 = (~w1454 & ~w1428) | (~w1454 & w8937) | (~w1428 & w8937);
assign w1456 = w1452 & w1455;
assign w1457 = ~w1453 & ~w1456;
assign w1458 = w267 & w271;
assign w1459 = ~w267 & ~w271;
assign w1460 = ~w1458 & ~w1459;
assign w1461 = w535 & w8938;
assign w1462 = pi568 & w535;
assign w1463 = w535 & w8939;
assign w1464 = pi563 & ~pi565;
assign w1465 = ~pi566 & w444;
assign w1466 = pi566 & ~w444;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = ~w449 & ~w463;
assign w1469 = pi568 & ~w535;
assign w1470 = ~w536 & w1468;
assign w1471 = w1470 & w8940;
assign w1472 = w1464 & w1471;
assign w1473 = w305 & w8942;
assign w1474 = (w1471 & w8943) | (w1471 & w8944) | (w8943 & w8944);
assign w1475 = ~w1473 & w1474;
assign w1476 = ~w1461 & ~w1463;
assign w1477 = ~w1475 & w1476;
assign w1478 = w535 & w8945;
assign w1479 = w535 & w8946;
assign w1480 = ~w348 & w8948;
assign w1481 = (w1471 & w8949) | (w1471 & w8950) | (w8949 & w8950);
assign w1482 = ~w1480 & w1481;
assign w1483 = ~w1478 & ~w1479;
assign w1484 = ~w1482 & w1483;
assign w1485 = w535 & w8951;
assign w1486 = w535 & w8952;
assign w1487 = pi563 & pi565;
assign w1488 = w1470 & w8953;
assign w1489 = w1487 & w1488;
assign w1490 = w305 & w8955;
assign w1491 = (w1488 & w8956) | (w1488 & w8957) | (w8956 & w8957);
assign w1492 = ~w1490 & w1491;
assign w1493 = ~w1485 & ~w1486;
assign w1494 = ~w1492 & w1493;
assign w1495 = w535 & w8958;
assign w1496 = w535 & w8959;
assign w1497 = ~w348 & w8961;
assign w1498 = (w1488 & w8962) | (w1488 & w8963) | (w8962 & w8963);
assign w1499 = ~w1497 & w1498;
assign w1500 = ~w1495 & ~w1496;
assign w1501 = ~w1499 & w1500;
assign w1502 = w535 & w8964;
assign w1503 = w535 & w8965;
assign w1504 = w1471 & w1487;
assign w1505 = w305 & w8967;
assign w1506 = (w1471 & w8968) | (w1471 & w8969) | (w8968 & w8969);
assign w1507 = ~w1505 & w1506;
assign w1508 = ~w1502 & ~w1503;
assign w1509 = ~w1507 & w1508;
assign w1510 = w535 & w8970;
assign w1511 = w535 & w8971;
assign w1512 = ~w348 & w8973;
assign w1513 = (w1471 & w8974) | (w1471 & w8975) | (w8974 & w8975);
assign w1514 = ~w1512 & w1513;
assign w1515 = ~w1510 & ~w1511;
assign w1516 = ~w1514 & w1515;
assign w1517 = w535 & w8976;
assign w1518 = w535 & w8977;
assign w1519 = w1464 & w1488;
assign w1520 = w305 & w8979;
assign w1521 = (w1488 & w8980) | (w1488 & w8981) | (w8980 & w8981);
assign w1522 = ~w1520 & w1521;
assign w1523 = ~w1517 & ~w1518;
assign w1524 = ~w1522 & w1523;
assign w1525 = w535 & w8982;
assign w1526 = w535 & w8983;
assign w1527 = ~w348 & w8985;
assign w1528 = (w1488 & w8986) | (w1488 & w8987) | (w8986 & w8987);
assign w1529 = ~w1527 & w1528;
assign w1530 = ~w1525 & ~w1526;
assign w1531 = ~w1529 & w1530;
assign w1532 = w535 & w8988;
assign w1533 = ~pi038 & pi673;
assign w1534 = w535 & w8989;
assign w1535 = pi565 & ~w1465;
assign w1536 = ~pi563 & ~w535;
assign w1537 = ~w1535 & w1536;
assign w1538 = w1471 & w1537;
assign w1539 = (~pi026 & ~w1471) | (~pi026 & w8991) | (~w1471 & w8991);
assign w1540 = ~w348 & w8992;
assign w1541 = ~w535 & ~w1539;
assign w1542 = ~w1540 & w1541;
assign w1543 = (~w351 & w8993) | (~w351 & w8994) | (w8993 & w8994);
assign w1544 = ~w1542 & w1543;
assign w1545 = w535 & w8995;
assign w1546 = ~pi039 & pi673;
assign w1547 = w535 & w8996;
assign w1548 = w305 & w8998;
assign w1549 = (~w535 & w1538) | (~w535 & w8999) | (w1538 & w8999);
assign w1550 = ~w1548 & w1549;
assign w1551 = (w305 & w9000) | (w305 & w9001) | (w9000 & w9001);
assign w1552 = ~w1550 & w1551;
assign w1553 = w535 & w9002;
assign w1554 = ~pi031 & pi673;
assign w1555 = ~pi041 & ~pi673;
assign w1556 = ~w1554 & ~w1555;
assign w1557 = w1462 & w1556;
assign w1558 = ~pi566 & ~w441;
assign w1559 = ~w441 & w9003;
assign w1560 = ~w444 & w1559;
assign w1561 = w1537 & w1560;
assign w1562 = (~pi028 & ~w1537) | (~pi028 & w9004) | (~w1537 & w9004);
assign w1563 = ~w348 & w9005;
assign w1564 = ~w535 & ~w1562;
assign w1565 = ~w1563 & w1564;
assign w1566 = ~w1553 & ~w1557;
assign w1567 = ~w1565 & w1566;
assign w1568 = w535 & w9006;
assign w1569 = ~pi030 & pi673;
assign w1570 = ~pi040 & ~pi673;
assign w1571 = ~w1569 & ~w1570;
assign w1572 = w1462 & w1571;
assign w1573 = (~pi029 & ~w1537) | (~pi029 & w9007) | (~w1537 & w9007);
assign w1574 = ~w535 & ~w1573;
assign w1575 = (w1574 & ~w305) | (w1574 & w9009) | (~w305 & w9009);
assign w1576 = ~w1568 & ~w1572;
assign w1577 = ~w1575 & w1576;
assign w1578 = w535 & w9010;
assign w1579 = ~pi034 & pi673;
assign w1580 = ~pi029 & ~pi673;
assign w1581 = ~w1579 & ~w1580;
assign w1582 = w1462 & w1581;
assign w1583 = ~w1462 & ~w1535;
assign w1584 = ~pi563 & ~w1583;
assign w1585 = ~w444 & w9011;
assign w1586 = ~w1583 & w9012;
assign w1587 = (~pi030 & w1583) | (~pi030 & w9013) | (w1583 & w9013);
assign w1588 = ~w535 & ~w1587;
assign w1589 = (w1588 & ~w305) | (w1588 & w9015) | (~w305 & w9015);
assign w1590 = ~w1578 & ~w1582;
assign w1591 = ~w1589 & w1590;
assign w1592 = w535 & w9016;
assign w1593 = ~pi035 & pi673;
assign w1594 = ~pi028 & ~pi673;
assign w1595 = ~w1593 & ~w1594;
assign w1596 = w1462 & w1595;
assign w1597 = (~pi031 & w1583) | (~pi031 & w9017) | (w1583 & w9017);
assign w1598 = ~w348 & w9018;
assign w1599 = ~w535 & ~w1597;
assign w1600 = ~w1598 & w1599;
assign w1601 = ~w1592 & ~w1596;
assign w1602 = ~w1600 & w1601;
assign w1603 = w535 & w9019;
assign w1604 = w1471 & w1584;
assign w1605 = w305 & w9020;
assign w1606 = (~w535 & w1604) | (~w535 & w9021) | (w1604 & w9021);
assign w1607 = ~w1605 & w1606;
assign w1608 = ~pi039 & ~pi673;
assign w1609 = w535 & w9023;
assign w1610 = (w1609 & ~w305) | (w1609 & w9024) | (~w305 & w9024);
assign w1611 = ~w1603 & ~w1607;
assign w1612 = ~w1610 & w1611;
assign w1613 = w535 & w9025;
assign w1614 = ~w348 & w9026;
assign w1615 = (~w535 & w1604) | (~w535 & w9027) | (w1604 & w9027);
assign w1616 = ~pi038 & ~pi673;
assign w1617 = ~w348 & w9028;
assign w1618 = w535 & w9029;
assign w1619 = ~w1617 & w1618;
assign w1620 = (~w1613 & w1614) | (~w1613 & w9030) | (w1614 & w9030);
assign w1621 = ~w1619 & w1620;
assign w1622 = w535 & w9031;
assign w1623 = ~pi040 & pi673;
assign w1624 = ~pi030 & ~pi673;
assign w1625 = ~w1623 & ~w1624;
assign w1626 = w1462 & w1625;
assign w1627 = ~w1583 & w9032;
assign w1628 = w305 & w9033;
assign w1629 = (~w535 & w1627) | (~w535 & w9034) | (w1627 & w9034);
assign w1630 = ~w1628 & w1629;
assign w1631 = ~w1622 & ~w1626;
assign w1632 = ~w1630 & w1631;
assign w1633 = w535 & w9035;
assign w1634 = ~pi041 & pi673;
assign w1635 = ~pi031 & ~pi673;
assign w1636 = ~w1634 & ~w1635;
assign w1637 = w1462 & w1636;
assign w1638 = ~w348 & w9036;
assign w1639 = (~w535 & w1627) | (~w535 & w9037) | (w1627 & w9037);
assign w1640 = ~w1638 & w1639;
assign w1641 = ~w1633 & ~w1637;
assign w1642 = ~w1640 & w1641;
assign w1643 = pi032 & ~pi673;
assign w1644 = pi027 & pi673;
assign w1645 = ~w1643 & ~w1644;
assign w1646 = w1462 & ~w1645;
assign w1647 = (pi036 & ~w535) | (pi036 & w9038) | (~w535 & w9038);
assign w1648 = ~w1646 & ~w1647;
assign w1649 = pi033 & ~pi673;
assign w1650 = pi026 & pi673;
assign w1651 = ~w1649 & ~w1650;
assign w1652 = w1462 & ~w1651;
assign w1653 = (pi037 & ~w535) | (pi037 & w9039) | (~w535 & w9039);
assign w1654 = ~w1652 & ~w1653;
assign w1655 = w535 & w9040;
assign w1656 = ~pi033 & pi673;
assign w1657 = ~pi026 & ~pi673;
assign w1658 = ~w1656 & ~w1657;
assign w1659 = w1462 & w1658;
assign w1660 = w1488 & w1537;
assign w1661 = (~pi038 & ~w1488) | (~pi038 & w9041) | (~w1488 & w9041);
assign w1662 = ~w348 & w9042;
assign w1663 = ~w535 & ~w1661;
assign w1664 = ~w1662 & w1663;
assign w1665 = ~w1655 & ~w1659;
assign w1666 = ~w1664 & w1665;
assign w1667 = w535 & w9043;
assign w1668 = ~pi032 & pi673;
assign w1669 = ~pi027 & ~pi673;
assign w1670 = ~w1668 & ~w1669;
assign w1671 = w1462 & w1670;
assign w1672 = (~pi039 & ~w1488) | (~pi039 & w9044) | (~w1488 & w9044);
assign w1673 = ~w535 & ~w1672;
assign w1674 = (w1673 & ~w305) | (w1673 & w9046) | (~w305 & w9046);
assign w1675 = ~w1667 & ~w1671;
assign w1676 = ~w1674 & w1675;
assign w1677 = w535 & w9047;
assign w1678 = ~pi029 & pi673;
assign w1679 = ~pi034 & ~pi673;
assign w1680 = ~w1678 & ~w1679;
assign w1681 = w1462 & w1680;
assign w1682 = ~w441 & w1585;
assign w1683 = w1537 & w1682;
assign w1684 = (~pi040 & ~w1537) | (~pi040 & w9048) | (~w1537 & w9048);
assign w1685 = ~w535 & ~w1684;
assign w1686 = (w1685 & ~w305) | (w1685 & w9050) | (~w305 & w9050);
assign w1687 = ~w1677 & ~w1681;
assign w1688 = ~w1686 & w1687;
assign w1689 = w535 & w9051;
assign w1690 = ~pi028 & pi673;
assign w1691 = ~pi035 & ~pi673;
assign w1692 = ~w1690 & ~w1691;
assign w1693 = w1462 & w1692;
assign w1694 = (~pi041 & ~w1537) | (~pi041 & w9052) | (~w1537 & w9052);
assign w1695 = ~w348 & w9053;
assign w1696 = ~w535 & ~w1694;
assign w1697 = ~w1695 & w1696;
assign w1698 = ~w1689 & ~w1693;
assign w1699 = ~w1697 & w1698;
assign w1700 = ~w1394 & w1409;
assign w1701 = w1394 & ~w1409;
assign w1702 = ~w1700 & ~w1701;
assign w1703 = w213 & w216;
assign w1704 = ~w213 & ~w216;
assign w1705 = ~w1703 & ~w1704;
assign w1706 = w1 & ~w1394;
assign w1707 = (~pi046 & ~w0) | (~pi046 & w9054) | (~w0 & w9054);
assign w1708 = (~w1707 & ~w1403) | (~w1707 & w9055) | (~w1403 & w9055);
assign w1709 = ~w1706 & w1708;
assign w1710 = ~w1394 & w9056;
assign w1711 = ~w1709 & ~w1710;
assign w1712 = w1 & ~w1432;
assign w1713 = (w1448 & w9057) | (w1448 & w9058) | (w9057 & w9058);
assign w1714 = w1 & w1432;
assign w1715 = (~w1448 & w9059) | (~w1448 & w9060) | (w9059 & w9060);
assign w1716 = ~w1713 & ~w1715;
assign w1717 = ~w1438 & ~w1716;
assign w1718 = (pi047 & ~w0) | (pi047 & w9061) | (~w0 & w9061);
assign w1719 = (~w1718 & ~w1438) | (~w1718 & w9062) | (~w1438 & w9062);
assign w1720 = w1716 & ~w1719;
assign w1721 = ~w1717 & ~w1720;
assign w1722 = w285 & w314;
assign w1723 = ~w285 & ~w314;
assign w1724 = ~w1722 & ~w1723;
assign w1725 = w332 & w358;
assign w1726 = ~w332 & ~w358;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = w1464 & w1559;
assign w1729 = (w1728 & ~w305) | (w1728 & w9063) | (~w305 & w9063);
assign w1730 = (pi050 & ~w1559) | (pi050 & w9064) | (~w1559 & w9064);
assign w1731 = ~w1729 & ~w1730;
assign w1732 = (w1728 & w348) | (w1728 & w9065) | (w348 & w9065);
assign w1733 = (pi051 & ~w1559) | (pi051 & w9066) | (~w1559 & w9066);
assign w1734 = ~w1732 & ~w1733;
assign w1735 = w1585 & w9067;
assign w1736 = (w1735 & ~w305) | (w1735 & w9068) | (~w305 & w9068);
assign w1737 = pi052 & ~w1735;
assign w1738 = ~w1736 & ~w1737;
assign w1739 = w1585 & w9069;
assign w1740 = (w1739 & w348) | (w1739 & w9070) | (w348 & w9070);
assign w1741 = pi053 & ~w1739;
assign w1742 = ~w1740 & ~w1741;
assign w1743 = (w1735 & w348) | (w1735 & w9071) | (w348 & w9071);
assign w1744 = pi054 & ~w1735;
assign w1745 = ~w1743 & ~w1744;
assign w1746 = (w1739 & ~w305) | (w1739 & w9072) | (~w305 & w9072);
assign w1747 = pi055 & ~w1739;
assign w1748 = ~w1746 & ~w1747;
assign w1749 = w1359 & w1368;
assign w1750 = ~w1359 & ~w1368;
assign w1751 = ~w1749 & ~w1750;
assign w1752 = w1365 & ~w1751;
assign w1753 = ~w1365 & w1751;
assign w1754 = ~w1752 & ~w1753;
assign w1755 = w400 & w403;
assign w1756 = ~w400 & ~w403;
assign w1757 = ~w1755 & ~w1756;
assign w1758 = w535 & w9073;
assign w1759 = w535 & w9074;
assign w1760 = w1359 & w1472;
assign w1761 = (w1471 & w9076) | (w1471 & w9077) | (w9076 & w9077);
assign w1762 = ~w1760 & w1761;
assign w1763 = ~w1758 & ~w1759;
assign w1764 = ~w1762 & w1763;
assign w1765 = w535 & w9078;
assign w1766 = w535 & w9079;
assign w1767 = w1359 & w1504;
assign w1768 = (w1471 & w9081) | (w1471 & w9082) | (w9081 & w9082);
assign w1769 = ~w1767 & w1768;
assign w1770 = ~w1765 & ~w1766;
assign w1771 = ~w1769 & w1770;
assign w1772 = w535 & w9083;
assign w1773 = w535 & w9084;
assign w1774 = w1359 & w1519;
assign w1775 = (w1488 & w9086) | (w1488 & w9087) | (w9086 & w9087);
assign w1776 = ~w1774 & w1775;
assign w1777 = ~w1772 & ~w1773;
assign w1778 = ~w1776 & w1777;
assign w1779 = w535 & w9088;
assign w1780 = w535 & w9089;
assign w1781 = w1359 & w1489;
assign w1782 = (w1488 & w9091) | (w1488 & w9092) | (w9091 & w9092);
assign w1783 = ~w1781 & w1782;
assign w1784 = ~w1779 & ~w1780;
assign w1785 = ~w1783 & w1784;
assign w1786 = ~pi067 & pi673;
assign w1787 = ~pi092 & ~pi673;
assign w1788 = ~w1786 & ~w1787;
assign w1789 = w1462 & ~w1788;
assign w1790 = (pi062 & ~w535) | (pi062 & w9093) | (~w535 & w9093);
assign w1791 = ~w1789 & ~w1790;
assign w1792 = w535 & w9094;
assign w1793 = ~pi064 & pi673;
assign w1794 = ~pi066 & ~pi673;
assign w1795 = ~w1793 & ~w1794;
assign w1796 = w1462 & w1795;
assign w1797 = (~pi063 & ~w1537) | (~pi063 & w9095) | (~w1537 & w9095);
assign w1798 = ~w535 & ~w1797;
assign w1799 = (w1798 & ~w1359) | (w1798 & w9096) | (~w1359 & w9096);
assign w1800 = ~w1792 & ~w1796;
assign w1801 = ~w1799 & w1800;
assign w1802 = w535 & w9097;
assign w1803 = ~pi068 & pi673;
assign w1804 = ~pi063 & ~pi673;
assign w1805 = ~w1803 & ~w1804;
assign w1806 = w1462 & w1805;
assign w1807 = (~pi064 & w1583) | (~pi064 & w9098) | (w1583 & w9098);
assign w1808 = ~w535 & ~w1807;
assign w1809 = (w1808 & ~w1359) | (w1808 & w9099) | (~w1359 & w9099);
assign w1810 = ~w1802 & ~w1806;
assign w1811 = ~w1809 & w1810;
assign w1812 = w535 & w9100;
assign w1813 = ~pi092 & pi673;
assign w1814 = ~pi067 & ~pi673;
assign w1815 = ~w1813 & ~w1814;
assign w1816 = w1462 & w1815;
assign w1817 = (~pi065 & ~w1488) | (~pi065 & w9101) | (~w1488 & w9101);
assign w1818 = ~w535 & ~w1817;
assign w1819 = (w1818 & ~w1359) | (w1818 & w9102) | (~w1359 & w9102);
assign w1820 = ~w1812 & ~w1816;
assign w1821 = ~w1819 & w1820;
assign w1822 = w535 & w9103;
assign w1823 = ~pi068 & ~pi673;
assign w1824 = ~pi063 & pi673;
assign w1825 = ~w1823 & ~w1824;
assign w1826 = w1462 & w1825;
assign w1827 = (~pi066 & ~w1537) | (~pi066 & w9104) | (~w1537 & w9104);
assign w1828 = ~w535 & ~w1827;
assign w1829 = (w1828 & ~w1359) | (w1828 & w9105) | (~w1359 & w9105);
assign w1830 = ~w1822 & ~w1826;
assign w1831 = ~w1829 & w1830;
assign w1832 = (~pi067 & ~w1471) | (~pi067 & w9106) | (~w1471 & w9106);
assign w1833 = ~w535 & ~w1832;
assign w1834 = (w1833 & ~w1359) | (w1833 & w9107) | (~w1359 & w9107);
assign w1835 = pi067 & w536;
assign w1836 = ~pi065 & pi673;
assign w1837 = w535 & w9108;
assign w1838 = (w1837 & ~w1359) | (w1837 & w9109) | (~w1359 & w9109);
assign w1839 = ~w1834 & ~w1835;
assign w1840 = ~w1838 & w1839;
assign w1841 = w535 & w9110;
assign w1842 = ~pi066 & pi673;
assign w1843 = ~pi064 & ~pi673;
assign w1844 = ~w1842 & ~w1843;
assign w1845 = w1462 & w1844;
assign w1846 = w1359 & w1627;
assign w1847 = (~w535 & w1627) | (~w535 & w9111) | (w1627 & w9111);
assign w1848 = ~w1846 & w1847;
assign w1849 = ~w1841 & ~w1845;
assign w1850 = ~w1848 & w1849;
assign w1851 = w1487 & w1559;
assign w1852 = (w1851 & ~w305) | (w1851 & w9112) | (~w305 & w9112);
assign w1853 = (pi069 & ~w1559) | (pi069 & w9113) | (~w1559 & w9113);
assign w1854 = ~w1852 & ~w1853;
assign w1855 = (w1851 & w348) | (w1851 & w9114) | (w348 & w9114);
assign w1856 = (pi070 & ~w1559) | (pi070 & w9115) | (~w1559 & w9115);
assign w1857 = ~w1855 & ~w1856;
assign w1858 = (w427 & ~w305) | (w427 & w9116) | (~w305 & w9116);
assign w1859 = (~pi071 & ~w101) | (~pi071 & w9117) | (~w101 & w9117);
assign w1860 = ~w1858 & ~w1859;
assign w1861 = (w427 & w348) | (w427 & w9118) | (w348 & w9118);
assign w1862 = (~pi072 & ~w101) | (~pi072 & w9119) | (~w101 & w9119);
assign w1863 = ~w1861 & ~w1862;
assign w1864 = w535 & w9120;
assign w1865 = w535 & w9121;
assign w1866 = w207 & w1472;
assign w1867 = (w1471 & w9123) | (w1471 & w9124) | (w9123 & w9124);
assign w1868 = ~w1866 & w1867;
assign w1869 = ~w1864 & ~w1865;
assign w1870 = ~w1868 & w1869;
assign w1871 = w535 & w9125;
assign w1872 = w535 & w9126;
assign w1873 = w255 & w1472;
assign w1874 = (w1471 & w9128) | (w1471 & w9129) | (w9128 & w9129);
assign w1875 = ~w1873 & w1874;
assign w1876 = ~w1871 & ~w1872;
assign w1877 = ~w1875 & w1876;
assign w1878 = w535 & w9130;
assign w1879 = w535 & w9131;
assign w1880 = (~w384 & w396) | (~w384 & w9133) | (w396 & w9133);
assign w1881 = ~w396 & w9134;
assign w1882 = ~w1880 & ~w1881;
assign w1883 = w1472 & ~w1882;
assign w1884 = (w1471 & w9135) | (w1471 & w9136) | (w9135 & w9136);
assign w1885 = ~w1883 & w1884;
assign w1886 = ~w1878 & ~w1879;
assign w1887 = ~w1885 & w1886;
assign w1888 = w535 & w9137;
assign w1889 = w535 & w9138;
assign w1890 = w207 & w1489;
assign w1891 = (w1488 & w9140) | (w1488 & w9141) | (w9140 & w9141);
assign w1892 = ~w1890 & w1891;
assign w1893 = ~w1888 & ~w1889;
assign w1894 = ~w1892 & w1893;
assign w1895 = w535 & w9142;
assign w1896 = w535 & w9143;
assign w1897 = w255 & w1489;
assign w1898 = (w1488 & w9145) | (w1488 & w9146) | (w9145 & w9146);
assign w1899 = ~w1897 & w1898;
assign w1900 = ~w1895 & ~w1896;
assign w1901 = ~w1899 & w1900;
assign w1902 = w535 & w9147;
assign w1903 = w535 & w9148;
assign w1904 = w1489 & ~w1882;
assign w1905 = (w1488 & w9150) | (w1488 & w9151) | (w9150 & w9151);
assign w1906 = ~w1904 & w1905;
assign w1907 = ~w1902 & ~w1903;
assign w1908 = ~w1906 & w1907;
assign w1909 = w535 & w9152;
assign w1910 = w535 & w9153;
assign w1911 = w255 & w1504;
assign w1912 = (w1471 & w9155) | (w1471 & w9156) | (w9155 & w9156);
assign w1913 = ~w1911 & w1912;
assign w1914 = ~w1909 & ~w1910;
assign w1915 = ~w1913 & w1914;
assign w1916 = w535 & w9157;
assign w1917 = w535 & w9158;
assign w1918 = w207 & w1504;
assign w1919 = (w1471 & w9160) | (w1471 & w9161) | (w9160 & w9161);
assign w1920 = ~w1918 & w1919;
assign w1921 = ~w1916 & ~w1917;
assign w1922 = ~w1920 & w1921;
assign w1923 = w535 & w9162;
assign w1924 = w535 & w9163;
assign w1925 = w1504 & ~w1882;
assign w1926 = (w1471 & w9165) | (w1471 & w9166) | (w9165 & w9166);
assign w1927 = ~w1925 & w1926;
assign w1928 = ~w1923 & ~w1924;
assign w1929 = ~w1927 & w1928;
assign w1930 = w535 & w9167;
assign w1931 = w535 & w9168;
assign w1932 = w207 & w1519;
assign w1933 = (w1488 & w9170) | (w1488 & w9171) | (w9170 & w9171);
assign w1934 = ~w1932 & w1933;
assign w1935 = ~w1930 & ~w1931;
assign w1936 = ~w1934 & w1935;
assign w1937 = w535 & w9172;
assign w1938 = w535 & w9173;
assign w1939 = w255 & w1519;
assign w1940 = (w1488 & w9175) | (w1488 & w9176) | (w9175 & w9176);
assign w1941 = ~w1939 & w1940;
assign w1942 = ~w1937 & ~w1938;
assign w1943 = ~w1941 & w1942;
assign w1944 = w535 & w9177;
assign w1945 = w535 & w9178;
assign w1946 = w1519 & ~w1882;
assign w1947 = (w1488 & w9180) | (w1488 & w9181) | (w9180 & w9181);
assign w1948 = ~w1946 & w1947;
assign w1949 = ~w1944 & ~w1945;
assign w1950 = ~w1948 & w1949;
assign w1951 = (~pi085 & ~w1471) | (~pi085 & w9182) | (~w1471 & w9182);
assign w1952 = ~w535 & ~w1951;
assign w1953 = (w1952 & w1882) | (w1952 & w9183) | (w1882 & w9183);
assign w1954 = pi085 & w536;
assign w1955 = ~pi102 & pi673;
assign w1956 = w535 & w9184;
assign w1957 = (w1956 & w1882) | (w1956 & w9185) | (w1882 & w9185);
assign w1958 = ~w1953 & ~w1954;
assign w1959 = ~w1957 & w1958;
assign w1960 = w535 & w9186;
assign w1961 = ~pi090 & pi673;
assign w1962 = ~pi104 & ~pi673;
assign w1963 = ~w1961 & ~w1962;
assign w1964 = w1462 & w1963;
assign w1965 = (~pi086 & ~w1537) | (~pi086 & w9187) | (~w1537 & w9187);
assign w1966 = ~w535 & ~w1965;
assign w1967 = (w1966 & ~w207) | (w1966 & w9188) | (~w207 & w9188);
assign w1968 = ~w1960 & ~w1964;
assign w1969 = ~w1967 & w1968;
assign w1970 = w535 & w9189;
assign w1971 = ~pi089 & pi673;
assign w1972 = ~pi103 & ~pi673;
assign w1973 = ~w1971 & ~w1972;
assign w1974 = w1462 & w1973;
assign w1975 = (~pi087 & ~w1537) | (~pi087 & w9190) | (~w1537 & w9190);
assign w1976 = ~w535 & ~w1975;
assign w1977 = (w1976 & ~w255) | (w1976 & w9191) | (~w255 & w9191);
assign w1978 = ~w1970 & ~w1974;
assign w1979 = ~w1977 & w1978;
assign w1980 = w535 & w9192;
assign w1981 = ~pi091 & pi673;
assign w1982 = ~pi105 & ~pi673;
assign w1983 = ~w1981 & ~w1982;
assign w1984 = w1462 & w1983;
assign w1985 = (~pi088 & ~w1537) | (~pi088 & w9193) | (~w1537 & w9193);
assign w1986 = ~w535 & ~w1985;
assign w1987 = (w1986 & w1882) | (w1986 & w9194) | (w1882 & w9194);
assign w1988 = ~w1980 & ~w1984;
assign w1989 = ~w1987 & w1988;
assign w1990 = w535 & w9195;
assign w1991 = ~pi095 & pi673;
assign w1992 = ~pi087 & ~pi673;
assign w1993 = ~w1991 & ~w1992;
assign w1994 = w1462 & w1993;
assign w1995 = (~pi089 & w1583) | (~pi089 & w9196) | (w1583 & w9196);
assign w1996 = ~w535 & ~w1995;
assign w1997 = (w1996 & ~w255) | (w1996 & w9197) | (~w255 & w9197);
assign w1998 = ~w1990 & ~w1994;
assign w1999 = ~w1997 & w1998;
assign w2000 = w535 & w9198;
assign w2001 = ~pi094 & pi673;
assign w2002 = ~pi086 & ~pi673;
assign w2003 = ~w2001 & ~w2002;
assign w2004 = w1462 & w2003;
assign w2005 = (~pi090 & w1583) | (~pi090 & w9199) | (w1583 & w9199);
assign w2006 = ~w535 & ~w2005;
assign w2007 = (w2006 & ~w207) | (w2006 & w9200) | (~w207 & w9200);
assign w2008 = ~w2000 & ~w2004;
assign w2009 = ~w2007 & w2008;
assign w2010 = w535 & w9201;
assign w2011 = ~pi096 & pi673;
assign w2012 = ~pi088 & ~pi673;
assign w2013 = ~w2011 & ~w2012;
assign w2014 = w1462 & w2013;
assign w2015 = (~pi091 & w1583) | (~pi091 & w9202) | (w1583 & w9202);
assign w2016 = ~w535 & ~w2015;
assign w2017 = (w2016 & w1882) | (w2016 & w9203) | (w1882 & w9203);
assign w2018 = ~w2010 & ~w2014;
assign w2019 = ~w2017 & w2018;
assign w2020 = w535 & w9204;
assign w2021 = ~pi065 & ~pi673;
assign w2022 = w535 & w9205;
assign w2023 = w1359 & w1604;
assign w2024 = (~w535 & w1604) | (~w535 & w9207) | (w1604 & w9207);
assign w2025 = ~w2023 & w2024;
assign w2026 = (w1359 & w9208) | (w1359 & w9209) | (w9208 & w9209);
assign w2027 = ~w2025 & w2026;
assign w2028 = pi112 & pi673;
assign w2029 = pi097 & ~pi673;
assign w2030 = ~w2028 & ~w2029;
assign w2031 = w1462 & ~w2030;
assign w2032 = (pi093 & ~w535) | (pi093 & w9210) | (~w535 & w9210);
assign w2033 = ~w2031 & ~w2032;
assign w2034 = w535 & w9211;
assign w2035 = ~pi104 & pi673;
assign w2036 = ~pi090 & ~pi673;
assign w2037 = ~w2035 & ~w2036;
assign w2038 = w1462 & w2037;
assign w2039 = w207 & w1627;
assign w2040 = (~w535 & w1627) | (~w535 & w9212) | (w1627 & w9212);
assign w2041 = ~w2039 & w2040;
assign w2042 = ~w2034 & ~w2038;
assign w2043 = ~w2041 & w2042;
assign w2044 = w535 & w9213;
assign w2045 = ~pi103 & pi673;
assign w2046 = ~pi089 & ~pi673;
assign w2047 = ~w2045 & ~w2046;
assign w2048 = w1462 & w2047;
assign w2049 = w255 & w1627;
assign w2050 = (~w535 & w1627) | (~w535 & w9214) | (w1627 & w9214);
assign w2051 = ~w2049 & w2050;
assign w2052 = ~w2044 & ~w2048;
assign w2053 = ~w2051 & w2052;
assign w2054 = w535 & w9215;
assign w2055 = ~pi105 & pi673;
assign w2056 = ~pi091 & ~pi673;
assign w2057 = ~w2055 & ~w2056;
assign w2058 = w1462 & w2057;
assign w2059 = w1627 & ~w1882;
assign w2060 = (~w535 & w1627) | (~w535 & w9216) | (w1627 & w9216);
assign w2061 = ~w2059 & w2060;
assign w2062 = ~w2054 & ~w2058;
assign w2063 = ~w2061 & w2062;
assign w2064 = w535 & w9217;
assign w2065 = w255 & w1604;
assign w2066 = (~w535 & w1604) | (~w535 & w9218) | (w1604 & w9218);
assign w2067 = ~w2065 & w2066;
assign w2068 = ~pi098 & ~pi673;
assign w2069 = w535 & w9219;
assign w2070 = (w2069 & ~w255) | (w2069 & w9220) | (~w255 & w9220);
assign w2071 = ~w2064 & ~w2067;
assign w2072 = ~w2070 & w2071;
assign w2073 = w535 & w9221;
assign w2074 = ~pi097 & pi673;
assign w2075 = ~pi112 & ~pi673;
assign w2076 = ~w2074 & ~w2075;
assign w2077 = w1462 & w2076;
assign w2078 = (~pi098 & ~w1488) | (~pi098 & w9222) | (~w1488 & w9222);
assign w2079 = ~w535 & ~w2078;
assign w2080 = (w2079 & ~w255) | (w2079 & w9223) | (~w255 & w9223);
assign w2081 = ~w2073 & ~w2077;
assign w2082 = ~w2080 & w2081;
assign w2083 = w535 & w9224;
assign w2084 = ~pi118 & ~pi673;
assign w2085 = ~pi115 & pi673;
assign w2086 = ~w2084 & ~w2085;
assign w2087 = w1462 & w2086;
assign w2088 = (~pi099 & ~w1488) | (~pi099 & w9225) | (~w1488 & w9225);
assign w2089 = ~w535 & ~w2088;
assign w2090 = (w2089 & ~w207) | (w2089 & w9226) | (~w207 & w9226);
assign w2091 = ~w2083 & ~w2087;
assign w2092 = ~w2090 & w2091;
assign w2093 = pi115 & ~pi673;
assign w2094 = pi118 & pi673;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = w1462 & ~w2095;
assign w2097 = (pi100 & ~w535) | (pi100 & w9227) | (~w535 & w9227);
assign w2098 = ~w2096 & ~w2097;
assign w2099 = pi116 & ~pi673;
assign w2100 = pi085 & pi673;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = w1462 & ~w2101;
assign w2103 = (pi101 & ~w535) | (pi101 & w9228) | (~w535 & w9228);
assign w2104 = ~w2102 & ~w2103;
assign w2105 = w535 & w9229;
assign w2106 = ~pi116 & pi673;
assign w2107 = ~pi085 & ~pi673;
assign w2108 = ~w2106 & ~w2107;
assign w2109 = w1462 & w2108;
assign w2110 = (~pi102 & ~w1488) | (~pi102 & w9230) | (~w1488 & w9230);
assign w2111 = ~w535 & ~w2110;
assign w2112 = (w2111 & w1882) | (w2111 & w9231) | (w1882 & w9231);
assign w2113 = ~w2105 & ~w2109;
assign w2114 = ~w2112 & w2113;
assign w2115 = w535 & w9232;
assign w2116 = ~pi087 & pi673;
assign w2117 = ~pi095 & ~pi673;
assign w2118 = ~w2116 & ~w2117;
assign w2119 = w1462 & w2118;
assign w2120 = (~pi103 & ~w1537) | (~pi103 & w9233) | (~w1537 & w9233);
assign w2121 = ~w535 & ~w2120;
assign w2122 = (w2121 & ~w255) | (w2121 & w9234) | (~w255 & w9234);
assign w2123 = ~w2115 & ~w2119;
assign w2124 = ~w2122 & w2123;
assign w2125 = w535 & w9235;
assign w2126 = ~pi086 & pi673;
assign w2127 = ~pi094 & ~pi673;
assign w2128 = ~w2126 & ~w2127;
assign w2129 = w1462 & w2128;
assign w2130 = (~pi104 & ~w1537) | (~pi104 & w9236) | (~w1537 & w9236);
assign w2131 = ~w535 & ~w2130;
assign w2132 = (w2131 & ~w207) | (w2131 & w9237) | (~w207 & w9237);
assign w2133 = ~w2125 & ~w2129;
assign w2134 = ~w2132 & w2133;
assign w2135 = w535 & w9238;
assign w2136 = ~pi088 & pi673;
assign w2137 = ~pi096 & ~pi673;
assign w2138 = ~w2136 & ~w2137;
assign w2139 = w1462 & w2138;
assign w2140 = (~pi105 & ~w1537) | (~pi105 & w9239) | (~w1537 & w9239);
assign w2141 = ~w535 & ~w2140;
assign w2142 = (w2141 & w1882) | (w2141 & w9240) | (w1882 & w9240);
assign w2143 = ~w2135 & ~w2139;
assign w2144 = ~w2142 & w2143;
assign w2145 = ~w1359 & w1728;
assign w2146 = (pi106 & ~w1559) | (pi106 & w9241) | (~w1559 & w9241);
assign w2147 = ~w2145 & ~w2146;
assign w2148 = ~w1359 & w1735;
assign w2149 = pi107 & ~w1735;
assign w2150 = ~w2148 & ~w2149;
assign w2151 = ~w1359 & w1851;
assign w2152 = (pi108 & ~w1559) | (pi108 & w9242) | (~w1559 & w9242);
assign w2153 = ~w2151 & ~w2152;
assign w2154 = ~w1359 & w1739;
assign w2155 = pi109 & ~w1739;
assign w2156 = ~w2154 & ~w2155;
assign w2157 = ~w1219 & ~w1235;
assign w2158 = ~w1346 & ~w2157;
assign w2159 = (w102 & w348) | (w102 & w9243) | (w348 & w9243);
assign w2160 = (~pi111 & ~w99) | (~pi111 & w9244) | (~w99 & w9244);
assign w2161 = ~w2159 & ~w2160;
assign w2162 = w535 & w9245;
assign w2163 = (~pi112 & ~w1471) | (~pi112 & w9246) | (~w1471 & w9246);
assign w2164 = ~w535 & ~w2163;
assign w2165 = (w2164 & ~w255) | (w2164 & w9247) | (~w255 & w9247);
assign w2166 = ~pi098 & pi673;
assign w2167 = w535 & w9248;
assign w2168 = (w2167 & ~w255) | (w2167 & w9249) | (~w255 & w9249);
assign w2169 = ~w2162 & ~w2165;
assign w2170 = ~w2168 & w2169;
assign w2171 = (w424 & w348) | (w424 & w9250) | (w348 & w9250);
assign w2172 = ~pi113 & ~w424;
assign w2173 = ~w2171 & ~w2172;
assign w2174 = (w424 & ~w305) | (w424 & w9251) | (~w305 & w9251);
assign w2175 = (~pi114 & ~w101) | (~pi114 & w9252) | (~w101 & w9252);
assign w2176 = ~w2174 & ~w2175;
assign w2177 = w535 & w9253;
assign w2178 = w207 & w1604;
assign w2179 = (~w535 & w1604) | (~w535 & w9254) | (w1604 & w9254);
assign w2180 = ~w2178 & w2179;
assign w2181 = ~pi099 & ~pi673;
assign w2182 = w535 & w9255;
assign w2183 = (w2182 & ~w207) | (w2182 & w9256) | (~w207 & w9256);
assign w2184 = ~w2177 & ~w2180;
assign w2185 = ~w2183 & w2184;
assign w2186 = ~pi102 & ~pi673;
assign w2187 = w535 & w9257;
assign w2188 = pi116 & w536;
assign w2189 = w1604 & ~w1882;
assign w2190 = (~w535 & w1604) | (~w535 & w9259) | (w1604 & w9259);
assign w2191 = ~w2189 & w2190;
assign w2192 = (~w1882 & w9260) | (~w1882 & w9261) | (w9260 & w9261);
assign w2193 = ~w2191 & w2192;
assign w2194 = (w102 & ~w305) | (w102 & w9262) | (~w305 & w9262);
assign w2195 = ~pi117 & ~w102;
assign w2196 = ~w2194 & ~w2195;
assign w2197 = w535 & w9263;
assign w2198 = (~pi118 & ~w1471) | (~pi118 & w9264) | (~w1471 & w9264);
assign w2199 = ~w535 & ~w2198;
assign w2200 = (w2199 & ~w207) | (w2199 & w9265) | (~w207 & w9265);
assign w2201 = ~pi099 & pi673;
assign w2202 = w535 & w9266;
assign w2203 = (w2202 & ~w207) | (w2202 & w9267) | (~w207 & w9267);
assign w2204 = ~w2197 & ~w2200;
assign w2205 = ~w2203 & w2204;
assign w2206 = ~w207 & w1728;
assign w2207 = (pi119 & ~w1559) | (pi119 & w9268) | (~w1559 & w9268);
assign w2208 = ~w2206 & ~w2207;
assign w2209 = (pi120 & ~w1559) | (pi120 & w9269) | (~w1559 & w9269);
assign w2210 = ~w255 & w1728;
assign w2211 = ~w2209 & ~w2210;
assign w2212 = w1728 & w1882;
assign w2213 = (pi121 & ~w1559) | (pi121 & w9270) | (~w1559 & w9270);
assign w2214 = ~w2212 & ~w2213;
assign w2215 = ~w207 & w1735;
assign w2216 = pi122 & ~w1735;
assign w2217 = ~w2215 & ~w2216;
assign w2218 = pi123 & ~w1735;
assign w2219 = ~w255 & w1735;
assign w2220 = ~w2218 & ~w2219;
assign w2221 = w1735 & w1882;
assign w2222 = pi124 & ~w1735;
assign w2223 = ~w2221 & ~w2222;
assign w2224 = ~w207 & w1851;
assign w2225 = (pi125 & ~w1559) | (pi125 & w9271) | (~w1559 & w9271);
assign w2226 = ~w2224 & ~w2225;
assign w2227 = (pi126 & ~w1559) | (pi126 & w9272) | (~w1559 & w9272);
assign w2228 = ~w255 & w1851;
assign w2229 = ~w2227 & ~w2228;
assign w2230 = w1851 & w1882;
assign w2231 = (pi127 & ~w1559) | (pi127 & w9273) | (~w1559 & w9273);
assign w2232 = ~w2230 & ~w2231;
assign w2233 = w1739 & w1882;
assign w2234 = pi128 & ~w1739;
assign w2235 = ~w2233 & ~w2234;
assign w2236 = ~w207 & w1739;
assign w2237 = pi129 & ~w1739;
assign w2238 = ~w2236 & ~w2237;
assign w2239 = pi130 & ~w1739;
assign w2240 = ~w255 & w1739;
assign w2241 = ~w2239 & ~w2240;
assign w2242 = w427 & w1359;
assign w2243 = (pi131 & ~w101) | (pi131 & w9274) | (~w101 & w9274);
assign w2244 = ~w2242 & ~w2243;
assign w2245 = w1 & ~w213;
assign w2246 = (pi133 & ~w0) | (pi133 & w9275) | (~w0 & w9275);
assign w2247 = ~w2245 & ~w2246;
assign w2248 = w1 & ~w261;
assign w2249 = (pi134 & ~w0) | (pi134 & w9276) | (~w0 & w9276);
assign w2250 = ~w2248 & ~w2249;
assign w2251 = w255 & w427;
assign w2252 = (pi135 & ~w101) | (pi135 & w9277) | (~w101 & w9277);
assign w2253 = ~w2251 & ~w2252;
assign w2254 = w1 & ~w1751;
assign w2255 = (~pi136 & ~w0) | (~pi136 & w9278) | (~w0 & w9278);
assign w2256 = ~w2254 & ~w2255;
assign w2257 = w427 & ~w1882;
assign w2258 = (pi137 & ~w101) | (pi137 & w9279) | (~w101 & w9279);
assign w2259 = ~w2257 & ~w2258;
assign w2260 = w207 & w427;
assign w2261 = (pi138 & ~w101) | (pi138 & w9280) | (~w101 & w9280);
assign w2262 = ~w2260 & ~w2261;
assign w2263 = ~w1394 & w1472;
assign w2264 = (w1471 & w9282) | (w1471 & w9283) | (w9282 & w9283);
assign w2265 = ~w2263 & w2264;
assign w2266 = w535 & w9284;
assign w2267 = w535 & w9285;
assign w2268 = ~w2266 & ~w2267;
assign w2269 = ~w2265 & w2268;
assign w2270 = ~w1394 & w1489;
assign w2271 = (w1488 & w9287) | (w1488 & w9288) | (w9287 & w9288);
assign w2272 = ~w2270 & w2271;
assign w2273 = w535 & w9289;
assign w2274 = w535 & w9290;
assign w2275 = ~w2273 & ~w2274;
assign w2276 = ~w2272 & w2275;
assign w2277 = ~w1394 & w1519;
assign w2278 = (w1488 & w9292) | (w1488 & w9293) | (w9292 & w9293);
assign w2279 = ~w2277 & w2278;
assign w2280 = w535 & w9294;
assign w2281 = w535 & w9295;
assign w2282 = ~w2280 & ~w2281;
assign w2283 = ~w2279 & w2282;
assign w2284 = ~w1394 & w1504;
assign w2285 = (w1471 & w9297) | (w1471 & w9298) | (w9297 & w9298);
assign w2286 = ~w2284 & w2285;
assign w2287 = w535 & w9299;
assign w2288 = w535 & w9300;
assign w2289 = ~w2287 & ~w2288;
assign w2290 = ~w2286 & w2289;
assign w2291 = (~pi143 & ~w1537) | (~pi143 & w9301) | (~w1537 & w9301);
assign w2292 = ~w535 & ~w2291;
assign w2293 = (w2292 & w1394) | (w2292 & w9302) | (w1394 & w9302);
assign w2294 = pi143 & w536;
assign w2295 = ~pi147 & pi673;
assign w2296 = ~pi151 & ~pi673;
assign w2297 = ~w2295 & ~w2296;
assign w2298 = w1462 & w2297;
assign w2299 = ~w2294 & ~w2298;
assign w2300 = ~w2293 & w2299;
assign w2301 = w102 & w1359;
assign w2302 = (pi144 & ~w99) | (pi144 & w9303) | (~w99 & w9303);
assign w2303 = ~w2301 & ~w2302;
assign w2304 = w207 & w424;
assign w2305 = (pi145 & ~w101) | (pi145 & w9304) | (~w101 & w9304);
assign w2306 = ~w2304 & ~w2305;
assign w2307 = w255 & w424;
assign w2308 = (pi146 & ~w101) | (pi146 & w9305) | (~w101 & w9305);
assign w2309 = ~w2307 & ~w2308;
assign w2310 = (~pi147 & w1583) | (~pi147 & w9306) | (w1583 & w9306);
assign w2311 = ~w535 & ~w2310;
assign w2312 = (w2311 & w1394) | (w2311 & w9307) | (w1394 & w9307);
assign w2313 = pi147 & w536;
assign w2314 = ~pi149 & pi673;
assign w2315 = ~pi143 & ~pi673;
assign w2316 = ~w2314 & ~w2315;
assign w2317 = w1462 & w2316;
assign w2318 = ~w2313 & ~w2317;
assign w2319 = ~w2312 & w2318;
assign w2320 = pi158 & ~pi673;
assign w2321 = pi152 & pi673;
assign w2322 = ~w2320 & ~w2321;
assign w2323 = w1462 & ~w2322;
assign w2324 = (pi148 & ~w535) | (pi148 & w9308) | (~w535 & w9308);
assign w2325 = ~w2323 & ~w2324;
assign w2326 = ~w1394 & w1627;
assign w2327 = (~w535 & w1627) | (~w535 & w9309) | (w1627 & w9309);
assign w2328 = ~w2326 & w2327;
assign w2329 = w535 & w9310;
assign w2330 = ~pi151 & pi673;
assign w2331 = ~pi147 & ~pi673;
assign w2332 = ~w2330 & ~w2331;
assign w2333 = w1462 & w2332;
assign w2334 = ~w2329 & ~w2333;
assign w2335 = ~w2328 & w2334;
assign w2336 = (~pi150 & ~w1488) | (~pi150 & w9311) | (~w1488 & w9311);
assign w2337 = ~w535 & ~w2336;
assign w2338 = (w2337 & w1394) | (w2337 & w9312) | (w1394 & w9312);
assign w2339 = pi150 & w536;
assign w2340 = ~pi152 & ~pi673;
assign w2341 = ~pi158 & pi673;
assign w2342 = ~w2340 & ~w2341;
assign w2343 = w1462 & w2342;
assign w2344 = ~w2339 & ~w2343;
assign w2345 = ~w2338 & w2344;
assign w2346 = (~pi151 & ~w1537) | (~pi151 & w9313) | (~w1537 & w9313);
assign w2347 = ~w535 & ~w2346;
assign w2348 = (w2347 & w1394) | (w2347 & w9314) | (w1394 & w9314);
assign w2349 = pi151 & w536;
assign w2350 = ~pi143 & pi673;
assign w2351 = ~pi149 & ~pi673;
assign w2352 = ~w2350 & ~w2351;
assign w2353 = w1462 & w2352;
assign w2354 = ~w2349 & ~w2353;
assign w2355 = ~w2348 & w2354;
assign w2356 = (~pi152 & ~w1471) | (~pi152 & w9315) | (~w1471 & w9315);
assign w2357 = ~w535 & ~w2356;
assign w2358 = (w2357 & w1394) | (w2357 & w9316) | (w1394 & w9316);
assign w2359 = pi152 & w536;
assign w2360 = ~pi150 & pi673;
assign w2361 = ~w164 & w1355;
assign w2362 = (~pi673 & w1355) | (~pi673 & w9317) | (w1355 & w9317);
assign w2363 = ~w2361 & w2362;
assign w2364 = w535 & w9318;
assign w2365 = (~w2359 & w2363) | (~w2359 & w9319) | (w2363 & w9319);
assign w2366 = ~w2358 & w2365;
assign w2367 = w424 & w1359;
assign w2368 = (pi153 & ~w101) | (pi153 & w9320) | (~w101 & w9320);
assign w2369 = ~w2367 & ~w2368;
assign w2370 = w102 & w255;
assign w2371 = (pi154 & ~w99) | (pi154 & w9321) | (~w99 & w9321);
assign w2372 = ~w2370 & ~w2371;
assign w2373 = w1 & w400;
assign w2374 = (pi155 & ~w0) | (pi155 & w9322) | (~w0 & w9322);
assign w2375 = ~w2373 & ~w2374;
assign w2376 = w102 & w207;
assign w2377 = (pi156 & ~w99) | (pi156 & w9323) | (~w99 & w9323);
assign w2378 = ~w2376 & ~w2377;
assign w2379 = w102 & ~w1882;
assign w2380 = (pi157 & ~w99) | (pi157 & w9324) | (~w99 & w9324);
assign w2381 = ~w2379 & ~w2380;
assign w2382 = w535 & w9325;
assign w2383 = ~w1604 & ~w2382;
assign w2384 = w1394 & ~w2383;
assign w2385 = (pi158 & ~w535) | (pi158 & w9326) | (~w535 & w9326);
assign w2386 = pi150 & ~pi673;
assign w2387 = w535 & w9327;
assign w2388 = (~w2387 & w1604) | (~w2387 & w9328) | (w1604 & w9328);
assign w2389 = ~w2384 & w2388;
assign w2390 = w424 & ~w1882;
assign w2391 = (pi159 & ~w101) | (pi159 & w9329) | (~w101 & w9329);
assign w2392 = ~w2390 & ~w2391;
assign w2393 = ~w1394 & w1728;
assign w2394 = (~pi160 & ~w1559) | (~pi160 & w9330) | (~w1559 & w9330);
assign w2395 = ~w2393 & ~w2394;
assign w2396 = ~w1394 & w1735;
assign w2397 = ~pi161 & ~w1735;
assign w2398 = ~w2396 & ~w2397;
assign w2399 = ~w1394 & w1851;
assign w2400 = (~pi162 & ~w1559) | (~pi162 & w9331) | (~w1559 & w9331);
assign w2401 = ~w2399 & ~w2400;
assign w2402 = ~w1394 & w1739;
assign w2403 = ~pi163 & ~w1739;
assign w2404 = ~w2402 & ~w2403;
assign w2405 = w1251 & w1339;
assign w2406 = ~w1251 & ~w1339;
assign w2407 = ~w2405 & ~w2406;
assign w2408 = w535 & w9332;
assign w2409 = w535 & w9333;
assign w2410 = (w1448 & w9335) | (w1448 & w9336) | (w9335 & w9336);
assign w2411 = (w1471 & w9337) | (w1471 & w9338) | (w9337 & w9338);
assign w2412 = ~w2410 & w2411;
assign w2413 = ~w2408 & ~w2409;
assign w2414 = ~w2412 & w2413;
assign w2415 = w535 & w9339;
assign w2416 = w535 & w9340;
assign w2417 = (w1448 & w9342) | (w1448 & w9343) | (w9342 & w9343);
assign w2418 = (w1471 & w9344) | (w1471 & w9345) | (w9344 & w9345);
assign w2419 = ~w2417 & w2418;
assign w2420 = ~w2415 & ~w2416;
assign w2421 = ~w2419 & w2420;
assign w2422 = w535 & w9346;
assign w2423 = w535 & w9347;
assign w2424 = (w1448 & w9349) | (w1448 & w9350) | (w9349 & w9350);
assign w2425 = (w1488 & w9351) | (w1488 & w9352) | (w9351 & w9352);
assign w2426 = ~w2424 & w2425;
assign w2427 = ~w2422 & ~w2423;
assign w2428 = ~w2426 & w2427;
assign w2429 = w535 & w9353;
assign w2430 = w535 & w9354;
assign w2431 = (w1448 & w9356) | (w1448 & w9357) | (w9356 & w9357);
assign w2432 = (w1488 & w9358) | (w1488 & w9359) | (w9358 & w9359);
assign w2433 = ~w2431 & w2432;
assign w2434 = ~w2429 & ~w2430;
assign w2435 = ~w2433 & w2434;
assign w2436 = w535 & w9360;
assign w2437 = ~pi180 & pi673;
assign w2438 = ~pi181 & ~pi673;
assign w2439 = ~w2437 & ~w2438;
assign w2440 = w1462 & w2439;
assign w2441 = (~pi172 & w1583) | (~pi172 & w9361) | (w1583 & w9361);
assign w2442 = ~w535 & ~w2441;
assign w2443 = (~w1448 & w9364) | (~w1448 & w9365) | (w9364 & w9365);
assign w2444 = ~w2436 & ~w2440;
assign w2445 = ~w2443 & w2444;
assign w2446 = ~pi175 & pi673;
assign w2447 = ~pi182 & ~pi673;
assign w2448 = ~w2446 & ~w2447;
assign w2449 = w1462 & ~w2448;
assign w2450 = (pi173 & ~w535) | (pi173 & w9366) | (~w535 & w9366);
assign w2451 = ~w2449 & ~w2450;
assign w2452 = w535 & w9367;
assign w2453 = ~pi175 & ~pi673;
assign w2454 = ~pi182 & pi673;
assign w2455 = ~w2453 & ~w2454;
assign w2456 = w1462 & w2455;
assign w2457 = (~pi174 & ~w1488) | (~pi174 & w9368) | (~w1488 & w9368);
assign w2458 = ~w535 & ~w2457;
assign w2459 = (~w1448 & w9371) | (~w1448 & w9372) | (w9371 & w9372);
assign w2460 = ~w2452 & ~w2456;
assign w2461 = ~w2459 & w2460;
assign w2462 = w535 & w9373;
assign w2463 = ~pi174 & pi673;
assign w2464 = w535 & w9374;
assign w2465 = (w1448 & w9376) | (w1448 & w9377) | (w9376 & w9377);
assign w2466 = (~w535 & w1538) | (~w535 & w9378) | (w1538 & w9378);
assign w2467 = ~w2465 & w2466;
assign w2468 = (w1448 & w9379) | (w1448 & w9380) | (w9379 & w9380);
assign w2469 = ~w2467 & w2468;
assign w2470 = (pi176 & ~w0) | (pi176 & w9381) | (~w0 & w9381);
assign w2471 = w1716 & ~w2470;
assign w2472 = w427 & ~w1394;
assign w2473 = (pi177 & ~w101) | (pi177 & w9382) | (~w101 & w9382);
assign w2474 = ~w2472 & ~w2473;
assign w2475 = w535 & w9383;
assign w2476 = ~pi181 & pi673;
assign w2477 = ~pi180 & ~pi673;
assign w2478 = ~w2476 & ~w2477;
assign w2479 = w1462 & w2478;
assign w2480 = (~pi179 & ~w1537) | (~pi179 & w9384) | (~w1537 & w9384);
assign w2481 = ~w535 & ~w2480;
assign w2482 = (~w1448 & w9387) | (~w1448 & w9388) | (w9387 & w9388);
assign w2483 = ~w2475 & ~w2479;
assign w2484 = ~w2482 & w2483;
assign w2485 = w535 & w9389;
assign w2486 = ~pi179 & pi673;
assign w2487 = ~pi172 & ~pi673;
assign w2488 = ~w2486 & ~w2487;
assign w2489 = w1462 & w2488;
assign w2490 = (w1448 & w9390) | (w1448 & w9391) | (w9390 & w9391);
assign w2491 = (~w535 & w1627) | (~w535 & w9392) | (w1627 & w9392);
assign w2492 = ~w2490 & w2491;
assign w2493 = ~w2485 & ~w2489;
assign w2494 = ~w2492 & w2493;
assign w2495 = w535 & w9393;
assign w2496 = ~pi172 & pi673;
assign w2497 = ~pi179 & ~pi673;
assign w2498 = ~w2496 & ~w2497;
assign w2499 = w1462 & w2498;
assign w2500 = (~pi181 & ~w1537) | (~pi181 & w9394) | (~w1537 & w9394);
assign w2501 = ~w535 & ~w2500;
assign w2502 = (~w1448 & w9397) | (~w1448 & w9398) | (w9397 & w9398);
assign w2503 = ~w2495 & ~w2499;
assign w2504 = ~w2502 & w2503;
assign w2505 = w535 & w9399;
assign w2506 = ~pi174 & ~pi673;
assign w2507 = w535 & w9402;
assign w2508 = (~w1448 & w9403) | (~w1448 & w9404) | (w9403 & w9404);
assign w2509 = (w1448 & w9405) | (w1448 & w9406) | (w9405 & w9406);
assign w2510 = (~w535 & w1604) | (~w535 & w9407) | (w1604 & w9407);
assign w2511 = ~w2509 & w2510;
assign w2512 = ~w2505 & ~w2508;
assign w2513 = ~w2511 & w2512;
assign w2514 = (~w1448 & w9408) | (~w1448 & w9409) | (w9408 & w9409);
assign w2515 = (~pi183 & ~w1559) | (~pi183 & w9410) | (~w1559 & w9410);
assign w2516 = ~w2514 & ~w2515;
assign w2517 = (~w1448 & w9411) | (~w1448 & w9412) | (w9411 & w9412);
assign w2518 = ~pi184 & ~w1739;
assign w2519 = ~w2517 & ~w2518;
assign w2520 = (~w1448 & w9413) | (~w1448 & w9414) | (w9413 & w9414);
assign w2521 = ~pi185 & ~w1735;
assign w2522 = ~w2520 & ~w2521;
assign w2523 = w102 & ~w1394;
assign w2524 = (pi186 & ~w99) | (pi186 & w9415) | (~w99 & w9415);
assign w2525 = ~w2523 & ~w2524;
assign w2526 = (~w1448 & w9416) | (~w1448 & w9417) | (w9416 & w9417);
assign w2527 = (~pi187 & ~w1559) | (~pi187 & w9418) | (~w1559 & w9418);
assign w2528 = ~w2526 & ~w2527;
assign w2529 = ~w1394 & w9419;
assign w2530 = w1 & w1397;
assign w2531 = (pi188 & ~w0) | (pi188 & w9420) | (~w0 & w9420);
assign w2532 = (~w2531 & ~w1394) | (~w2531 & w9421) | (~w1394 & w9421);
assign w2533 = ~w2529 & w2532;
assign w2534 = w424 & ~w1394;
assign w2535 = (pi189 & ~w101) | (pi189 & w9422) | (~w101 & w9422);
assign w2536 = ~w2534 & ~w2535;
assign w2537 = (~w1448 & w9423) | (~w1448 & w9424) | (w9423 & w9424);
assign w2538 = (~pi191 & ~w101) | (~pi191 & w9425) | (~w101 & w9425);
assign w2539 = ~w2537 & ~w2538;
assign w2540 = w1022 & ~w1244;
assign w2541 = ~w1321 & ~w2540;
assign w2542 = (~w1448 & w9426) | (~w1448 & w9427) | (w9426 & w9427);
assign w2543 = (~pi193 & ~w99) | (~pi193 & w9428) | (~w99 & w9428);
assign w2544 = ~w2542 & ~w2543;
assign w2545 = (~w1448 & w9429) | (~w1448 & w9430) | (w9429 & w9430);
assign w2546 = (~pi194 & ~w101) | (~pi194 & w9431) | (~w101 & w9431);
assign w2547 = ~w2545 & ~w2546;
assign w2548 = (pi196 & ~w0) | (pi196 & w9432) | (~w0 & w9432);
assign w2549 = pi551 & w418;
assign w2550 = pi390 & pi665;
assign w2551 = pi550 & w2550;
assign w2552 = w2550 & w9433;
assign w2553 = pi665 & w18;
assign w2554 = (~w18 & w9435) | (~w18 & w9436) | (w9435 & w9436);
assign w2555 = ~pi551 & w2552;
assign w2556 = ~w18 & w2555;
assign w2557 = ~w2554 & ~w2556;
assign w2558 = ~pi559 & ~w2557;
assign w2559 = ~w2549 & ~w2558;
assign w2560 = pi552 & w418;
assign w2561 = (~pi552 & ~w2550) | (~pi552 & w9437) | (~w2550 & w9437);
assign w2562 = ~pi559 & ~w2561;
assign w2563 = (~w18 & w9438) | (~w18 & w9439) | (w9438 & w9439);
assign w2564 = ~w2560 & ~w2563;
assign w2565 = w2559 & ~w2564;
assign w2566 = ~w2559 & w2564;
assign w2567 = ~w2565 & ~w2566;
assign w2568 = pi559 & w22;
assign w2569 = ~w18 & w9440;
assign w2570 = pi390 & ~w2569;
assign w2571 = (~pi390 & w18) | (~pi390 & w9441) | (w18 & w9441);
assign w2572 = (~pi559 & w2571) | (~pi559 & w9442) | (w2571 & w9442);
assign w2573 = ~w418 & ~w2572;
assign w2574 = ~w2570 & ~w2573;
assign w2575 = pi550 & w418;
assign w2576 = ~pi550 & ~w2550;
assign w2577 = (~pi559 & ~w18) | (~pi559 & w9443) | (~w18 & w9443);
assign w2578 = ~w2551 & ~w2576;
assign w2579 = (~w18 & w9444) | (~w18 & w9445) | (w9444 & w9445);
assign w2580 = ~w2575 & ~w2579;
assign w2581 = ~w2574 & w2580;
assign w2582 = w2574 & ~w2580;
assign w2583 = w2574 & w9446;
assign w2584 = ~w2581 & ~w2583;
assign w2585 = ~w2567 & ~w2584;
assign w2586 = ~w19 & w9447;
assign w2587 = (~pi288 & w19) | (~pi288 & w9448) | (w19 & w9448);
assign w2588 = ~w2586 & ~w2587;
assign w2589 = pi154 & ~w2588;
assign w2590 = ~pi154 & w2588;
assign w2591 = ~w2589 & ~w2590;
assign w2592 = w2585 & w2591;
assign w2593 = ~w2585 & ~w2591;
assign w2594 = ~w2592 & ~w2593;
assign w2595 = (pi228 & w19) | (pi228 & w9449) | (w19 & w9449);
assign w2596 = ~w19 & w9450;
assign w2597 = ~w2595 & ~w2596;
assign w2598 = w2594 & w2597;
assign w2599 = ~w2594 & ~w2597;
assign w2600 = ~w2598 & ~w2599;
assign w2601 = (pi204 & w19) | (pi204 & w9451) | (w19 & w9451);
assign w2602 = ~w19 & w9452;
assign w2603 = ~w2601 & ~w2602;
assign w2604 = w2600 & ~w2603;
assign w2605 = ~w2600 & w2603;
assign w2606 = ~w2604 & ~w2605;
assign w2607 = w623 & w2606;
assign w2608 = (w1 & w2606) | (w1 & w9453) | (w2606 & w9453);
assign w2609 = ~w2607 & w2608;
assign w2610 = ~w2548 & ~w2609;
assign w2611 = (pi238 & w19) | (pi238 & w9454) | (w19 & w9454);
assign w2612 = ~w19 & w9455;
assign w2613 = ~w2611 & ~w2612;
assign w2614 = w2574 & w2580;
assign w2615 = w2565 & w2614;
assign w2616 = w2566 & w2581;
assign w2617 = ~w2615 & ~w2616;
assign w2618 = pi156 & ~w2617;
assign w2619 = ~pi156 & w2617;
assign w2620 = ~w2618 & ~w2619;
assign w2621 = ~w19 & w9456;
assign w2622 = (~pi333 & w19) | (~pi333 & w9457) | (w19 & w9457);
assign w2623 = ~w2621 & ~w2622;
assign w2624 = w2620 & ~w2623;
assign w2625 = ~w2620 & w2623;
assign w2626 = ~w2624 & ~w2625;
assign w2627 = w2613 & w2626;
assign w2628 = ~w2613 & ~w2626;
assign w2629 = ~w2627 & ~w2628;
assign w2630 = (pi215 & w19) | (pi215 & w9458) | (w19 & w9458);
assign w2631 = ~w19 & w9459;
assign w2632 = ~w2630 & ~w2631;
assign w2633 = w2629 & w2632;
assign w2634 = ~w2629 & ~w2632;
assign w2635 = ~w2633 & ~w2634;
assign w2636 = w1123 & ~w2635;
assign w2637 = ~w1123 & w2635;
assign w2638 = ~w2636 & ~w2637;
assign w2639 = w1 & ~w2638;
assign w2640 = (pi197 & ~w0) | (pi197 & w9460) | (~w0 & w9460);
assign w2641 = ~w2639 & ~w2640;
assign w2642 = (~pi198 & ~w0) | (~pi198 & w9461) | (~w0 & w9461);
assign w2643 = ~w2567 & w2582;
assign w2644 = (pi332 & w19) | (pi332 & w9462) | (w19 & w9462);
assign w2645 = ~w19 & w9463;
assign w2646 = ~w2644 & ~w2645;
assign w2647 = pi117 & ~w2646;
assign w2648 = ~pi117 & w2646;
assign w2649 = ~w2647 & ~w2648;
assign w2650 = ~w2567 & w9464;
assign w2651 = (~w2649 & w2567) | (~w2649 & w9465) | (w2567 & w9465);
assign w2652 = ~w2650 & ~w2651;
assign w2653 = (pi239 & w19) | (pi239 & w9466) | (w19 & w9466);
assign w2654 = ~w19 & w9467;
assign w2655 = ~w2653 & ~w2654;
assign w2656 = w2652 & ~w2655;
assign w2657 = ~w2652 & w2655;
assign w2658 = ~w2656 & ~w2657;
assign w2659 = (pi214 & w19) | (pi214 & w9468) | (w19 & w9468);
assign w2660 = ~w19 & w9469;
assign w2661 = ~w2659 & ~w2660;
assign w2662 = w2658 & w2661;
assign w2663 = ~w2658 & ~w2661;
assign w2664 = ~w2662 & ~w2663;
assign w2665 = w931 & w2664;
assign w2666 = (w1 & w2664) | (w1 & w9470) | (w2664 & w9470);
assign w2667 = ~w2665 & w2666;
assign w2668 = ~w2642 & ~w2667;
assign w2669 = (pi199 & ~w0) | (pi199 & w9471) | (~w0 & w9471);
assign w2670 = w2559 & ~w2580;
assign w2671 = ~w2574 & w2670;
assign w2672 = w2670 & w9472;
assign w2673 = pi111 & ~w2672;
assign w2674 = ~pi111 & w2672;
assign w2675 = ~w2673 & ~w2674;
assign w2676 = ~w19 & w9473;
assign w2677 = (~pi394 & w19) | (~pi394 & w9474) | (w19 & w9474);
assign w2678 = ~w2676 & ~w2677;
assign w2679 = w2675 & ~w2678;
assign w2680 = ~w2675 & w2678;
assign w2681 = ~w2679 & ~w2680;
assign w2682 = ~w19 & w9475;
assign w2683 = (~pi249 & w19) | (~pi249 & w9476) | (w19 & w9476);
assign w2684 = ~w2682 & ~w2683;
assign w2685 = w2681 & ~w2684;
assign w2686 = ~w2681 & w2684;
assign w2687 = ~w2685 & ~w2686;
assign w2688 = (pi226 & w19) | (pi226 & w9477) | (w19 & w9477);
assign w2689 = ~w19 & w9478;
assign w2690 = ~w2688 & ~w2689;
assign w2691 = ~w2687 & w2690;
assign w2692 = w2687 & ~w2690;
assign w2693 = ~w2691 & ~w2692;
assign w2694 = w1 & ~w2693;
assign w2695 = w1 & ~w422;
assign w2696 = (w2695 & w2693) | (w2695 & w9480) | (w2693 & w9480);
assign w2697 = (~w2669 & w2693) | (~w2669 & w9481) | (w2693 & w9481);
assign w2698 = ~w2696 & w2697;
assign w2699 = (pi200 & ~w0) | (pi200 & w9482) | (~w0 & w9482);
assign w2700 = ~w2574 & w9483;
assign w2701 = pi144 & ~w2700;
assign w2702 = ~pi144 & w2700;
assign w2703 = ~w2701 & ~w2702;
assign w2704 = ~w19 & w9484;
assign w2705 = (~pi387 & w19) | (~pi387 & w9485) | (w19 & w9485);
assign w2706 = ~w2704 & ~w2705;
assign w2707 = w2703 & ~w2706;
assign w2708 = ~w2703 & w2706;
assign w2709 = ~w2707 & ~w2708;
assign w2710 = ~w19 & w9486;
assign w2711 = (~pi248 & w19) | (~pi248 & w9487) | (w19 & w9487);
assign w2712 = ~w2710 & ~w2711;
assign w2713 = w2709 & ~w2712;
assign w2714 = ~w2709 & w2712;
assign w2715 = ~w2713 & ~w2714;
assign w2716 = (pi227 & w19) | (pi227 & w9488) | (w19 & w9488);
assign w2717 = ~w19 & w9489;
assign w2718 = ~w2716 & ~w2717;
assign w2719 = w2715 & ~w2718;
assign w2720 = ~w2715 & w2718;
assign w2721 = ~w2719 & ~w2720;
assign w2722 = w1100 & w2721;
assign w2723 = (w1 & w2721) | (w1 & w9490) | (w2721 & w9490);
assign w2724 = ~w2722 & w2723;
assign w2725 = ~w2699 & ~w2724;
assign w2726 = (pi201 & ~w0) | (pi201 & w9491) | (~w0 & w9491);
assign w2727 = w2566 & w2614;
assign w2728 = pi157 & ~w2727;
assign w2729 = ~pi157 & w2727;
assign w2730 = ~w2728 & ~w2729;
assign w2731 = ~w19 & w9492;
assign w2732 = (~pi389 & w19) | (~pi389 & w9493) | (w19 & w9493);
assign w2733 = ~w2731 & ~w2732;
assign w2734 = w2730 & ~w2733;
assign w2735 = ~w2730 & w2733;
assign w2736 = ~w2734 & ~w2735;
assign w2737 = ~w19 & w9494;
assign w2738 = (~pi250 & w19) | (~pi250 & w9495) | (w19 & w9495);
assign w2739 = ~w2737 & ~w2738;
assign w2740 = w2736 & ~w2739;
assign w2741 = ~w2736 & w2739;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = (pi225 & w19) | (pi225 & w9496) | (w19 & w9496);
assign w2744 = ~w19 & w9497;
assign w2745 = ~w2743 & ~w2744;
assign w2746 = ~w2742 & w2745;
assign w2747 = w2742 & ~w2745;
assign w2748 = ~w2746 & ~w2747;
assign w2749 = w1 & ~w2748;
assign w2750 = w1 & ~w811;
assign w2751 = (w2750 & w2748) | (w2750 & w9499) | (w2748 & w9499);
assign w2752 = (~w2726 & w2748) | (~w2726 & w9500) | (w2748 & w9500);
assign w2753 = ~w2751 & w2752;
assign w2754 = (~pi202 & ~w0) | (~pi202 & w9501) | (~w0 & w9501);
assign w2755 = (pi251 & w19) | (pi251 & w9502) | (w19 & w9502);
assign w2756 = ~w19 & w9503;
assign w2757 = ~w2755 & ~w2756;
assign w2758 = (pi193 & w2616) | (pi193 & w9504) | (w2616 & w9504);
assign w2759 = ~w2616 & w9505;
assign w2760 = ~w2758 & ~w2759;
assign w2761 = ~w19 & w9506;
assign w2762 = (~pi388 & w19) | (~pi388 & w9507) | (w19 & w9507);
assign w2763 = ~w2761 & ~w2762;
assign w2764 = w2760 & ~w2763;
assign w2765 = ~w2760 & w2763;
assign w2766 = ~w2764 & ~w2765;
assign w2767 = w2757 & w2766;
assign w2768 = ~w2757 & ~w2766;
assign w2769 = ~w2767 & ~w2768;
assign w2770 = (pi223 & w19) | (pi223 & w9508) | (w19 & w9508);
assign w2771 = ~w19 & w9509;
assign w2772 = ~w2770 & ~w2771;
assign w2773 = w2769 & w2772;
assign w2774 = ~w2769 & ~w2772;
assign w2775 = ~w2773 & ~w2774;
assign w2776 = w1 & w2775;
assign w2777 = w1 & ~w717;
assign w2778 = (~w2754 & w717) | (~w2754 & w9510) | (w717 & w9510);
assign w2779 = (w2778 & ~w2775) | (w2778 & w9511) | (~w2775 & w9511);
assign w2780 = w2775 & w2777;
assign w2781 = ~w2779 & ~w2780;
assign w2782 = (~pi203 & ~w0) | (~pi203 & w9512) | (~w0 & w9512);
assign w2783 = (w2564 & w2643) | (w2564 & w9513) | (w2643 & w9513);
assign w2784 = ~pi924 & w27;
assign w2785 = (~pi396 & w19) | (~pi396 & w9514) | (w19 & w9514);
assign w2786 = (pi186 & w2784) | (pi186 & w9515) | (w2784 & w9515);
assign w2787 = ~w2784 & w9516;
assign w2788 = ~w2786 & ~w2787;
assign w2789 = w2783 & w2788;
assign w2790 = ~w2783 & ~w2788;
assign w2791 = ~w2789 & ~w2790;
assign w2792 = (pi247 & w19) | (pi247 & w9517) | (w19 & w9517);
assign w2793 = ~w19 & w9518;
assign w2794 = ~w2792 & ~w2793;
assign w2795 = w2791 & w2794;
assign w2796 = ~w2791 & ~w2794;
assign w2797 = ~w2795 & ~w2796;
assign w2798 = (pi224 & w19) | (pi224 & w9519) | (w19 & w9519);
assign w2799 = ~w19 & w9520;
assign w2800 = ~w2798 & ~w2799;
assign w2801 = ~w2797 & ~w2800;
assign w2802 = w2797 & w2800;
assign w2803 = ~w2801 & ~w2802;
assign w2804 = w1 & ~w2803;
assign w2805 = (~w2782 & w911) | (~w2782 & w9521) | (w911 & w9521);
assign w2806 = ~w2804 & w2805;
assign w2807 = ~w2803 & w9522;
assign w2808 = ~w2806 & ~w2807;
assign w2809 = w1 & w2606;
assign w2810 = (pi204 & ~w0) | (pi204 & w9523) | (~w0 & w9523);
assign w2811 = ~w2809 & ~w2810;
assign w2812 = (~pi205 & ~w0) | (~pi205 & w9524) | (~w0 & w9524);
assign w2813 = ~w19 & w9525;
assign w2814 = (~pi414 & w19) | (~pi414 & w9526) | (w19 & w9526);
assign w2815 = ~w2813 & ~w2814;
assign w2816 = pi189 & ~w2815;
assign w2817 = ~pi189 & w2815;
assign w2818 = ~w2816 & ~w2817;
assign w2819 = ~w19 & w9527;
assign w2820 = (~pi292 & w19) | (~pi292 & w9528) | (w19 & w9528);
assign w2821 = ~w2819 & ~w2820;
assign w2822 = w2818 & ~w2821;
assign w2823 = ~w2818 & w2821;
assign w2824 = ~w2822 & ~w2823;
assign w2825 = (pi231 & w19) | (pi231 & w9529) | (w19 & w9529);
assign w2826 = ~w19 & w9530;
assign w2827 = ~w2825 & ~w2826;
assign w2828 = w2824 & ~w2827;
assign w2829 = ~w2824 & w2827;
assign w2830 = ~w2828 & ~w2829;
assign w2831 = (pi205 & w19) | (pi205 & w9531) | (w19 & w9531);
assign w2832 = ~w19 & w9532;
assign w2833 = ~w2831 & ~w2832;
assign w2834 = w2830 & w2833;
assign w2835 = (w1 & w2830) | (w1 & w9533) | (w2830 & w9533);
assign w2836 = ~w2834 & w2835;
assign w2837 = ~w2812 & ~w2836;
assign w2838 = (~pi206 & ~w0) | (~pi206 & w9534) | (~w0 & w9534);
assign w2839 = ~w19 & w9535;
assign w2840 = (~pi437 & w19) | (~pi437 & w9536) | (w19 & w9536);
assign w2841 = ~w2839 & ~w2840;
assign w2842 = pi145 & ~w2841;
assign w2843 = ~pi145 & w2841;
assign w2844 = ~w2842 & ~w2843;
assign w2845 = ~w19 & w9537;
assign w2846 = (~pi291 & w19) | (~pi291 & w9538) | (w19 & w9538);
assign w2847 = ~w2845 & ~w2846;
assign w2848 = w2844 & ~w2847;
assign w2849 = ~w2844 & w2847;
assign w2850 = ~w2848 & ~w2849;
assign w2851 = (pi232 & w19) | (pi232 & w9539) | (w19 & w9539);
assign w2852 = ~w19 & w9540;
assign w2853 = ~w2851 & ~w2852;
assign w2854 = w2850 & ~w2853;
assign w2855 = ~w2850 & w2853;
assign w2856 = ~w2854 & ~w2855;
assign w2857 = (pi206 & w19) | (pi206 & w9541) | (w19 & w9541);
assign w2858 = ~w19 & w9542;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = w2856 & w2859;
assign w2861 = (w1 & w2856) | (w1 & w9543) | (w2856 & w9543);
assign w2862 = ~w2860 & w2861;
assign w2863 = ~w2838 & ~w2862;
assign w2864 = (~pi207 & ~w0) | (~pi207 & w9544) | (~w0 & w9544);
assign w2865 = ~w19 & w9545;
assign w2866 = (~pi415 & w19) | (~pi415 & w9546) | (w19 & w9546);
assign w2867 = ~w2865 & ~w2866;
assign w2868 = pi146 & ~w2867;
assign w2869 = ~pi146 & w2867;
assign w2870 = ~w2868 & ~w2869;
assign w2871 = ~pi870 & w27;
assign w2872 = ~pi293 & ~w27;
assign w2873 = ~w2871 & ~w2872;
assign w2874 = w2870 & ~w2873;
assign w2875 = ~w2870 & w2873;
assign w2876 = ~w2874 & ~w2875;
assign w2877 = pi233 & ~w27;
assign w2878 = ~pi838 & w27;
assign w2879 = ~w2877 & ~w2878;
assign w2880 = w2876 & ~w2879;
assign w2881 = ~w2876 & w2879;
assign w2882 = ~w2880 & ~w2881;
assign w2883 = pi207 & ~w27;
assign w2884 = pi806 & w27;
assign w2885 = ~w2883 & ~w2884;
assign w2886 = ~w2882 & ~w2885;
assign w2887 = w2882 & w2885;
assign w2888 = w1 & ~w2886;
assign w2889 = ~w2887 & w2888;
assign w2890 = ~w2864 & ~w2889;
assign w2891 = pi208 & ~w1;
assign w2892 = ~pi903 & w27;
assign w2893 = ~pi416 & ~w27;
assign w2894 = ~w2892 & ~w2893;
assign w2895 = pi114 & ~w2894;
assign w2896 = ~pi114 & w2894;
assign w2897 = ~w2895 & ~w2896;
assign w2898 = ~pi871 & w27;
assign w2899 = ~pi252 & ~w27;
assign w2900 = ~w2898 & ~w2899;
assign w2901 = w2897 & ~w2900;
assign w2902 = ~w2897 & w2900;
assign w2903 = ~w2901 & ~w2902;
assign w2904 = pi237 & ~w27;
assign w2905 = ~pi839 & w27;
assign w2906 = ~w2904 & ~w2905;
assign w2907 = w2903 & ~w2906;
assign w2908 = ~w2903 & w2906;
assign w2909 = ~w2907 & ~w2908;
assign w2910 = w1 & ~w2909;
assign w2911 = pi208 & ~w27;
assign w2912 = pi807 & w27;
assign w2913 = ~w2911 & ~w2912;
assign w2914 = w2910 & ~w2913;
assign w2915 = w1 & w2913;
assign w2916 = w2909 & w2915;
assign w2917 = ~w2891 & ~w2916;
assign w2918 = ~w2914 & w2917;
assign w2919 = pi209 & ~w1;
assign w2920 = ~pi904 & w27;
assign w2921 = ~pi417 & ~w27;
assign w2922 = ~w2920 & ~w2921;
assign w2923 = pi113 & ~w2922;
assign w2924 = ~pi113 & w2922;
assign w2925 = ~w2923 & ~w2924;
assign w2926 = ~pi872 & w27;
assign w2927 = ~pi294 & ~w27;
assign w2928 = ~w2926 & ~w2927;
assign w2929 = w2925 & ~w2928;
assign w2930 = ~w2925 & w2928;
assign w2931 = ~w2929 & ~w2930;
assign w2932 = pi234 & ~w27;
assign w2933 = ~pi840 & w27;
assign w2934 = ~w2932 & ~w2933;
assign w2935 = w2931 & ~w2934;
assign w2936 = ~w2931 & w2934;
assign w2937 = ~w2935 & ~w2936;
assign w2938 = pi209 & ~w27;
assign w2939 = pi808 & w27;
assign w2940 = ~w2938 & ~w2939;
assign w2941 = w2937 & ~w2940;
assign w2942 = ~w2937 & w2940;
assign w2943 = w1 & ~w2941;
assign w2944 = ~w2942 & w2943;
assign w2945 = ~w2919 & ~w2944;
assign w2946 = ~pi210 & ~w1;
assign w2947 = ~pi898 & w27;
assign w2948 = ~pi413 & ~w27;
assign w2949 = ~w2947 & ~w2948;
assign w2950 = pi153 & ~w2949;
assign w2951 = ~pi153 & w2949;
assign w2952 = ~w2950 & ~w2951;
assign w2953 = ~pi866 & w27;
assign w2954 = ~pi289 & ~w27;
assign w2955 = ~w2953 & ~w2954;
assign w2956 = w2952 & ~w2955;
assign w2957 = ~w2952 & w2955;
assign w2958 = ~w2956 & ~w2957;
assign w2959 = pi229 & ~w27;
assign w2960 = ~pi834 & w27;
assign w2961 = ~w2959 & ~w2960;
assign w2962 = w2958 & ~w2961;
assign w2963 = ~w2958 & w2961;
assign w2964 = ~w2962 & ~w2963;
assign w2965 = pi210 & ~w27;
assign w2966 = pi802 & w27;
assign w2967 = ~w2965 & ~w2966;
assign w2968 = ~w2964 & ~w2967;
assign w2969 = w2964 & w2967;
assign w2970 = w1 & ~w2968;
assign w2971 = ~w2969 & w2970;
assign w2972 = ~w2946 & ~w2971;
assign w2973 = ~pi211 & ~w1;
assign w2974 = ~pi899 & w27;
assign w2975 = ~pi409 & ~w27;
assign w2976 = ~w2974 & ~w2975;
assign w2977 = pi194 & ~w2976;
assign w2978 = ~pi194 & w2976;
assign w2979 = ~w2977 & ~w2978;
assign w2980 = ~pi867 & w27;
assign w2981 = ~pi290 & ~w27;
assign w2982 = ~w2980 & ~w2981;
assign w2983 = w2979 & ~w2982;
assign w2984 = ~w2979 & w2982;
assign w2985 = ~w2983 & ~w2984;
assign w2986 = pi230 & ~w27;
assign w2987 = ~pi835 & w27;
assign w2988 = ~w2986 & ~w2987;
assign w2989 = w2985 & ~w2988;
assign w2990 = ~w2985 & w2988;
assign w2991 = ~w2989 & ~w2990;
assign w2992 = pi211 & ~w27;
assign w2993 = pi803 & w27;
assign w2994 = ~w2992 & ~w2993;
assign w2995 = ~w2991 & ~w2994;
assign w2996 = w2991 & w2994;
assign w2997 = w1 & ~w2995;
assign w2998 = ~w2996 & w2997;
assign w2999 = ~w2973 & ~w2998;
assign w3000 = ~pi212 & ~w1;
assign w3001 = ~pi921 & w27;
assign w3002 = ~pi419 & ~w27;
assign w3003 = ~w3001 & ~w3002;
assign w3004 = pi137 & ~w3003;
assign w3005 = ~pi137 & w3003;
assign w3006 = ~w3004 & ~w3005;
assign w3007 = ~pi889 & w27;
assign w3008 = ~pi296 & ~w27;
assign w3009 = ~w3007 & ~w3008;
assign w3010 = w3006 & ~w3009;
assign w3011 = ~w3006 & w3009;
assign w3012 = ~w3010 & ~w3011;
assign w3013 = pi236 & ~w27;
assign w3014 = ~pi857 & w27;
assign w3015 = ~w3013 & ~w3014;
assign w3016 = w3012 & ~w3015;
assign w3017 = ~w3012 & w3015;
assign w3018 = ~w3016 & ~w3017;
assign w3019 = pi212 & ~w27;
assign w3020 = pi825 & w27;
assign w3021 = ~w3019 & ~w3020;
assign w3022 = ~w3018 & ~w3021;
assign w3023 = w3018 & w3021;
assign w3024 = w1 & ~w3022;
assign w3025 = ~w3023 & w3024;
assign w3026 = ~w3000 & ~w3025;
assign w3027 = pi213 & ~w1;
assign w3028 = ~pi905 & w27;
assign w3029 = ~pi418 & ~w27;
assign w3030 = ~w3028 & ~w3029;
assign w3031 = pi159 & ~w3030;
assign w3032 = ~pi159 & w3030;
assign w3033 = ~w3031 & ~w3032;
assign w3034 = ~pi873 & w27;
assign w3035 = ~pi295 & ~w27;
assign w3036 = ~w3034 & ~w3035;
assign w3037 = w3033 & ~w3036;
assign w3038 = ~w3033 & w3036;
assign w3039 = ~w3037 & ~w3038;
assign w3040 = pi235 & ~w27;
assign w3041 = ~pi841 & w27;
assign w3042 = ~w3040 & ~w3041;
assign w3043 = w3039 & ~w3042;
assign w3044 = ~w3039 & w3042;
assign w3045 = ~w3043 & ~w3044;
assign w3046 = pi213 & ~w27;
assign w3047 = pi809 & w27;
assign w3048 = ~w3046 & ~w3047;
assign w3049 = w3045 & ~w3048;
assign w3050 = ~w3045 & w3048;
assign w3051 = w1 & ~w3049;
assign w3052 = ~w3050 & w3051;
assign w3053 = ~w3027 & ~w3052;
assign w3054 = pi214 & ~w1;
assign w3055 = w1 & ~w2664;
assign w3056 = ~w3054 & ~w3055;
assign w3057 = w1 & w2635;
assign w3058 = pi215 & ~w1;
assign w3059 = ~w3057 & ~w3058;
assign w3060 = ~pi216 & ~w1;
assign w3061 = ~pi915 & w27;
assign w3062 = ~pi421 & ~w27;
assign w3063 = ~w3061 & ~w3062;
assign w3064 = pi191 & ~w3063;
assign w3065 = ~pi191 & w3063;
assign w3066 = ~w3064 & ~w3065;
assign w3067 = ~pi883 & w27;
assign w3068 = ~pi298 & ~w27;
assign w3069 = ~w3067 & ~w3068;
assign w3070 = w3066 & ~w3069;
assign w3071 = ~w3066 & w3069;
assign w3072 = ~w3070 & ~w3071;
assign w3073 = pi240 & ~w27;
assign w3074 = ~pi851 & w27;
assign w3075 = ~w3073 & ~w3074;
assign w3076 = w3072 & ~w3075;
assign w3077 = ~w3072 & w3075;
assign w3078 = ~w3076 & ~w3077;
assign w3079 = pi216 & ~w27;
assign w3080 = pi819 & w27;
assign w3081 = ~w3079 & ~w3080;
assign w3082 = ~w3078 & ~w3081;
assign w3083 = w3078 & w3081;
assign w3084 = w1 & ~w3082;
assign w3085 = ~w3083 & w3084;
assign w3086 = ~w3060 & ~w3085;
assign w3087 = ~pi217 & ~w1;
assign w3088 = ~pi914 & w27;
assign w3089 = ~pi430 & ~w27;
assign w3090 = ~w3088 & ~w3089;
assign w3091 = pi131 & ~w3090;
assign w3092 = ~pi131 & w3090;
assign w3093 = ~w3091 & ~w3092;
assign w3094 = ~pi882 & w27;
assign w3095 = ~pi334 & ~w27;
assign w3096 = ~w3094 & ~w3095;
assign w3097 = w3093 & ~w3096;
assign w3098 = ~w3093 & w3096;
assign w3099 = ~w3097 & ~w3098;
assign w3100 = pi245 & ~w27;
assign w3101 = ~pi850 & w27;
assign w3102 = ~w3100 & ~w3101;
assign w3103 = w3099 & ~w3102;
assign w3104 = ~w3099 & w3102;
assign w3105 = ~w3103 & ~w3104;
assign w3106 = pi217 & ~w27;
assign w3107 = pi818 & w27;
assign w3108 = ~w3106 & ~w3107;
assign w3109 = ~w3105 & ~w3108;
assign w3110 = w3105 & w3108;
assign w3111 = w1 & ~w3109;
assign w3112 = ~w3110 & w3111;
assign w3113 = ~w3087 & ~w3112;
assign w3114 = ~pi218 & ~w1;
assign w3115 = ~pi917 & w27;
assign w3116 = ~pi431 & ~w27;
assign w3117 = ~w3115 & ~w3116;
assign w3118 = pi138 & ~w3117;
assign w3119 = ~pi138 & w3117;
assign w3120 = ~w3118 & ~w3119;
assign w3121 = ~pi885 & w27;
assign w3122 = ~pi335 & ~w27;
assign w3123 = ~w3121 & ~w3122;
assign w3124 = w3120 & ~w3123;
assign w3125 = ~w3120 & w3123;
assign w3126 = ~w3124 & ~w3125;
assign w3127 = pi242 & ~w27;
assign w3128 = ~pi853 & w27;
assign w3129 = ~w3127 & ~w3128;
assign w3130 = w3126 & ~w3129;
assign w3131 = ~w3126 & w3129;
assign w3132 = ~w3130 & ~w3131;
assign w3133 = pi218 & ~w27;
assign w3134 = pi821 & w27;
assign w3135 = ~w3133 & ~w3134;
assign w3136 = ~w3132 & ~w3135;
assign w3137 = w3132 & w3135;
assign w3138 = w1 & ~w3136;
assign w3139 = ~w3137 & w3138;
assign w3140 = ~w3114 & ~w3139;
assign w3141 = ~pi219 & ~w1;
assign w3142 = ~pi916 & w27;
assign w3143 = ~pi433 & ~w27;
assign w3144 = ~w3142 & ~w3143;
assign w3145 = pi177 & ~w3144;
assign w3146 = ~pi177 & w3144;
assign w3147 = ~w3145 & ~w3146;
assign w3148 = ~pi884 & w27;
assign w3149 = ~pi338 & ~w27;
assign w3150 = ~w3148 & ~w3149;
assign w3151 = w3147 & ~w3150;
assign w3152 = ~w3147 & w3150;
assign w3153 = ~w3151 & ~w3152;
assign w3154 = pi241 & ~w27;
assign w3155 = ~pi852 & w27;
assign w3156 = ~w3154 & ~w3155;
assign w3157 = w3153 & ~w3156;
assign w3158 = ~w3153 & w3156;
assign w3159 = ~w3157 & ~w3158;
assign w3160 = pi219 & ~w27;
assign w3161 = pi820 & w27;
assign w3162 = ~w3160 & ~w3161;
assign w3163 = ~w3159 & ~w3162;
assign w3164 = w3159 & w3162;
assign w3165 = w1 & ~w3163;
assign w3166 = ~w3164 & w3165;
assign w3167 = ~w3141 & ~w3166;
assign w3168 = ~pi220 & ~w1;
assign w3169 = ~pi919 & w27;
assign w3170 = ~pi436 & ~w27;
assign w3171 = ~w3169 & ~w3170;
assign w3172 = pi071 & ~w3171;
assign w3173 = ~pi071 & w3171;
assign w3174 = ~w3172 & ~w3173;
assign w3175 = ~pi887 & w27;
assign w3176 = ~pi337 & ~w27;
assign w3177 = ~w3175 & ~w3176;
assign w3178 = w3174 & ~w3177;
assign w3179 = ~w3174 & w3177;
assign w3180 = ~w3178 & ~w3179;
assign w3181 = pi246 & ~w27;
assign w3182 = ~pi855 & w27;
assign w3183 = ~w3181 & ~w3182;
assign w3184 = w3180 & ~w3183;
assign w3185 = ~w3180 & w3183;
assign w3186 = ~w3184 & ~w3185;
assign w3187 = pi220 & ~w27;
assign w3188 = pi823 & w27;
assign w3189 = ~w3187 & ~w3188;
assign w3190 = ~w3186 & ~w3189;
assign w3191 = w3186 & w3189;
assign w3192 = w1 & ~w3190;
assign w3193 = ~w3191 & w3192;
assign w3194 = ~w3168 & ~w3193;
assign w3195 = ~pi221 & ~w1;
assign w3196 = ~pi920 & w27;
assign w3197 = ~pi434 & ~w27;
assign w3198 = ~w3196 & ~w3197;
assign w3199 = pi072 & ~w3198;
assign w3200 = ~pi072 & w3198;
assign w3201 = ~w3199 & ~w3200;
assign w3202 = ~pi888 & w27;
assign w3203 = ~pi339 & ~w27;
assign w3204 = ~w3202 & ~w3203;
assign w3205 = w3201 & ~w3204;
assign w3206 = ~w3201 & w3204;
assign w3207 = ~w3205 & ~w3206;
assign w3208 = pi244 & ~w27;
assign w3209 = ~pi856 & w27;
assign w3210 = ~w3208 & ~w3209;
assign w3211 = w3207 & ~w3210;
assign w3212 = ~w3207 & w3210;
assign w3213 = ~w3211 & ~w3212;
assign w3214 = pi221 & ~w27;
assign w3215 = pi824 & w27;
assign w3216 = ~w3214 & ~w3215;
assign w3217 = ~w3213 & ~w3216;
assign w3218 = w3213 & w3216;
assign w3219 = w1 & ~w3217;
assign w3220 = ~w3218 & w3219;
assign w3221 = ~w3195 & ~w3220;
assign w3222 = ~pi222 & ~w1;
assign w3223 = ~pi918 & w27;
assign w3224 = ~pi432 & ~w27;
assign w3225 = ~w3223 & ~w3224;
assign w3226 = pi135 & ~w3225;
assign w3227 = ~pi135 & w3225;
assign w3228 = ~w3226 & ~w3227;
assign w3229 = ~pi886 & w27;
assign w3230 = ~pi336 & ~w27;
assign w3231 = ~w3229 & ~w3230;
assign w3232 = w3228 & ~w3231;
assign w3233 = ~w3228 & w3231;
assign w3234 = ~w3232 & ~w3233;
assign w3235 = pi243 & ~w27;
assign w3236 = ~pi854 & w27;
assign w3237 = ~w3235 & ~w3236;
assign w3238 = w3234 & ~w3237;
assign w3239 = ~w3234 & w3237;
assign w3240 = ~w3238 & ~w3239;
assign w3241 = pi222 & ~w27;
assign w3242 = pi822 & w27;
assign w3243 = ~w3241 & ~w3242;
assign w3244 = ~w3240 & ~w3243;
assign w3245 = w3240 & w3243;
assign w3246 = w1 & ~w3244;
assign w3247 = ~w3245 & w3246;
assign w3248 = ~w3222 & ~w3247;
assign w3249 = pi223 & ~w1;
assign w3250 = ~w2776 & ~w3249;
assign w3251 = pi224 & ~w1;
assign w3252 = ~w2804 & ~w3251;
assign w3253 = ~pi225 & ~w1;
assign w3254 = ~w2749 & ~w3253;
assign w3255 = ~pi226 & ~w1;
assign w3256 = ~w2694 & ~w3255;
assign w3257 = w1 & w2721;
assign w3258 = pi227 & ~w1;
assign w3259 = ~w3257 & ~w3258;
assign w3260 = pi228 & ~w1;
assign w3261 = w1 & ~w2600;
assign w3262 = ~w3260 & ~w3261;
assign w3263 = pi229 & ~w1;
assign w3264 = w1 & ~w2964;
assign w3265 = ~w3263 & ~w3264;
assign w3266 = pi230 & ~w1;
assign w3267 = w1 & ~w2991;
assign w3268 = ~w3266 & ~w3267;
assign w3269 = pi231 & ~w1;
assign w3270 = w1 & ~w2830;
assign w3271 = ~w3269 & ~w3270;
assign w3272 = pi232 & ~w1;
assign w3273 = w1 & ~w2856;
assign w3274 = ~w3272 & ~w3273;
assign w3275 = pi233 & ~w1;
assign w3276 = w1 & ~w2882;
assign w3277 = ~w3275 & ~w3276;
assign w3278 = pi234 & ~w1;
assign w3279 = w1 & ~w2937;
assign w3280 = ~w3278 & ~w3279;
assign w3281 = pi235 & ~w1;
assign w3282 = w1 & ~w3045;
assign w3283 = ~w3281 & ~w3282;
assign w3284 = pi236 & ~w1;
assign w3285 = w1 & ~w3018;
assign w3286 = ~w3284 & ~w3285;
assign w3287 = pi237 & ~w1;
assign w3288 = ~w2910 & ~w3287;
assign w3289 = w1 & ~w2629;
assign w3290 = pi238 & ~w1;
assign w3291 = ~w3289 & ~w3290;
assign w3292 = pi239 & ~w1;
assign w3293 = w1 & ~w2658;
assign w3294 = ~w3292 & ~w3293;
assign w3295 = pi240 & ~w1;
assign w3296 = w1 & ~w3078;
assign w3297 = ~w3295 & ~w3296;
assign w3298 = pi241 & ~w1;
assign w3299 = w1 & ~w3159;
assign w3300 = ~w3298 & ~w3299;
assign w3301 = pi242 & ~w1;
assign w3302 = w1 & ~w3132;
assign w3303 = ~w3301 & ~w3302;
assign w3304 = pi243 & ~w1;
assign w3305 = w1 & ~w3240;
assign w3306 = ~w3304 & ~w3305;
assign w3307 = pi244 & ~w1;
assign w3308 = w1 & ~w3213;
assign w3309 = ~w3307 & ~w3308;
assign w3310 = pi245 & ~w1;
assign w3311 = w1 & ~w3105;
assign w3312 = ~w3310 & ~w3311;
assign w3313 = pi246 & ~w1;
assign w3314 = w1 & ~w3186;
assign w3315 = ~w3313 & ~w3314;
assign w3316 = pi247 & ~w1;
assign w3317 = w1 & ~w2797;
assign w3318 = ~w3316 & ~w3317;
assign w3319 = w1 & w2715;
assign w3320 = pi248 & ~w1;
assign w3321 = ~w3319 & ~w3320;
assign w3322 = w1 & w2687;
assign w3323 = pi249 & ~w1;
assign w3324 = ~w3322 & ~w3323;
assign w3325 = w1 & w2742;
assign w3326 = pi250 & ~w1;
assign w3327 = ~w3325 & ~w3326;
assign w3328 = w1 & ~w2769;
assign w3329 = pi251 & ~w1;
assign w3330 = ~w3328 & ~w3329;
assign w3331 = w1 & ~w2903;
assign w3332 = pi252 & ~w1;
assign w3333 = ~w3331 & ~w3332;
assign w3334 = ~pi669 & pi673;
assign w3335 = pi673 & w22;
assign w3336 = ~pi555 & pi557;
assign w3337 = w525 & w3336;
assign w3338 = ~w3335 & ~w3337;
assign w3339 = ~pi669 & ~w3338;
assign w3340 = pi666 & ~pi673;
assign w3341 = ~w3339 & ~w3340;
assign w3342 = ~w3334 & w3341;
assign w3343 = ~pi562 & ~w3342;
assign w3344 = w528 & ~w3343;
assign w3345 = ~pi673 & ~w22;
assign w3346 = pi656 & w3345;
assign w3347 = pi126 & w469;
assign w3348 = ~w469 & ~w3345;
assign w3349 = pi734 & w3348;
assign w3350 = ~w3346 & ~w3347;
assign w3351 = ~w3349 & w3350;
assign w3352 = w3344 & ~w3351;
assign w3353 = ~pi673 & w468;
assign w3354 = ~w3335 & ~w3353;
assign w3355 = ~w3339 & w3354;
assign w3356 = ~w3334 & w3355;
assign w3357 = pi126 & ~w3356;
assign w3358 = w3340 & w3355;
assign w3359 = pi656 & w3358;
assign w3360 = ~w3357 & ~w3359;
assign w3361 = ~pi562 & ~w3360;
assign w3362 = ~w3352 & ~w3361;
assign w3363 = pi862 & ~w3362;
assign w3364 = ~pi862 & w3362;
assign w3365 = w2568 & ~w3363;
assign w3366 = ~w3364 & w3365;
assign w3367 = ~w23 & w2553;
assign w3368 = ~pi253 & ~w3367;
assign w3369 = ~pi204 & ~w3362;
assign w3370 = pi204 & w3362;
assign w3371 = ~w3369 & ~w3370;
assign w3372 = w3367 & ~w3371;
assign w3373 = ~w2568 & ~w3368;
assign w3374 = ~w3372 & w3373;
assign w3375 = ~w3366 & ~w3374;
assign w3376 = pi075 & w469;
assign w3377 = pi649 & w3345;
assign w3378 = pi785 & w3348;
assign w3379 = ~w3376 & ~w3377;
assign w3380 = ~w3378 & w3379;
assign w3381 = w3344 & ~w3380;
assign w3382 = pi075 & ~w3356;
assign w3383 = pi649 & w3358;
assign w3384 = ~w3382 & ~w3383;
assign w3385 = ~pi562 & ~w3384;
assign w3386 = ~w3381 & ~w3385;
assign w3387 = pi913 & ~w3386;
assign w3388 = ~pi913 & w3386;
assign w3389 = w2568 & ~w3387;
assign w3390 = ~w3388 & w3389;
assign w3391 = ~pi254 & ~w3367;
assign w3392 = ~pi155 & ~w3386;
assign w3393 = pi155 & w3386;
assign w3394 = ~w3392 & ~w3393;
assign w3395 = w3367 & ~w3394;
assign w3396 = ~w2568 & ~w3391;
assign w3397 = ~w3395 & w3396;
assign w3398 = ~w3390 & ~w3397;
assign w3399 = pi646 & w3345;
assign w3400 = pi127 & w469;
assign w3401 = pi737 & w3348;
assign w3402 = ~w3399 & ~w3400;
assign w3403 = ~w3401 & w3402;
assign w3404 = w3344 & ~w3403;
assign w3405 = pi127 & ~w3356;
assign w3406 = pi646 & w3358;
assign w3407 = ~w3405 & ~w3406;
assign w3408 = ~pi562 & ~w3407;
assign w3409 = ~w3404 & ~w3408;
assign w3410 = pi865 & ~w3409;
assign w3411 = ~pi865 & w3409;
assign w3412 = w2568 & ~w3410;
assign w3413 = ~w3411 & w3412;
assign w3414 = ~pi255 & ~w3367;
assign w3415 = ~pi225 & ~w3409;
assign w3416 = pi225 & w3409;
assign w3417 = ~w3415 & ~w3416;
assign w3418 = w3367 & ~w3417;
assign w3419 = ~w2568 & ~w3414;
assign w3420 = ~w3418 & w3419;
assign w3421 = ~w3413 & ~w3420;
assign w3422 = pi037 & w469;
assign w3423 = pi538 & w3345;
assign w3424 = pi680 & w3348;
assign w3425 = ~w3422 & ~w3423;
assign w3426 = ~w3424 & w3425;
assign w3427 = w3344 & ~w3426;
assign w3428 = pi037 & ~w3356;
assign w3429 = pi538 & w3358;
assign w3430 = ~w3428 & ~w3429;
assign w3431 = ~pi562 & ~w3430;
assign w3432 = ~w3427 & ~w3431;
assign w3433 = pi808 & ~w3432;
assign w3434 = ~pi808 & w3432;
assign w3435 = w2568 & ~w3433;
assign w3436 = ~w3434 & w3435;
assign w3437 = ~pi256 & ~w3367;
assign w3438 = pi209 & ~w3432;
assign w3439 = ~pi209 & w3432;
assign w3440 = ~w3438 & ~w3439;
assign w3441 = w3367 & ~w3440;
assign w3442 = ~w2568 & ~w3437;
assign w3443 = ~w3441 & w3442;
assign w3444 = ~w3436 & ~w3443;
assign w3445 = pi608 & w3345;
assign w3446 = pi083 & w469;
assign w3447 = pi750 & w3348;
assign w3448 = ~w3445 & ~w3446;
assign w3449 = ~w3447 & w3448;
assign w3450 = w3344 & ~w3449;
assign w3451 = pi083 & ~w3356;
assign w3452 = pi608 & w3358;
assign w3453 = ~w3451 & ~w3452;
assign w3454 = ~pi562 & ~w3453;
assign w3455 = ~w3450 & ~w3454;
assign w3456 = pi878 & ~w3455;
assign w3457 = ~pi878 & w3455;
assign w3458 = w2568 & ~w3456;
assign w3459 = ~w3457 & w3458;
assign w3460 = ~pi257 & ~w3367;
assign w3461 = pi044 & ~w3455;
assign w3462 = ~pi044 & w3455;
assign w3463 = ~w3461 & ~w3462;
assign w3464 = w3367 & ~w3463;
assign w3465 = ~w2568 & ~w3460;
assign w3466 = ~w3464 & w3465;
assign w3467 = ~w3459 & ~w3466;
assign w3468 = ~pi185 & w469;
assign w3469 = pi521 & w3345;
assign w3470 = pi699 & w3348;
assign w3471 = ~w3468 & ~w3469;
assign w3472 = ~w3470 & w3471;
assign w3473 = w3344 & ~w3472;
assign w3474 = ~pi185 & ~w3356;
assign w3475 = pi521 & w3358;
assign w3476 = ~w3474 & ~w3475;
assign w3477 = ~pi562 & ~w3476;
assign w3478 = ~w3473 & ~w3477;
assign w3479 = pi827 & ~w3478;
assign w3480 = ~pi827 & w3478;
assign w3481 = w2568 & ~w3479;
assign w3482 = ~w3480 & w3481;
assign w3483 = ~pi258 & ~w3367;
assign w3484 = pi202 & ~w3478;
assign w3485 = ~pi202 & w3478;
assign w3486 = ~w3484 & ~w3485;
assign w3487 = w3367 & ~w3486;
assign w3488 = ~w2568 & ~w3483;
assign w3489 = ~w3487 & w3488;
assign w3490 = ~w3482 & ~w3489;
assign w3491 = pi024 & w469;
assign w3492 = pi592 & w3345;
assign w3493 = pi751 & w3348;
assign w3494 = ~w3491 & ~w3492;
assign w3495 = ~w3493 & w3494;
assign w3496 = w3344 & ~w3495;
assign w3497 = pi024 & ~w3356;
assign w3498 = pi592 & w3358;
assign w3499 = ~w3497 & ~w3498;
assign w3500 = ~pi562 & ~w3499;
assign w3501 = ~w3496 & ~w3500;
assign w3502 = pi879 & ~w3501;
assign w3503 = ~pi879 & w3501;
assign w3504 = w2568 & ~w3502;
assign w3505 = ~w3503 & w3504;
assign w3506 = ~pi259 & ~w3367;
assign w3507 = pi048 & ~w3501;
assign w3508 = ~pi048 & w3501;
assign w3509 = ~w3507 & ~w3508;
assign w3510 = w3367 & ~w3509;
assign w3511 = ~w2568 & ~w3506;
assign w3512 = ~w3510 & w3511;
assign w3513 = ~w3505 & ~w3512;
assign w3514 = pi025 & w469;
assign w3515 = pi593 & w3345;
assign w3516 = pi752 & w3348;
assign w3517 = ~w3514 & ~w3515;
assign w3518 = ~w3516 & w3517;
assign w3519 = w3344 & ~w3518;
assign w3520 = pi025 & ~w3356;
assign w3521 = pi593 & w3358;
assign w3522 = ~w3520 & ~w3521;
assign w3523 = ~pi562 & ~w3522;
assign w3524 = ~w3519 & ~w3523;
assign w3525 = pi880 & ~w3524;
assign w3526 = ~pi880 & w3524;
assign w3527 = w2568 & ~w3525;
assign w3528 = ~w3526 & w3527;
assign w3529 = ~pi260 & ~w3367;
assign w3530 = pi049 & ~w3524;
assign w3531 = ~pi049 & w3524;
assign w3532 = ~w3530 & ~w3531;
assign w3533 = w3367 & ~w3532;
assign w3534 = ~w2568 & ~w3529;
assign w3535 = ~w3533 & w3534;
assign w3536 = ~w3528 & ~w3535;
assign w3537 = pi662 & w3345;
assign w3538 = pi084 & w469;
assign w3539 = pi753 & w3348;
assign w3540 = ~w3537 & ~w3538;
assign w3541 = ~w3539 & w3540;
assign w3542 = w3344 & ~w3541;
assign w3543 = pi084 & ~w3356;
assign w3544 = pi662 & w3358;
assign w3545 = ~w3543 & ~w3544;
assign w3546 = ~pi562 & ~w3545;
assign w3547 = ~w3542 & ~w3546;
assign w3548 = pi881 & ~w3547;
assign w3549 = ~pi881 & w3547;
assign w3550 = w2568 & ~w3548;
assign w3551 = ~w3549 & w3550;
assign w3552 = ~pi261 & ~w3367;
assign w3553 = pi057 & ~w3547;
assign w3554 = ~pi057 & w3547;
assign w3555 = ~w3553 & ~w3554;
assign w3556 = w3367 & ~w3555;
assign w3557 = ~w2568 & ~w3552;
assign w3558 = ~w3556 & w3557;
assign w3559 = ~w3551 & ~w3558;
assign w3560 = pi522 & w3345;
assign w3561 = pi161 & w469;
assign w3562 = pi700 & w3348;
assign w3563 = ~w3560 & ~w3561;
assign w3564 = ~w3562 & w3563;
assign w3565 = w3344 & ~w3564;
assign w3566 = pi161 & ~w3356;
assign w3567 = pi522 & w3358;
assign w3568 = ~w3566 & ~w3567;
assign w3569 = ~pi562 & ~w3568;
assign w3570 = ~w3565 & ~w3569;
assign w3571 = pi828 & ~w3570;
assign w3572 = ~pi828 & w3570;
assign w3573 = w2568 & ~w3571;
assign w3574 = ~w3572 & w3573;
assign w3575 = ~pi262 & ~w3367;
assign w3576 = pi203 & ~w3570;
assign w3577 = ~pi203 & w3570;
assign w3578 = ~w3576 & ~w3577;
assign w3579 = w3367 & ~w3578;
assign w3580 = ~w2568 & ~w3575;
assign w3581 = ~w3579 & w3580;
assign w3582 = ~w3574 & ~w3581;
assign w3583 = pi543 & w3345;
assign w3584 = pi052 & w469;
assign w3585 = pi703 & w3348;
assign w3586 = ~w3583 & ~w3584;
assign w3587 = ~w3585 & w3586;
assign w3588 = w3344 & ~w3587;
assign w3589 = pi052 & ~w3356;
assign w3590 = pi543 & w3358;
assign w3591 = ~w3589 & ~w3590;
assign w3592 = ~pi562 & ~w3591;
assign w3593 = ~w3588 & ~w3592;
assign w3594 = pi831 & ~w3593;
assign w3595 = ~pi831 & w3593;
assign w3596 = w2568 & ~w3594;
assign w3597 = ~w3595 & w3596;
assign w3598 = ~pi263 & ~w3367;
assign w3599 = pi198 & ~w3593;
assign w3600 = ~pi198 & w3593;
assign w3601 = ~w3599 & ~w3600;
assign w3602 = w3367 & ~w3601;
assign w3603 = ~w2568 & ~w3598;
assign w3604 = ~w3602 & w3603;
assign w3605 = ~w3597 & ~w3604;
assign w3606 = pi061 & w469;
assign w3607 = pi527 & w3345;
assign w3608 = pi682 & w3348;
assign w3609 = ~w3606 & ~w3607;
assign w3610 = ~w3608 & w3609;
assign w3611 = w3344 & ~w3610;
assign w3612 = pi061 & ~w3356;
assign w3613 = pi527 & w3358;
assign w3614 = ~w3612 & ~w3613;
assign w3615 = ~pi562 & ~w3614;
assign w3616 = ~w3611 & ~w3615;
assign w3617 = pi810 & ~w3616;
assign w3618 = ~pi810 & w3616;
assign w3619 = w2568 & ~w3617;
assign w3620 = ~w3618 & w3619;
assign w3621 = ~pi264 & ~w3367;
assign w3622 = pi009 & ~w3616;
assign w3623 = ~pi009 & w3616;
assign w3624 = ~w3622 & ~w3623;
assign w3625 = w3367 & ~w3624;
assign w3626 = ~w2568 & ~w3621;
assign w3627 = ~w3625 & w3626;
assign w3628 = ~w3620 & ~w3627;
assign w3629 = pi168 & w469;
assign w3630 = pi571 & w3345;
assign w3631 = pi779 & w3348;
assign w3632 = ~w3629 & ~w3630;
assign w3633 = ~w3631 & w3632;
assign w3634 = w3344 & ~w3633;
assign w3635 = pi168 & ~w3356;
assign w3636 = pi571 & w3358;
assign w3637 = ~w3635 & ~w3636;
assign w3638 = ~pi562 & ~w3637;
assign w3639 = ~w3634 & ~w3638;
assign w3640 = pi907 & ~w3639;
assign w3641 = ~pi907 & w3639;
assign w3642 = w2568 & ~w3640;
assign w3643 = ~w3641 & w3642;
assign w3644 = ~pi265 & ~w3367;
assign w3645 = ~pi176 & ~w3639;
assign w3646 = pi176 & w3639;
assign w3647 = ~w3645 & ~w3646;
assign w3648 = w3367 & ~w3647;
assign w3649 = ~w2568 & ~w3644;
assign w3650 = ~w3648 & w3649;
assign w3651 = ~w3643 & ~w3650;
assign w3652 = ~pi062 & w469;
assign w3653 = pi540 & w3345;
assign w3654 = pi674 & w3348;
assign w3655 = ~w3652 & ~w3653;
assign w3656 = ~w3654 & w3655;
assign w3657 = w3344 & ~w3656;
assign w3658 = ~pi062 & ~w3356;
assign w3659 = pi540 & w3358;
assign w3660 = ~w3658 & ~w3659;
assign w3661 = ~pi562 & ~w3660;
assign w3662 = ~w3657 & ~w3661;
assign w3663 = pi802 & ~w3662;
assign w3664 = ~pi802 & w3662;
assign w3665 = w2568 & ~w3663;
assign w3666 = ~w3664 & w3665;
assign w3667 = ~pi266 & ~w3367;
assign w3668 = pi210 & ~w3662;
assign w3669 = ~pi210 & w3662;
assign w3670 = ~w3668 & ~w3669;
assign w3671 = w3367 & ~w3670;
assign w3672 = ~w2568 & ~w3667;
assign w3673 = ~w3671 & w3672;
assign w3674 = ~w3666 & ~w3673;
assign w3675 = pi139 & w469;
assign w3676 = pi591 & w3345;
assign w3677 = pi780 & w3348;
assign w3678 = ~w3675 & ~w3676;
assign w3679 = ~w3677 & w3678;
assign w3680 = w3344 & ~w3679;
assign w3681 = pi139 & ~w3356;
assign w3682 = pi591 & w3358;
assign w3683 = ~w3681 & ~w3682;
assign w3684 = ~pi562 & ~w3683;
assign w3685 = ~w3680 & ~w3684;
assign w3686 = pi908 & ~w3685;
assign w3687 = ~pi908 & w3685;
assign w3688 = w2568 & ~w3686;
assign w3689 = ~w3687 & w3688;
assign w3690 = ~pi267 & ~w3367;
assign w3691 = ~pi188 & ~w3685;
assign w3692 = pi188 & w3685;
assign w3693 = ~w3691 & ~w3692;
assign w3694 = w3367 & ~w3693;
assign w3695 = ~w2568 & ~w3690;
assign w3696 = ~w3694 & w3695;
assign w3697 = ~w3689 & ~w3696;
assign w3698 = pi636 & w3345;
assign w3699 = pi073 & w469;
assign w3700 = pi781 & w3348;
assign w3701 = ~w3698 & ~w3699;
assign w3702 = ~w3700 & w3701;
assign w3703 = w3344 & ~w3702;
assign w3704 = pi073 & ~w3356;
assign w3705 = pi636 & w3358;
assign w3706 = ~w3704 & ~w3705;
assign w3707 = ~pi562 & ~w3706;
assign w3708 = ~w3703 & ~w3707;
assign w3709 = pi909 & ~w3708;
assign w3710 = ~pi909 & w3708;
assign w3711 = w2568 & ~w3709;
assign w3712 = ~w3710 & w3711;
assign w3713 = ~pi268 & ~w3367;
assign w3714 = ~pi133 & ~w3708;
assign w3715 = pi133 & w3708;
assign w3716 = ~w3714 & ~w3715;
assign w3717 = w3367 & ~w3716;
assign w3718 = ~w2568 & ~w3713;
assign w3719 = ~w3717 & w3718;
assign w3720 = ~w3712 & ~w3719;
assign w3721 = pi594 & w3345;
assign w3722 = pi160 & w469;
assign w3723 = pi796 & w3348;
assign w3724 = ~w3721 & ~w3722;
assign w3725 = ~w3723 & w3724;
assign w3726 = w3344 & ~w3725;
assign w3727 = pi160 & ~w3356;
assign w3728 = pi594 & w3358;
assign w3729 = ~w3727 & ~w3728;
assign w3730 = ~pi562 & ~w3729;
assign w3731 = ~w3726 & ~w3730;
assign w3732 = pi924 & ~w3731;
assign w3733 = ~pi924 & w3731;
assign w3734 = w2568 & ~w3732;
assign w3735 = ~w3733 & w3734;
assign w3736 = ~pi269 & ~w3367;
assign w3737 = pi396 & ~w3731;
assign w3738 = ~pi396 & w3731;
assign w3739 = ~w3737 & ~w3738;
assign w3740 = w3367 & ~w3739;
assign w3741 = ~w2568 & ~w3736;
assign w3742 = ~w3740 & w3741;
assign w3743 = ~w3735 & ~w3742;
assign w3744 = pi100 & w469;
assign w3745 = pi493 & w3345;
assign w3746 = pi677 & w3348;
assign w3747 = ~w3744 & ~w3745;
assign w3748 = ~w3746 & w3747;
assign w3749 = w3344 & ~w3748;
assign w3750 = pi100 & ~w3356;
assign w3751 = pi493 & w3358;
assign w3752 = ~w3750 & ~w3751;
assign w3753 = ~pi562 & ~w3752;
assign w3754 = ~w3749 & ~w3753;
assign w3755 = pi805 & ~w3754;
assign w3756 = ~pi805 & w3754;
assign w3757 = w2568 & ~w3755;
assign w3758 = ~w3756 & w3757;
assign w3759 = ~pi270 & ~w3367;
assign w3760 = pi206 & ~w3754;
assign w3761 = ~pi206 & w3754;
assign w3762 = ~w3760 & ~w3761;
assign w3763 = w3367 & ~w3762;
assign w3764 = ~w2568 & ~w3759;
assign w3765 = ~w3763 & w3764;
assign w3766 = ~w3758 & ~w3765;
assign w3767 = pi169 & w469;
assign w3768 = pi652 & w3345;
assign w3769 = pi715 & w3348;
assign w3770 = ~w3767 & ~w3768;
assign w3771 = ~w3769 & w3770;
assign w3772 = w3344 & ~w3771;
assign w3773 = pi169 & ~w3356;
assign w3774 = pi652 & w3358;
assign w3775 = ~w3773 & ~w3774;
assign w3776 = ~pi562 & ~w3775;
assign w3777 = ~w3772 & ~w3776;
assign w3778 = pi843 & ~w3777;
assign w3779 = ~pi843 & w3777;
assign w3780 = w2568 & ~w3778;
assign w3781 = ~w3779 & w3780;
assign w3782 = ~pi271 & ~w3367;
assign w3783 = pi043 & ~w3777;
assign w3784 = ~pi043 & w3777;
assign w3785 = ~w3783 & ~w3784;
assign w3786 = w3367 & ~w3785;
assign w3787 = ~w2568 & ~w3782;
assign w3788 = ~w3786 & w3787;
assign w3789 = ~w3781 & ~w3788;
assign w3790 = pi119 & w469;
assign w3791 = pi624 & w3345;
assign w3792 = pi797 & w3348;
assign w3793 = ~w3790 & ~w3791;
assign w3794 = ~w3792 & w3793;
assign w3795 = w3344 & ~w3794;
assign w3796 = pi119 & ~w3356;
assign w3797 = pi624 & w3358;
assign w3798 = ~w3796 & ~w3797;
assign w3799 = ~pi562 & ~w3798;
assign w3800 = ~w3795 & ~w3799;
assign w3801 = pi925 & ~w3800;
assign w3802 = ~pi925 & w3800;
assign w3803 = w2568 & ~w3801;
assign w3804 = ~w3802 & w3803;
assign w3805 = ~pi272 & ~w3367;
assign w3806 = pi333 & ~w3800;
assign w3807 = ~pi333 & w3800;
assign w3808 = ~w3806 & ~w3807;
assign w3809 = w3367 & ~w3808;
assign w3810 = ~w2568 & ~w3805;
assign w3811 = ~w3809 & w3810;
assign w3812 = ~w3804 & ~w3811;
assign w3813 = pi638 & w3345;
assign w3814 = pi142 & w469;
assign w3815 = pi716 & w3348;
assign w3816 = ~w3813 & ~w3814;
assign w3817 = ~w3815 & w3816;
assign w3818 = w3344 & ~w3817;
assign w3819 = pi142 & ~w3356;
assign w3820 = pi638 & w3358;
assign w3821 = ~w3819 & ~w3820;
assign w3822 = ~pi562 & ~w3821;
assign w3823 = ~w3818 & ~w3822;
assign w3824 = pi844 & ~w3823;
assign w3825 = ~pi844 & w3823;
assign w3826 = w2568 & ~w3824;
assign w3827 = ~w3825 & w3826;
assign w3828 = ~pi273 & ~w3367;
assign w3829 = pi042 & ~w3823;
assign w3830 = ~pi042 & w3823;
assign w3831 = ~w3829 & ~w3830;
assign w3832 = w3367 & ~w3831;
assign w3833 = ~w2568 & ~w3828;
assign w3834 = ~w3832 & w3833;
assign w3835 = ~w3827 & ~w3834;
assign w3836 = pi607 & w3345;
assign w3837 = pi080 & w469;
assign w3838 = pi717 & w3348;
assign w3839 = ~w3836 & ~w3837;
assign w3840 = ~w3838 & w3839;
assign w3841 = w3344 & ~w3840;
assign w3842 = pi080 & ~w3356;
assign w3843 = pi607 & w3358;
assign w3844 = ~w3842 & ~w3843;
assign w3845 = ~pi562 & ~w3844;
assign w3846 = ~w3841 & ~w3845;
assign w3847 = pi845 & ~w3846;
assign w3848 = ~pi845 & w3846;
assign w3849 = w2568 & ~w3847;
assign w3850 = ~w3848 & w3849;
assign w3851 = ~pi274 & ~w3367;
assign w3852 = pi012 & ~w3846;
assign w3853 = ~pi012 & w3846;
assign w3854 = ~w3852 & ~w3853;
assign w3855 = w3367 & ~w3854;
assign w3856 = ~w2568 & ~w3851;
assign w3857 = ~w3855 & w3856;
assign w3858 = ~w3850 & ~w3857;
assign w3859 = pi637 & w3345;
assign w3860 = pi079 & w469;
assign w3861 = pi718 & w3348;
assign w3862 = ~w3859 & ~w3860;
assign w3863 = ~w3861 & w3862;
assign w3864 = w3344 & ~w3863;
assign w3865 = pi079 & ~w3356;
assign w3866 = pi637 & w3358;
assign w3867 = ~w3865 & ~w3866;
assign w3868 = ~pi562 & ~w3867;
assign w3869 = ~w3864 & ~w3868;
assign w3870 = pi846 & ~w3869;
assign w3871 = ~pi846 & w3869;
assign w3872 = w2568 & ~w3870;
assign w3873 = ~w3871 & w3872;
assign w3874 = ~pi275 & ~w3367;
assign w3875 = pi013 & ~w3869;
assign w3876 = ~pi013 & w3869;
assign w3877 = ~w3875 & ~w3876;
assign w3878 = w3367 & ~w3877;
assign w3879 = ~w2568 & ~w3874;
assign w3880 = ~w3878 & w3879;
assign w3881 = ~w3873 & ~w3880;
assign w3882 = pi074 & w469;
assign w3883 = pi572 & w3345;
assign w3884 = pi782 & w3348;
assign w3885 = ~w3882 & ~w3883;
assign w3886 = ~w3884 & w3885;
assign w3887 = w3344 & ~w3886;
assign w3888 = pi074 & ~w3356;
assign w3889 = pi572 & w3358;
assign w3890 = ~w3888 & ~w3889;
assign w3891 = ~pi562 & ~w3890;
assign w3892 = ~w3887 & ~w3891;
assign w3893 = pi910 & ~w3892;
assign w3894 = ~pi910 & w3892;
assign w3895 = w2568 & ~w3893;
assign w3896 = ~w3894 & w3895;
assign w3897 = ~pi276 & ~w3367;
assign w3898 = ~pi134 & ~w3892;
assign w3899 = pi134 & w3892;
assign w3900 = ~w3898 & ~w3899;
assign w3901 = w3367 & ~w3900;
assign w3902 = ~w2568 & ~w3897;
assign w3903 = ~w3901 & w3902;
assign w3904 = ~w3896 & ~w3903;
assign w3905 = pi615 & w3345;
assign w3906 = pi050 & w469;
assign w3907 = pi799 & w3348;
assign w3908 = ~w3905 & ~w3906;
assign w3909 = ~w3907 & w3908;
assign w3910 = w3344 & ~w3909;
assign w3911 = pi050 & ~w3356;
assign w3912 = pi615 & w3358;
assign w3913 = ~w3911 & ~w3912;
assign w3914 = ~pi562 & ~w3913;
assign w3915 = ~w3910 & ~w3914;
assign w3916 = pi927 & ~w3915;
assign w3917 = ~pi927 & w3915;
assign w3918 = w2568 & ~w3916;
assign w3919 = ~w3917 & w3918;
assign w3920 = ~pi277 & ~w3367;
assign w3921 = pi332 & ~w3915;
assign w3922 = ~pi332 & w3915;
assign w3923 = ~w3921 & ~w3922;
assign w3924 = w3367 & ~w3923;
assign w3925 = ~w2568 & ~w3920;
assign w3926 = ~w3924 & w3925;
assign w3927 = ~w3919 & ~w3926;
assign w3928 = pi622 & w3345;
assign w3929 = pi023 & w469;
assign w3930 = pi720 & w3348;
assign w3931 = ~w3928 & ~w3929;
assign w3932 = ~w3930 & w3931;
assign w3933 = w3344 & ~w3932;
assign w3934 = pi023 & ~w3356;
assign w3935 = pi622 & w3358;
assign w3936 = ~w3934 & ~w3935;
assign w3937 = ~pi562 & ~w3936;
assign w3938 = ~w3933 & ~w3937;
assign w3939 = pi848 & ~w3938;
assign w3940 = ~pi848 & w3938;
assign w3941 = w2568 & ~w3939;
assign w3942 = ~w3940 & w3941;
assign w3943 = ~pi278 & ~w3367;
assign w3944 = pi015 & ~w3938;
assign w3945 = ~pi015 & w3938;
assign w3946 = ~w3944 & ~w3945;
assign w3947 = w3367 & ~w3946;
assign w3948 = ~w2568 & ~w3943;
assign w3949 = ~w3947 & w3948;
assign w3950 = ~w3942 & ~w3949;
assign w3951 = pi605 & w3345;
assign w3952 = pi081 & w469;
assign w3953 = pi721 & w3348;
assign w3954 = ~w3951 & ~w3952;
assign w3955 = ~w3953 & w3954;
assign w3956 = w3344 & ~w3955;
assign w3957 = pi081 & ~w3356;
assign w3958 = pi605 & w3358;
assign w3959 = ~w3957 & ~w3958;
assign w3960 = ~pi562 & ~w3959;
assign w3961 = ~w3956 & ~w3960;
assign w3962 = pi849 & ~w3961;
assign w3963 = ~pi849 & w3961;
assign w3964 = w2568 & ~w3962;
assign w3965 = ~w3963 & w3964;
assign w3966 = ~pi279 & ~w3367;
assign w3967 = pi016 & ~w3961;
assign w3968 = ~pi016 & w3961;
assign w3969 = ~w3967 & ~w3968;
assign w3970 = w3367 & ~w3969;
assign w3971 = ~w2568 & ~w3966;
assign w3972 = ~w3970 & w3971;
assign w3973 = ~w3965 & ~w3972;
assign w3974 = pi601 & w3345;
assign w3975 = pi051 & w469;
assign w3976 = pi800 & w3348;
assign w3977 = ~w3974 & ~w3975;
assign w3978 = ~w3976 & w3977;
assign w3979 = w3344 & ~w3978;
assign w3980 = pi051 & ~w3356;
assign w3981 = pi601 & w3358;
assign w3982 = ~w3980 & ~w3981;
assign w3983 = ~pi562 & ~w3982;
assign w3984 = ~w3979 & ~w3983;
assign w3985 = pi928 & ~w3984;
assign w3986 = ~pi928 & w3984;
assign w3987 = w2568 & ~w3985;
assign w3988 = ~w3986 & w3987;
assign w3989 = ~pi280 & ~w3367;
assign w3990 = pi394 & ~w3984;
assign w3991 = ~pi394 & w3984;
assign w3992 = ~w3990 & ~w3991;
assign w3993 = w3367 & ~w3992;
assign w3994 = ~w2568 & ~w3989;
assign w3995 = ~w3993 & w3994;
assign w3996 = ~w3988 & ~w3995;
assign w3997 = pi660 & w3345;
assign w3998 = pi121 & w469;
assign w3999 = pi801 & w3348;
assign w4000 = ~w3997 & ~w3998;
assign w4001 = ~w3999 & w4000;
assign w4002 = w3344 & ~w4001;
assign w4003 = pi121 & ~w3356;
assign w4004 = pi660 & w3358;
assign w4005 = ~w4003 & ~w4004;
assign w4006 = ~pi562 & ~w4005;
assign w4007 = ~w4002 & ~w4006;
assign w4008 = pi929 & ~w4007;
assign w4009 = ~pi929 & w4007;
assign w4010 = w2568 & ~w4008;
assign w4011 = ~w4009 & w4010;
assign w4012 = ~pi281 & ~w3367;
assign w4013 = pi389 & ~w4007;
assign w4014 = ~pi389 & w4007;
assign w4015 = ~w4013 & ~w4014;
assign w4016 = w3367 & ~w4015;
assign w4017 = ~w2568 & ~w4012;
assign w4018 = ~w4016 & w4017;
assign w4019 = ~w4011 & ~w4018;
assign w4020 = pi525 & w3345;
assign w4021 = pi140 & w469;
assign w4022 = pi684 & w3348;
assign w4023 = ~w4020 & ~w4021;
assign w4024 = ~w4022 & w4023;
assign w4025 = w3344 & ~w4024;
assign w4026 = pi140 & ~w3356;
assign w4027 = pi525 & w3358;
assign w4028 = ~w4026 & ~w4027;
assign w4029 = ~pi562 & ~w4028;
assign w4030 = ~w4025 & ~w4029;
assign w4031 = pi812 & ~w4030;
assign w4032 = ~pi812 & w4030;
assign w4033 = w2568 & ~w4031;
assign w4034 = ~w4032 & w4033;
assign w4035 = ~pi282 & ~w3367;
assign w4036 = pi010 & ~w4030;
assign w4037 = ~pi010 & w4030;
assign w4038 = ~w4036 & ~w4037;
assign w4039 = w3367 & ~w4038;
assign w4040 = ~w2568 & ~w4035;
assign w4041 = ~w4039 & w4040;
assign w4042 = ~w4034 & ~w4041;
assign w4043 = pi530 & w3345;
assign w4044 = pi020 & w469;
assign w4045 = pi687 & w3348;
assign w4046 = ~w4043 & ~w4044;
assign w4047 = ~w4045 & w4046;
assign w4048 = w3344 & ~w4047;
assign w4049 = pi020 & ~w3356;
assign w4050 = pi530 & w3358;
assign w4051 = ~w4049 & ~w4050;
assign w4052 = ~pi562 & ~w4051;
assign w4053 = ~w4048 & ~w4052;
assign w4054 = pi815 & ~w4053;
assign w4055 = ~pi815 & w4053;
assign w4056 = w2568 & ~w4054;
assign w4057 = ~w4055 & w4056;
assign w4058 = ~pi283 & ~w3367;
assign w4059 = pi002 & ~w4053;
assign w4060 = ~pi002 & w4053;
assign w4061 = ~w4059 & ~w4060;
assign w4062 = w3367 & ~w4061;
assign w4063 = ~w2568 & ~w4058;
assign w4064 = ~w4062 & w4063;
assign w4065 = ~w4057 & ~w4064;
assign w4066 = pi573 & w3345;
assign w4067 = pi019 & w469;
assign w4068 = pi784 & w3348;
assign w4069 = ~w4066 & ~w4067;
assign w4070 = ~w4068 & w4069;
assign w4071 = w3344 & ~w4070;
assign w4072 = pi019 & ~w3356;
assign w4073 = pi573 & w3358;
assign w4074 = ~w4072 & ~w4073;
assign w4075 = ~pi562 & ~w4074;
assign w4076 = ~w4071 & ~w4075;
assign w4077 = pi912 & ~w4076;
assign w4078 = ~pi912 & w4076;
assign w4079 = w2568 & ~w4077;
assign w4080 = ~w4078 & w4079;
assign w4081 = ~pi284 & ~w3367;
assign w4082 = pi166 & ~w4076;
assign w4083 = ~pi166 & w4076;
assign w4084 = ~w4082 & ~w4083;
assign w4085 = w3367 & ~w4084;
assign w4086 = ~w2568 & ~w4081;
assign w4087 = ~w4085 & w4086;
assign w4088 = ~w4080 & ~w4087;
assign w4089 = pi626 & w3345;
assign w4090 = pi162 & w469;
assign w4091 = pi732 & w3348;
assign w4092 = ~w4089 & ~w4090;
assign w4093 = ~w4091 & w4092;
assign w4094 = w3344 & ~w4093;
assign w4095 = pi162 & ~w3356;
assign w4096 = pi626 & w3358;
assign w4097 = ~w4095 & ~w4096;
assign w4098 = ~pi562 & ~w4097;
assign w4099 = ~w4094 & ~w4098;
assign w4100 = pi860 & ~w4099;
assign w4101 = ~pi860 & w4099;
assign w4102 = w2568 & ~w4100;
assign w4103 = ~w4101 & w4102;
assign w4104 = ~pi285 & ~w3367;
assign w4105 = ~pi224 & ~w4099;
assign w4106 = pi224 & w4099;
assign w4107 = ~w4105 & ~w4106;
assign w4108 = w3367 & ~w4107;
assign w4109 = ~w2568 & ~w4104;
assign w4110 = ~w4108 & w4109;
assign w4111 = ~w4103 & ~w4110;
assign w4112 = ~pi183 & w469;
assign w4113 = pi586 & w3345;
assign w4114 = pi731 & w3348;
assign w4115 = ~w4112 & ~w4113;
assign w4116 = ~w4114 & w4115;
assign w4117 = w3344 & ~w4116;
assign w4118 = ~pi183 & ~w3356;
assign w4119 = pi586 & w3358;
assign w4120 = ~w4118 & ~w4119;
assign w4121 = ~pi562 & ~w4120;
assign w4122 = ~w4117 & ~w4121;
assign w4123 = pi859 & ~w4122;
assign w4124 = ~pi859 & w4122;
assign w4125 = w2568 & ~w4123;
assign w4126 = ~w4124 & w4125;
assign w4127 = ~pi286 & ~w3367;
assign w4128 = ~pi223 & ~w4122;
assign w4129 = pi223 & w4122;
assign w4130 = ~w4128 & ~w4129;
assign w4131 = w3367 & ~w4130;
assign w4132 = ~w2568 & ~w4127;
assign w4133 = ~w4131 & w4132;
assign w4134 = ~w4126 & ~w4133;
assign w4135 = pi631 & w3345;
assign w4136 = pi125 & w469;
assign w4137 = pi733 & w3348;
assign w4138 = ~w4135 & ~w4136;
assign w4139 = ~w4137 & w4138;
assign w4140 = w3344 & ~w4139;
assign w4141 = pi125 & ~w3356;
assign w4142 = pi631 & w3358;
assign w4143 = ~w4141 & ~w4142;
assign w4144 = ~pi562 & ~w4143;
assign w4145 = ~w4140 & ~w4144;
assign w4146 = pi861 & ~w4145;
assign w4147 = ~pi861 & w4145;
assign w4148 = w2568 & ~w4146;
assign w4149 = ~w4147 & w4148;
assign w4150 = ~pi287 & ~w3367;
assign w4151 = ~pi215 & ~w4145;
assign w4152 = pi215 & w4145;
assign w4153 = ~w4151 & ~w4152;
assign w4154 = w3367 & ~w4153;
assign w4155 = ~w2568 & ~w4150;
assign w4156 = ~w4154 & w4155;
assign w4157 = ~w4149 & ~w4156;
assign w4158 = w1 & w2594;
assign w4159 = pi288 & ~w1;
assign w4160 = ~w4158 & ~w4159;
assign w4161 = w1 & ~w2958;
assign w4162 = pi289 & ~w1;
assign w4163 = ~w4161 & ~w4162;
assign w4164 = w1 & ~w2985;
assign w4165 = pi290 & ~w1;
assign w4166 = ~w4164 & ~w4165;
assign w4167 = w1 & ~w2850;
assign w4168 = pi291 & ~w1;
assign w4169 = ~w4167 & ~w4168;
assign w4170 = w1 & ~w2824;
assign w4171 = pi292 & ~w1;
assign w4172 = ~w4170 & ~w4171;
assign w4173 = w1 & ~w2876;
assign w4174 = pi293 & ~w1;
assign w4175 = ~w4173 & ~w4174;
assign w4176 = w1 & ~w2931;
assign w4177 = pi294 & ~w1;
assign w4178 = ~w4176 & ~w4177;
assign w4179 = w1 & ~w3039;
assign w4180 = pi295 & ~w1;
assign w4181 = ~w4179 & ~w4180;
assign w4182 = w1 & ~w3012;
assign w4183 = pi296 & ~w1;
assign w4184 = ~w4182 & ~w4183;
assign w4185 = pi544 & w3345;
assign w4186 = pi036 & w469;
assign w4187 = pi679 & w3348;
assign w4188 = ~w4185 & ~w4186;
assign w4189 = ~w4187 & w4188;
assign w4190 = w3344 & ~w4189;
assign w4191 = pi036 & ~w3356;
assign w4192 = pi544 & w3358;
assign w4193 = ~w4191 & ~w4192;
assign w4194 = ~pi562 & ~w4193;
assign w4195 = ~w4190 & ~w4194;
assign w4196 = pi807 & ~w4195;
assign w4197 = ~pi807 & w4195;
assign w4198 = w2568 & ~w4196;
assign w4199 = ~w4197 & w4198;
assign w4200 = ~pi297 & ~w3367;
assign w4201 = pi208 & ~w4195;
assign w4202 = ~pi208 & w4195;
assign w4203 = ~w4201 & ~w4202;
assign w4204 = w3367 & ~w4203;
assign w4205 = ~w2568 & ~w4200;
assign w4206 = ~w4204 & w4205;
assign w4207 = ~w4199 & ~w4206;
assign w4208 = w1 & ~w3072;
assign w4209 = pi298 & ~w1;
assign w4210 = ~w4208 & ~w4209;
assign w4211 = pi059 & w469;
assign w4212 = pi648 & w3345;
assign w4213 = pi714 & w3348;
assign w4214 = ~w4211 & ~w4212;
assign w4215 = ~w4213 & w4214;
assign w4216 = w3344 & ~w4215;
assign w4217 = pi059 & ~w3356;
assign w4218 = pi648 & w3358;
assign w4219 = ~w4217 & ~w4218;
assign w4220 = ~pi562 & ~w4219;
assign w4221 = ~w4216 & ~w4220;
assign w4222 = pi842 & ~w4221;
assign w4223 = ~pi842 & w4221;
assign w4224 = w2568 & ~w4222;
assign w4225 = ~w4223 & w4224;
assign w4226 = ~pi299 & ~w3367;
assign w4227 = pi017 & ~w4221;
assign w4228 = ~pi017 & w4221;
assign w4229 = ~w4227 & ~w4228;
assign w4230 = w3367 & ~w4229;
assign w4231 = ~w2568 & ~w4226;
assign w4232 = ~w4230 & w4231;
assign w4233 = ~w4225 & ~w4232;
assign w4234 = pi120 & w469;
assign w4235 = pi642 & w3345;
assign w4236 = pi798 & w3348;
assign w4237 = ~w4234 & ~w4235;
assign w4238 = ~w4236 & w4237;
assign w4239 = w3344 & ~w4238;
assign w4240 = pi120 & ~w3356;
assign w4241 = pi642 & w3358;
assign w4242 = ~w4240 & ~w4241;
assign w4243 = ~pi562 & ~w4242;
assign w4244 = ~w4239 & ~w4243;
assign w4245 = pi926 & ~w4244;
assign w4246 = ~pi926 & w4244;
assign w4247 = w2568 & ~w4245;
assign w4248 = ~w4246 & w4247;
assign w4249 = ~pi300 & ~w3367;
assign w4250 = pi288 & ~w4244;
assign w4251 = ~pi288 & w4244;
assign w4252 = ~w4250 & ~w4251;
assign w4253 = w3367 & ~w4252;
assign w4254 = ~w2568 & ~w4249;
assign w4255 = ~w4253 & w4254;
assign w4256 = ~w4248 & ~w4255;
assign w4257 = pi069 & w469;
assign w4258 = pi645 & w3345;
assign w4259 = pi735 & w3348;
assign w4260 = ~w4257 & ~w4258;
assign w4261 = ~w4259 & w4260;
assign w4262 = w3344 & ~w4261;
assign w4263 = pi069 & ~w3356;
assign w4264 = pi645 & w3358;
assign w4265 = ~w4263 & ~w4264;
assign w4266 = ~pi562 & ~w4265;
assign w4267 = ~w4262 & ~w4266;
assign w4268 = pi863 & ~w4267;
assign w4269 = ~pi863 & w4267;
assign w4270 = w2568 & ~w4268;
assign w4271 = ~w4269 & w4270;
assign w4272 = ~pi301 & ~w3367;
assign w4273 = ~pi214 & ~w4267;
assign w4274 = pi214 & w4267;
assign w4275 = ~w4273 & ~w4274;
assign w4276 = w3367 & ~w4275;
assign w4277 = ~w2568 & ~w4272;
assign w4278 = ~w4276 & w4277;
assign w4279 = ~w4271 & ~w4278;
assign w4280 = pi070 & w469;
assign w4281 = pi619 & w3345;
assign w4282 = pi736 & w3348;
assign w4283 = ~w4280 & ~w4281;
assign w4284 = ~w4282 & w4283;
assign w4285 = w3344 & ~w4284;
assign w4286 = pi070 & ~w3356;
assign w4287 = pi619 & w3358;
assign w4288 = ~w4286 & ~w4287;
assign w4289 = ~pi562 & ~w4288;
assign w4290 = ~w4285 & ~w4289;
assign w4291 = pi864 & ~w4290;
assign w4292 = ~pi864 & w4290;
assign w4293 = w2568 & ~w4291;
assign w4294 = ~w4292 & w4293;
assign w4295 = ~pi302 & ~w3367;
assign w4296 = ~pi226 & ~w4290;
assign w4297 = pi226 & w4290;
assign w4298 = ~w4296 & ~w4297;
assign w4299 = w3367 & ~w4298;
assign w4300 = ~w2568 & ~w4295;
assign w4301 = ~w4299 & w4300;
assign w4302 = ~w4294 & ~w4301;
assign w4303 = ~pi173 & w469;
assign w4304 = pi520 & w3345;
assign w4305 = pi675 & w3348;
assign w4306 = ~w4303 & ~w4304;
assign w4307 = ~w4305 & w4306;
assign w4308 = w3344 & ~w4307;
assign w4309 = ~pi173 & ~w3356;
assign w4310 = pi520 & w3358;
assign w4311 = ~w4309 & ~w4310;
assign w4312 = ~pi562 & ~w4311;
assign w4313 = ~w4308 & ~w4312;
assign w4314 = pi803 & ~w4313;
assign w4315 = ~pi803 & w4313;
assign w4316 = w2568 & ~w4314;
assign w4317 = ~w4315 & w4316;
assign w4318 = ~pi303 & ~w3367;
assign w4319 = pi211 & ~w4313;
assign w4320 = ~pi211 & w4313;
assign w4321 = ~w4319 & ~w4320;
assign w4322 = w3367 & ~w4321;
assign w4323 = ~w2568 & ~w4318;
assign w4324 = ~w4322 & w4323;
assign w4325 = ~w4317 & ~w4324;
assign w4326 = pi170 & w469;
assign w4327 = pi659 & w3345;
assign w4328 = pi747 & w3348;
assign w4329 = ~w4326 & ~w4327;
assign w4330 = ~w4328 & w4329;
assign w4331 = w3344 & ~w4330;
assign w4332 = pi170 & ~w3356;
assign w4333 = pi659 & w3358;
assign w4334 = ~w4332 & ~w4333;
assign w4335 = ~pi562 & ~w4334;
assign w4336 = ~w4331 & ~w4335;
assign w4337 = pi875 & ~w4336;
assign w4338 = ~pi875 & w4336;
assign w4339 = w2568 & ~w4337;
assign w4340 = ~w4338 & w4339;
assign w4341 = ~pi304 & ~w3367;
assign w4342 = ~pi047 & ~w4336;
assign w4343 = pi047 & w4336;
assign w4344 = ~w4342 & ~w4343;
assign w4345 = w3367 & ~w4344;
assign w4346 = ~w2568 & ~w4341;
assign w4347 = ~w4345 & w4346;
assign w4348 = ~w4340 & ~w4347;
assign w4349 = pi141 & w469;
assign w4350 = pi603 & w3345;
assign w4351 = pi748 & w3348;
assign w4352 = ~w4349 & ~w4350;
assign w4353 = ~w4351 & w4352;
assign w4354 = w3344 & ~w4353;
assign w4355 = pi141 & ~w3356;
assign w4356 = pi603 & w3358;
assign w4357 = ~w4355 & ~w4356;
assign w4358 = ~pi562 & ~w4357;
assign w4359 = ~w4354 & ~w4358;
assign w4360 = pi876 & ~w4359;
assign w4361 = ~pi876 & w4359;
assign w4362 = w2568 & ~w4360;
assign w4363 = ~w4361 & w4362;
assign w4364 = ~pi305 & ~w3367;
assign w4365 = ~pi046 & ~w4359;
assign w4366 = pi046 & w4359;
assign w4367 = ~w4365 & ~w4366;
assign w4368 = w3367 & ~w4367;
assign w4369 = ~w2568 & ~w4364;
assign w4370 = ~w4368 & w4369;
assign w4371 = ~w4363 & ~w4370;
assign w4372 = pi107 & w469;
assign w4373 = pi541 & w3345;
assign w4374 = pi698 & w3348;
assign w4375 = ~w4372 & ~w4373;
assign w4376 = ~w4374 & w4375;
assign w4377 = w3344 & ~w4376;
assign w4378 = pi107 & ~w3356;
assign w4379 = pi541 & w3358;
assign w4380 = ~w4378 & ~w4379;
assign w4381 = ~pi562 & ~w4380;
assign w4382 = ~w4377 & ~w4381;
assign w4383 = pi826 & ~w4382;
assign w4384 = ~pi826 & w4382;
assign w4385 = w2568 & ~w4383;
assign w4386 = ~w4384 & w4385;
assign w4387 = ~pi306 & ~w3367;
assign w4388 = pi200 & ~w4382;
assign w4389 = ~pi200 & w4382;
assign w4390 = ~w4388 & ~w4389;
assign w4391 = w3367 & ~w4390;
assign w4392 = ~w2568 & ~w4387;
assign w4393 = ~w4391 & w4392;
assign w4394 = ~w4386 & ~w4393;
assign w4395 = pi582 & w3345;
assign w4396 = pi060 & w469;
assign w4397 = pi746 & w3348;
assign w4398 = ~w4395 & ~w4396;
assign w4399 = ~w4397 & w4398;
assign w4400 = w3344 & ~w4399;
assign w4401 = pi060 & ~w3356;
assign w4402 = pi582 & w3358;
assign w4403 = ~w4401 & ~w4402;
assign w4404 = ~pi562 & ~w4403;
assign w4405 = ~w4400 & ~w4404;
assign w4406 = pi874 & ~w4405;
assign w4407 = ~pi874 & w4405;
assign w4408 = w2568 & ~w4406;
assign w4409 = ~w4407 & w4408;
assign w4410 = ~pi307 & ~w3367;
assign w4411 = pi056 & ~w4405;
assign w4412 = ~pi056 & w4405;
assign w4413 = ~w4411 & ~w4412;
assign w4414 = w3367 & ~w4413;
assign w4415 = ~w2568 & ~w4410;
assign w4416 = ~w4414 & w4415;
assign w4417 = ~w4409 & ~w4416;
assign w4418 = pi101 & w469;
assign w4419 = pi546 & w3345;
assign w4420 = pi681 & w3348;
assign w4421 = ~w4418 & ~w4419;
assign w4422 = ~w4420 & w4421;
assign w4423 = w3344 & ~w4422;
assign w4424 = pi101 & ~w3356;
assign w4425 = pi546 & w3358;
assign w4426 = ~w4424 & ~w4425;
assign w4427 = ~pi562 & ~w4426;
assign w4428 = ~w4423 & ~w4427;
assign w4429 = pi809 & ~w4428;
assign w4430 = ~pi809 & w4428;
assign w4431 = w2568 & ~w4429;
assign w4432 = ~w4430 & w4431;
assign w4433 = ~pi308 & ~w3367;
assign w4434 = pi213 & ~w4428;
assign w4435 = ~pi213 & w4428;
assign w4436 = ~w4434 & ~w4435;
assign w4437 = w3367 & ~w4436;
assign w4438 = ~w2568 & ~w4433;
assign w4439 = ~w4437 & w4438;
assign w4440 = ~w4432 & ~w4439;
assign w4441 = pi123 & w469;
assign w4442 = pi468 & w3345;
assign w4443 = pi702 & w3348;
assign w4444 = ~w4441 & ~w4442;
assign w4445 = ~w4443 & w4444;
assign w4446 = w3344 & ~w4445;
assign w4447 = pi123 & ~w3356;
assign w4448 = pi468 & w3358;
assign w4449 = ~w4447 & ~w4448;
assign w4450 = ~pi562 & ~w4449;
assign w4451 = ~w4446 & ~w4450;
assign w4452 = pi830 & ~w4451;
assign w4453 = ~pi830 & w4451;
assign w4454 = w2568 & ~w4452;
assign w4455 = ~w4453 & w4454;
assign w4456 = ~pi309 & ~w3367;
assign w4457 = pi196 & ~w4451;
assign w4458 = ~pi196 & w4451;
assign w4459 = ~w4457 & ~w4458;
assign w4460 = w3367 & ~w4459;
assign w4461 = ~w2568 & ~w4456;
assign w4462 = ~w4460 & w4461;
assign w4463 = ~w4455 & ~w4462;
assign w4464 = pi569 & w3345;
assign w4465 = pi058 & w469;
assign w4466 = pi778 & w3348;
assign w4467 = ~w4464 & ~w4465;
assign w4468 = ~w4466 & w4467;
assign w4469 = w3344 & ~w4468;
assign w4470 = pi058 & ~w3356;
assign w4471 = pi569 & w3358;
assign w4472 = ~w4470 & ~w4471;
assign w4473 = ~pi562 & ~w4472;
assign w4474 = ~w4469 & ~w4473;
assign w4475 = pi906 & ~w4474;
assign w4476 = ~pi906 & w4474;
assign w4477 = w2568 & ~w4475;
assign w4478 = ~w4476 & w4477;
assign w4479 = ~pi310 & ~w3367;
assign w4480 = ~pi136 & ~w4474;
assign w4481 = pi136 & w4474;
assign w4482 = ~w4480 & ~w4481;
assign w4483 = w3367 & ~w4482;
assign w4484 = ~w2568 & ~w4479;
assign w4485 = ~w4483 & w4484;
assign w4486 = ~w4478 & ~w4485;
assign w4487 = pi534 & w3345;
assign w4488 = pi054 & w469;
assign w4489 = pi704 & w3348;
assign w4490 = ~w4487 & ~w4488;
assign w4491 = ~w4489 & w4490;
assign w4492 = w3344 & ~w4491;
assign w4493 = pi054 & ~w3356;
assign w4494 = pi534 & w3358;
assign w4495 = ~w4493 & ~w4494;
assign w4496 = ~pi562 & ~w4495;
assign w4497 = ~w4492 & ~w4496;
assign w4498 = pi832 & ~w4497;
assign w4499 = ~pi832 & w4497;
assign w4500 = w2568 & ~w4498;
assign w4501 = ~w4499 & w4500;
assign w4502 = ~pi311 & ~w3367;
assign w4503 = pi199 & ~w4497;
assign w4504 = ~pi199 & w4497;
assign w4505 = ~w4503 & ~w4504;
assign w4506 = w3367 & ~w4505;
assign w4507 = ~w2568 & ~w4502;
assign w4508 = ~w4506 & w4507;
assign w4509 = ~w4501 & ~w4508;
assign w4510 = pi524 & w3345;
assign w4511 = pi148 & w469;
assign w4512 = pi676 & w3348;
assign w4513 = ~w4510 & ~w4511;
assign w4514 = ~w4512 & w4513;
assign w4515 = w3344 & ~w4514;
assign w4516 = pi148 & ~w3356;
assign w4517 = pi524 & w3358;
assign w4518 = ~w4516 & ~w4517;
assign w4519 = ~pi562 & ~w4518;
assign w4520 = ~w4515 & ~w4519;
assign w4521 = pi804 & ~w4520;
assign w4522 = ~pi804 & w4520;
assign w4523 = w2568 & ~w4521;
assign w4524 = ~w4522 & w4523;
assign w4525 = ~pi312 & ~w3367;
assign w4526 = pi205 & ~w4520;
assign w4527 = ~pi205 & w4520;
assign w4528 = ~w4526 & ~w4527;
assign w4529 = w3367 & ~w4528;
assign w4530 = ~w2568 & ~w4525;
assign w4531 = ~w4529 & w4530;
assign w4532 = ~w4524 & ~w4531;
assign w4533 = pi548 & w3345;
assign w4534 = pi124 & w469;
assign w4535 = pi705 & w3348;
assign w4536 = ~w4533 & ~w4534;
assign w4537 = ~w4535 & w4536;
assign w4538 = w3344 & ~w4537;
assign w4539 = pi124 & ~w3356;
assign w4540 = pi548 & w3358;
assign w4541 = ~w4539 & ~w4540;
assign w4542 = ~pi562 & ~w4541;
assign w4543 = ~w4538 & ~w4542;
assign w4544 = pi833 & ~w4543;
assign w4545 = ~pi833 & w4543;
assign w4546 = w2568 & ~w4544;
assign w4547 = ~w4545 & w4546;
assign w4548 = ~pi313 & ~w3367;
assign w4549 = pi201 & ~w4543;
assign w4550 = ~pi201 & w4543;
assign w4551 = ~w4549 & ~w4550;
assign w4552 = w3367 & ~w4551;
assign w4553 = ~w2568 & ~w4548;
assign w4554 = ~w4552 & w4553;
assign w4555 = ~w4547 & ~w4554;
assign w4556 = pi602 & w3345;
assign w4557 = pi163 & w469;
assign w4558 = pi764 & w3348;
assign w4559 = ~w4556 & ~w4557;
assign w4560 = ~w4558 & w4559;
assign w4561 = w3344 & ~w4560;
assign w4562 = pi163 & ~w3356;
assign w4563 = pi602 & w3358;
assign w4564 = ~w4562 & ~w4563;
assign w4565 = ~pi562 & ~w4564;
assign w4566 = ~w4561 & ~w4565;
assign w4567 = pi892 & ~w4566;
assign w4568 = ~pi892 & w4566;
assign w4569 = w2568 & ~w4567;
assign w4570 = ~w4568 & w4569;
assign w4571 = ~pi314 & ~w3367;
assign w4572 = ~pi247 & ~w4566;
assign w4573 = pi247 & w4566;
assign w4574 = ~w4572 & ~w4573;
assign w4575 = w3367 & ~w4574;
assign w4576 = ~w2568 & ~w4571;
assign w4577 = ~w4575 & w4576;
assign w4578 = ~w4570 & ~w4577;
assign w4579 = pi584 & w3345;
assign w4580 = pi129 & w469;
assign w4581 = pi765 & w3348;
assign w4582 = ~w4579 & ~w4580;
assign w4583 = ~w4581 & w4582;
assign w4584 = w3344 & ~w4583;
assign w4585 = pi129 & ~w3356;
assign w4586 = pi584 & w3358;
assign w4587 = ~w4585 & ~w4586;
assign w4588 = ~pi562 & ~w4587;
assign w4589 = ~w4584 & ~w4588;
assign w4590 = pi893 & ~w4589;
assign w4591 = ~pi893 & w4589;
assign w4592 = w2568 & ~w4590;
assign w4593 = ~w4591 & w4592;
assign w4594 = ~pi315 & ~w3367;
assign w4595 = pi238 & ~w4589;
assign w4596 = ~pi238 & w4589;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = w3367 & ~w4597;
assign w4599 = ~w2568 & ~w4594;
assign w4600 = ~w4598 & w4599;
assign w4601 = ~w4593 & ~w4600;
assign w4602 = pi130 & w469;
assign w4603 = pi654 & w3345;
assign w4604 = pi766 & w3348;
assign w4605 = ~w4602 & ~w4603;
assign w4606 = ~w4604 & w4605;
assign w4607 = w3344 & ~w4606;
assign w4608 = pi130 & ~w3356;
assign w4609 = pi654 & w3358;
assign w4610 = ~w4608 & ~w4609;
assign w4611 = ~pi562 & ~w4610;
assign w4612 = ~w4607 & ~w4611;
assign w4613 = pi894 & ~w4612;
assign w4614 = ~pi894 & w4612;
assign w4615 = w2568 & ~w4613;
assign w4616 = ~w4614 & w4615;
assign w4617 = ~pi316 & ~w3367;
assign w4618 = ~pi228 & ~w4612;
assign w4619 = pi228 & w4612;
assign w4620 = ~w4618 & ~w4619;
assign w4621 = w3367 & ~w4620;
assign w4622 = ~w2568 & ~w4617;
assign w4623 = ~w4621 & w4622;
assign w4624 = ~w4616 & ~w4623;
assign w4625 = ~pi158 & ~w3356;
assign w4626 = ~pi650 & w3358;
assign w4627 = ~w4625 & ~w4626;
assign w4628 = ~pi562 & ~w4627;
assign w4629 = pi650 & w3345;
assign w4630 = pi158 & w469;
assign w4631 = pi708 & w3348;
assign w4632 = ~w4629 & ~w4630;
assign w4633 = ~w4631 & w4632;
assign w4634 = w3344 & w4633;
assign w4635 = ~w4628 & ~w4634;
assign w4636 = ~pi836 & ~w4635;
assign w4637 = pi836 & w4635;
assign w4638 = w2568 & ~w4636;
assign w4639 = ~w4637 & w4638;
assign w4640 = ~pi317 & ~w3367;
assign w4641 = pi231 & ~w4635;
assign w4642 = ~pi231 & w4635;
assign w4643 = ~w4641 & ~w4642;
assign w4644 = w3367 & ~w4643;
assign w4645 = ~w2568 & ~w4640;
assign w4646 = ~w4644 & w4645;
assign w4647 = ~w4639 & ~w4646;
assign w4648 = pi055 & w469;
assign w4649 = pi590 & w3345;
assign w4650 = pi767 & w3348;
assign w4651 = ~w4648 & ~w4649;
assign w4652 = ~w4650 & w4651;
assign w4653 = w3344 & ~w4652;
assign w4654 = pi055 & ~w3356;
assign w4655 = pi590 & w3358;
assign w4656 = ~w4654 & ~w4655;
assign w4657 = ~pi562 & ~w4656;
assign w4658 = ~w4653 & ~w4657;
assign w4659 = pi895 & ~w4658;
assign w4660 = ~pi895 & w4658;
assign w4661 = w2568 & ~w4659;
assign w4662 = ~w4660 & w4661;
assign w4663 = ~pi318 & ~w3367;
assign w4664 = ~pi239 & ~w4658;
assign w4665 = pi239 & w4658;
assign w4666 = ~w4664 & ~w4665;
assign w4667 = w3367 & ~w4666;
assign w4668 = ~w2568 & ~w4663;
assign w4669 = ~w4667 & w4668;
assign w4670 = ~w4662 & ~w4669;
assign w4671 = pi510 & w3345;
assign w4672 = pi076 & w469;
assign w4673 = pi685 & w3348;
assign w4674 = ~w4671 & ~w4672;
assign w4675 = ~w4673 & w4674;
assign w4676 = w3344 & ~w4675;
assign w4677 = pi076 & ~w3356;
assign w4678 = pi510 & w3358;
assign w4679 = ~w4677 & ~w4678;
assign w4680 = ~pi562 & ~w4679;
assign w4681 = ~w4676 & ~w4680;
assign w4682 = pi813 & ~w4681;
assign w4683 = ~pi813 & w4681;
assign w4684 = w2568 & ~w4682;
assign w4685 = ~w4683 & w4684;
assign w4686 = ~pi319 & ~w3367;
assign w4687 = pi000 & ~w4681;
assign w4688 = ~pi000 & w4681;
assign w4689 = ~w4687 & ~w4688;
assign w4690 = w3367 & ~w4689;
assign w4691 = ~w2568 & ~w4686;
assign w4692 = ~w4690 & w4691;
assign w4693 = ~w4685 & ~w4692;
assign w4694 = pi053 & w469;
assign w4695 = pi639 & w3345;
assign w4696 = pi768 & w3348;
assign w4697 = ~w4694 & ~w4695;
assign w4698 = ~w4696 & w4697;
assign w4699 = w3344 & ~w4698;
assign w4700 = pi053 & ~w3356;
assign w4701 = pi639 & w3358;
assign w4702 = ~w4700 & ~w4701;
assign w4703 = ~pi562 & ~w4702;
assign w4704 = ~w4699 & ~w4703;
assign w4705 = pi896 & ~w4704;
assign w4706 = ~pi896 & w4704;
assign w4707 = w2568 & ~w4705;
assign w4708 = ~w4706 & w4707;
assign w4709 = ~pi320 & ~w3367;
assign w4710 = pi249 & ~w4704;
assign w4711 = ~pi249 & w4704;
assign w4712 = ~w4710 & ~w4711;
assign w4713 = w3367 & ~w4712;
assign w4714 = ~w2568 & ~w4709;
assign w4715 = ~w4713 & w4714;
assign w4716 = ~w4708 & ~w4715;
assign w4717 = pi661 & w3345;
assign w4718 = pi128 & w469;
assign w4719 = pi769 & w3348;
assign w4720 = ~w4717 & ~w4718;
assign w4721 = ~w4719 & w4720;
assign w4722 = w3344 & ~w4721;
assign w4723 = pi128 & ~w3356;
assign w4724 = pi661 & w3358;
assign w4725 = ~w4723 & ~w4724;
assign w4726 = ~pi562 & ~w4725;
assign w4727 = ~w4722 & ~w4726;
assign w4728 = pi897 & ~w4727;
assign w4729 = ~pi897 & w4727;
assign w4730 = w2568 & ~w4728;
assign w4731 = ~w4729 & w4730;
assign w4732 = ~pi321 & ~w3367;
assign w4733 = pi250 & ~w4727;
assign w4734 = ~pi250 & w4727;
assign w4735 = ~w4733 & ~w4734;
assign w4736 = w3367 & ~w4735;
assign w4737 = ~w2568 & ~w4732;
assign w4738 = ~w4736 & w4737;
assign w4739 = ~w4731 & ~w4738;
assign w4740 = pi647 & w3345;
assign w4741 = pi106 & w469;
assign w4742 = pi794 & w3348;
assign w4743 = ~w4740 & ~w4741;
assign w4744 = ~w4742 & w4743;
assign w4745 = w3344 & ~w4744;
assign w4746 = pi106 & ~w3356;
assign w4747 = pi647 & w3358;
assign w4748 = ~w4746 & ~w4747;
assign w4749 = ~pi562 & ~w4748;
assign w4750 = ~w4745 & ~w4749;
assign w4751 = pi922 & ~w4750;
assign w4752 = ~pi922 & w4750;
assign w4753 = w2568 & ~w4751;
assign w4754 = ~w4752 & w4753;
assign w4755 = ~pi322 & ~w3367;
assign w4756 = pi387 & ~w4750;
assign w4757 = ~pi387 & w4750;
assign w4758 = ~w4756 & ~w4757;
assign w4759 = w3367 & ~w4758;
assign w4760 = ~w2568 & ~w4755;
assign w4761 = ~w4759 & w4760;
assign w4762 = ~w4754 & ~w4761;
assign w4763 = pi523 & w3345;
assign w4764 = pi171 & w469;
assign w4765 = pi683 & w3348;
assign w4766 = ~w4763 & ~w4764;
assign w4767 = ~w4765 & w4766;
assign w4768 = w3344 & ~w4767;
assign w4769 = pi171 & ~w3356;
assign w4770 = pi523 & w3358;
assign w4771 = ~w4769 & ~w4770;
assign w4772 = ~pi562 & ~w4771;
assign w4773 = ~w4768 & ~w4772;
assign w4774 = pi811 & ~w4773;
assign w4775 = ~pi811 & w4773;
assign w4776 = w2568 & ~w4774;
assign w4777 = ~w4775 & w4776;
assign w4778 = ~pi323 & ~w3367;
assign w4779 = pi011 & ~w4773;
assign w4780 = ~pi011 & w4773;
assign w4781 = ~w4779 & ~w4780;
assign w4782 = w3367 & ~w4781;
assign w4783 = ~w2568 & ~w4778;
assign w4784 = ~w4782 & w4783;
assign w4785 = ~w4777 & ~w4784;
assign w4786 = pi653 & w3345;
assign w4787 = ~pi187 & w469;
assign w4788 = pi795 & w3348;
assign w4789 = ~w4786 & ~w4787;
assign w4790 = ~w4788 & w4789;
assign w4791 = w3344 & ~w4790;
assign w4792 = ~pi187 & ~w3356;
assign w4793 = pi653 & w3358;
assign w4794 = ~w4792 & ~w4793;
assign w4795 = ~pi562 & ~w4794;
assign w4796 = ~w4791 & ~w4795;
assign w4797 = pi923 & ~w4796;
assign w4798 = ~pi923 & w4796;
assign w4799 = w2568 & ~w4797;
assign w4800 = ~w4798 & w4799;
assign w4801 = ~pi324 & ~w3367;
assign w4802 = pi388 & ~w4796;
assign w4803 = ~pi388 & w4796;
assign w4804 = ~w4802 & ~w4803;
assign w4805 = w3367 & ~w4804;
assign w4806 = ~w2568 & ~w4801;
assign w4807 = ~w4805 & w4806;
assign w4808 = ~w4800 & ~w4807;
assign w4809 = pi022 & w469;
assign w4810 = pi575 & w3345;
assign w4811 = pi719 & w3348;
assign w4812 = ~w4809 & ~w4810;
assign w4813 = ~w4811 & w4812;
assign w4814 = w3344 & ~w4813;
assign w4815 = pi022 & ~w3356;
assign w4816 = pi575 & w3358;
assign w4817 = ~w4815 & ~w4816;
assign w4818 = ~pi562 & ~w4817;
assign w4819 = ~w4814 & ~w4818;
assign w4820 = pi847 & ~w4819;
assign w4821 = ~pi847 & w4819;
assign w4822 = w2568 & ~w4820;
assign w4823 = ~w4821 & w4822;
assign w4824 = ~pi325 & ~w3367;
assign w4825 = pi014 & ~w4819;
assign w4826 = ~pi014 & w4819;
assign w4827 = ~w4825 & ~w4826;
assign w4828 = w3367 & ~w4827;
assign w4829 = ~w2568 & ~w4824;
assign w4830 = ~w4828 & w4829;
assign w4831 = ~w4823 & ~w4830;
assign w4832 = pi093 & w469;
assign w4833 = pi469 & w3345;
assign w4834 = pi678 & w3348;
assign w4835 = ~w4832 & ~w4833;
assign w4836 = ~w4834 & w4835;
assign w4837 = w3344 & ~w4836;
assign w4838 = pi093 & ~w3356;
assign w4839 = pi469 & w3358;
assign w4840 = ~w4838 & ~w4839;
assign w4841 = ~pi562 & ~w4840;
assign w4842 = ~w4837 & ~w4841;
assign w4843 = pi806 & ~w4842;
assign w4844 = ~pi806 & w4842;
assign w4845 = w2568 & ~w4843;
assign w4846 = ~w4844 & w4845;
assign w4847 = ~pi326 & ~w3367;
assign w4848 = pi207 & ~w4842;
assign w4849 = ~pi207 & w4842;
assign w4850 = ~w4848 & ~w4849;
assign w4851 = w3367 & ~w4850;
assign w4852 = ~w2568 & ~w4847;
assign w4853 = ~w4851 & w4852;
assign w4854 = ~w4846 & ~w4853;
assign w4855 = pi466 & w3345;
assign w4856 = pi077 & w469;
assign w4857 = pi686 & w3348;
assign w4858 = ~w4855 & ~w4856;
assign w4859 = ~w4857 & w4858;
assign w4860 = w3344 & ~w4859;
assign w4861 = pi077 & ~w3356;
assign w4862 = pi466 & w3358;
assign w4863 = ~w4861 & ~w4862;
assign w4864 = ~pi562 & ~w4863;
assign w4865 = ~w4860 & ~w4864;
assign w4866 = pi814 & ~w4865;
assign w4867 = ~pi814 & w4865;
assign w4868 = w2568 & ~w4866;
assign w4869 = ~w4867 & w4868;
assign w4870 = ~pi327 & ~w3367;
assign w4871 = pi001 & ~w4865;
assign w4872 = ~pi001 & w4865;
assign w4873 = ~w4871 & ~w4872;
assign w4874 = w3367 & ~w4873;
assign w4875 = ~w2568 & ~w4870;
assign w4876 = ~w4874 & w4875;
assign w4877 = ~w4869 & ~w4876;
assign w4878 = pi612 & w3345;
assign w4879 = pi018 & w469;
assign w4880 = pi783 & w3348;
assign w4881 = ~w4878 & ~w4879;
assign w4882 = ~w4880 & w4881;
assign w4883 = w3344 & ~w4882;
assign w4884 = pi018 & ~w3356;
assign w4885 = pi612 & w3358;
assign w4886 = ~w4884 & ~w4885;
assign w4887 = ~pi562 & ~w4886;
assign w4888 = ~w4883 & ~w4887;
assign w4889 = pi911 & ~w4888;
assign w4890 = ~pi911 & w4888;
assign w4891 = w2568 & ~w4889;
assign w4892 = ~w4890 & w4891;
assign w4893 = ~pi328 & ~w3367;
assign w4894 = pi167 & ~w4888;
assign w4895 = ~pi167 & w4888;
assign w4896 = ~w4894 & ~w4895;
assign w4897 = w3367 & ~w4896;
assign w4898 = ~w2568 & ~w4893;
assign w4899 = ~w4897 & w4898;
assign w4900 = ~w4892 & ~w4899;
assign w4901 = pi021 & w469;
assign w4902 = pi539 & w3345;
assign w4903 = pi688 & w3348;
assign w4904 = ~w4901 & ~w4902;
assign w4905 = ~w4903 & w4904;
assign w4906 = w3344 & ~w4905;
assign w4907 = pi021 & ~w3356;
assign w4908 = pi539 & w3358;
assign w4909 = ~w4907 & ~w4908;
assign w4910 = ~pi562 & ~w4909;
assign w4911 = ~w4906 & ~w4910;
assign w4912 = pi816 & ~w4911;
assign w4913 = ~pi816 & w4911;
assign w4914 = w2568 & ~w4912;
assign w4915 = ~w4913 & w4914;
assign w4916 = ~pi329 & ~w3367;
assign w4917 = pi003 & ~w4911;
assign w4918 = ~pi003 & w4911;
assign w4919 = ~w4917 & ~w4918;
assign w4920 = w3367 & ~w4919;
assign w4921 = ~w2568 & ~w4916;
assign w4922 = ~w4920 & w4921;
assign w4923 = ~w4915 & ~w4922;
assign w4924 = pi108 & w469;
assign w4925 = pi604 & w3345;
assign w4926 = pi730 & w3348;
assign w4927 = ~w4924 & ~w4925;
assign w4928 = ~w4926 & w4927;
assign w4929 = w3344 & ~w4928;
assign w4930 = pi108 & ~w3356;
assign w4931 = pi604 & w3358;
assign w4932 = ~w4930 & ~w4931;
assign w4933 = ~pi562 & ~w4932;
assign w4934 = ~w4929 & ~w4933;
assign w4935 = pi858 & ~w4934;
assign w4936 = ~pi858 & w4934;
assign w4937 = w2568 & ~w4935;
assign w4938 = ~w4936 & w4937;
assign w4939 = ~pi330 & ~w3367;
assign w4940 = ~pi227 & ~w4934;
assign w4941 = pi227 & w4934;
assign w4942 = ~w4940 & ~w4941;
assign w4943 = w3367 & ~w4942;
assign w4944 = ~w2568 & ~w4939;
assign w4945 = ~w4943 & w4944;
assign w4946 = ~w4938 & ~w4945;
assign w4947 = pi549 & w3345;
assign w4948 = pi078 & w469;
assign w4949 = pi689 & w3348;
assign w4950 = ~w4947 & ~w4948;
assign w4951 = ~w4949 & w4950;
assign w4952 = w3344 & ~w4951;
assign w4953 = pi078 & ~w3356;
assign w4954 = pi549 & w3358;
assign w4955 = ~w4953 & ~w4954;
assign w4956 = ~pi562 & ~w4955;
assign w4957 = ~w4952 & ~w4956;
assign w4958 = pi817 & ~w4957;
assign w4959 = ~pi817 & w4957;
assign w4960 = w2568 & ~w4958;
assign w4961 = ~w4959 & w4960;
assign w4962 = ~pi331 & ~w3367;
assign w4963 = pi004 & ~w4957;
assign w4964 = ~pi004 & w4957;
assign w4965 = ~w4963 & ~w4964;
assign w4966 = w3367 & ~w4965;
assign w4967 = ~w2568 & ~w4962;
assign w4968 = ~w4966 & w4967;
assign w4969 = ~w4961 & ~w4968;
assign w4970 = pi332 & ~w1;
assign w4971 = w1 & ~w2652;
assign w4972 = ~w4970 & ~w4971;
assign w4973 = w1 & w2626;
assign w4974 = pi333 & ~w1;
assign w4975 = ~w4973 & ~w4974;
assign w4976 = w1 & ~w3099;
assign w4977 = pi334 & ~w1;
assign w4978 = ~w4976 & ~w4977;
assign w4979 = w1 & ~w3126;
assign w4980 = pi335 & ~w1;
assign w4981 = ~w4979 & ~w4980;
assign w4982 = w1 & ~w3234;
assign w4983 = pi336 & ~w1;
assign w4984 = ~w4982 & ~w4983;
assign w4985 = w1 & ~w3180;
assign w4986 = pi337 & ~w1;
assign w4987 = ~w4985 & ~w4986;
assign w4988 = w1 & ~w3153;
assign w4989 = pi338 & ~w1;
assign w4990 = ~w4988 & ~w4989;
assign w4991 = w1 & ~w3207;
assign w4992 = pi339 & ~w1;
assign w4993 = ~w4991 & ~w4992;
assign w4994 = pi122 & w469;
assign w4995 = pi509 & w3345;
assign w4996 = pi701 & w3348;
assign w4997 = ~w4994 & ~w4995;
assign w4998 = ~w4996 & w4997;
assign w4999 = w3344 & ~w4998;
assign w5000 = pi122 & ~w3356;
assign w5001 = pi509 & w3358;
assign w5002 = ~w5000 & ~w5001;
assign w5003 = ~pi562 & ~w5002;
assign w5004 = ~w4999 & ~w5003;
assign w5005 = pi829 & ~w5004;
assign w5006 = ~pi829 & w5004;
assign w5007 = w2568 & ~w5005;
assign w5008 = ~w5006 & w5007;
assign w5009 = ~pi340 & ~w3367;
assign w5010 = pi197 & ~w5004;
assign w5011 = ~pi197 & w5004;
assign w5012 = ~w5010 & ~w5011;
assign w5013 = w3367 & ~w5012;
assign w5014 = ~w2568 & ~w5009;
assign w5015 = ~w5013 & w5014;
assign w5016 = ~w5008 & ~w5015;
assign w5017 = pi644 & w3345;
assign w5018 = pi082 & w469;
assign w5019 = pi749 & w3348;
assign w5020 = ~w5017 & ~w5018;
assign w5021 = ~w5019 & w5020;
assign w5022 = w3344 & ~w5021;
assign w5023 = pi082 & ~w3356;
assign w5024 = pi644 & w3358;
assign w5025 = ~w5023 & ~w5024;
assign w5026 = ~pi562 & ~w5025;
assign w5027 = ~w5022 & ~w5026;
assign w5028 = pi877 & ~w5027;
assign w5029 = ~pi877 & w5027;
assign w5030 = w2568 & ~w5028;
assign w5031 = ~w5029 & w5030;
assign w5032 = ~pi341 & ~w3367;
assign w5033 = pi045 & ~w5027;
assign w5034 = ~pi045 & w5027;
assign w5035 = ~w5033 & ~w5034;
assign w5036 = w3367 & ~w5035;
assign w5037 = ~w2568 & ~w5032;
assign w5038 = ~w5036 & w5037;
assign w5039 = ~w5031 & ~w5038;
assign w5040 = pi112 & ~w3356;
assign w5041 = pi664 & w3358;
assign w5042 = ~w5040 & ~w5041;
assign w5043 = ~pi562 & ~w5042;
assign w5044 = pi774 & w3348;
assign w5045 = pi664 & w3345;
assign w5046 = ~w468 & w2028;
assign w5047 = ~w5045 & ~w5046;
assign w5048 = ~w5044 & w5047;
assign w5049 = w3344 & ~w5048;
assign w5050 = ~w5043 & ~w5049;
assign w5051 = pi902 & ~w5050;
assign w5052 = ~pi902 & w5050;
assign w5053 = w2568 & ~w5051;
assign w5054 = ~w5052 & w5053;
assign w5055 = ~pi342 & ~w3367;
assign w5056 = pi415 & ~w5050;
assign w5057 = ~pi415 & w5050;
assign w5058 = ~w5056 & ~w5057;
assign w5059 = w3367 & ~w5058;
assign w5060 = ~w2568 & ~w5055;
assign w5061 = ~w5059 & w5060;
assign w5062 = ~w5054 & ~w5061;
assign w5063 = ~pi182 & ~w3356;
assign w5064 = ~pi587 & w3358;
assign w5065 = ~w5063 & ~w5064;
assign w5066 = ~pi562 & ~w5065;
assign w5067 = pi587 & w3345;
assign w5068 = pi182 & w469;
assign w5069 = pi707 & w3348;
assign w5070 = ~w5067 & ~w5068;
assign w5071 = ~w5069 & w5070;
assign w5072 = w3344 & w5071;
assign w5073 = ~w5066 & ~w5072;
assign w5074 = ~pi835 & ~w5073;
assign w5075 = pi835 & w5073;
assign w5076 = w2568 & ~w5074;
assign w5077 = ~w5075 & w5076;
assign w5078 = ~pi343 & ~w3367;
assign w5079 = pi230 & ~w5073;
assign w5080 = ~pi230 & w5073;
assign w5081 = ~w5079 & ~w5080;
assign w5082 = w3367 & ~w5081;
assign w5083 = ~w2568 & ~w5078;
assign w5084 = ~w5082 & w5083;
assign w5085 = ~w5077 & ~w5084;
assign w5086 = pi085 & w469;
assign w5087 = pi611 & w3345;
assign w5088 = pi777 & w3348;
assign w5089 = ~w5086 & ~w5087;
assign w5090 = ~w5088 & w5089;
assign w5091 = w3344 & ~w5090;
assign w5092 = pi085 & ~w3356;
assign w5093 = pi611 & w3358;
assign w5094 = ~w5092 & ~w5093;
assign w5095 = ~pi562 & ~w5094;
assign w5096 = ~w5091 & ~w5095;
assign w5097 = pi905 & ~w5096;
assign w5098 = ~pi905 & w5096;
assign w5099 = w2568 & ~w5097;
assign w5100 = ~w5098 & w5099;
assign w5101 = ~pi344 & ~w3367;
assign w5102 = pi418 & ~w5096;
assign w5103 = ~pi418 & w5096;
assign w5104 = ~w5102 & ~w5103;
assign w5105 = w3367 & ~w5104;
assign w5106 = ~w2568 & ~w5101;
assign w5107 = ~w5105 & w5106;
assign w5108 = ~w5100 & ~w5107;
assign w5109 = pi152 & w469;
assign w5110 = pi579 & w3345;
assign w5111 = pi772 & w3348;
assign w5112 = ~w5109 & ~w5110;
assign w5113 = ~w5111 & w5112;
assign w5114 = w3344 & ~w5113;
assign w5115 = pi152 & ~w3356;
assign w5116 = pi579 & w3358;
assign w5117 = ~w5115 & ~w5116;
assign w5118 = ~pi562 & ~w5117;
assign w5119 = ~w5114 & ~w5118;
assign w5120 = pi900 & ~w5119;
assign w5121 = ~pi900 & w5119;
assign w5122 = w2568 & ~w5120;
assign w5123 = ~w5121 & w5122;
assign w5124 = ~pi345 & ~w3367;
assign w5125 = pi414 & ~w5119;
assign w5126 = ~pi414 & w5119;
assign w5127 = ~w5125 & ~w5126;
assign w5128 = w3367 & ~w5127;
assign w5129 = ~w2568 & ~w5124;
assign w5130 = ~w5128 & w5129;
assign w5131 = ~w5123 & ~w5130;
assign w5132 = ~pi115 & ~w3356;
assign w5133 = ~pi663 & w3358;
assign w5134 = ~w5132 & ~w5133;
assign w5135 = ~pi562 & ~w5134;
assign w5136 = pi663 & w3345;
assign w5137 = pi115 & w469;
assign w5138 = pi709 & w3348;
assign w5139 = ~w5136 & ~w5137;
assign w5140 = ~w5138 & w5139;
assign w5141 = w3344 & w5140;
assign w5142 = ~w5135 & ~w5141;
assign w5143 = ~pi837 & ~w5142;
assign w5144 = pi837 & w5142;
assign w5145 = w2568 & ~w5143;
assign w5146 = ~w5144 & w5145;
assign w5147 = ~pi346 & ~w3367;
assign w5148 = pi232 & ~w5142;
assign w5149 = ~pi232 & w5142;
assign w5150 = ~w5148 & ~w5149;
assign w5151 = w3367 & ~w5150;
assign w5152 = ~w2568 & ~w5147;
assign w5153 = ~w5151 & w5152;
assign w5154 = ~w5146 & ~w5153;
assign w5155 = ~pi669 & ~pi673;
assign w5156 = pi435 & w469;
assign w5157 = ~w5155 & ~w5156;
assign w5158 = ~pi562 & ~w3338;
assign w5159 = ~pi560 & ~pi561;
assign w5160 = ~w5157 & w5159;
assign w5161 = ~w5158 & w5160;
assign w5162 = pi560 & pi561;
assign w5163 = pi407 & w5162;
assign w5164 = ~pi560 & pi561;
assign w5165 = pi406 & w5164;
assign w5166 = pi560 & ~pi561;
assign w5167 = pi395 & w5166;
assign w5168 = pi397 & w5161;
assign w5169 = ~w5163 & ~w5165;
assign w5170 = ~w5167 & w5169;
assign w5171 = w469 & w5170;
assign w5172 = ~w5168 & w5171;
assign w5173 = pi151 & w5166;
assign w5174 = pi149 & w5164;
assign w5175 = pi147 & w5162;
assign w5176 = pi143 & w5161;
assign w5177 = ~w5173 & ~w5174;
assign w5178 = ~w5175 & w5177;
assign w5179 = ~w469 & w5178;
assign w5180 = ~w5176 & w5179;
assign w5181 = ~w5172 & ~w5180;
assign w5182 = pi323 & w5162;
assign w5183 = pi271 & w5164;
assign w5184 = pi304 & w5166;
assign w5185 = pi265 & w5161;
assign w5186 = ~w5182 & ~w5183;
assign w5187 = ~w5184 & w5186;
assign w5188 = w469 & w5187;
assign w5189 = ~w5185 & w5188;
assign w5190 = pi171 & w5162;
assign w5191 = pi169 & w5164;
assign w5192 = pi170 & w5166;
assign w5193 = pi168 & w5161;
assign w5194 = ~w5190 & ~w5191;
assign w5195 = ~w5192 & w5194;
assign w5196 = ~w469 & w5195;
assign w5197 = ~w5193 & w5196;
assign w5198 = ~w5189 & ~w5197;
assign w5199 = pi303 & w5162;
assign w5200 = pi343 & w5164;
assign w5201 = pi354 & w5166;
assign w5202 = pi377 & w5161;
assign w5203 = ~w5199 & ~w5200;
assign w5204 = ~w5201 & w5203;
assign w5205 = w469 & w5204;
assign w5206 = ~w5202 & w5205;
assign w5207 = ~pi173 & w5162;
assign w5208 = pi174 & w5166;
assign w5209 = pi182 & w5164;
assign w5210 = pi175 & w5161;
assign w5211 = ~w5207 & ~w5208;
assign w5212 = ~w5209 & w5211;
assign w5213 = ~w469 & w5212;
assign w5214 = ~w5210 & w5213;
assign w5215 = ~w5206 & ~w5214;
assign w5216 = ~w5198 & ~w5215;
assign w5217 = w5198 & w5215;
assign w5218 = ~w5216 & ~w5217;
assign w5219 = ~w5181 & ~w5218;
assign w5220 = w5181 & w5218;
assign w5221 = ~w5219 & ~w5220;
assign w5222 = pi367 & w5166;
assign w5223 = pi383 & w5164;
assign w5224 = pi386 & w5162;
assign w5225 = pi403 & w5161;
assign w5226 = ~w5222 & ~w5223;
assign w5227 = ~w5224 & w5226;
assign w5228 = w469 & w5227;
assign w5229 = ~w5225 & w5228;
assign w5230 = pi172 & w5162;
assign w5231 = pi180 & w5164;
assign w5232 = pi179 & w5166;
assign w5233 = pi181 & w5161;
assign w5234 = ~w5230 & ~w5231;
assign w5235 = ~w5232 & w5234;
assign w5236 = ~w469 & w5235;
assign w5237 = ~w5233 & w5236;
assign w5238 = ~w5229 & ~w5237;
assign w5239 = pi356 & w5166;
assign w5240 = pi317 & w5164;
assign w5241 = pi312 & w5162;
assign w5242 = pi345 & w5161;
assign w5243 = ~w5239 & ~w5240;
assign w5244 = ~w5241 & w5243;
assign w5245 = w469 & w5244;
assign w5246 = ~w5242 & w5245;
assign w5247 = pi148 & w5162;
assign w5248 = pi150 & w5166;
assign w5249 = pi158 & w5164;
assign w5250 = pi152 & w5161;
assign w5251 = ~w5247 & ~w5248;
assign w5252 = ~w5249 & w5251;
assign w5253 = ~w469 & w5252;
assign w5254 = ~w5250 & w5253;
assign w5255 = ~w5246 & ~w5254;
assign w5256 = pi258 & w5162;
assign w5257 = pi286 & w5164;
assign w5258 = pi392 & w5166;
assign w5259 = pi324 & w5161;
assign w5260 = ~w5256 & ~w5257;
assign w5261 = ~w5258 & w5260;
assign w5262 = w469 & w5261;
assign w5263 = ~w5259 & w5262;
assign w5264 = ~pi183 & w5164;
assign w5265 = ~pi185 & w5162;
assign w5266 = ~pi184 & w5166;
assign w5267 = ~pi187 & w5161;
assign w5268 = ~w5264 & ~w5265;
assign w5269 = ~w5266 & w5268;
assign w5270 = ~w469 & w5269;
assign w5271 = ~w5267 & w5270;
assign w5272 = ~w5263 & ~w5271;
assign w5273 = w5255 & ~w5272;
assign w5274 = ~w5255 & w5272;
assign w5275 = ~w5273 & ~w5274;
assign w5276 = w5238 & w5275;
assign w5277 = ~w5238 & ~w5275;
assign w5278 = ~w5276 & ~w5277;
assign w5279 = ~w5221 & ~w5278;
assign w5280 = w5221 & w5278;
assign w5281 = ~w5279 & ~w5280;
assign w5282 = ~pi673 & ~w5281;
assign w5283 = pi359 & w5166;
assign w5284 = pi380 & w5164;
assign w5285 = pi297 & w5162;
assign w5286 = pi351 & w5161;
assign w5287 = ~w5283 & ~w5284;
assign w5288 = ~w5285 & w5287;
assign w5289 = w469 & w5288;
assign w5290 = ~w5286 & w5289;
assign w5291 = pi036 & w5162;
assign w5292 = pi032 & w5164;
assign w5293 = pi039 & w5166;
assign w5294 = pi027 & w5161;
assign w5295 = ~w5291 & ~w5292;
assign w5296 = ~w5293 & w5295;
assign w5297 = ~w469 & w5296;
assign w5298 = ~w5294 & w5297;
assign w5299 = ~w5290 & ~w5298;
assign w5300 = pi362 & w5161;
assign w5301 = pi361 & w5166;
assign w5302 = pi381 & w5164;
assign w5303 = pi256 & w5162;
assign w5304 = ~w5301 & ~w5302;
assign w5305 = ~w5303 & w5304;
assign w5306 = w469 & w5305;
assign w5307 = ~w5300 & w5306;
assign w5308 = pi026 & w5161;
assign w5309 = pi033 & w5164;
assign w5310 = pi037 & w5162;
assign w5311 = pi038 & w5166;
assign w5312 = ~w5309 & ~w5310;
assign w5313 = ~w5311 & w5312;
assign w5314 = ~w469 & w5313;
assign w5315 = ~w5308 & w5314;
assign w5316 = ~w5307 & ~w5315;
assign w5317 = pi391 & w5161;
assign w5318 = pi370 & w5166;
assign w5319 = pi398 & w5164;
assign w5320 = pi360 & w5162;
assign w5321 = ~w5318 & ~w5319;
assign w5322 = ~w5320 & w5321;
assign w5323 = w469 & w5322;
assign w5324 = ~w5317 & w5323;
assign w5325 = pi028 & w5161;
assign w5326 = pi041 & w5166;
assign w5327 = pi031 & w5162;
assign w5328 = pi035 & w5164;
assign w5329 = ~w5326 & ~w5327;
assign w5330 = ~w5328 & w5329;
assign w5331 = ~w469 & w5330;
assign w5332 = ~w5325 & w5331;
assign w5333 = ~w5324 & ~w5332;
assign w5334 = ~w5316 & ~w5333;
assign w5335 = w5316 & w5333;
assign w5336 = ~w5334 & ~w5335;
assign w5337 = ~w5299 & ~w5336;
assign w5338 = w5299 & w5336;
assign w5339 = ~w5337 & ~w5338;
assign w5340 = pi358 & w5162;
assign w5341 = pi402 & w5164;
assign w5342 = pi369 & w5166;
assign w5343 = pi393 & w5161;
assign w5344 = ~w5340 & ~w5341;
assign w5345 = ~w5342 & w5344;
assign w5346 = w469 & w5345;
assign w5347 = ~w5343 & w5346;
assign w5348 = pi030 & w5162;
assign w5349 = pi034 & w5164;
assign w5350 = pi040 & w5166;
assign w5351 = pi029 & w5161;
assign w5352 = ~w5348 & ~w5349;
assign w5353 = ~w5350 & w5352;
assign w5354 = ~w469 & w5353;
assign w5355 = ~w5351 & w5354;
assign w5356 = ~w5347 & ~w5355;
assign w5357 = pi328 & w5161;
assign w5358 = pi259 & w5166;
assign w5359 = pi325 & w5164;
assign w5360 = pi283 & w5162;
assign w5361 = ~w5358 & ~w5359;
assign w5362 = ~w5360 & w5361;
assign w5363 = w469 & w5362;
assign w5364 = ~w5357 & w5363;
assign w5365 = pi018 & w5161;
assign w5366 = pi024 & w5166;
assign w5367 = pi020 & w5162;
assign w5368 = pi022 & w5164;
assign w5369 = ~w5366 & ~w5367;
assign w5370 = ~w5368 & w5369;
assign w5371 = ~w469 & w5370;
assign w5372 = ~w5365 & w5371;
assign w5373 = ~w5364 & ~w5372;
assign w5374 = pi277 & w5161;
assign w5375 = pi318 & w5166;
assign w5376 = pi301 & w5164;
assign w5377 = pi263 & w5162;
assign w5378 = ~w5375 & ~w5376;
assign w5379 = ~w5377 & w5378;
assign w5380 = w469 & w5379;
assign w5381 = ~w5374 & w5380;
assign w5382 = pi050 & w5161;
assign w5383 = pi069 & w5164;
assign w5384 = pi052 & w5162;
assign w5385 = pi055 & w5166;
assign w5386 = ~w5383 & ~w5384;
assign w5387 = ~w5385 & w5386;
assign w5388 = ~w469 & w5387;
assign w5389 = ~w5382 & w5388;
assign w5390 = ~w5381 & ~w5389;
assign w5391 = ~w5373 & ~w5390;
assign w5392 = w5373 & w5390;
assign w5393 = ~w5391 & ~w5392;
assign w5394 = ~w5356 & ~w5393;
assign w5395 = w5356 & w5393;
assign w5396 = ~w5394 & ~w5395;
assign w5397 = w5339 & ~w5396;
assign w5398 = ~w5339 & w5396;
assign w5399 = ~w5397 & ~w5398;
assign w5400 = pi085 & w5161;
assign w5401 = pi102 & w5166;
assign w5402 = pi101 & w5162;
assign w5403 = pi116 & w5164;
assign w5404 = ~w5401 & ~w5402;
assign w5405 = ~w5403 & w5404;
assign w5406 = ~w469 & w5405;
assign w5407 = ~w5400 & w5406;
assign w5408 = pi344 & w5161;
assign w5409 = pi308 & w5162;
assign w5410 = pi382 & w5164;
assign w5411 = pi399 & w5166;
assign w5412 = ~w5409 & ~w5410;
assign w5413 = ~w5411 & w5412;
assign w5414 = w469 & w5413;
assign w5415 = ~w5408 & w5414;
assign w5416 = ~w5407 & ~w5415;
assign w5417 = pi375 & w5161;
assign w5418 = pi363 & w5162;
assign w5419 = pi385 & w5164;
assign w5420 = pi372 & w5166;
assign w5421 = ~w5418 & ~w5419;
assign w5422 = ~w5420 & w5421;
assign w5423 = w469 & w5422;
assign w5424 = ~w5417 & w5423;
assign w5425 = pi088 & w5161;
assign w5426 = pi096 & w5164;
assign w5427 = pi091 & w5162;
assign w5428 = pi105 & w5166;
assign w5429 = ~w5426 & ~w5427;
assign w5430 = ~w5428 & w5429;
assign w5431 = ~w469 & w5430;
assign w5432 = ~w5425 & w5431;
assign w5433 = ~w5424 & ~w5432;
assign w5434 = ~w5416 & ~w5433;
assign w5435 = w5416 & w5433;
assign w5436 = ~w5434 & ~w5435;
assign w5437 = pi284 & w5161;
assign w5438 = pi329 & w5162;
assign w5439 = pi260 & w5166;
assign w5440 = pi278 & w5164;
assign w5441 = ~w5438 & ~w5439;
assign w5442 = ~w5440 & w5441;
assign w5443 = w469 & w5442;
assign w5444 = ~w5437 & w5443;
assign w5445 = pi019 & w5161;
assign w5446 = pi023 & w5164;
assign w5447 = pi021 & w5162;
assign w5448 = pi025 & w5166;
assign w5449 = ~w5446 & ~w5447;
assign w5450 = ~w5448 & w5449;
assign w5451 = ~w469 & w5450;
assign w5452 = ~w5445 & w5451;
assign w5453 = ~w5444 & ~w5452;
assign w5454 = pi280 & w5161;
assign w5455 = pi311 & w5162;
assign w5456 = pi320 & w5166;
assign w5457 = pi302 & w5164;
assign w5458 = ~w5455 & ~w5456;
assign w5459 = ~w5457 & w5458;
assign w5460 = w469 & w5459;
assign w5461 = ~w5454 & w5460;
assign w5462 = pi051 & w5161;
assign w5463 = pi053 & w5166;
assign w5464 = pi054 & w5162;
assign w5465 = pi070 & w5164;
assign w5466 = ~w5463 & ~w5464;
assign w5467 = ~w5465 & w5466;
assign w5468 = ~w469 & w5467;
assign w5469 = ~w5462 & w5468;
assign w5470 = ~w5461 & ~w5469;
assign w5471 = ~w5453 & ~w5470;
assign w5472 = w5453 & w5470;
assign w5473 = ~w5471 & ~w5472;
assign w5474 = w5336 & ~w5473;
assign w5475 = ~w5336 & w5473;
assign w5476 = ~w5474 & ~w5475;
assign w5477 = w5436 & w5476;
assign w5478 = ~w5436 & ~w5476;
assign w5479 = ~w5477 & ~w5478;
assign w5480 = w5399 & w5479;
assign w5481 = ~w5399 & ~w5479;
assign w5482 = pi673 & ~w5480;
assign w5483 = ~w5481 & w5482;
assign w5484 = ~w5282 & ~w5483;
assign w5485 = pi257 & w5166;
assign w5486 = pi275 & w5164;
assign w5487 = pi327 & w5162;
assign w5488 = pi276 & w5161;
assign w5489 = ~w5485 & ~w5486;
assign w5490 = ~w5487 & w5489;
assign w5491 = w469 & w5490;
assign w5492 = ~w5488 & w5491;
assign w5493 = pi077 & w5162;
assign w5494 = pi079 & w5164;
assign w5495 = pi083 & w5166;
assign w5496 = pi074 & w5161;
assign w5497 = ~w5493 & ~w5494;
assign w5498 = ~w5495 & w5497;
assign w5499 = ~w469 & w5498;
assign w5500 = ~w5496 & w5499;
assign w5501 = ~w5492 & ~w5500;
assign w5502 = ~w5281 & w5501;
assign w5503 = w5281 & ~w5501;
assign w5504 = ~w5502 & ~w5503;
assign w5505 = w5484 & w5504;
assign w5506 = ~w5484 & ~w5504;
assign w5507 = ~w5505 & ~w5506;
assign w5508 = pi316 & w5166;
assign w5509 = pi253 & w5164;
assign w5510 = pi309 & w5162;
assign w5511 = pi300 & w5161;
assign w5512 = ~w5508 & ~w5509;
assign w5513 = ~w5510 & w5512;
assign w5514 = w469 & w5513;
assign w5515 = ~w5511 & w5514;
assign w5516 = pi123 & w5162;
assign w5517 = pi130 & w5166;
assign w5518 = pi126 & w5164;
assign w5519 = pi120 & w5161;
assign w5520 = ~w5516 & ~w5517;
assign w5521 = ~w5518 & w5520;
assign w5522 = ~w469 & w5521;
assign w5523 = ~w5519 & w5522;
assign w5524 = ~w5515 & ~w5523;
assign w5525 = pi384 & w5164;
assign w5526 = pi355 & w5162;
assign w5527 = pi371 & w5166;
assign w5528 = pi365 & w5161;
assign w5529 = ~w5525 & ~w5526;
assign w5530 = ~w5527 & w5529;
assign w5531 = w469 & w5530;
assign w5532 = ~w5528 & w5531;
assign w5533 = pi095 & w5164;
assign w5534 = pi103 & w5166;
assign w5535 = pi089 & w5162;
assign w5536 = pi087 & w5161;
assign w5537 = ~w5533 & ~w5534;
assign w5538 = ~w5535 & w5537;
assign w5539 = ~w469 & w5538;
assign w5540 = ~w5536 & w5539;
assign w5541 = ~w5532 & ~w5540;
assign w5542 = ~w5524 & ~w5541;
assign w5543 = w5524 & w5541;
assign w5544 = ~w5542 & ~w5543;
assign w5545 = pi121 & w5161;
assign w5546 = pi128 & w5166;
assign w5547 = pi124 & w5162;
assign w5548 = pi127 & w5164;
assign w5549 = ~w5546 & ~w5547;
assign w5550 = ~w5548 & w5549;
assign w5551 = ~w469 & w5550;
assign w5552 = ~w5545 & w5551;
assign w5553 = pi281 & w5161;
assign w5554 = pi313 & w5162;
assign w5555 = pi255 & w5164;
assign w5556 = pi321 & w5166;
assign w5557 = ~w5554 & ~w5555;
assign w5558 = ~w5556 & w5557;
assign w5559 = w469 & w5558;
assign w5560 = ~w5553 & w5559;
assign w5561 = ~w5552 & ~w5560;
assign w5562 = ~w5416 & ~w5561;
assign w5563 = w5416 & w5561;
assign w5564 = ~w5562 & ~w5563;
assign w5565 = pi357 & w5166;
assign w5566 = pi346 & w5164;
assign w5567 = pi270 & w5162;
assign w5568 = pi379 & w5161;
assign w5569 = ~w5565 & ~w5566;
assign w5570 = ~w5567 & w5569;
assign w5571 = w469 & w5570;
assign w5572 = ~w5568 & w5571;
assign w5573 = pi100 & w5162;
assign w5574 = pi115 & w5164;
assign w5575 = pi099 & w5166;
assign w5576 = pi118 & w5161;
assign w5577 = ~w5573 & ~w5574;
assign w5578 = ~w5575 & w5577;
assign w5579 = ~w469 & w5578;
assign w5580 = ~w5576 & w5579;
assign w5581 = ~w5572 & ~w5580;
assign w5582 = pi315 & w5166;
assign w5583 = pi287 & w5164;
assign w5584 = pi340 & w5162;
assign w5585 = pi272 & w5161;
assign w5586 = ~w5582 & ~w5583;
assign w5587 = ~w5584 & w5586;
assign w5588 = w469 & w5587;
assign w5589 = ~w5585 & w5588;
assign w5590 = pi122 & w5162;
assign w5591 = pi129 & w5166;
assign w5592 = pi125 & w5164;
assign w5593 = pi119 & w5161;
assign w5594 = ~w5590 & ~w5591;
assign w5595 = ~w5592 & w5594;
assign w5596 = ~w469 & w5595;
assign w5597 = ~w5593 & w5596;
assign w5598 = ~w5589 & ~w5597;
assign w5599 = ~w5581 & ~w5598;
assign w5600 = w5581 & w5598;
assign w5601 = ~w5599 & ~w5600;
assign w5602 = w5564 & ~w5601;
assign w5603 = ~w5564 & w5601;
assign w5604 = ~w5602 & ~w5603;
assign w5605 = w5544 & w5604;
assign w5606 = ~w5544 & ~w5604;
assign w5607 = ~w5605 & ~w5606;
assign w5608 = ~w5507 & ~w5607;
assign w5609 = w5161 & w5608;
assign w5610 = w5161 & w5607;
assign w5611 = w5507 & w5610;
assign w5612 = pi347 & ~w5161;
assign w5613 = ~w5611 & ~w5612;
assign w5614 = ~w5609 & w5613;
assign w5615 = w5524 & ~w5581;
assign w5616 = ~w5524 & w5581;
assign w5617 = ~w5615 & ~w5616;
assign w5618 = pi319 & w5162;
assign w5619 = pi274 & w5164;
assign w5620 = pi341 & w5166;
assign w5621 = pi268 & w5161;
assign w5622 = ~w5618 & ~w5619;
assign w5623 = ~w5620 & w5622;
assign w5624 = w469 & w5623;
assign w5625 = ~w5621 & w5624;
assign w5626 = pi082 & w5166;
assign w5627 = pi080 & w5164;
assign w5628 = pi076 & w5162;
assign w5629 = pi073 & w5161;
assign w5630 = ~w5626 & ~w5627;
assign w5631 = ~w5628 & w5630;
assign w5632 = ~w469 & w5631;
assign w5633 = ~w5629 & w5632;
assign w5634 = ~w5625 & ~w5633;
assign w5635 = pi254 & w5161;
assign w5636 = pi331 & w5162;
assign w5637 = pi279 & w5164;
assign w5638 = pi261 & w5166;
assign w5639 = ~w5636 & ~w5637;
assign w5640 = ~w5638 & w5639;
assign w5641 = w469 & w5640;
assign w5642 = ~w5635 & w5641;
assign w5643 = pi075 & w5161;
assign w5644 = pi081 & w5164;
assign w5645 = pi078 & w5162;
assign w5646 = pi084 & w5166;
assign w5647 = ~w5644 & ~w5645;
assign w5648 = ~w5646 & w5647;
assign w5649 = ~w469 & w5648;
assign w5650 = ~w5643 & w5649;
assign w5651 = ~w5642 & ~w5650;
assign w5652 = ~w5416 & ~w5651;
assign w5653 = w5416 & w5651;
assign w5654 = ~w5652 & ~w5653;
assign w5655 = w5634 & ~w5654;
assign w5656 = ~w5634 & w5654;
assign w5657 = ~w5655 & ~w5656;
assign w5658 = w5617 & w5657;
assign w5659 = ~w5617 & ~w5657;
assign w5660 = ~w5658 & ~w5659;
assign w5661 = pi305 & w5166;
assign w5662 = pi273 & w5164;
assign w5663 = pi282 & w5162;
assign w5664 = pi267 & w5161;
assign w5665 = ~w5661 & ~w5662;
assign w5666 = ~w5663 & w5665;
assign w5667 = w469 & w5666;
assign w5668 = ~w5664 & w5667;
assign w5669 = pi140 & w5162;
assign w5670 = pi142 & w5164;
assign w5671 = pi141 & w5166;
assign w5672 = pi139 & w5161;
assign w5673 = ~w5669 & ~w5670;
assign w5674 = ~w5671 & w5673;
assign w5675 = ~w469 & w5674;
assign w5676 = ~w5672 & w5675;
assign w5677 = ~w5668 & ~w5676;
assign w5678 = ~w5215 & ~w5272;
assign w5679 = w5215 & w5272;
assign w5680 = ~w5678 & ~w5679;
assign w5681 = ~w5677 & ~w5680;
assign w5682 = w5677 & w5680;
assign w5683 = ~w5681 & ~w5682;
assign w5684 = pi314 & w5166;
assign w5685 = pi285 & w5164;
assign w5686 = pi262 & w5162;
assign w5687 = pi269 & w5161;
assign w5688 = ~w5684 & ~w5685;
assign w5689 = ~w5686 & w5688;
assign w5690 = w469 & w5689;
assign w5691 = ~w5687 & w5690;
assign w5692 = pi161 & w5162;
assign w5693 = pi163 & w5166;
assign w5694 = pi162 & w5164;
assign w5695 = pi160 & w5161;
assign w5696 = ~w5692 & ~w5693;
assign w5697 = ~w5694 & w5696;
assign w5698 = ~w469 & w5697;
assign w5699 = ~w5695 & w5698;
assign w5700 = ~w5691 & ~w5699;
assign w5701 = w5238 & ~w5700;
assign w5702 = ~w5238 & w5700;
assign w5703 = ~w5701 & ~w5702;
assign w5704 = w5198 & w5703;
assign w5705 = ~w5198 & ~w5703;
assign w5706 = ~w5704 & ~w5705;
assign w5707 = ~w5683 & ~w5706;
assign w5708 = w5683 & w5706;
assign w5709 = ~w5707 & ~w5708;
assign w5710 = ~pi673 & ~w5709;
assign w5711 = ~w5299 & ~w5473;
assign w5712 = w5299 & w5473;
assign w5713 = ~w5711 & ~w5712;
assign w5714 = w5396 & ~w5713;
assign w5715 = ~w5396 & w5713;
assign w5716 = ~w5714 & ~w5715;
assign w5717 = ~w5561 & ~w5651;
assign w5718 = w5561 & w5651;
assign w5719 = ~w5717 & ~w5718;
assign w5720 = w5476 & w5719;
assign w5721 = ~w5476 & ~w5719;
assign w5722 = ~w5720 & ~w5721;
assign w5723 = w5716 & w5722;
assign w5724 = ~w5716 & ~w5722;
assign w5725 = pi673 & ~w5723;
assign w5726 = ~w5724 & w5725;
assign w5727 = ~w5710 & ~w5726;
assign w5728 = pi401 & w5166;
assign w5729 = pi326 & w5162;
assign w5730 = pi378 & w5164;
assign w5731 = pi342 & w5161;
assign w5732 = ~w5728 & ~w5729;
assign w5733 = ~w5730 & w5732;
assign w5734 = w469 & w5733;
assign w5735 = ~w5731 & w5734;
assign w5736 = pi093 & w5162;
assign w5737 = pi098 & w5166;
assign w5738 = pi097 & w5164;
assign w5739 = pi112 & w5161;
assign w5740 = ~w5736 & ~w5737;
assign w5741 = ~w5738 & w5740;
assign w5742 = ~w469 & w5741;
assign w5743 = ~w5739 & w5742;
assign w5744 = ~w5735 & ~w5743;
assign w5745 = ~w5541 & ~w5744;
assign w5746 = w5541 & w5744;
assign w5747 = ~w5745 & ~w5746;
assign w5748 = w5709 & ~w5747;
assign w5749 = ~w5709 & w5747;
assign w5750 = ~w5748 & ~w5749;
assign w5751 = w5727 & w5750;
assign w5752 = ~w5727 & ~w5750;
assign w5753 = ~w5751 & ~w5752;
assign w5754 = w5660 & ~w5753;
assign w5755 = w5161 & w5754;
assign w5756 = w5161 & ~w5660;
assign w5757 = w5753 & w5756;
assign w5758 = pi348 & ~w5161;
assign w5759 = ~w5757 & ~w5758;
assign w5760 = ~w5755 & w5759;
assign w5761 = ~w5524 & ~w5744;
assign w5762 = w5524 & w5744;
assign w5763 = ~w5761 & ~w5762;
assign w5764 = ~w5433 & ~w5651;
assign w5765 = w5433 & w5651;
assign w5766 = ~w5764 & ~w5765;
assign w5767 = pi404 & w5162;
assign w5768 = pi405 & w5164;
assign w5769 = pi368 & w5166;
assign w5770 = pi364 & w5161;
assign w5771 = ~w5767 & ~w5768;
assign w5772 = ~w5769 & w5771;
assign w5773 = w469 & w5772;
assign w5774 = ~w5770 & w5773;
assign w5775 = pi104 & w5166;
assign w5776 = pi094 & w5164;
assign w5777 = pi090 & w5162;
assign w5778 = pi086 & w5161;
assign w5779 = ~w5775 & ~w5776;
assign w5780 = ~w5777 & w5779;
assign w5781 = ~w469 & w5780;
assign w5782 = ~w5778 & w5781;
assign w5783 = ~w5774 & ~w5782;
assign w5784 = w5634 & ~w5783;
assign w5785 = ~w5634 & w5783;
assign w5786 = ~w5784 & ~w5785;
assign w5787 = w5766 & w5786;
assign w5788 = ~w5766 & ~w5786;
assign w5789 = ~w5787 & ~w5788;
assign w5790 = w5763 & w5789;
assign w5791 = ~w5763 & ~w5789;
assign w5792 = ~w5790 & ~w5791;
assign w5793 = ~w5507 & ~w5792;
assign w5794 = w5161 & w5793;
assign w5795 = w5161 & w5792;
assign w5796 = w5507 & w5795;
assign w5797 = pi349 & ~w5161;
assign w5798 = ~w5796 & ~w5797;
assign w5799 = ~w5794 & w5798;
assign w5800 = ~w5433 & ~w5561;
assign w5801 = w5433 & w5561;
assign w5802 = ~w5800 & ~w5801;
assign w5803 = w5501 & ~w5802;
assign w5804 = ~w5501 & w5802;
assign w5805 = ~w5803 & ~w5804;
assign w5806 = w5598 & ~w5805;
assign w5807 = ~w5598 & w5805;
assign w5808 = ~w5806 & ~w5807;
assign w5809 = w5783 & w5808;
assign w5810 = ~w5783 & ~w5808;
assign w5811 = ~w5809 & ~w5810;
assign w5812 = w5753 & ~w5811;
assign w5813 = w5161 & w5812;
assign w5814 = w5161 & w5811;
assign w5815 = ~w5753 & w5814;
assign w5816 = pi350 & ~w5161;
assign w5817 = ~w5815 & ~w5816;
assign w5818 = ~w5813 & w5817;
assign w5819 = pi027 & w469;
assign w5820 = pi628 & w3345;
assign w5821 = pi775 & w3348;
assign w5822 = ~w5819 & ~w5820;
assign w5823 = ~w5821 & w5822;
assign w5824 = w3344 & ~w5823;
assign w5825 = pi027 & ~w3356;
assign w5826 = pi628 & w3358;
assign w5827 = ~w5825 & ~w5826;
assign w5828 = ~pi562 & ~w5827;
assign w5829 = ~w5824 & ~w5828;
assign w5830 = pi903 & ~w5829;
assign w5831 = ~pi903 & w5829;
assign w5832 = w2568 & ~w5830;
assign w5833 = ~w5831 & w5832;
assign w5834 = ~pi351 & ~w3367;
assign w5835 = pi416 & ~w5829;
assign w5836 = ~pi416 & w5829;
assign w5837 = ~w5835 & ~w5836;
assign w5838 = w3367 & ~w5837;
assign w5839 = ~w2568 & ~w5834;
assign w5840 = ~w5838 & w5839;
assign w5841 = ~w5833 & ~w5840;
assign w5842 = ~pi063 & ~w3356;
assign w5843 = ~pi574 & w3358;
assign w5844 = ~w5842 & ~w5843;
assign w5845 = ~pi562 & ~w5844;
assign w5846 = pi574 & w3345;
assign w5847 = pi063 & w469;
assign w5848 = pi786 & w3348;
assign w5849 = ~w5846 & ~w5847;
assign w5850 = ~w5848 & w5849;
assign w5851 = w3344 & w5850;
assign w5852 = ~w5845 & ~w5851;
assign w5853 = ~pi914 & ~w5852;
assign w5854 = pi914 & w5852;
assign w5855 = w2568 & ~w5853;
assign w5856 = ~w5854 & w5855;
assign w5857 = ~pi352 & ~w3367;
assign w5858 = ~pi430 & ~w5852;
assign w5859 = pi430 & w5852;
assign w5860 = ~w5858 & ~w5859;
assign w5861 = w3367 & ~w5860;
assign w5862 = ~w2568 & ~w5857;
assign w5863 = ~w5861 & w5862;
assign w5864 = ~w5856 & ~w5863;
assign w5865 = pi595 & w3345;
assign w5866 = pi065 & w469;
assign w5867 = pi738 & w3348;
assign w5868 = ~w5865 & ~w5866;
assign w5869 = ~w5867 & w5868;
assign w5870 = pi562 & ~w5869;
assign w5871 = ~pi065 & ~w3355;
assign w5872 = ~w3334 & ~w3340;
assign w5873 = ~w1836 & ~w5872;
assign w5874 = ~w3334 & ~w5869;
assign w5875 = w3355 & ~w5873;
assign w5876 = ~w5874 & w5875;
assign w5877 = ~pi595 & w3358;
assign w5878 = ~pi562 & ~w5871;
assign w5879 = ~w5876 & w5878;
assign w5880 = ~w5877 & w5879;
assign w5881 = ~w5870 & ~w5880;
assign w5882 = pi866 & ~w5881;
assign w5883 = ~pi866 & w5881;
assign w5884 = w2568 & ~w5882;
assign w5885 = ~w5883 & w5884;
assign w5886 = ~pi353 & ~w3367;
assign w5887 = pi289 & ~w5881;
assign w5888 = ~pi289 & w5881;
assign w5889 = ~w5887 & ~w5888;
assign w5890 = w3367 & ~w5889;
assign w5891 = ~w2568 & ~w5886;
assign w5892 = ~w5890 & w5891;
assign w5893 = ~w5885 & ~w5892;
assign w5894 = pi588 & w3345;
assign w5895 = pi174 & w469;
assign w5896 = pi739 & w3348;
assign w5897 = ~w5894 & ~w5895;
assign w5898 = ~w5896 & w5897;
assign w5899 = pi562 & ~w5898;
assign w5900 = ~pi174 & ~w3355;
assign w5901 = ~w2463 & ~w5872;
assign w5902 = ~w3334 & ~w5898;
assign w5903 = w3355 & ~w5901;
assign w5904 = ~w5902 & w5903;
assign w5905 = ~pi588 & w3358;
assign w5906 = ~pi562 & ~w5900;
assign w5907 = ~w5904 & w5906;
assign w5908 = ~w5905 & w5907;
assign w5909 = ~w5899 & ~w5908;
assign w5910 = pi867 & ~w5909;
assign w5911 = ~pi867 & w5909;
assign w5912 = w2568 & ~w5910;
assign w5913 = ~w5911 & w5912;
assign w5914 = ~pi354 & ~w3367;
assign w5915 = pi290 & ~w5909;
assign w5916 = ~pi290 & w5909;
assign w5917 = ~w5915 & ~w5916;
assign w5918 = w3367 & ~w5917;
assign w5919 = ~w2568 & ~w5914;
assign w5920 = ~w5918 & w5919;
assign w5921 = ~w5913 & ~w5920;
assign w5922 = pi089 & w469;
assign w5923 = pi467 & w3345;
assign w5924 = pi694 & w3348;
assign w5925 = ~w5922 & ~w5923;
assign w5926 = ~w5924 & w5925;
assign w5927 = pi562 & ~w5926;
assign w5928 = ~pi089 & ~w3355;
assign w5929 = ~w1971 & ~w5872;
assign w5930 = ~w3334 & ~w5926;
assign w5931 = w3355 & ~w5929;
assign w5932 = ~w5930 & w5931;
assign w5933 = ~pi467 & w3358;
assign w5934 = ~pi562 & ~w5928;
assign w5935 = ~w5932 & w5934;
assign w5936 = ~w5933 & w5935;
assign w5937 = ~w5927 & ~w5936;
assign w5938 = pi822 & ~w5937;
assign w5939 = ~pi822 & w5937;
assign w5940 = w2568 & ~w5938;
assign w5941 = ~w5939 & w5940;
assign w5942 = ~pi355 & ~w3367;
assign w5943 = pi222 & ~w5937;
assign w5944 = ~pi222 & w5937;
assign w5945 = ~w5943 & ~w5944;
assign w5946 = w3367 & ~w5945;
assign w5947 = ~w2568 & ~w5942;
assign w5948 = ~w5946 & w5947;
assign w5949 = ~w5941 & ~w5948;
assign w5950 = pi150 & w469;
assign w5951 = pi634 & w3345;
assign w5952 = pi740 & w3348;
assign w5953 = ~w5950 & ~w5951;
assign w5954 = ~w5952 & w5953;
assign w5955 = pi562 & ~w5954;
assign w5956 = ~pi150 & ~w3355;
assign w5957 = ~w2360 & ~w5872;
assign w5958 = ~w3334 & ~w5954;
assign w5959 = w3355 & ~w5957;
assign w5960 = ~w5958 & w5959;
assign w5961 = ~pi634 & w3358;
assign w5962 = ~pi562 & ~w5956;
assign w5963 = ~w5960 & w5962;
assign w5964 = ~w5961 & w5963;
assign w5965 = ~w5955 & ~w5964;
assign w5966 = pi868 & ~w5965;
assign w5967 = ~pi868 & w5965;
assign w5968 = w2568 & ~w5966;
assign w5969 = ~w5967 & w5968;
assign w5970 = ~pi356 & ~w3367;
assign w5971 = pi292 & ~w5965;
assign w5972 = ~pi292 & w5965;
assign w5973 = ~w5971 & ~w5972;
assign w5974 = w3367 & ~w5973;
assign w5975 = ~w2568 & ~w5970;
assign w5976 = ~w5974 & w5975;
assign w5977 = ~w5969 & ~w5976;
assign w5978 = pi576 & w3345;
assign w5979 = pi099 & w469;
assign w5980 = pi741 & w3348;
assign w5981 = ~w5978 & ~w5979;
assign w5982 = ~w5980 & w5981;
assign w5983 = pi562 & ~w5982;
assign w5984 = ~pi099 & ~w3355;
assign w5985 = ~w2201 & ~w5872;
assign w5986 = ~w3334 & ~w5982;
assign w5987 = w3355 & ~w5985;
assign w5988 = ~w5986 & w5987;
assign w5989 = ~pi576 & w3358;
assign w5990 = ~pi562 & ~w5984;
assign w5991 = ~w5988 & w5990;
assign w5992 = ~w5989 & w5991;
assign w5993 = ~w5983 & ~w5992;
assign w5994 = pi869 & ~w5993;
assign w5995 = ~pi869 & w5993;
assign w5996 = w2568 & ~w5994;
assign w5997 = ~w5995 & w5996;
assign w5998 = ~pi357 & ~w3367;
assign w5999 = pi291 & ~w5993;
assign w6000 = ~pi291 & w5993;
assign w6001 = ~w5999 & ~w6000;
assign w6002 = w3367 & ~w6001;
assign w6003 = ~w2568 & ~w5998;
assign w6004 = ~w6002 & w6003;
assign w6005 = ~w5997 & ~w6004;
assign w6006 = pi531 & w3345;
assign w6007 = pi030 & w469;
assign w6008 = pi695 & w3348;
assign w6009 = ~w6006 & ~w6007;
assign w6010 = ~w6008 & w6009;
assign w6011 = pi562 & ~w6010;
assign w6012 = ~pi030 & ~w3355;
assign w6013 = ~w1569 & ~w5872;
assign w6014 = ~w3334 & ~w6010;
assign w6015 = w3355 & ~w6013;
assign w6016 = ~w6014 & w6015;
assign w6017 = ~pi531 & w3358;
assign w6018 = ~pi562 & ~w6012;
assign w6019 = ~w6016 & w6018;
assign w6020 = ~w6017 & w6019;
assign w6021 = ~w6011 & ~w6020;
assign w6022 = pi823 & ~w6021;
assign w6023 = ~pi823 & w6021;
assign w6024 = w2568 & ~w6022;
assign w6025 = ~w6023 & w6024;
assign w6026 = ~pi358 & ~w3367;
assign w6027 = pi220 & ~w6021;
assign w6028 = ~pi220 & w6021;
assign w6029 = ~w6027 & ~w6028;
assign w6030 = w3367 & ~w6029;
assign w6031 = ~w2568 & ~w6026;
assign w6032 = ~w6030 & w6031;
assign w6033 = ~w6025 & ~w6032;
assign w6034 = pi039 & w469;
assign w6035 = pi585 & w3345;
assign w6036 = pi743 & w3348;
assign w6037 = ~w6034 & ~w6035;
assign w6038 = ~w6036 & w6037;
assign w6039 = pi562 & ~w6038;
assign w6040 = ~pi039 & ~w3355;
assign w6041 = ~w1546 & ~w5872;
assign w6042 = ~w3334 & ~w6038;
assign w6043 = w3355 & ~w6041;
assign w6044 = ~w6042 & w6043;
assign w6045 = ~pi585 & w3358;
assign w6046 = ~pi562 & ~w6040;
assign w6047 = ~w6044 & w6046;
assign w6048 = ~w6045 & w6047;
assign w6049 = ~w6039 & ~w6048;
assign w6050 = pi871 & ~w6049;
assign w6051 = ~pi871 & w6049;
assign w6052 = w2568 & ~w6050;
assign w6053 = ~w6051 & w6052;
assign w6054 = ~pi359 & ~w3367;
assign w6055 = pi252 & ~w6049;
assign w6056 = ~pi252 & w6049;
assign w6057 = ~w6055 & ~w6056;
assign w6058 = w3367 & ~w6057;
assign w6059 = ~w2568 & ~w6054;
assign w6060 = ~w6058 & w6059;
assign w6061 = ~w6053 & ~w6060;
assign w6062 = pi533 & w3345;
assign w6063 = pi031 & w469;
assign w6064 = pi696 & w3348;
assign w6065 = ~w6062 & ~w6063;
assign w6066 = ~w6064 & w6065;
assign w6067 = pi562 & ~w6066;
assign w6068 = ~pi031 & ~w3355;
assign w6069 = ~w1554 & ~w5872;
assign w6070 = ~w3334 & ~w6066;
assign w6071 = w3355 & ~w6069;
assign w6072 = ~w6070 & w6071;
assign w6073 = ~pi533 & w3358;
assign w6074 = ~pi562 & ~w6068;
assign w6075 = ~w6072 & w6074;
assign w6076 = ~w6073 & w6075;
assign w6077 = ~w6067 & ~w6076;
assign w6078 = pi824 & ~w6077;
assign w6079 = ~pi824 & w6077;
assign w6080 = w2568 & ~w6078;
assign w6081 = ~w6079 & w6080;
assign w6082 = ~pi360 & ~w3367;
assign w6083 = pi221 & ~w6077;
assign w6084 = ~pi221 & w6077;
assign w6085 = ~w6083 & ~w6084;
assign w6086 = w3367 & ~w6085;
assign w6087 = ~w2568 & ~w6082;
assign w6088 = ~w6086 & w6087;
assign w6089 = ~w6081 & ~w6088;
assign w6090 = pi577 & w3345;
assign w6091 = pi038 & w469;
assign w6092 = pi744 & w3348;
assign w6093 = ~w6090 & ~w6091;
assign w6094 = ~w6092 & w6093;
assign w6095 = pi562 & ~w6094;
assign w6096 = ~pi038 & ~w3355;
assign w6097 = ~w1533 & ~w5872;
assign w6098 = ~w3334 & ~w6094;
assign w6099 = w3355 & ~w6097;
assign w6100 = ~w6098 & w6099;
assign w6101 = ~pi577 & w3358;
assign w6102 = ~pi562 & ~w6096;
assign w6103 = ~w6100 & w6102;
assign w6104 = ~w6101 & w6103;
assign w6105 = ~w6095 & ~w6104;
assign w6106 = pi872 & ~w6105;
assign w6107 = ~pi872 & w6105;
assign w6108 = w2568 & ~w6106;
assign w6109 = ~w6107 & w6108;
assign w6110 = ~pi361 & ~w3367;
assign w6111 = pi294 & ~w6105;
assign w6112 = ~pi294 & w6105;
assign w6113 = ~w6111 & ~w6112;
assign w6114 = w3367 & ~w6113;
assign w6115 = ~w2568 & ~w6110;
assign w6116 = ~w6114 & w6115;
assign w6117 = ~w6109 & ~w6116;
assign w6118 = pi026 & w469;
assign w6119 = pi570 & w3345;
assign w6120 = pi776 & w3348;
assign w6121 = ~w6118 & ~w6119;
assign w6122 = ~w6120 & w6121;
assign w6123 = pi562 & ~w6122;
assign w6124 = ~pi026 & ~w3355;
assign w6125 = pi026 & ~w3356;
assign w6126 = ~w3340 & w6122;
assign w6127 = ~w3334 & ~w6126;
assign w6128 = ~w6125 & ~w6127;
assign w6129 = ~pi570 & w3358;
assign w6130 = ~pi562 & ~w6124;
assign w6131 = ~w6129 & w6130;
assign w6132 = ~w6128 & w6131;
assign w6133 = ~w6123 & ~w6132;
assign w6134 = pi904 & ~w6133;
assign w6135 = ~pi904 & w6133;
assign w6136 = w2568 & ~w6134;
assign w6137 = ~w6135 & w6136;
assign w6138 = ~pi362 & ~w3367;
assign w6139 = pi417 & ~w6133;
assign w6140 = ~pi417 & w6133;
assign w6141 = ~w6139 & ~w6140;
assign w6142 = w3367 & ~w6141;
assign w6143 = ~w2568 & ~w6138;
assign w6144 = ~w6142 & w6143;
assign w6145 = ~w6137 & ~w6144;
assign w6146 = pi091 & w469;
assign w6147 = pi547 & w3345;
assign w6148 = pi697 & w3348;
assign w6149 = ~w6146 & ~w6147;
assign w6150 = ~w6148 & w6149;
assign w6151 = pi562 & ~w6150;
assign w6152 = ~pi091 & ~w3355;
assign w6153 = ~w1981 & ~w5872;
assign w6154 = ~w3334 & ~w6150;
assign w6155 = w3355 & ~w6153;
assign w6156 = ~w6154 & w6155;
assign w6157 = ~pi547 & w3358;
assign w6158 = ~pi562 & ~w6152;
assign w6159 = ~w6156 & w6158;
assign w6160 = ~w6157 & w6159;
assign w6161 = ~w6151 & ~w6160;
assign w6162 = pi825 & ~w6161;
assign w6163 = ~pi825 & w6161;
assign w6164 = w2568 & ~w6162;
assign w6165 = ~w6163 & w6164;
assign w6166 = ~pi363 & ~w3367;
assign w6167 = pi212 & ~w6161;
assign w6168 = ~pi212 & w6161;
assign w6169 = ~w6167 & ~w6168;
assign w6170 = w3367 & ~w6169;
assign w6171 = ~w2568 & ~w6166;
assign w6172 = ~w6170 & w6171;
assign w6173 = ~w6165 & ~w6172;
assign w6174 = pi621 & w3345;
assign w6175 = pi086 & w469;
assign w6176 = pi789 & w3348;
assign w6177 = ~w6174 & ~w6175;
assign w6178 = ~w6176 & w6177;
assign w6179 = pi562 & ~w6178;
assign w6180 = ~pi086 & ~w3355;
assign w6181 = ~w2126 & ~w5872;
assign w6182 = ~w3334 & ~w6178;
assign w6183 = w3355 & ~w6181;
assign w6184 = ~w6182 & w6183;
assign w6185 = ~pi621 & w3358;
assign w6186 = ~pi562 & ~w6180;
assign w6187 = ~w6184 & w6186;
assign w6188 = ~w6185 & w6187;
assign w6189 = ~w6179 & ~w6188;
assign w6190 = pi917 & ~w6189;
assign w6191 = ~pi917 & w6189;
assign w6192 = w2568 & ~w6190;
assign w6193 = ~w6191 & w6192;
assign w6194 = ~pi364 & ~w3367;
assign w6195 = pi431 & ~w6189;
assign w6196 = ~pi431 & w6189;
assign w6197 = ~w6195 & ~w6196;
assign w6198 = w3367 & ~w6197;
assign w6199 = ~w2568 & ~w6194;
assign w6200 = ~w6198 & w6199;
assign w6201 = ~w6193 & ~w6200;
assign w6202 = pi087 & w469;
assign w6203 = pi597 & w3345;
assign w6204 = pi790 & w3348;
assign w6205 = ~w6202 & ~w6203;
assign w6206 = ~w6204 & w6205;
assign w6207 = pi562 & ~w6206;
assign w6208 = ~pi087 & ~w3355;
assign w6209 = ~w2116 & ~w5872;
assign w6210 = ~w3334 & ~w6206;
assign w6211 = w3355 & ~w6209;
assign w6212 = ~w6210 & w6211;
assign w6213 = ~pi597 & w3358;
assign w6214 = ~pi562 & ~w6208;
assign w6215 = ~w6212 & w6214;
assign w6216 = ~w6213 & w6215;
assign w6217 = ~w6207 & ~w6216;
assign w6218 = pi918 & ~w6217;
assign w6219 = ~pi918 & w6217;
assign w6220 = w2568 & ~w6218;
assign w6221 = ~w6219 & w6220;
assign w6222 = ~pi365 & ~w3367;
assign w6223 = pi432 & ~w6217;
assign w6224 = ~pi432 & w6217;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = w3367 & ~w6225;
assign w6227 = ~w2568 & ~w6222;
assign w6228 = ~w6226 & w6227;
assign w6229 = ~w6221 & ~w6228;
assign w6230 = pi066 & w469;
assign w6231 = pi623 & w3345;
assign w6232 = pi754 & w3348;
assign w6233 = ~w6230 & ~w6231;
assign w6234 = ~w6232 & w6233;
assign w6235 = pi562 & ~w6234;
assign w6236 = ~pi066 & ~w3355;
assign w6237 = ~w1842 & ~w5872;
assign w6238 = ~w3334 & ~w6234;
assign w6239 = w3355 & ~w6237;
assign w6240 = ~w6238 & w6239;
assign w6241 = ~pi623 & w3358;
assign w6242 = ~pi562 & ~w6236;
assign w6243 = ~w6240 & w6242;
assign w6244 = ~w6241 & w6243;
assign w6245 = ~w6235 & ~w6244;
assign w6246 = pi882 & ~w6245;
assign w6247 = ~pi882 & w6245;
assign w6248 = w2568 & ~w6246;
assign w6249 = ~w6247 & w6248;
assign w6250 = ~pi366 & ~w3367;
assign w6251 = pi334 & ~w6245;
assign w6252 = ~pi334 & w6245;
assign w6253 = ~w6251 & ~w6252;
assign w6254 = w3367 & ~w6253;
assign w6255 = ~w2568 & ~w6250;
assign w6256 = ~w6254 & w6255;
assign w6257 = ~w6249 & ~w6256;
assign w6258 = pi179 & w469;
assign w6259 = pi635 & w3345;
assign w6260 = pi755 & w3348;
assign w6261 = ~w6258 & ~w6259;
assign w6262 = ~w6260 & w6261;
assign w6263 = pi562 & ~w6262;
assign w6264 = ~pi179 & ~w3355;
assign w6265 = ~w2486 & ~w5872;
assign w6266 = ~w3334 & ~w6262;
assign w6267 = w3355 & ~w6265;
assign w6268 = ~w6266 & w6267;
assign w6269 = ~pi635 & w3358;
assign w6270 = ~pi562 & ~w6264;
assign w6271 = ~w6268 & w6270;
assign w6272 = ~w6269 & w6271;
assign w6273 = ~w6263 & ~w6272;
assign w6274 = pi883 & ~w6273;
assign w6275 = ~pi883 & w6273;
assign w6276 = w2568 & ~w6274;
assign w6277 = ~w6275 & w6276;
assign w6278 = ~pi367 & ~w3367;
assign w6279 = pi298 & ~w6273;
assign w6280 = ~pi298 & w6273;
assign w6281 = ~w6279 & ~w6280;
assign w6282 = w3367 & ~w6281;
assign w6283 = ~w2568 & ~w6278;
assign w6284 = ~w6282 & w6283;
assign w6285 = ~w6277 & ~w6284;
assign w6286 = pi625 & w3345;
assign w6287 = pi104 & w469;
assign w6288 = pi757 & w3348;
assign w6289 = ~w6286 & ~w6287;
assign w6290 = ~w6288 & w6289;
assign w6291 = pi562 & ~w6290;
assign w6292 = ~pi104 & ~w3355;
assign w6293 = ~w2035 & ~w5872;
assign w6294 = ~w3334 & ~w6290;
assign w6295 = w3355 & ~w6293;
assign w6296 = ~w6294 & w6295;
assign w6297 = ~pi625 & w3358;
assign w6298 = ~pi562 & ~w6292;
assign w6299 = ~w6296 & w6298;
assign w6300 = ~w6297 & w6299;
assign w6301 = ~w6291 & ~w6300;
assign w6302 = pi885 & ~w6301;
assign w6303 = ~pi885 & w6301;
assign w6304 = w2568 & ~w6302;
assign w6305 = ~w6303 & w6304;
assign w6306 = ~pi368 & ~w3367;
assign w6307 = pi335 & ~w6301;
assign w6308 = ~pi335 & w6301;
assign w6309 = ~w6307 & ~w6308;
assign w6310 = w3367 & ~w6309;
assign w6311 = ~w2568 & ~w6306;
assign w6312 = ~w6310 & w6311;
assign w6313 = ~w6305 & ~w6312;
assign w6314 = pi578 & w3345;
assign w6315 = pi040 & w469;
assign w6316 = pi759 & w3348;
assign w6317 = ~w6314 & ~w6315;
assign w6318 = ~w6316 & w6317;
assign w6319 = pi562 & ~w6318;
assign w6320 = ~pi040 & ~w3355;
assign w6321 = ~w1623 & ~w5872;
assign w6322 = ~w3334 & ~w6318;
assign w6323 = w3355 & ~w6321;
assign w6324 = ~w6322 & w6323;
assign w6325 = ~pi578 & w3358;
assign w6326 = ~pi562 & ~w6320;
assign w6327 = ~w6324 & w6326;
assign w6328 = ~w6325 & w6327;
assign w6329 = ~w6319 & ~w6328;
assign w6330 = pi887 & ~w6329;
assign w6331 = ~pi887 & w6329;
assign w6332 = w2568 & ~w6330;
assign w6333 = ~w6331 & w6332;
assign w6334 = ~pi369 & ~w3367;
assign w6335 = pi337 & ~w6329;
assign w6336 = ~pi337 & w6329;
assign w6337 = ~w6335 & ~w6336;
assign w6338 = w3367 & ~w6337;
assign w6339 = ~w2568 & ~w6334;
assign w6340 = ~w6338 & w6339;
assign w6341 = ~w6333 & ~w6340;
assign w6342 = pi598 & w3345;
assign w6343 = pi041 & w469;
assign w6344 = pi760 & w3348;
assign w6345 = ~w6342 & ~w6343;
assign w6346 = ~w6344 & w6345;
assign w6347 = pi562 & ~w6346;
assign w6348 = ~pi041 & ~w3355;
assign w6349 = ~w1634 & ~w5872;
assign w6350 = ~w3334 & ~w6346;
assign w6351 = w3355 & ~w6349;
assign w6352 = ~w6350 & w6351;
assign w6353 = ~pi598 & w3358;
assign w6354 = ~pi562 & ~w6348;
assign w6355 = ~w6352 & w6354;
assign w6356 = ~w6353 & w6355;
assign w6357 = ~w6347 & ~w6356;
assign w6358 = pi888 & ~w6357;
assign w6359 = ~pi888 & w6357;
assign w6360 = w2568 & ~w6358;
assign w6361 = ~w6359 & w6360;
assign w6362 = ~pi370 & ~w3367;
assign w6363 = pi339 & ~w6357;
assign w6364 = ~pi339 & w6357;
assign w6365 = ~w6363 & ~w6364;
assign w6366 = w3367 & ~w6365;
assign w6367 = ~w2568 & ~w6362;
assign w6368 = ~w6366 & w6367;
assign w6369 = ~w6361 & ~w6368;
assign w6370 = pi610 & w3345;
assign w6371 = pi103 & w469;
assign w6372 = pi758 & w3348;
assign w6373 = ~w6370 & ~w6371;
assign w6374 = ~w6372 & w6373;
assign w6375 = pi562 & ~w6374;
assign w6376 = ~pi103 & ~w3355;
assign w6377 = ~w2045 & ~w5872;
assign w6378 = ~w3334 & ~w6374;
assign w6379 = w3355 & ~w6377;
assign w6380 = ~w6378 & w6379;
assign w6381 = ~pi610 & w3358;
assign w6382 = ~pi562 & ~w6376;
assign w6383 = ~w6380 & w6382;
assign w6384 = ~w6381 & w6383;
assign w6385 = ~w6375 & ~w6384;
assign w6386 = pi886 & ~w6385;
assign w6387 = ~pi886 & w6385;
assign w6388 = w2568 & ~w6386;
assign w6389 = ~w6387 & w6388;
assign w6390 = ~pi371 & ~w3367;
assign w6391 = pi336 & ~w6385;
assign w6392 = ~pi336 & w6385;
assign w6393 = ~w6391 & ~w6392;
assign w6394 = w3367 & ~w6393;
assign w6395 = ~w2568 & ~w6390;
assign w6396 = ~w6394 & w6395;
assign w6397 = ~w6389 & ~w6396;
assign w6398 = pi632 & w3345;
assign w6399 = pi105 & w469;
assign w6400 = pi761 & w3348;
assign w6401 = ~w6398 & ~w6399;
assign w6402 = ~w6400 & w6401;
assign w6403 = pi562 & ~w6402;
assign w6404 = ~pi105 & ~w3355;
assign w6405 = ~w2055 & ~w5872;
assign w6406 = ~w3334 & ~w6402;
assign w6407 = w3355 & ~w6405;
assign w6408 = ~w6406 & w6407;
assign w6409 = ~pi632 & w3358;
assign w6410 = ~pi562 & ~w6404;
assign w6411 = ~w6408 & w6410;
assign w6412 = ~w6409 & w6411;
assign w6413 = ~w6403 & ~w6412;
assign w6414 = pi889 & ~w6413;
assign w6415 = ~pi889 & w6413;
assign w6416 = w2568 & ~w6414;
assign w6417 = ~w6415 & w6416;
assign w6418 = ~pi372 & ~w3367;
assign w6419 = pi296 & ~w6413;
assign w6420 = ~pi296 & w6413;
assign w6421 = ~w6419 & ~w6420;
assign w6422 = w3367 & ~w6421;
assign w6423 = ~w2568 & ~w6418;
assign w6424 = ~w6422 & w6423;
assign w6425 = ~w6417 & ~w6424;
assign w6426 = pi109 & w469;
assign w6427 = pi599 & w3345;
assign w6428 = pi762 & w3348;
assign w6429 = ~w6426 & ~w6427;
assign w6430 = ~w6428 & w6429;
assign w6431 = w3344 & ~w6430;
assign w6432 = pi109 & ~w3356;
assign w6433 = pi599 & w3358;
assign w6434 = ~w6432 & ~w6433;
assign w6435 = ~pi562 & ~w6434;
assign w6436 = ~w6431 & ~w6435;
assign w6437 = pi890 & ~w6436;
assign w6438 = ~pi890 & w6436;
assign w6439 = w2568 & ~w6437;
assign w6440 = ~w6438 & w6439;
assign w6441 = ~pi373 & ~w3367;
assign w6442 = pi248 & ~w6436;
assign w6443 = ~pi248 & w6436;
assign w6444 = ~w6442 & ~w6443;
assign w6445 = w3367 & ~w6444;
assign w6446 = ~w2568 & ~w6441;
assign w6447 = ~w6445 & w6446;
assign w6448 = ~w6440 & ~w6447;
assign w6449 = pi092 & w469;
assign w6450 = pi643 & w3345;
assign w6451 = pi706 & w3348;
assign w6452 = ~w6449 & ~w6450;
assign w6453 = ~w6451 & w6452;
assign w6454 = pi562 & ~w6453;
assign w6455 = ~pi092 & ~w3355;
assign w6456 = ~w1813 & ~w5872;
assign w6457 = ~w3334 & ~w6453;
assign w6458 = w3355 & ~w6456;
assign w6459 = ~w6457 & w6458;
assign w6460 = ~pi643 & w3358;
assign w6461 = ~pi562 & ~w6455;
assign w6462 = ~w6459 & w6461;
assign w6463 = ~w6460 & w6462;
assign w6464 = ~w6454 & ~w6463;
assign w6465 = pi834 & ~w6464;
assign w6466 = ~pi834 & w6464;
assign w6467 = w2568 & ~w6465;
assign w6468 = ~w6466 & w6467;
assign w6469 = ~pi374 & ~w3367;
assign w6470 = ~pi229 & ~w6464;
assign w6471 = pi229 & w6464;
assign w6472 = ~w6470 & ~w6471;
assign w6473 = w3367 & ~w6472;
assign w6474 = ~w2568 & ~w6469;
assign w6475 = ~w6473 & w6474;
assign w6476 = ~w6468 & ~w6475;
assign w6477 = pi088 & w469;
assign w6478 = pi614 & w3345;
assign w6479 = pi793 & w3348;
assign w6480 = ~w6477 & ~w6478;
assign w6481 = ~w6479 & w6480;
assign w6482 = pi562 & ~w6481;
assign w6483 = ~pi088 & ~w3355;
assign w6484 = ~w2136 & ~w5872;
assign w6485 = ~w3334 & ~w6481;
assign w6486 = w3355 & ~w6484;
assign w6487 = ~w6485 & w6486;
assign w6488 = ~pi614 & w3358;
assign w6489 = ~pi562 & ~w6483;
assign w6490 = ~w6487 & w6489;
assign w6491 = ~w6488 & w6490;
assign w6492 = ~w6482 & ~w6491;
assign w6493 = pi921 & ~w6492;
assign w6494 = ~pi921 & w6492;
assign w6495 = w2568 & ~w6493;
assign w6496 = ~w6494 & w6495;
assign w6497 = ~pi375 & ~w3367;
assign w6498 = pi419 & ~w6492;
assign w6499 = ~pi419 & w6492;
assign w6500 = ~w6498 & ~w6499;
assign w6501 = w3367 & ~w6500;
assign w6502 = ~w2568 & ~w6497;
assign w6503 = ~w6501 & w6502;
assign w6504 = ~w6496 & ~w6503;
assign w6505 = ~pi067 & w469;
assign w6506 = ~pi620 & w3345;
assign w6507 = ~pi770 & w3348;
assign w6508 = ~w6505 & ~w6506;
assign w6509 = ~w6507 & w6508;
assign w6510 = pi562 & w6509;
assign w6511 = ~pi067 & ~w3355;
assign w6512 = ~w1786 & ~w5872;
assign w6513 = ~w3334 & w6509;
assign w6514 = w3355 & ~w6512;
assign w6515 = ~w6513 & w6514;
assign w6516 = ~pi620 & w3358;
assign w6517 = ~pi562 & ~w6511;
assign w6518 = ~w6515 & w6517;
assign w6519 = ~w6516 & w6518;
assign w6520 = ~w6510 & ~w6519;
assign w6521 = pi898 & ~w6520;
assign w6522 = ~pi898 & w6520;
assign w6523 = w2568 & ~w6521;
assign w6524 = ~w6522 & w6523;
assign w6525 = ~pi376 & ~w3367;
assign w6526 = pi413 & ~w6520;
assign w6527 = ~pi413 & w6520;
assign w6528 = ~w6526 & ~w6527;
assign w6529 = w3367 & ~w6528;
assign w6530 = ~w2568 & ~w6525;
assign w6531 = ~w6529 & w6530;
assign w6532 = ~w6524 & ~w6531;
assign w6533 = ~pi175 & ~w3355;
assign w6534 = ~w468 & w2446;
assign w6535 = ~pi771 & w3348;
assign w6536 = ~pi606 & w3345;
assign w6537 = ~w6534 & ~w6536;
assign w6538 = ~w6535 & w6537;
assign w6539 = ~w3334 & w6538;
assign w6540 = ~w2446 & ~w5872;
assign w6541 = ~w6539 & ~w6540;
assign w6542 = ~pi606 & w3340;
assign w6543 = ~w6541 & ~w6542;
assign w6544 = w3355 & ~w6543;
assign w6545 = ~w6533 & ~w6544;
assign w6546 = ~pi562 & ~w6545;
assign w6547 = pi562 & ~w6538;
assign w6548 = ~w6546 & ~w6547;
assign w6549 = ~pi899 & ~w6548;
assign w6550 = pi899 & w6548;
assign w6551 = w2568 & ~w6549;
assign w6552 = ~w6550 & w6551;
assign w6553 = ~pi377 & ~w3367;
assign w6554 = ~pi409 & ~w6548;
assign w6555 = pi409 & w6548;
assign w6556 = ~w6554 & ~w6555;
assign w6557 = w3367 & ~w6556;
assign w6558 = ~w2568 & ~w6553;
assign w6559 = ~w6557 & w6558;
assign w6560 = ~w6552 & ~w6559;
assign w6561 = pi616 & w3345;
assign w6562 = pi097 & w469;
assign w6563 = pi710 & w3348;
assign w6564 = ~w6561 & ~w6562;
assign w6565 = ~w6563 & w6564;
assign w6566 = pi562 & ~w6565;
assign w6567 = ~pi097 & ~w3355;
assign w6568 = ~w2074 & ~w5872;
assign w6569 = ~w3334 & ~w6565;
assign w6570 = w3355 & ~w6568;
assign w6571 = ~w6569 & w6570;
assign w6572 = ~pi616 & w3358;
assign w6573 = ~pi562 & ~w6567;
assign w6574 = ~w6571 & w6573;
assign w6575 = ~w6572 & w6574;
assign w6576 = ~w6566 & ~w6575;
assign w6577 = pi838 & ~w6576;
assign w6578 = ~pi838 & w6576;
assign w6579 = w2568 & ~w6577;
assign w6580 = ~w6578 & w6579;
assign w6581 = ~pi378 & ~w3367;
assign w6582 = ~pi233 & ~w6576;
assign w6583 = pi233 & w6576;
assign w6584 = ~w6582 & ~w6583;
assign w6585 = w3367 & ~w6584;
assign w6586 = ~w2568 & ~w6581;
assign w6587 = ~w6585 & w6586;
assign w6588 = ~w6580 & ~w6587;
assign w6589 = pi118 & w469;
assign w6590 = pi581 & w3345;
assign w6591 = pi773 & w3348;
assign w6592 = ~w6589 & ~w6590;
assign w6593 = ~w6591 & w6592;
assign w6594 = pi562 & ~w6593;
assign w6595 = ~pi118 & ~w3355;
assign w6596 = pi118 & ~w3356;
assign w6597 = ~w3340 & w6593;
assign w6598 = ~w3334 & ~w6597;
assign w6599 = ~w6596 & ~w6598;
assign w6600 = ~pi581 & w3358;
assign w6601 = ~pi562 & ~w6595;
assign w6602 = ~w6600 & w6601;
assign w6603 = ~w6599 & w6602;
assign w6604 = ~w6594 & ~w6603;
assign w6605 = pi901 & ~w6604;
assign w6606 = ~pi901 & w6604;
assign w6607 = w2568 & ~w6605;
assign w6608 = ~w6606 & w6607;
assign w6609 = ~pi379 & ~w3367;
assign w6610 = pi437 & ~w6604;
assign w6611 = ~pi437 & w6604;
assign w6612 = ~w6610 & ~w6611;
assign w6613 = w3367 & ~w6612;
assign w6614 = ~w2568 & ~w6609;
assign w6615 = ~w6613 & w6614;
assign w6616 = ~w6608 & ~w6615;
assign w6617 = pi609 & w3345;
assign w6618 = pi032 & w469;
assign w6619 = pi711 & w3348;
assign w6620 = ~w6617 & ~w6618;
assign w6621 = ~w6619 & w6620;
assign w6622 = pi562 & ~w6621;
assign w6623 = ~pi032 & ~w3355;
assign w6624 = ~w1668 & ~w5872;
assign w6625 = ~w3334 & ~w6621;
assign w6626 = w3355 & ~w6624;
assign w6627 = ~w6625 & w6626;
assign w6628 = ~pi609 & w3358;
assign w6629 = ~pi562 & ~w6623;
assign w6630 = ~w6627 & w6629;
assign w6631 = ~w6628 & w6630;
assign w6632 = ~w6622 & ~w6631;
assign w6633 = pi839 & ~w6632;
assign w6634 = ~pi839 & w6632;
assign w6635 = w2568 & ~w6633;
assign w6636 = ~w6634 & w6635;
assign w6637 = ~pi380 & ~w3367;
assign w6638 = ~pi237 & ~w6632;
assign w6639 = pi237 & w6632;
assign w6640 = ~w6638 & ~w6639;
assign w6641 = w3367 & ~w6640;
assign w6642 = ~w2568 & ~w6637;
assign w6643 = ~w6641 & w6642;
assign w6644 = ~w6636 & ~w6643;
assign w6645 = pi658 & w3345;
assign w6646 = pi033 & w469;
assign w6647 = pi712 & w3348;
assign w6648 = ~w6645 & ~w6646;
assign w6649 = ~w6647 & w6648;
assign w6650 = pi562 & ~w6649;
assign w6651 = ~pi033 & ~w3355;
assign w6652 = ~w1656 & ~w5872;
assign w6653 = ~w3334 & ~w6649;
assign w6654 = w3355 & ~w6652;
assign w6655 = ~w6653 & w6654;
assign w6656 = ~pi658 & w3358;
assign w6657 = ~pi562 & ~w6651;
assign w6658 = ~w6655 & w6657;
assign w6659 = ~w6656 & w6658;
assign w6660 = ~w6650 & ~w6659;
assign w6661 = pi840 & ~w6660;
assign w6662 = ~pi840 & w6660;
assign w6663 = w2568 & ~w6661;
assign w6664 = ~w6662 & w6663;
assign w6665 = ~pi381 & ~w3367;
assign w6666 = ~pi234 & ~w6660;
assign w6667 = pi234 & w6660;
assign w6668 = ~w6666 & ~w6667;
assign w6669 = w3367 & ~w6668;
assign w6670 = ~w2568 & ~w6665;
assign w6671 = ~w6669 & w6670;
assign w6672 = ~w6664 & ~w6671;
assign w6673 = pi116 & w469;
assign w6674 = pi617 & w3345;
assign w6675 = pi713 & w3348;
assign w6676 = ~w6673 & ~w6674;
assign w6677 = ~w6675 & w6676;
assign w6678 = pi562 & ~w6677;
assign w6679 = ~pi116 & ~w3355;
assign w6680 = ~w2106 & ~w5872;
assign w6681 = ~w3334 & ~w6677;
assign w6682 = w3355 & ~w6680;
assign w6683 = ~w6681 & w6682;
assign w6684 = ~pi617 & w3358;
assign w6685 = ~pi562 & ~w6679;
assign w6686 = ~w6683 & w6685;
assign w6687 = ~w6684 & w6686;
assign w6688 = ~w6678 & ~w6687;
assign w6689 = pi841 & ~w6688;
assign w6690 = ~pi841 & w6688;
assign w6691 = w2568 & ~w6689;
assign w6692 = ~w6690 & w6691;
assign w6693 = ~pi382 & ~w3367;
assign w6694 = ~pi235 & ~w6688;
assign w6695 = pi235 & w6688;
assign w6696 = ~w6694 & ~w6695;
assign w6697 = w3367 & ~w6696;
assign w6698 = ~w2568 & ~w6693;
assign w6699 = ~w6697 & w6698;
assign w6700 = ~w6692 & ~w6699;
assign w6701 = pi180 & w469;
assign w6702 = pi596 & w3345;
assign w6703 = pi723 & w3348;
assign w6704 = ~w6701 & ~w6702;
assign w6705 = ~w6703 & w6704;
assign w6706 = pi562 & ~w6705;
assign w6707 = ~pi180 & ~w3355;
assign w6708 = ~w2437 & ~w5872;
assign w6709 = ~w3334 & ~w6705;
assign w6710 = w3355 & ~w6708;
assign w6711 = ~w6709 & w6710;
assign w6712 = ~pi596 & w3358;
assign w6713 = ~pi562 & ~w6707;
assign w6714 = ~w6711 & w6713;
assign w6715 = ~w6712 & w6714;
assign w6716 = ~w6706 & ~w6715;
assign w6717 = pi851 & ~w6716;
assign w6718 = ~pi851 & w6716;
assign w6719 = w2568 & ~w6717;
assign w6720 = ~w6718 & w6719;
assign w6721 = ~pi383 & ~w3367;
assign w6722 = ~pi240 & ~w6716;
assign w6723 = pi240 & w6716;
assign w6724 = ~w6722 & ~w6723;
assign w6725 = w3367 & ~w6724;
assign w6726 = ~w2568 & ~w6721;
assign w6727 = ~w6725 & w6726;
assign w6728 = ~w6720 & ~w6727;
assign w6729 = pi095 & w469;
assign w6730 = pi630 & w3345;
assign w6731 = pi726 & w3348;
assign w6732 = ~w6729 & ~w6730;
assign w6733 = ~w6731 & w6732;
assign w6734 = pi562 & ~w6733;
assign w6735 = ~pi095 & ~w3355;
assign w6736 = ~w1991 & ~w5872;
assign w6737 = ~w3334 & ~w6733;
assign w6738 = w3355 & ~w6736;
assign w6739 = ~w6737 & w6738;
assign w6740 = ~pi630 & w3358;
assign w6741 = ~pi562 & ~w6735;
assign w6742 = ~w6739 & w6741;
assign w6743 = ~w6740 & w6742;
assign w6744 = ~w6734 & ~w6743;
assign w6745 = pi854 & ~w6744;
assign w6746 = ~pi854 & w6744;
assign w6747 = w2568 & ~w6745;
assign w6748 = ~w6746 & w6747;
assign w6749 = ~pi384 & ~w3367;
assign w6750 = ~pi243 & ~w6744;
assign w6751 = pi243 & w6744;
assign w6752 = ~w6750 & ~w6751;
assign w6753 = w3367 & ~w6752;
assign w6754 = ~w2568 & ~w6749;
assign w6755 = ~w6753 & w6754;
assign w6756 = ~w6748 & ~w6755;
assign w6757 = pi618 & w3345;
assign w6758 = pi096 & w469;
assign w6759 = pi729 & w3348;
assign w6760 = ~w6757 & ~w6758;
assign w6761 = ~w6759 & w6760;
assign w6762 = pi562 & ~w6761;
assign w6763 = ~pi096 & ~w3355;
assign w6764 = ~w2011 & ~w5872;
assign w6765 = ~w3334 & ~w6761;
assign w6766 = w3355 & ~w6764;
assign w6767 = ~w6765 & w6766;
assign w6768 = ~pi618 & w3358;
assign w6769 = ~pi562 & ~w6763;
assign w6770 = ~w6767 & w6769;
assign w6771 = ~w6768 & w6770;
assign w6772 = ~w6762 & ~w6771;
assign w6773 = pi857 & ~w6772;
assign w6774 = ~pi857 & w6772;
assign w6775 = w2568 & ~w6773;
assign w6776 = ~w6774 & w6775;
assign w6777 = ~pi385 & ~w3367;
assign w6778 = ~pi236 & ~w6772;
assign w6779 = pi236 & w6772;
assign w6780 = ~w6778 & ~w6779;
assign w6781 = w3367 & ~w6780;
assign w6782 = ~w2568 & ~w6777;
assign w6783 = ~w6781 & w6782;
assign w6784 = ~w6776 & ~w6783;
assign w6785 = pi172 & w469;
assign w6786 = pi518 & w3345;
assign w6787 = pi691 & w3348;
assign w6788 = ~w6785 & ~w6786;
assign w6789 = ~w6787 & w6788;
assign w6790 = pi562 & ~w6789;
assign w6791 = ~pi172 & ~w3355;
assign w6792 = ~w2496 & ~w5872;
assign w6793 = ~w3334 & ~w6789;
assign w6794 = w3355 & ~w6792;
assign w6795 = ~w6793 & w6794;
assign w6796 = ~pi518 & w3358;
assign w6797 = ~pi562 & ~w6791;
assign w6798 = ~w6795 & w6797;
assign w6799 = ~w6796 & w6798;
assign w6800 = ~w6790 & ~w6799;
assign w6801 = pi819 & ~w6800;
assign w6802 = ~pi819 & w6800;
assign w6803 = w2568 & ~w6801;
assign w6804 = ~w6802 & w6803;
assign w6805 = ~pi386 & ~w3367;
assign w6806 = pi216 & ~w6800;
assign w6807 = ~pi216 & w6800;
assign w6808 = ~w6806 & ~w6807;
assign w6809 = w3367 & ~w6808;
assign w6810 = ~w2568 & ~w6805;
assign w6811 = ~w6809 & w6810;
assign w6812 = ~w6804 & ~w6811;
assign w6813 = w1 & ~w2709;
assign w6814 = pi387 & ~w1;
assign w6815 = ~w6813 & ~w6814;
assign w6816 = w1 & w2766;
assign w6817 = pi388 & ~w1;
assign w6818 = ~w6816 & ~w6817;
assign w6819 = w1 & ~w2736;
assign w6820 = pi389 & ~w1;
assign w6821 = ~w6819 & ~w6820;
assign w6822 = ~w2572 & ~w2574;
assign w6823 = pi028 & w469;
assign w6824 = pi629 & w3345;
assign w6825 = pi792 & w3348;
assign w6826 = ~w6823 & ~w6824;
assign w6827 = ~w6825 & w6826;
assign w6828 = pi562 & ~w6827;
assign w6829 = ~pi028 & ~w3355;
assign w6830 = ~w1690 & ~w5872;
assign w6831 = ~w3334 & ~w6827;
assign w6832 = w3355 & ~w6830;
assign w6833 = ~w6831 & w6832;
assign w6834 = ~pi629 & w3358;
assign w6835 = ~pi562 & ~w6829;
assign w6836 = ~w6833 & w6835;
assign w6837 = ~w6834 & w6836;
assign w6838 = ~w6828 & ~w6837;
assign w6839 = pi920 & ~w6838;
assign w6840 = ~pi920 & w6838;
assign w6841 = w2568 & ~w6839;
assign w6842 = ~w6840 & w6841;
assign w6843 = ~pi391 & ~w3367;
assign w6844 = pi434 & ~w6838;
assign w6845 = ~pi434 & w6838;
assign w6846 = ~w6844 & ~w6845;
assign w6847 = w3367 & ~w6846;
assign w6848 = ~w2568 & ~w6843;
assign w6849 = ~w6847 & w6848;
assign w6850 = ~w6842 & ~w6849;
assign w6851 = ~pi184 & w469;
assign w6852 = pi600 & w3345;
assign w6853 = pi763 & w3348;
assign w6854 = ~w6851 & ~w6852;
assign w6855 = ~w6853 & w6854;
assign w6856 = w3344 & ~w6855;
assign w6857 = ~pi184 & ~w3356;
assign w6858 = pi600 & w3358;
assign w6859 = ~w6857 & ~w6858;
assign w6860 = ~pi562 & ~w6859;
assign w6861 = ~w6856 & ~w6860;
assign w6862 = pi891 & ~w6861;
assign w6863 = ~pi891 & w6861;
assign w6864 = w2568 & ~w6862;
assign w6865 = ~w6863 & w6864;
assign w6866 = ~pi392 & ~w3367;
assign w6867 = pi251 & ~w6861;
assign w6868 = ~pi251 & w6861;
assign w6869 = ~w6867 & ~w6868;
assign w6870 = w3367 & ~w6869;
assign w6871 = ~w2568 & ~w6866;
assign w6872 = ~w6870 & w6871;
assign w6873 = ~w6865 & ~w6872;
assign w6874 = pi029 & w469;
assign w6875 = pi655 & w3345;
assign w6876 = pi791 & w3348;
assign w6877 = ~w6874 & ~w6875;
assign w6878 = ~w6876 & w6877;
assign w6879 = pi562 & ~w6878;
assign w6880 = ~pi029 & ~w3355;
assign w6881 = ~w1678 & ~w5872;
assign w6882 = ~w3334 & ~w6878;
assign w6883 = w3355 & ~w6881;
assign w6884 = ~w6882 & w6883;
assign w6885 = ~pi655 & w3358;
assign w6886 = ~pi562 & ~w6880;
assign w6887 = ~w6884 & w6886;
assign w6888 = ~w6885 & w6887;
assign w6889 = ~w6879 & ~w6888;
assign w6890 = pi919 & ~w6889;
assign w6891 = ~pi919 & w6889;
assign w6892 = w2568 & ~w6890;
assign w6893 = ~w6891 & w6892;
assign w6894 = ~pi393 & ~w3367;
assign w6895 = pi436 & ~w6889;
assign w6896 = ~pi436 & w6889;
assign w6897 = ~w6895 & ~w6896;
assign w6898 = w3367 & ~w6897;
assign w6899 = ~w2568 & ~w6894;
assign w6900 = ~w6898 & w6899;
assign w6901 = ~w6893 & ~w6900;
assign w6902 = w1 & ~w2681;
assign w6903 = pi394 & ~w1;
assign w6904 = ~w6902 & ~w6903;
assign w6905 = pi151 & w469;
assign w6906 = pi580 & w3345;
assign w6907 = pi756 & w3348;
assign w6908 = ~w6905 & ~w6906;
assign w6909 = ~w6907 & w6908;
assign w6910 = pi562 & ~w6909;
assign w6911 = ~pi151 & ~w3355;
assign w6912 = ~w2330 & ~w5872;
assign w6913 = ~w3334 & ~w6909;
assign w6914 = w3355 & ~w6912;
assign w6915 = ~w6913 & w6914;
assign w6916 = ~pi580 & w3358;
assign w6917 = ~pi562 & ~w6911;
assign w6918 = ~w6915 & w6917;
assign w6919 = ~w6916 & w6918;
assign w6920 = ~w6910 & ~w6919;
assign w6921 = pi884 & ~w6920;
assign w6922 = ~pi884 & w6920;
assign w6923 = w2568 & ~w6921;
assign w6924 = ~w6922 & w6923;
assign w6925 = ~pi395 & ~w3367;
assign w6926 = pi338 & ~w6920;
assign w6927 = ~pi338 & w6920;
assign w6928 = ~w6926 & ~w6927;
assign w6929 = w3367 & ~w6928;
assign w6930 = ~w2568 & ~w6925;
assign w6931 = ~w6929 & w6930;
assign w6932 = ~w6924 & ~w6931;
assign w6933 = w1 & w2791;
assign w6934 = pi396 & ~w1;
assign w6935 = ~w6933 & ~w6934;
assign w6936 = pi143 & w469;
assign w6937 = pi657 & w3345;
assign w6938 = pi788 & w3348;
assign w6939 = ~w6936 & ~w6937;
assign w6940 = ~w6938 & w6939;
assign w6941 = pi562 & ~w6940;
assign w6942 = ~pi143 & ~w3355;
assign w6943 = ~w2350 & ~w5872;
assign w6944 = ~w3334 & ~w6940;
assign w6945 = w3355 & ~w6943;
assign w6946 = ~w6944 & w6945;
assign w6947 = ~pi657 & w3358;
assign w6948 = ~pi562 & ~w6942;
assign w6949 = ~w6946 & w6948;
assign w6950 = ~w6947 & w6949;
assign w6951 = ~w6941 & ~w6950;
assign w6952 = pi916 & ~w6951;
assign w6953 = ~pi916 & w6951;
assign w6954 = w2568 & ~w6952;
assign w6955 = ~w6953 & w6954;
assign w6956 = ~pi397 & ~w3367;
assign w6957 = pi433 & ~w6951;
assign w6958 = ~pi433 & w6951;
assign w6959 = ~w6957 & ~w6958;
assign w6960 = w3367 & ~w6959;
assign w6961 = ~w2568 & ~w6956;
assign w6962 = ~w6960 & w6961;
assign w6963 = ~w6955 & ~w6962;
assign w6964 = pi035 & w469;
assign w6965 = pi640 & w3345;
assign w6966 = pi728 & w3348;
assign w6967 = ~w6964 & ~w6965;
assign w6968 = ~w6966 & w6967;
assign w6969 = pi562 & ~w6968;
assign w6970 = ~pi035 & ~w3355;
assign w6971 = ~w1593 & ~w5872;
assign w6972 = ~w3334 & ~w6968;
assign w6973 = w3355 & ~w6971;
assign w6974 = ~w6972 & w6973;
assign w6975 = ~pi640 & w3358;
assign w6976 = ~pi562 & ~w6970;
assign w6977 = ~w6974 & w6976;
assign w6978 = ~w6975 & w6977;
assign w6979 = ~w6969 & ~w6978;
assign w6980 = pi856 & ~w6979;
assign w6981 = ~pi856 & w6979;
assign w6982 = w2568 & ~w6980;
assign w6983 = ~w6981 & w6982;
assign w6984 = ~pi398 & ~w3367;
assign w6985 = ~pi244 & ~w6979;
assign w6986 = pi244 & w6979;
assign w6987 = ~w6985 & ~w6986;
assign w6988 = w3367 & ~w6987;
assign w6989 = ~w2568 & ~w6984;
assign w6990 = ~w6988 & w6989;
assign w6991 = ~w6983 & ~w6990;
assign w6992 = pi589 & w3345;
assign w6993 = pi102 & w469;
assign w6994 = pi745 & w3348;
assign w6995 = ~w6992 & ~w6993;
assign w6996 = ~w6994 & w6995;
assign w6997 = pi562 & ~w6996;
assign w6998 = ~pi102 & ~w3355;
assign w6999 = ~w1955 & ~w5872;
assign w7000 = ~w3334 & ~w6996;
assign w7001 = w3355 & ~w6999;
assign w7002 = ~w7000 & w7001;
assign w7003 = ~pi589 & w3358;
assign w7004 = ~pi562 & ~w6998;
assign w7005 = ~w7002 & w7004;
assign w7006 = ~w7003 & w7005;
assign w7007 = ~w6997 & ~w7006;
assign w7008 = pi873 & ~w7007;
assign w7009 = ~pi873 & w7007;
assign w7010 = w2568 & ~w7008;
assign w7011 = ~w7009 & w7010;
assign w7012 = ~pi399 & ~w3367;
assign w7013 = pi295 & ~w7007;
assign w7014 = ~pi295 & w7007;
assign w7015 = ~w7013 & ~w7014;
assign w7016 = w3367 & ~w7015;
assign w7017 = ~w2568 & ~w7012;
assign w7018 = ~w7016 & w7017;
assign w7019 = ~w7011 & ~w7018;
assign w7020 = pi535 & w3345;
assign w7021 = pi064 & w469;
assign w7022 = pi690 & w3348;
assign w7023 = ~w7020 & ~w7021;
assign w7024 = ~w7022 & w7023;
assign w7025 = pi562 & ~w7024;
assign w7026 = ~pi064 & ~w3355;
assign w7027 = ~w1793 & ~w5872;
assign w7028 = ~w3334 & ~w7024;
assign w7029 = w3355 & ~w7027;
assign w7030 = ~w7028 & w7029;
assign w7031 = ~pi535 & w3358;
assign w7032 = ~pi562 & ~w7026;
assign w7033 = ~w7030 & w7032;
assign w7034 = ~w7031 & w7033;
assign w7035 = ~w7025 & ~w7034;
assign w7036 = pi818 & ~w7035;
assign w7037 = ~pi818 & w7035;
assign w7038 = w2568 & ~w7036;
assign w7039 = ~w7037 & w7038;
assign w7040 = ~pi400 & ~w3367;
assign w7041 = pi217 & ~w7035;
assign w7042 = ~pi217 & w7035;
assign w7043 = ~w7041 & ~w7042;
assign w7044 = w3367 & ~w7043;
assign w7045 = ~w2568 & ~w7040;
assign w7046 = ~w7044 & w7045;
assign w7047 = ~w7039 & ~w7046;
assign w7048 = pi627 & w3345;
assign w7049 = pi098 & w469;
assign w7050 = pi742 & w3348;
assign w7051 = ~w7048 & ~w7049;
assign w7052 = ~w7050 & w7051;
assign w7053 = pi562 & ~w7052;
assign w7054 = ~pi098 & ~w3355;
assign w7055 = ~w2166 & ~w5872;
assign w7056 = ~w3334 & ~w7052;
assign w7057 = w3355 & ~w7055;
assign w7058 = ~w7056 & w7057;
assign w7059 = ~pi627 & w3358;
assign w7060 = ~pi562 & ~w7054;
assign w7061 = ~w7058 & w7060;
assign w7062 = ~w7059 & w7061;
assign w7063 = ~w7053 & ~w7062;
assign w7064 = pi870 & ~w7063;
assign w7065 = ~pi870 & w7063;
assign w7066 = w2568 & ~w7064;
assign w7067 = ~w7065 & w7066;
assign w7068 = ~pi401 & ~w3367;
assign w7069 = pi293 & ~w7063;
assign w7070 = ~pi293 & w7063;
assign w7071 = ~w7069 & ~w7070;
assign w7072 = w3367 & ~w7071;
assign w7073 = ~w2568 & ~w7068;
assign w7074 = ~w7072 & w7073;
assign w7075 = ~w7067 & ~w7074;
assign w7076 = pi034 & w469;
assign w7077 = pi613 & w3345;
assign w7078 = pi727 & w3348;
assign w7079 = ~w7076 & ~w7077;
assign w7080 = ~w7078 & w7079;
assign w7081 = pi562 & ~w7080;
assign w7082 = ~pi034 & ~w3355;
assign w7083 = ~w1579 & ~w5872;
assign w7084 = ~w3334 & ~w7080;
assign w7085 = w3355 & ~w7083;
assign w7086 = ~w7084 & w7085;
assign w7087 = ~pi613 & w3358;
assign w7088 = ~pi562 & ~w7082;
assign w7089 = ~w7086 & w7088;
assign w7090 = ~w7087 & w7089;
assign w7091 = ~w7081 & ~w7090;
assign w7092 = pi855 & ~w7091;
assign w7093 = ~pi855 & w7091;
assign w7094 = w2568 & ~w7092;
assign w7095 = ~w7093 & w7094;
assign w7096 = ~pi402 & ~w3367;
assign w7097 = ~pi246 & ~w7091;
assign w7098 = pi246 & w7091;
assign w7099 = ~w7097 & ~w7098;
assign w7100 = w3367 & ~w7099;
assign w7101 = ~w2568 & ~w7096;
assign w7102 = ~w7100 & w7101;
assign w7103 = ~w7095 & ~w7102;
assign w7104 = pi181 & w469;
assign w7105 = pi651 & w3345;
assign w7106 = pi787 & w3348;
assign w7107 = ~w7104 & ~w7105;
assign w7108 = ~w7106 & w7107;
assign w7109 = pi562 & ~w7108;
assign w7110 = ~pi181 & ~w3355;
assign w7111 = ~w2476 & ~w5872;
assign w7112 = ~w3334 & ~w7108;
assign w7113 = w3355 & ~w7111;
assign w7114 = ~w7112 & w7113;
assign w7115 = ~pi651 & w3358;
assign w7116 = ~pi562 & ~w7110;
assign w7117 = ~w7114 & w7116;
assign w7118 = ~w7115 & w7117;
assign w7119 = ~w7109 & ~w7118;
assign w7120 = pi915 & ~w7119;
assign w7121 = ~pi915 & w7119;
assign w7122 = w2568 & ~w7120;
assign w7123 = ~w7121 & w7122;
assign w7124 = ~pi403 & ~w3367;
assign w7125 = pi421 & ~w7119;
assign w7126 = ~pi421 & w7119;
assign w7127 = ~w7125 & ~w7126;
assign w7128 = w3367 & ~w7127;
assign w7129 = ~w2568 & ~w7124;
assign w7130 = ~w7128 & w7129;
assign w7131 = ~w7123 & ~w7130;
assign w7132 = pi090 & w469;
assign w7133 = pi511 & w3345;
assign w7134 = pi693 & w3348;
assign w7135 = ~w7132 & ~w7133;
assign w7136 = ~w7134 & w7135;
assign w7137 = pi562 & ~w7136;
assign w7138 = ~pi090 & ~w3355;
assign w7139 = ~w1961 & ~w5872;
assign w7140 = ~w3334 & ~w7136;
assign w7141 = w3355 & ~w7139;
assign w7142 = ~w7140 & w7141;
assign w7143 = ~pi511 & w3358;
assign w7144 = ~pi562 & ~w7138;
assign w7145 = ~w7142 & w7144;
assign w7146 = ~w7143 & w7145;
assign w7147 = ~w7137 & ~w7146;
assign w7148 = pi821 & ~w7147;
assign w7149 = ~pi821 & w7147;
assign w7150 = w2568 & ~w7148;
assign w7151 = ~w7149 & w7150;
assign w7152 = ~pi404 & ~w3367;
assign w7153 = pi218 & ~w7147;
assign w7154 = ~pi218 & w7147;
assign w7155 = ~w7153 & ~w7154;
assign w7156 = w3367 & ~w7155;
assign w7157 = ~w2568 & ~w7152;
assign w7158 = ~w7156 & w7157;
assign w7159 = ~w7151 & ~w7158;
assign w7160 = pi094 & w469;
assign w7161 = pi633 & w3345;
assign w7162 = pi725 & w3348;
assign w7163 = ~w7160 & ~w7161;
assign w7164 = ~w7162 & w7163;
assign w7165 = pi562 & ~w7164;
assign w7166 = ~pi094 & ~w3355;
assign w7167 = ~w2001 & ~w5872;
assign w7168 = ~w3334 & ~w7164;
assign w7169 = w3355 & ~w7167;
assign w7170 = ~w7168 & w7169;
assign w7171 = ~pi633 & w3358;
assign w7172 = ~pi562 & ~w7166;
assign w7173 = ~w7170 & w7172;
assign w7174 = ~w7171 & w7173;
assign w7175 = ~w7165 & ~w7174;
assign w7176 = pi853 & ~w7175;
assign w7177 = ~pi853 & w7175;
assign w7178 = w2568 & ~w7176;
assign w7179 = ~w7177 & w7178;
assign w7180 = ~pi405 & ~w3367;
assign w7181 = ~pi242 & ~w7175;
assign w7182 = pi242 & w7175;
assign w7183 = ~w7181 & ~w7182;
assign w7184 = w3367 & ~w7183;
assign w7185 = ~w2568 & ~w7180;
assign w7186 = ~w7184 & w7185;
assign w7187 = ~w7179 & ~w7186;
assign w7188 = pi149 & w469;
assign w7189 = pi641 & w3345;
assign w7190 = pi724 & w3348;
assign w7191 = ~w7188 & ~w7189;
assign w7192 = ~w7190 & w7191;
assign w7193 = pi562 & ~w7192;
assign w7194 = ~pi149 & ~w3355;
assign w7195 = ~w2314 & ~w5872;
assign w7196 = ~w3334 & ~w7192;
assign w7197 = w3355 & ~w7195;
assign w7198 = ~w7196 & w7197;
assign w7199 = ~pi641 & w3358;
assign w7200 = ~pi562 & ~w7194;
assign w7201 = ~w7198 & w7200;
assign w7202 = ~w7199 & w7201;
assign w7203 = ~w7193 & ~w7202;
assign w7204 = pi852 & ~w7203;
assign w7205 = ~pi852 & w7203;
assign w7206 = w2568 & ~w7204;
assign w7207 = ~w7205 & w7206;
assign w7208 = ~pi406 & ~w3367;
assign w7209 = ~pi241 & ~w7203;
assign w7210 = pi241 & w7203;
assign w7211 = ~w7209 & ~w7210;
assign w7212 = w3367 & ~w7211;
assign w7213 = ~w2568 & ~w7208;
assign w7214 = ~w7212 & w7213;
assign w7215 = ~w7207 & ~w7214;
assign w7216 = pi147 & w469;
assign w7217 = pi519 & w3345;
assign w7218 = pi692 & w3348;
assign w7219 = ~w7216 & ~w7217;
assign w7220 = ~w7218 & w7219;
assign w7221 = pi562 & ~w7220;
assign w7222 = ~pi147 & ~w3355;
assign w7223 = ~w2295 & ~w5872;
assign w7224 = ~w3334 & ~w7220;
assign w7225 = w3355 & ~w7223;
assign w7226 = ~w7224 & w7225;
assign w7227 = ~pi519 & w3358;
assign w7228 = ~pi562 & ~w7222;
assign w7229 = ~w7226 & w7228;
assign w7230 = ~w7227 & w7229;
assign w7231 = ~w7221 & ~w7230;
assign w7232 = pi820 & ~w7231;
assign w7233 = ~pi820 & w7231;
assign w7234 = w2568 & ~w7232;
assign w7235 = ~w7233 & w7234;
assign w7236 = ~pi407 & ~w3367;
assign w7237 = pi219 & ~w7231;
assign w7238 = ~pi219 & w7231;
assign w7239 = ~w7237 & ~w7238;
assign w7240 = w3367 & ~w7239;
assign w7241 = ~w2568 & ~w7236;
assign w7242 = ~w7240 & w7241;
assign w7243 = ~w7235 & ~w7242;
assign w7244 = pi068 & w469;
assign w7245 = pi583 & w3345;
assign w7246 = pi722 & w3348;
assign w7247 = ~w7244 & ~w7245;
assign w7248 = ~w7246 & w7247;
assign w7249 = pi562 & ~w7248;
assign w7250 = ~pi068 & ~w3355;
assign w7251 = ~w1803 & ~w5872;
assign w7252 = ~w3334 & ~w7248;
assign w7253 = w3355 & ~w7251;
assign w7254 = ~w7252 & w7253;
assign w7255 = ~pi583 & w3358;
assign w7256 = ~pi562 & ~w7250;
assign w7257 = ~w7254 & w7256;
assign w7258 = ~w7255 & w7257;
assign w7259 = ~w7249 & ~w7258;
assign w7260 = pi850 & ~w7259;
assign w7261 = ~pi850 & w7259;
assign w7262 = w2568 & ~w7260;
assign w7263 = ~w7261 & w7262;
assign w7264 = ~pi408 & ~w3367;
assign w7265 = ~pi245 & ~w7259;
assign w7266 = pi245 & w7259;
assign w7267 = ~w7265 & ~w7266;
assign w7268 = w3367 & ~w7267;
assign w7269 = ~w2568 & ~w7264;
assign w7270 = ~w7268 & w7269;
assign w7271 = ~w7263 & ~w7270;
assign w7272 = w1 & w2979;
assign w7273 = pi409 & ~w1;
assign w7274 = ~w7272 & ~w7273;
assign w7275 = ~w5255 & ~w5677;
assign w7276 = w5255 & w5677;
assign w7277 = ~w7275 & ~w7276;
assign w7278 = w5598 & ~w5654;
assign w7279 = ~w5598 & w5654;
assign w7280 = ~w7278 & ~w7279;
assign w7281 = ~w7277 & ~w7280;
assign w7282 = w7277 & w7280;
assign w7283 = ~w7281 & ~w7282;
assign w7284 = ~w5581 & ~w5783;
assign w7285 = w5581 & w5783;
assign w7286 = ~w7284 & ~w7285;
assign w7287 = pi266 & w5162;
assign w7288 = pi374 & w5164;
assign w7289 = pi353 & w5166;
assign w7290 = pi376 & w5161;
assign w7291 = ~w7287 & ~w7288;
assign w7292 = ~w7289 & w7291;
assign w7293 = w469 & w7292;
assign w7294 = ~w7290 & w7293;
assign w7295 = pi065 & w5166;
assign w7296 = pi092 & w5164;
assign w7297 = ~pi062 & w5162;
assign w7298 = pi067 & w5161;
assign w7299 = ~w7295 & ~w7296;
assign w7300 = ~w7297 & w7299;
assign w7301 = ~w469 & w7300;
assign w7302 = ~w7298 & w7301;
assign w7303 = ~w7294 & ~w7302;
assign w7304 = pi373 & w5166;
assign w7305 = pi330 & w5164;
assign w7306 = pi306 & w5162;
assign w7307 = pi322 & w5161;
assign w7308 = ~w7304 & ~w7305;
assign w7309 = ~w7306 & w7308;
assign w7310 = w469 & w7309;
assign w7311 = ~w7307 & w7310;
assign w7312 = pi109 & w5166;
assign w7313 = pi108 & w5164;
assign w7314 = pi107 & w5162;
assign w7315 = pi106 & w5161;
assign w7316 = ~w7312 & ~w7313;
assign w7317 = ~w7314 & w7316;
assign w7318 = ~w469 & w7317;
assign w7319 = ~w7315 & w7318;
assign w7320 = ~w7311 & ~w7319;
assign w7321 = ~w7303 & ~w7320;
assign w7322 = w7303 & w7320;
assign w7323 = ~w7321 & ~w7322;
assign w7324 = w5564 & ~w7323;
assign w7325 = ~w5564 & w7323;
assign w7326 = ~w7324 & ~w7325;
assign w7327 = pi408 & w5164;
assign w7328 = pi400 & w5162;
assign w7329 = pi366 & w5166;
assign w7330 = pi352 & w5161;
assign w7331 = ~w7327 & ~w7328;
assign w7332 = ~w7329 & w7331;
assign w7333 = w469 & w7332;
assign w7334 = ~w7330 & w7333;
assign w7335 = pi068 & w5164;
assign w7336 = pi066 & w5166;
assign w7337 = pi064 & w5162;
assign w7338 = pi063 & w5161;
assign w7339 = ~w7335 & ~w7336;
assign w7340 = ~w7337 & w7339;
assign w7341 = ~w469 & w7340;
assign w7342 = ~w7338 & w7341;
assign w7343 = ~w7334 & ~w7342;
assign w7344 = pi307 & w5166;
assign w7345 = pi299 & w5164;
assign w7346 = pi264 & w5162;
assign w7347 = pi310 & w5161;
assign w7348 = ~w7344 & ~w7345;
assign w7349 = ~w7346 & w7348;
assign w7350 = w469 & w7349;
assign w7351 = ~w7347 & w7350;
assign w7352 = pi061 & w5162;
assign w7353 = pi060 & w5166;
assign w7354 = pi059 & w5164;
assign w7355 = pi058 & w5161;
assign w7356 = ~w7352 & ~w7353;
assign w7357 = ~w7354 & w7356;
assign w7358 = ~w469 & w7357;
assign w7359 = ~w7355 & w7358;
assign w7360 = ~w7351 & ~w7359;
assign w7361 = ~w5766 & ~w7360;
assign w7362 = w5766 & w7360;
assign w7363 = ~w7361 & ~w7362;
assign w7364 = ~w7343 & ~w7363;
assign w7365 = w7343 & w7363;
assign w7366 = ~w7364 & ~w7365;
assign w7367 = w7326 & w7366;
assign w7368 = ~w7326 & ~w7366;
assign w7369 = ~w7367 & ~w7368;
assign w7370 = ~w5198 & ~w5272;
assign w7371 = w5198 & w5272;
assign w7372 = ~w7370 & ~w7371;
assign w7373 = w5716 & w7372;
assign w7374 = ~w5716 & ~w7372;
assign w7375 = ~w7373 & ~w7374;
assign w7376 = w7369 & w7375;
assign w7377 = ~w7369 & ~w7375;
assign w7378 = pi673 & ~w7376;
assign w7379 = ~w7377 & w7378;
assign w7380 = w7286 & w7379;
assign w7381 = ~w7286 & ~w7379;
assign w7382 = ~w7380 & ~w7381;
assign w7383 = w5161 & ~w7283;
assign w7384 = w7382 & w7383;
assign w7385 = w5161 & w7283;
assign w7386 = w7380 & w7385;
assign w7387 = ~w7286 & w7385;
assign w7388 = ~w7379 & w7387;
assign w7389 = pi410 & ~w5161;
assign w7390 = ~w7388 & ~w7389;
assign w7391 = ~w7386 & w7390;
assign w7392 = ~w7384 & w7391;
assign w7393 = ~w5215 & w5238;
assign w7394 = w5215 & ~w5238;
assign w7395 = ~w7393 & ~w7394;
assign w7396 = w5399 & w7395;
assign w7397 = ~w5399 & ~w7395;
assign w7398 = ~w7396 & ~w7397;
assign w7399 = ~w7369 & w7398;
assign w7400 = w7369 & ~w7398;
assign w7401 = pi673 & ~w7399;
assign w7402 = ~w7400 & w7401;
assign w7403 = ~w5634 & w7402;
assign w7404 = w5634 & ~w7402;
assign w7405 = ~w7403 & ~w7404;
assign w7406 = ~w5181 & ~w5677;
assign w7407 = w5181 & w5677;
assign w7408 = ~w7406 & ~w7407;
assign w7409 = w5766 & ~w7408;
assign w7410 = ~w5766 & w7408;
assign w7411 = ~w7409 & ~w7410;
assign w7412 = w5601 & w7411;
assign w7413 = ~w5601 & ~w7411;
assign w7414 = ~w7412 & ~w7413;
assign w7415 = w5161 & w7414;
assign w7416 = w7405 & w7415;
assign w7417 = w5161 & ~w7414;
assign w7418 = w7403 & w7417;
assign w7419 = pi411 & ~w5161;
assign w7420 = w5634 & w7417;
assign w7421 = ~w7402 & w7420;
assign w7422 = ~w7419 & ~w7421;
assign w7423 = ~w7418 & w7422;
assign w7424 = ~w7416 & w7423;
assign w7425 = ~w5255 & ~w5700;
assign w7426 = w5255 & w5700;
assign w7427 = ~w7425 & ~w7426;
assign w7428 = ~w5564 & w5783;
assign w7429 = w5564 & ~w5783;
assign w7430 = ~w7428 & ~w7429;
assign w7431 = ~w7427 & ~w7430;
assign w7432 = w7427 & w7430;
assign w7433 = ~w7431 & ~w7432;
assign w7434 = w5598 & w7433;
assign w7435 = ~w5598 & ~w7433;
assign w7436 = ~w7434 & ~w7435;
assign w7437 = w5161 & w7436;
assign w7438 = w7405 & w7437;
assign w7439 = w5161 & ~w7436;
assign w7440 = w7403 & w7439;
assign w7441 = pi412 & ~w5161;
assign w7442 = w5634 & w7439;
assign w7443 = ~w7402 & w7442;
assign w7444 = ~w7441 & ~w7443;
assign w7445 = ~w7440 & w7444;
assign w7446 = ~w7438 & w7445;
assign w7447 = w1 & w2952;
assign w7448 = pi413 & ~w1;
assign w7449 = ~w7447 & ~w7448;
assign w7450 = w1 & w2818;
assign w7451 = pi414 & ~w1;
assign w7452 = ~w7450 & ~w7451;
assign w7453 = w1 & w2870;
assign w7454 = pi415 & ~w1;
assign w7455 = ~w7453 & ~w7454;
assign w7456 = w1 & w2897;
assign w7457 = pi416 & ~w1;
assign w7458 = ~w7456 & ~w7457;
assign w7459 = w1 & w2925;
assign w7460 = pi417 & ~w1;
assign w7461 = ~w7459 & ~w7460;
assign w7462 = w1 & w3033;
assign w7463 = pi418 & ~w1;
assign w7464 = ~w7462 & ~w7463;
assign w7465 = w1 & w3006;
assign w7466 = pi419 & ~w1;
assign w7467 = ~w7465 & ~w7466;
assign w7468 = ~w5181 & ~w5700;
assign w7469 = w5181 & w5700;
assign w7470 = ~w7468 & ~w7469;
assign w7471 = w5802 & ~w7470;
assign w7472 = ~w5802 & w7470;
assign w7473 = ~w7471 & ~w7472;
assign w7474 = ~w5634 & ~w7473;
assign w7475 = w5634 & w7473;
assign w7476 = ~w7474 & ~w7475;
assign w7477 = w5161 & w7476;
assign w7478 = ~w7382 & w7477;
assign w7479 = ~w7286 & w7379;
assign w7480 = w5161 & ~w7476;
assign w7481 = w7479 & w7480;
assign w7482 = pi420 & ~w5161;
assign w7483 = w7286 & w7480;
assign w7484 = ~w7379 & w7483;
assign w7485 = ~w7482 & ~w7484;
assign w7486 = ~w7481 & w7485;
assign w7487 = ~w7478 & w7486;
assign w7488 = w1 & w3066;
assign w7489 = pi421 & ~w1;
assign w7490 = ~w7488 & ~w7489;
assign w7491 = w5164 & w5608;
assign w7492 = w5164 & w5607;
assign w7493 = w5507 & w7492;
assign w7494 = pi422 & ~w5164;
assign w7495 = ~w7493 & ~w7494;
assign w7496 = ~w7491 & w7495;
assign w7497 = w5164 & w5754;
assign w7498 = w5164 & ~w5660;
assign w7499 = w5753 & w7498;
assign w7500 = pi423 & ~w5164;
assign w7501 = ~w7499 & ~w7500;
assign w7502 = ~w7497 & w7501;
assign w7503 = w5164 & w5812;
assign w7504 = w5164 & w5811;
assign w7505 = ~w5753 & w7504;
assign w7506 = pi424 & ~w5164;
assign w7507 = ~w7505 & ~w7506;
assign w7508 = ~w7503 & w7507;
assign w7509 = w5166 & w5608;
assign w7510 = w5166 & w5607;
assign w7511 = w5507 & w7510;
assign w7512 = pi425 & ~w5166;
assign w7513 = ~w7511 & ~w7512;
assign w7514 = ~w7509 & w7513;
assign w7515 = w5164 & w5793;
assign w7516 = w5164 & w5792;
assign w7517 = w5507 & w7516;
assign w7518 = pi426 & ~w5164;
assign w7519 = ~w7517 & ~w7518;
assign w7520 = ~w7515 & w7519;
assign w7521 = w5166 & w5793;
assign w7522 = w5166 & w5792;
assign w7523 = w5507 & w7522;
assign w7524 = pi427 & ~w5166;
assign w7525 = ~w7523 & ~w7524;
assign w7526 = ~w7521 & w7525;
assign w7527 = w5166 & w5754;
assign w7528 = w5166 & ~w5660;
assign w7529 = w5753 & w7528;
assign w7530 = pi428 & ~w5166;
assign w7531 = ~w7529 & ~w7530;
assign w7532 = ~w7527 & w7531;
assign w7533 = w5166 & w5812;
assign w7534 = w5166 & w5811;
assign w7535 = ~w5753 & w7534;
assign w7536 = pi429 & ~w5166;
assign w7537 = ~w7535 & ~w7536;
assign w7538 = ~w7533 & w7537;
assign w7539 = w1 & w3093;
assign w7540 = pi430 & ~w1;
assign w7541 = ~w7539 & ~w7540;
assign w7542 = w1 & w3120;
assign w7543 = pi431 & ~w1;
assign w7544 = ~w7542 & ~w7543;
assign w7545 = w1 & w3228;
assign w7546 = pi432 & ~w1;
assign w7547 = ~w7545 & ~w7546;
assign w7548 = w1 & w3147;
assign w7549 = pi433 & ~w1;
assign w7550 = ~w7548 & ~w7549;
assign w7551 = w1 & w3201;
assign w7552 = pi434 & ~w1;
assign w7553 = ~w7551 & ~w7552;
assign w7554 = ~w23 & ~w2577;
assign w7555 = w1 & w3174;
assign w7556 = pi436 & ~w1;
assign w7557 = ~w7555 & ~w7556;
assign w7558 = w1 & w2844;
assign w7559 = pi437 & ~w1;
assign w7560 = ~w7558 & ~w7559;
assign w7561 = ~w5238 & ~w5726;
assign w7562 = w5238 & w5726;
assign w7563 = ~w7561 & ~w7562;
assign w7564 = ~w5680 & ~w7360;
assign w7565 = w5680 & w7360;
assign w7566 = ~w7564 & ~w7565;
assign w7567 = ~w7563 & ~w7566;
assign w7568 = w7563 & w7566;
assign w7569 = ~w7567 & ~w7568;
assign w7570 = ~w5654 & ~w7303;
assign w7571 = w5654 & w7303;
assign w7572 = ~w7570 & ~w7571;
assign w7573 = w5161 & w7572;
assign w7574 = w7569 & w7573;
assign w7575 = w5161 & ~w7572;
assign w7576 = w7568 & w7575;
assign w7577 = ~w7566 & w7575;
assign w7578 = ~w7563 & w7577;
assign w7579 = pi438 & ~w5161;
assign w7580 = ~w7578 & ~w7579;
assign w7581 = ~w7576 & w7580;
assign w7582 = ~w7574 & w7581;
assign w7583 = ~w5564 & ~w7360;
assign w7584 = w5564 & w7360;
assign w7585 = ~w7583 & ~w7584;
assign w7586 = ~w7320 & ~w7585;
assign w7587 = w7320 & w7585;
assign w7588 = ~w7586 & ~w7587;
assign w7589 = w5476 & w5802;
assign w7590 = ~w5476 & ~w5802;
assign w7591 = ~w7589 & ~w7590;
assign w7592 = ~w7588 & w7591;
assign w7593 = w7588 & ~w7591;
assign w7594 = pi673 & ~w7592;
assign w7595 = ~w7593 & w7594;
assign w7596 = w5221 & ~w7427;
assign w7597 = ~w5221 & w7427;
assign w7598 = ~w7596 & ~w7597;
assign w7599 = w7595 & w7598;
assign w7600 = ~w7595 & ~w7598;
assign w7601 = ~w7599 & ~w7600;
assign w7602 = w5161 & w7601;
assign w7603 = pi439 & ~w5161;
assign w7604 = ~w7602 & ~w7603;
assign w7605 = ~w5483 & ~w7372;
assign w7606 = w5483 & w7372;
assign w7607 = ~w7605 & ~w7606;
assign w7608 = ~w5215 & ~w7607;
assign w7609 = w5215 & w7607;
assign w7610 = ~w7608 & ~w7609;
assign w7611 = w5161 & w7366;
assign w7612 = w7610 & w7611;
assign w7613 = w5161 & ~w7366;
assign w7614 = w7609 & w7613;
assign w7615 = ~w5215 & w7613;
assign w7616 = ~w7607 & w7615;
assign w7617 = pi440 & ~w5161;
assign w7618 = ~w7616 & ~w7617;
assign w7619 = ~w7614 & w7618;
assign w7620 = ~w7612 & w7619;
assign w7621 = ~w5802 & w7303;
assign w7622 = w5802 & ~w7303;
assign w7623 = ~w7621 & ~w7622;
assign w7624 = w7343 & w7623;
assign w7625 = ~w7343 & ~w7623;
assign w7626 = ~w7624 & ~w7625;
assign w7627 = w5654 & w7626;
assign w7628 = ~w5654 & ~w7626;
assign w7629 = ~w7627 & ~w7628;
assign w7630 = ~w5479 & ~w7629;
assign w7631 = w5479 & w7629;
assign w7632 = pi673 & ~w7630;
assign w7633 = ~w7631 & w7632;
assign w7634 = ~w5706 & w7277;
assign w7635 = w5706 & ~w7277;
assign w7636 = ~w7634 & ~w7635;
assign w7637 = w7633 & w7636;
assign w7638 = ~w7633 & ~w7636;
assign w7639 = ~w7637 & ~w7638;
assign w7640 = w5161 & ~w7639;
assign w7641 = pi441 & ~w5161;
assign w7642 = ~w7640 & ~w7641;
assign w7643 = ~w7320 & ~w7343;
assign w7644 = w7320 & w7343;
assign w7645 = ~w7643 & ~w7644;
assign w7646 = w5218 & ~w7645;
assign w7647 = ~w5218 & w7645;
assign w7648 = ~w7646 & ~w7647;
assign w7649 = w5802 & ~w7648;
assign w7650 = ~w5802 & w7648;
assign w7651 = ~w7649 & ~w7650;
assign w7652 = w7563 & w7651;
assign w7653 = ~w7563 & ~w7651;
assign w7654 = ~w7652 & ~w7653;
assign w7655 = w5161 & ~w7654;
assign w7656 = pi442 & ~w5161;
assign w7657 = ~w7655 & ~w7656;
assign w7658 = ~w7408 & w7595;
assign w7659 = w7408 & ~w7595;
assign w7660 = ~w7658 & ~w7659;
assign w7661 = w5278 & w7660;
assign w7662 = ~w5278 & ~w7660;
assign w7663 = ~w7661 & ~w7662;
assign w7664 = w5161 & ~w7663;
assign w7665 = pi443 & ~w5161;
assign w7666 = ~w7664 & ~w7665;
assign w7667 = w5164 & w7436;
assign w7668 = w7405 & w7667;
assign w7669 = w5164 & ~w7436;
assign w7670 = w7403 & w7669;
assign w7671 = pi444 & ~w5164;
assign w7672 = w5634 & w7669;
assign w7673 = ~w7402 & w7672;
assign w7674 = ~w7671 & ~w7673;
assign w7675 = ~w7670 & w7674;
assign w7676 = ~w7668 & w7675;
assign w7677 = w5164 & ~w7283;
assign w7678 = w7382 & w7677;
assign w7679 = w5164 & w7283;
assign w7680 = w7380 & w7679;
assign w7681 = ~w7286 & w7679;
assign w7682 = ~w7379 & w7681;
assign w7683 = pi445 & ~w5164;
assign w7684 = ~w7682 & ~w7683;
assign w7685 = ~w7680 & w7684;
assign w7686 = ~w7678 & w7685;
assign w7687 = w5164 & w7414;
assign w7688 = w7405 & w7687;
assign w7689 = w5164 & ~w7414;
assign w7690 = w7403 & w7689;
assign w7691 = pi446 & ~w5164;
assign w7692 = w5634 & w7689;
assign w7693 = ~w7402 & w7692;
assign w7694 = ~w7691 & ~w7693;
assign w7695 = ~w7690 & w7694;
assign w7696 = ~w7688 & w7695;
assign w7697 = w5164 & w7476;
assign w7698 = ~w7382 & w7697;
assign w7699 = w5164 & ~w7476;
assign w7700 = w7479 & w7699;
assign w7701 = pi447 & ~w5164;
assign w7702 = w7286 & w7699;
assign w7703 = ~w7379 & w7702;
assign w7704 = ~w7701 & ~w7703;
assign w7705 = ~w7700 & w7704;
assign w7706 = ~w7698 & w7705;
assign w7707 = w5166 & w7436;
assign w7708 = w7405 & w7707;
assign w7709 = w5166 & ~w7436;
assign w7710 = w7403 & w7709;
assign w7711 = pi448 & ~w5166;
assign w7712 = w5634 & w7709;
assign w7713 = ~w7402 & w7712;
assign w7714 = ~w7711 & ~w7713;
assign w7715 = ~w7710 & w7714;
assign w7716 = ~w7708 & w7715;
assign w7717 = w5166 & ~w7283;
assign w7718 = w7382 & w7717;
assign w7719 = w5166 & w7283;
assign w7720 = w7380 & w7719;
assign w7721 = ~w7286 & w7719;
assign w7722 = ~w7379 & w7721;
assign w7723 = pi449 & ~w5166;
assign w7724 = ~w7722 & ~w7723;
assign w7725 = ~w7720 & w7724;
assign w7726 = ~w7718 & w7725;
assign w7727 = ~w5238 & w7607;
assign w7728 = w5238 & ~w7607;
assign w7729 = ~w7727 & ~w7728;
assign w7730 = w5161 & w7326;
assign w7731 = w7729 & w7730;
assign w7732 = w5161 & ~w7326;
assign w7733 = w7727 & w7732;
assign w7734 = pi450 & ~w5161;
assign w7735 = w5238 & w7732;
assign w7736 = ~w7607 & w7735;
assign w7737 = ~w7734 & ~w7736;
assign w7738 = ~w7733 & w7737;
assign w7739 = ~w7731 & w7738;
assign w7740 = w5683 & ~w7470;
assign w7741 = ~w5683 & w7470;
assign w7742 = ~w7740 & ~w7741;
assign w7743 = w7633 & w7742;
assign w7744 = ~w7633 & ~w7742;
assign w7745 = ~w7743 & ~w7744;
assign w7746 = w5161 & ~w7745;
assign w7747 = ~pi451 & ~w5161;
assign w7748 = ~w7746 & ~w7747;
assign w7749 = w5166 & w7476;
assign w7750 = ~w7382 & w7749;
assign w7751 = w5166 & ~w7476;
assign w7752 = w7479 & w7751;
assign w7753 = pi452 & ~w5166;
assign w7754 = w7286 & w7751;
assign w7755 = ~w7379 & w7754;
assign w7756 = ~w7753 & ~w7755;
assign w7757 = ~w7752 & w7756;
assign w7758 = ~w7750 & w7757;
assign w7759 = w5166 & w7414;
assign w7760 = w7405 & w7759;
assign w7761 = w5166 & ~w7414;
assign w7762 = w7403 & w7761;
assign w7763 = pi453 & ~w5166;
assign w7764 = w5634 & w7761;
assign w7765 = ~w7402 & w7764;
assign w7766 = ~w7763 & ~w7765;
assign w7767 = ~w7762 & w7766;
assign w7768 = ~w7760 & w7767;
assign w7769 = pi673 & ~w5716;
assign w7770 = w7360 & ~w7626;
assign w7771 = ~w7360 & w7626;
assign w7772 = ~w7770 & ~w7771;
assign w7773 = w7769 & w7772;
assign w7774 = ~w7769 & ~w7772;
assign w7775 = ~w7773 & ~w7774;
assign w7776 = w5161 & ~w7775;
assign w7777 = pi454 & ~w5161;
assign w7778 = ~w7776 & ~w7777;
assign w7779 = ~w7411 & ~w7433;
assign w7780 = w7411 & w7433;
assign w7781 = ~w7779 & ~w7780;
assign w7782 = w5479 & w5581;
assign w7783 = ~w5479 & ~w5581;
assign w7784 = ~w7782 & ~w7783;
assign w7785 = w7781 & ~w7784;
assign w7786 = ~w7781 & w7784;
assign w7787 = pi673 & ~w7785;
assign w7788 = ~w7786 & w7787;
assign w7789 = ~w5393 & w5501;
assign w7790 = w5393 & ~w5501;
assign w7791 = ~w7789 & ~w7790;
assign w7792 = w5541 & w7791;
assign w7793 = ~w5541 & ~w7791;
assign w7794 = ~w7792 & ~w7793;
assign w7795 = w5299 & ~w7794;
assign w7796 = ~w5299 & w7794;
assign w7797 = ~w7795 & ~w7796;
assign w7798 = w7788 & w7797;
assign w7799 = ~w7788 & ~w7797;
assign w7800 = ~w7798 & ~w7799;
assign w7801 = w5161 & ~w7800;
assign w7802 = pi455 & ~w5161;
assign w7803 = ~w7801 & ~w7802;
assign w7804 = ~w7283 & ~w7473;
assign w7805 = w7283 & w7473;
assign w7806 = ~w7804 & ~w7805;
assign w7807 = w5634 & w5722;
assign w7808 = ~w5634 & ~w5722;
assign w7809 = ~w7807 & ~w7808;
assign w7810 = ~w7806 & w7809;
assign w7811 = w7806 & ~w7809;
assign w7812 = pi673 & ~w7810;
assign w7813 = ~w7811 & w7812;
assign w7814 = ~w5299 & ~w5356;
assign w7815 = w5299 & w5356;
assign w7816 = ~w7814 & ~w7815;
assign w7817 = w5373 & ~w7816;
assign w7818 = ~w5373 & w7816;
assign w7819 = ~w7817 & ~w7818;
assign w7820 = w5544 & ~w7819;
assign w7821 = ~w5544 & w7819;
assign w7822 = ~w7820 & ~w7821;
assign w7823 = w7813 & w7822;
assign w7824 = ~w7813 & ~w7822;
assign w7825 = ~w7823 & ~w7824;
assign w7826 = w5161 & ~w7825;
assign w7827 = pi456 & ~w5161;
assign w7828 = ~w7826 & ~w7827;
assign w7829 = w5604 & w5747;
assign w7830 = ~w5604 & ~w5747;
assign w7831 = ~w7829 & ~w7830;
assign w7832 = w5789 & w7831;
assign w7833 = ~w5789 & ~w7831;
assign w7834 = pi673 & ~w7832;
assign w7835 = ~w7833 & w7834;
assign w7836 = ~w5373 & ~w5470;
assign w7837 = w5373 & w5470;
assign w7838 = ~w7836 & ~w7837;
assign w7839 = w5316 & ~w5453;
assign w7840 = ~w5316 & w5453;
assign w7841 = ~w7839 & ~w7840;
assign w7842 = w5356 & w7841;
assign w7843 = ~w5356 & ~w7841;
assign w7844 = ~w7842 & ~w7843;
assign w7845 = w7838 & ~w7844;
assign w7846 = ~w7838 & w7844;
assign w7847 = ~w7845 & ~w7846;
assign w7848 = w7835 & w7847;
assign w7849 = ~w7835 & ~w7847;
assign w7850 = ~w7848 & ~w7849;
assign w7851 = w5161 & ~w7850;
assign w7852 = pi457 & ~w5161;
assign w7853 = ~w7851 & ~w7852;
assign w7854 = w7572 & ~w7645;
assign w7855 = ~w7572 & w7645;
assign w7856 = ~w7854 & ~w7855;
assign w7857 = w7769 & w7856;
assign w7858 = ~w7769 & ~w7856;
assign w7859 = ~w7857 & ~w7858;
assign w7860 = w5161 & w7859;
assign w7861 = pi458 & ~w5161;
assign w7862 = ~w7860 & ~w7861;
assign w7863 = pi673 & ~w5399;
assign w7864 = w7323 & ~w7363;
assign w7865 = ~w7323 & w7363;
assign w7866 = ~w7864 & ~w7865;
assign w7867 = w7863 & w7866;
assign w7868 = ~w7863 & ~w7866;
assign w7869 = ~w7867 & ~w7868;
assign w7870 = w5161 & w7869;
assign w7871 = pi459 & ~w5161;
assign w7872 = ~w7870 & ~w7871;
assign w7873 = w7585 & ~w7645;
assign w7874 = ~w7585 & w7645;
assign w7875 = ~w7873 & ~w7874;
assign w7876 = w7863 & w7875;
assign w7877 = ~w7863 & ~w7875;
assign w7878 = ~w7876 & ~w7877;
assign w7879 = w5161 & w7878;
assign w7880 = pi460 & ~w5161;
assign w7881 = ~w7879 & ~w7880;
assign w7882 = w5660 & w5811;
assign w7883 = ~w5660 & ~w5811;
assign w7884 = pi673 & ~w7882;
assign w7885 = ~w7883 & w7884;
assign w7886 = ~w5333 & ~w5390;
assign w7887 = w5333 & w5390;
assign w7888 = ~w7886 & ~w7887;
assign w7889 = ~w7844 & w7888;
assign w7890 = w7844 & ~w7888;
assign w7891 = ~w7889 & ~w7890;
assign w7892 = w7885 & w7891;
assign w7893 = ~w7885 & ~w7891;
assign w7894 = ~w7892 & ~w7893;
assign w7895 = w5161 & ~w7894;
assign w7896 = pi461 & ~w5161;
assign w7897 = ~w7895 & ~w7896;
assign w7898 = w5339 & ~w7838;
assign w7899 = ~w5339 & w7838;
assign w7900 = ~w7898 & ~w7899;
assign w7901 = w7885 & w7900;
assign w7902 = ~w7885 & ~w7900;
assign w7903 = ~w7901 & ~w7902;
assign w7904 = w5161 & ~w7903;
assign w7905 = ~pi462 & ~w5161;
assign w7906 = ~w7904 & ~w7905;
assign w7907 = w5713 & ~w7888;
assign w7908 = ~w5713 & w7888;
assign w7909 = ~w7907 & ~w7908;
assign w7910 = w7835 & w7909;
assign w7911 = ~w7835 & ~w7909;
assign w7912 = ~w7910 & ~w7911;
assign w7913 = w5161 & ~w7912;
assign w7914 = ~pi463 & ~w5161;
assign w7915 = ~w7913 & ~w7914;
assign w7916 = pi464 & ~w5161;
assign w7917 = w5501 & ~w5744;
assign w7918 = ~w5501 & w5744;
assign w7919 = ~w7917 & ~w7918;
assign w7920 = w7816 & w7919;
assign w7921 = ~w7816 & ~w7919;
assign w7922 = ~w7920 & ~w7921;
assign w7923 = w5390 & ~w7922;
assign w7924 = ~w5390 & w7922;
assign w7925 = ~w7923 & ~w7924;
assign w7926 = w7813 & w7925;
assign w7927 = ~w7813 & ~w7925;
assign w7928 = ~w7926 & ~w7927;
assign w7929 = w5161 & ~w7928;
assign w7930 = ~w7916 & ~w7929;
assign w7931 = w5396 & ~w5763;
assign w7932 = ~w5396 & w5763;
assign w7933 = ~w7931 & ~w7932;
assign w7934 = w7788 & w7933;
assign w7935 = ~w7788 & ~w7933;
assign w7936 = ~w7934 & ~w7935;
assign w7937 = w5161 & ~w7936;
assign w7938 = ~pi465 & ~w5161;
assign w7939 = ~w7937 & ~w7938;
assign w7940 = w5162 & w5753;
assign w7941 = w5162 & w5660;
assign w7942 = ~pi466 & ~w5162;
assign w7943 = ~w7941 & ~w7942;
assign w7944 = ~w7940 & w7943;
assign w7945 = w5753 & w7941;
assign w7946 = ~w7944 & ~w7945;
assign w7947 = w5162 & w5507;
assign w7948 = ~w5792 & w7947;
assign w7949 = w5162 & w5792;
assign w7950 = ~w5507 & w7949;
assign w7951 = pi467 & ~w5162;
assign w7952 = ~w7950 & ~w7951;
assign w7953 = ~w7948 & w7952;
assign w7954 = ~pi468 & ~w5162;
assign w7955 = w5162 & w5811;
assign w7956 = ~w7954 & ~w7955;
assign w7957 = ~w7940 & ~w7956;
assign w7958 = ~w5811 & w7940;
assign w7959 = ~w7957 & ~w7958;
assign w7960 = ~w5607 & w7947;
assign w7961 = w5162 & w5607;
assign w7962 = ~w5507 & w7961;
assign w7963 = pi469 & ~w5162;
assign w7964 = ~w7962 & ~w7963;
assign w7965 = ~w7960 & w7964;
assign w7966 = w5164 & w7326;
assign w7967 = w7729 & w7966;
assign w7968 = w5164 & ~w7326;
assign w7969 = w7727 & w7968;
assign w7970 = pi470 & ~w5164;
assign w7971 = w5238 & w7968;
assign w7972 = ~w7607 & w7971;
assign w7973 = ~w7970 & ~w7972;
assign w7974 = ~w7969 & w7973;
assign w7975 = ~w7967 & w7974;
assign w7976 = w5164 & ~w7745;
assign w7977 = ~pi471 & ~w5164;
assign w7978 = ~w7976 & ~w7977;
assign w7979 = w5164 & w7601;
assign w7980 = pi472 & ~w5164;
assign w7981 = ~w7979 & ~w7980;
assign w7982 = w5164 & w7572;
assign w7983 = w7569 & w7982;
assign w7984 = w5164 & ~w7572;
assign w7985 = w7568 & w7984;
assign w7986 = ~w7566 & w7984;
assign w7987 = ~w7563 & w7986;
assign w7988 = pi473 & ~w5164;
assign w7989 = ~w7987 & ~w7988;
assign w7990 = ~w7985 & w7989;
assign w7991 = ~w7983 & w7990;
assign w7992 = w5164 & w7366;
assign w7993 = w7610 & w7992;
assign w7994 = w5164 & ~w7366;
assign w7995 = w7609 & w7994;
assign w7996 = ~w5215 & w7994;
assign w7997 = ~w7607 & w7996;
assign w7998 = pi474 & ~w5164;
assign w7999 = ~w7997 & ~w7998;
assign w8000 = ~w7995 & w7999;
assign w8001 = ~w7993 & w8000;
assign w8002 = w5164 & ~w7639;
assign w8003 = pi475 & ~w5164;
assign w8004 = ~w8002 & ~w8003;
assign w8005 = w5164 & ~w7654;
assign w8006 = pi476 & ~w5164;
assign w8007 = ~w8005 & ~w8006;
assign w8008 = w5164 & ~w7663;
assign w8009 = pi477 & ~w5164;
assign w8010 = ~w8008 & ~w8009;
assign w8011 = w5166 & w7326;
assign w8012 = w7729 & w8011;
assign w8013 = w5166 & ~w7326;
assign w8014 = w7727 & w8013;
assign w8015 = pi478 & ~w5166;
assign w8016 = w5238 & w8013;
assign w8017 = ~w7607 & w8016;
assign w8018 = ~w8015 & ~w8017;
assign w8019 = ~w8014 & w8018;
assign w8020 = ~w8012 & w8019;
assign w8021 = w5166 & ~w7745;
assign w8022 = ~pi479 & ~w5166;
assign w8023 = ~w8021 & ~w8022;
assign w8024 = w5166 & w7601;
assign w8025 = pi480 & ~w5166;
assign w8026 = ~w8024 & ~w8025;
assign w8027 = w5166 & w7572;
assign w8028 = w7569 & w8027;
assign w8029 = w5166 & ~w7572;
assign w8030 = w7568 & w8029;
assign w8031 = ~w7566 & w8029;
assign w8032 = ~w7563 & w8031;
assign w8033 = pi481 & ~w5166;
assign w8034 = ~w8032 & ~w8033;
assign w8035 = ~w8030 & w8034;
assign w8036 = ~w8028 & w8035;
assign w8037 = w5166 & w7366;
assign w8038 = w7610 & w8037;
assign w8039 = w5166 & ~w7366;
assign w8040 = w7609 & w8039;
assign w8041 = ~w5215 & w8039;
assign w8042 = ~w7607 & w8041;
assign w8043 = pi482 & ~w5166;
assign w8044 = ~w8042 & ~w8043;
assign w8045 = ~w8040 & w8044;
assign w8046 = ~w8038 & w8045;
assign w8047 = w5166 & ~w7639;
assign w8048 = pi483 & ~w5166;
assign w8049 = ~w8047 & ~w8048;
assign w8050 = w5166 & ~w7654;
assign w8051 = pi484 & ~w5166;
assign w8052 = ~w8050 & ~w8051;
assign w8053 = w5166 & ~w7663;
assign w8054 = pi485 & ~w5166;
assign w8055 = ~w8053 & ~w8054;
assign w8056 = w5164 & ~w7825;
assign w8057 = pi486 & ~w5164;
assign w8058 = ~w8056 & ~w8057;
assign w8059 = w5164 & ~w7894;
assign w8060 = pi487 & ~w5164;
assign w8061 = ~w8059 & ~w8060;
assign w8062 = w5166 & ~w7936;
assign w8063 = ~pi488 & ~w5166;
assign w8064 = ~w8062 & ~w8063;
assign w8065 = pi489 & ~w5164;
assign w8066 = w5164 & ~w7928;
assign w8067 = ~w8065 & ~w8066;
assign w8068 = w5164 & ~w7936;
assign w8069 = ~pi490 & ~w5164;
assign w8070 = ~w8068 & ~w8069;
assign w8071 = w5164 & ~w7800;
assign w8072 = pi491 & ~w5164;
assign w8073 = ~w8071 & ~w8072;
assign w8074 = pi492 & ~w5166;
assign w8075 = w5166 & ~w7928;
assign w8076 = ~w8074 & ~w8075;
assign w8077 = w5162 & w7436;
assign w8078 = w7405 & w8077;
assign w8079 = w5162 & ~w7436;
assign w8080 = w7403 & w8079;
assign w8081 = ~pi493 & ~w5162;
assign w8082 = w5634 & w8079;
assign w8083 = ~w7402 & w8082;
assign w8084 = ~w8081 & ~w8083;
assign w8085 = ~w8080 & w8084;
assign w8086 = ~w8078 & w8085;
assign w8087 = w5164 & ~w7912;
assign w8088 = ~pi494 & ~w5164;
assign w8089 = ~w8087 & ~w8088;
assign w8090 = w5164 & ~w7903;
assign w8091 = ~pi495 & ~w5164;
assign w8092 = ~w8090 & ~w8091;
assign w8093 = w5164 & ~w7850;
assign w8094 = pi496 & ~w5164;
assign w8095 = ~w8093 & ~w8094;
assign w8096 = w5166 & ~w7912;
assign w8097 = ~pi497 & ~w5166;
assign w8098 = ~w8096 & ~w8097;
assign w8099 = w5166 & ~w7903;
assign w8100 = ~pi498 & ~w5166;
assign w8101 = ~w8099 & ~w8100;
assign w8102 = w5166 & ~w7850;
assign w8103 = pi499 & ~w5166;
assign w8104 = ~w8102 & ~w8103;
assign w8105 = w5166 & ~w7894;
assign w8106 = pi500 & ~w5166;
assign w8107 = ~w8105 & ~w8106;
assign w8108 = w5164 & w7878;
assign w8109 = pi501 & ~w5164;
assign w8110 = ~w8108 & ~w8109;
assign w8111 = w5164 & w7869;
assign w8112 = pi502 & ~w5164;
assign w8113 = ~w8111 & ~w8112;
assign w8114 = w5164 & ~w7775;
assign w8115 = pi503 & ~w5164;
assign w8116 = ~w8114 & ~w8115;
assign w8117 = w5166 & w7878;
assign w8118 = pi504 & ~w5166;
assign w8119 = ~w8117 & ~w8118;
assign w8120 = w5166 & ~w7775;
assign w8121 = pi505 & ~w5166;
assign w8122 = ~w8120 & ~w8121;
assign w8123 = w5166 & w7869;
assign w8124 = pi506 & ~w5166;
assign w8125 = ~w8123 & ~w8124;
assign w8126 = w5166 & w7859;
assign w8127 = pi507 & ~w5166;
assign w8128 = ~w8126 & ~w8127;
assign w8129 = w5164 & w7859;
assign w8130 = pi508 & ~w5164;
assign w8131 = ~w8129 & ~w8130;
assign w8132 = w5162 & w7286;
assign w8133 = ~w7379 & w8132;
assign w8134 = w5162 & ~w7286;
assign w8135 = w7379 & w8134;
assign w8136 = ~w8133 & ~w8135;
assign w8137 = w7476 & ~w8136;
assign w8138 = ~w7476 & w8132;
assign w8139 = w7379 & w8138;
assign w8140 = pi509 & ~w5162;
assign w8141 = ~w7476 & w8134;
assign w8142 = ~w7379 & w8141;
assign w8143 = ~w8139 & ~w8140;
assign w8144 = ~w8142 & w8143;
assign w8145 = ~w8137 & w8144;
assign w8146 = w5162 & w7283;
assign w8147 = w7382 & w8146;
assign w8148 = ~pi510 & ~w5162;
assign w8149 = ~w8146 & ~w8148;
assign w8150 = w8136 & w8149;
assign w8151 = ~w8147 & ~w8150;
assign w8152 = w5162 & w7414;
assign w8153 = w7405 & w8152;
assign w8154 = w5162 & ~w7414;
assign w8155 = w7403 & w8154;
assign w8156 = ~pi511 & ~w5162;
assign w8157 = w5634 & w8154;
assign w8158 = ~w7402 & w8157;
assign w8159 = ~w8156 & ~w8158;
assign w8160 = ~w8155 & w8159;
assign w8161 = ~w8153 & w8160;
assign w8162 = w5166 & ~w7800;
assign w8163 = pi512 & ~w5166;
assign w8164 = ~w8162 & ~w8163;
assign w8165 = w5166 & ~w7825;
assign w8166 = pi513 & ~w5166;
assign w8167 = ~w8165 & ~w8166;
assign w8168 = w5544 & ~w7922;
assign w8169 = ~w5544 & w7922;
assign w8170 = pi673 & ~w8168;
assign w8171 = ~w8169 & w8170;
assign w8172 = w5470 & ~w5719;
assign w8173 = ~w5470 & w5719;
assign w8174 = ~w8172 & ~w8173;
assign w8175 = ~w5316 & ~w5433;
assign w8176 = w5316 & w5433;
assign w8177 = ~w8175 & ~w8176;
assign w8178 = w8174 & ~w8177;
assign w8179 = ~w8174 & w8177;
assign w8180 = ~w8178 & ~w8179;
assign w8181 = w8171 & w8180;
assign w8182 = ~w8171 & ~w8180;
assign w8183 = ~w8181 & ~w8182;
assign w8184 = w5161 & ~w8183;
assign w8185 = pi514 & ~w5161;
assign w8186 = ~w8184 & ~w8185;
assign w8187 = w5763 & ~w7794;
assign w8188 = ~w5763 & w7794;
assign w8189 = pi673 & ~w8187;
assign w8190 = ~w8188 & w8189;
assign w8191 = ~w5453 & ~w5564;
assign w8192 = w5453 & w5564;
assign w8193 = ~w8191 & ~w8192;
assign w8194 = w8177 & ~w8193;
assign w8195 = ~w8177 & w8193;
assign w8196 = ~w8194 & ~w8195;
assign w8197 = w8190 & w8196;
assign w8198 = ~w8190 & ~w8196;
assign w8199 = ~w8197 & ~w8198;
assign w8200 = w5161 & w8199;
assign w8201 = pi515 & ~w5161;
assign w8202 = ~w8200 & ~w8201;
assign w8203 = ~w5333 & ~w5651;
assign w8204 = w5333 & w5651;
assign w8205 = ~w8203 & ~w8204;
assign w8206 = ~w5436 & ~w8205;
assign w8207 = w5436 & w8205;
assign w8208 = ~w8206 & ~w8207;
assign w8209 = w5470 & ~w8208;
assign w8210 = ~w5470 & w8208;
assign w8211 = ~w8209 & ~w8210;
assign w8212 = w8190 & w8211;
assign w8213 = ~w8190 & ~w8211;
assign w8214 = ~w8212 & ~w8213;
assign w8215 = w5161 & w8214;
assign w8216 = pi516 & ~w5161;
assign w8217 = ~w8215 & ~w8216;
assign w8218 = w8193 & ~w8205;
assign w8219 = ~w8193 & w8205;
assign w8220 = ~w8218 & ~w8219;
assign w8221 = w8171 & w8220;
assign w8222 = ~w8171 & ~w8220;
assign w8223 = ~w8221 & ~w8222;
assign w8224 = w5161 & w8223;
assign w8225 = pi517 & ~w5161;
assign w8226 = ~w8224 & ~w8225;
assign w8227 = w5162 & w7366;
assign w8228 = ~pi518 & ~w5162;
assign w8229 = ~w8227 & ~w8228;
assign w8230 = w7610 & ~w8229;
assign w8231 = pi518 & ~w5162;
assign w8232 = ~w8227 & ~w8231;
assign w8233 = ~w7610 & w8232;
assign w8234 = ~w8230 & ~w8233;
assign w8235 = w5162 & w7639;
assign w8236 = pi519 & ~w5162;
assign w8237 = ~w8235 & ~w8236;
assign w8238 = w5162 & w7326;
assign w8239 = w7729 & w8238;
assign w8240 = w5162 & ~w7326;
assign w8241 = w7727 & w8240;
assign w8242 = ~pi520 & ~w5162;
assign w8243 = w5238 & w8240;
assign w8244 = ~w7607 & w8243;
assign w8245 = ~w8242 & ~w8244;
assign w8246 = ~w8241 & w8245;
assign w8247 = ~w8239 & w8246;
assign w8248 = w5162 & ~w7654;
assign w8249 = ~pi521 & ~w5162;
assign w8250 = ~w8248 & ~w8249;
assign w8251 = w5162 & w7663;
assign w8252 = pi522 & ~w5162;
assign w8253 = ~w8251 & ~w8252;
assign w8254 = ~pi523 & ~w5162;
assign w8255 = w5162 & ~w7572;
assign w8256 = ~w8254 & ~w8255;
assign w8257 = ~w7569 & ~w8256;
assign w8258 = w5162 & w7572;
assign w8259 = ~w8254 & ~w8258;
assign w8260 = w7569 & ~w8259;
assign w8261 = ~w8257 & ~w8260;
assign w8262 = w5162 & ~w7745;
assign w8263 = pi524 & ~w5162;
assign w8264 = ~w8262 & ~w8263;
assign w8265 = w5162 & ~w7601;
assign w8266 = pi525 & ~w5162;
assign w8267 = ~w8265 & ~w8266;
assign w8268 = w5166 & w8199;
assign w8269 = pi526 & ~w5166;
assign w8270 = ~w8268 & ~w8269;
assign w8271 = w5162 & ~w7859;
assign w8272 = pi527 & ~w5162;
assign w8273 = ~w8271 & ~w8272;
assign w8274 = w5164 & w8223;
assign w8275 = pi528 & ~w5164;
assign w8276 = ~w8274 & ~w8275;
assign w8277 = w5166 & ~w8183;
assign w8278 = pi529 & ~w5166;
assign w8279 = ~w8277 & ~w8278;
assign w8280 = w5162 & w7928;
assign w8281 = pi530 & ~w5162;
assign w8282 = ~w8280 & ~w8281;
assign w8283 = w5162 & w7800;
assign w8284 = pi531 & ~w5162;
assign w8285 = ~w8283 & ~w8284;
assign w8286 = w5164 & w8214;
assign w8287 = pi532 & ~w5164;
assign w8288 = ~w8286 & ~w8287;
assign w8289 = w5162 & w7850;
assign w8290 = pi533 & ~w5162;
assign w8291 = ~w8289 & ~w8290;
assign w8292 = w5162 & w7894;
assign w8293 = pi534 & ~w5162;
assign w8294 = ~w8292 & ~w8293;
assign w8295 = w5162 & ~w7869;
assign w8296 = pi535 & ~w5162;
assign w8297 = ~w8295 & ~w8296;
assign w8298 = w5164 & w8199;
assign w8299 = pi536 & ~w5164;
assign w8300 = ~w8298 & ~w8299;
assign w8301 = w5164 & ~w8183;
assign w8302 = pi537 & ~w5164;
assign w8303 = ~w8301 & ~w8302;
assign w8304 = w5162 & ~w7912;
assign w8305 = pi538 & ~w5162;
assign w8306 = ~w8304 & ~w8305;
assign w8307 = w5162 & ~w7903;
assign w8308 = pi539 & ~w5162;
assign w8309 = ~w8307 & ~w8308;
assign w8310 = w5162 & ~w7878;
assign w8311 = pi540 & ~w5162;
assign w8312 = ~w8310 & ~w8311;
assign w8313 = w5162 & w7775;
assign w8314 = pi541 & ~w5162;
assign w8315 = ~w8313 & ~w8314;
assign w8316 = w5166 & w8214;
assign w8317 = pi542 & ~w5166;
assign w8318 = ~w8316 & ~w8317;
assign w8319 = w5162 & w7825;
assign w8320 = pi543 & ~w5162;
assign w8321 = ~w8319 & ~w8320;
assign w8322 = w5162 & ~w7936;
assign w8323 = pi544 & ~w5162;
assign w8324 = ~w8322 & ~w8323;
assign w8325 = w5166 & w8223;
assign w8326 = pi545 & ~w5166;
assign w8327 = ~w8325 & ~w8326;
assign w8328 = w5162 & ~w8183;
assign w8329 = ~pi546 & ~w5162;
assign w8330 = ~w8328 & ~w8329;
assign w8331 = w5162 & ~w8223;
assign w8332 = pi547 & ~w5162;
assign w8333 = ~w8331 & ~w8332;
assign w8334 = pi548 & ~w5162;
assign w8335 = w5162 & ~w8214;
assign w8336 = ~w8334 & ~w8335;
assign w8337 = w5162 & ~w8199;
assign w8338 = pi549 & ~w5162;
assign w8339 = ~w8337 & ~w8338;
assign w8340 = pi550 & w2568;
assign w8341 = ~w2579 & ~w8340;
assign w8342 = pi551 & w2568;
assign w8343 = ~w2558 & ~w8342;
assign w8344 = pi552 & w2568;
assign w8345 = ~w2563 & ~w8344;
assign w8346 = ~w102 & ~w419;
assign w8347 = pi562 & pi672;
assign w8348 = pi673 & w8347;
assign w8349 = pi562 & ~pi672;
assign w8350 = pi555 & w8349;
assign w8351 = pi435 & ~w528;
assign w8352 = ~pi562 & ~w8351;
assign w8353 = ~pi557 & ~w3334;
assign w8354 = w3341 & ~w8353;
assign w8355 = ~w467 & ~w3336;
assign w8356 = w8354 & ~w8355;
assign w8357 = ~w8354 & w8355;
assign w8358 = w8352 & ~w8356;
assign w8359 = ~w8357 & w8358;
assign w8360 = ~w8348 & ~w8350;
assign w8361 = ~w8359 & w8360;
assign w8362 = pi556 & w8349;
assign w8363 = pi555 & pi557;
assign w8364 = ~w3341 & w8363;
assign w8365 = pi556 & w8364;
assign w8366 = w20 & w3334;
assign w8367 = w466 & w8366;
assign w8368 = pi556 & ~w8366;
assign w8369 = ~w8367 & ~w8368;
assign w8370 = ~w8364 & w8369;
assign w8371 = w8352 & ~w8365;
assign w8372 = ~w8370 & w8371;
assign w8373 = ~w8362 & ~w8372;
assign w8374 = ~w3343 & ~w8347;
assign w8375 = pi557 & ~w8374;
assign w8376 = ~w3342 & w8352;
assign w8377 = ~pi557 & ~w8376;
assign w8378 = ~w8375 & ~w8377;
assign w8379 = pi558 & w8349;
assign w8380 = ~pi558 & ~w8365;
assign w8381 = pi558 & w8365;
assign w8382 = w8352 & ~w8367;
assign w8383 = ~w8380 & w8382;
assign w8384 = ~w8381 & w8383;
assign w8385 = ~w8348 & ~w8379;
assign w8386 = ~w8384 & w8385;
assign w8387 = pi669 & w5158;
assign w8388 = pi667 & ~w3343;
assign w8389 = ~w8351 & ~w8387;
assign w8390 = ~w8388 & w8389;
assign w8391 = ~w5161 & ~w5164;
assign w8392 = ~w5164 & ~w5166;
assign w8393 = ~w8349 & ~w8351;
assign w8394 = ~w537 & ~w1536;
assign w8395 = pi566 & w441;
assign w8396 = pi565 & ~w8395;
assign w8397 = ~w456 & ~w8396;
assign w8398 = ~w1558 & ~w8395;
assign w8399 = ~w452 & w1469;
assign w8400 = ~w1489 & ~w8399;
assign w8401 = pi569 & ~w5162;
assign w8402 = ~pi458 & w5162;
assign w8403 = ~w8401 & ~w8402;
assign w8404 = pi570 & ~w5162;
assign w8405 = ~pi463 & w5162;
assign w8406 = ~w8404 & ~w8405;
assign w8407 = pi571 & ~w5162;
assign w8408 = ~pi438 & w5162;
assign w8409 = ~w8407 & ~w8408;
assign w8410 = pi572 & ~w5162;
assign w8411 = ~pi348 & w5162;
assign w8412 = ~w8410 & ~w8411;
assign w8413 = pi573 & ~w5162;
assign w8414 = ~pi462 & w5162;
assign w8415 = ~w8413 & ~w8414;
assign w8416 = pi574 & ~w5162;
assign w8417 = ~pi459 & w5162;
assign w8418 = ~w8416 & ~w8417;
assign w8419 = pi575 & ~w5162;
assign w8420 = ~pi489 & w5162;
assign w8421 = ~w8419 & ~w8420;
assign w8422 = pi576 & ~w5162;
assign w8423 = ~pi448 & w5162;
assign w8424 = ~w8422 & ~w8423;
assign w8425 = pi577 & ~w5162;
assign w8426 = ~pi497 & w5162;
assign w8427 = ~w8425 & ~w8426;
assign w8428 = pi578 & ~w5162;
assign w8429 = ~pi512 & w5162;
assign w8430 = ~w8428 & ~w8429;
assign w8431 = pi579 & ~w5162;
assign w8432 = ~pi451 & w5162;
assign w8433 = ~w8431 & ~w8432;
assign w8434 = pi580 & ~w5162;
assign w8435 = ~pi483 & w5162;
assign w8436 = ~w8434 & ~w8435;
assign w8437 = pi581 & ~w5162;
assign w8438 = ~pi412 & w5162;
assign w8439 = ~w8437 & ~w8438;
assign w8440 = pi582 & ~w5162;
assign w8441 = ~pi507 & w5162;
assign w8442 = ~w8440 & ~w8441;
assign w8443 = pi583 & ~w5162;
assign w8444 = ~pi502 & w5162;
assign w8445 = ~w8443 & ~w8444;
assign w8446 = pi584 & ~w5162;
assign w8447 = ~pi452 & w5162;
assign w8448 = ~w8446 & ~w8447;
assign w8449 = pi585 & ~w5162;
assign w8450 = ~pi488 & w5162;
assign w8451 = ~w8449 & ~w8450;
assign w8452 = pi586 & ~w5162;
assign w8453 = ~pi476 & w5162;
assign w8454 = ~w8452 & ~w8453;
assign w8455 = pi587 & ~w5162;
assign w8456 = ~pi470 & w5162;
assign w8457 = ~w8455 & ~w8456;
assign w8458 = pi588 & ~w5162;
assign w8459 = ~pi478 & w5162;
assign w8460 = ~w8458 & ~w8459;
assign w8461 = pi589 & ~w5162;
assign w8462 = ~pi529 & w5162;
assign w8463 = ~w8461 & ~w8462;
assign w8464 = pi590 & ~w5162;
assign w8465 = ~pi513 & w5162;
assign w8466 = ~w8464 & ~w8465;
assign w8467 = pi591 & ~w5162;
assign w8468 = ~pi439 & w5162;
assign w8469 = ~w8467 & ~w8468;
assign w8470 = pi592 & ~w5162;
assign w8471 = ~pi492 & w5162;
assign w8472 = ~w8470 & ~w8471;
assign w8473 = pi593 & ~w5162;
assign w8474 = ~pi498 & w5162;
assign w8475 = ~w8473 & ~w8474;
assign w8476 = pi594 & ~w5162;
assign w8477 = ~pi443 & w5162;
assign w8478 = ~w8476 & ~w8477;
assign w8479 = pi595 & ~w5162;
assign w8480 = ~pi504 & w5162;
assign w8481 = ~w8479 & ~w8480;
assign w8482 = pi596 & ~w5162;
assign w8483 = ~pi474 & w5162;
assign w8484 = ~w8482 & ~w8483;
assign w8485 = pi597 & ~w5162;
assign w8486 = ~pi349 & w5162;
assign w8487 = ~w8485 & ~w8486;
assign w8488 = pi598 & ~w5162;
assign w8489 = ~pi499 & w5162;
assign w8490 = ~w8488 & ~w8489;
assign w8491 = pi599 & ~w5162;
assign w8492 = ~pi505 & w5162;
assign w8493 = ~w8491 & ~w8492;
assign w8494 = pi600 & ~w5162;
assign w8495 = ~pi484 & w5162;
assign w8496 = ~w8494 & ~w8495;
assign w8497 = pi601 & ~w5162;
assign w8498 = ~pi461 & w5162;
assign w8499 = ~w8497 & ~w8498;
assign w8500 = pi602 & ~w5162;
assign w8501 = ~pi485 & w5162;
assign w8502 = ~w8500 & ~w8501;
assign w8503 = pi603 & ~w5162;
assign w8504 = ~pi480 & w5162;
assign w8505 = ~w8503 & ~w8504;
assign w8506 = pi604 & ~w5162;
assign w8507 = ~pi503 & w5162;
assign w8508 = ~w8506 & ~w8507;
assign w8509 = pi605 & ~w5162;
assign w8510 = ~pi536 & w5162;
assign w8511 = ~w8509 & ~w8510;
assign w8512 = pi606 & ~w5162;
assign w8513 = ~pi450 & w5162;
assign w8514 = ~w8512 & ~w8513;
assign w8515 = pi607 & ~w5162;
assign w8516 = ~pi445 & w5162;
assign w8517 = ~w8515 & ~w8516;
assign w8518 = pi608 & ~w5162;
assign w8519 = ~pi428 & w5162;
assign w8520 = ~w8518 & ~w8519;
assign w8521 = pi609 & ~w5162;
assign w8522 = ~pi490 & w5162;
assign w8523 = ~w8521 & ~w8522;
assign w8524 = pi610 & ~w5162;
assign w8525 = ~pi427 & w5162;
assign w8526 = ~w8524 & ~w8525;
assign w8527 = pi611 & ~w5162;
assign w8528 = ~pi514 & w5162;
assign w8529 = ~w8527 & ~w8528;
assign w8530 = pi612 & ~w5162;
assign w8531 = ~pi464 & w5162;
assign w8532 = ~w8530 & ~w8531;
assign w8533 = pi613 & ~w5162;
assign w8534 = ~pi491 & w5162;
assign w8535 = ~w8533 & ~w8534;
assign w8536 = pi614 & ~w5162;
assign w8537 = ~pi517 & w5162;
assign w8538 = ~w8536 & ~w8537;
assign w8539 = pi615 & ~w5162;
assign w8540 = ~pi456 & w5162;
assign w8541 = ~w8539 & ~w8540;
assign w8542 = pi616 & ~w5162;
assign w8543 = ~pi422 & w5162;
assign w8544 = ~w8542 & ~w8543;
assign w8545 = pi617 & ~w5162;
assign w8546 = ~pi537 & w5162;
assign w8547 = ~w8545 & ~w8546;
assign w8548 = pi618 & ~w5162;
assign w8549 = ~pi528 & w5162;
assign w8550 = ~w8548 & ~w8549;
assign w8551 = pi619 & ~w5162;
assign w8552 = ~pi487 & w5162;
assign w8553 = ~w8551 & ~w8552;
assign w8554 = pi620 & ~w5162;
assign w8555 = ~pi460 & w5162;
assign w8556 = ~w8554 & ~w8555;
assign w8557 = pi621 & ~w5162;
assign w8558 = ~pi411 & w5162;
assign w8559 = ~w8557 & ~w8558;
assign w8560 = pi622 & ~w5162;
assign w8561 = ~pi495 & w5162;
assign w8562 = ~w8560 & ~w8561;
assign w8563 = pi623 & ~w5162;
assign w8564 = ~pi506 & w5162;
assign w8565 = ~w8563 & ~w8564;
assign w8566 = pi624 & ~w5162;
assign w8567 = ~pi420 & w5162;
assign w8568 = ~w8566 & ~w8567;
assign w8569 = pi625 & ~w5162;
assign w8570 = ~pi453 & w5162;
assign w8571 = ~w8569 & ~w8570;
assign w8572 = pi626 & ~w5162;
assign w8573 = ~pi477 & w5162;
assign w8574 = ~w8572 & ~w8573;
assign w8575 = pi627 & ~w5162;
assign w8576 = ~pi425 & w5162;
assign w8577 = ~w8575 & ~w8576;
assign w8578 = pi628 & ~w5162;
assign w8579 = ~pi465 & w5162;
assign w8580 = ~w8578 & ~w8579;
assign w8581 = pi629 & ~w5162;
assign w8582 = ~pi457 & w5162;
assign w8583 = ~w8581 & ~w8582;
assign w8584 = pi630 & ~w5162;
assign w8585 = ~pi426 & w5162;
assign w8586 = ~w8584 & ~w8585;
assign w8587 = pi631 & ~w5162;
assign w8588 = ~pi447 & w5162;
assign w8589 = ~w8587 & ~w8588;
assign w8590 = pi632 & ~w5162;
assign w8591 = ~pi545 & w5162;
assign w8592 = ~w8590 & ~w8591;
assign w8593 = pi633 & ~w5162;
assign w8594 = ~pi446 & w5162;
assign w8595 = ~w8593 & ~w8594;
assign w8596 = pi634 & ~w5162;
assign w8597 = ~pi479 & w5162;
assign w8598 = ~w8596 & ~w8597;
assign w8599 = pi635 & ~w5162;
assign w8600 = ~pi482 & w5162;
assign w8601 = ~w8599 & ~w8600;
assign w8602 = pi636 & ~w5162;
assign w8603 = ~pi410 & w5162;
assign w8604 = ~w8602 & ~w8603;
assign w8605 = pi637 & ~w5162;
assign w8606 = ~pi423 & w5162;
assign w8607 = ~w8605 & ~w8606;
assign w8608 = pi638 & ~w5162;
assign w8609 = ~pi472 & w5162;
assign w8610 = ~w8608 & ~w8609;
assign w8611 = pi639 & ~w5162;
assign w8612 = ~pi500 & w5162;
assign w8613 = ~w8611 & ~w8612;
assign w8614 = pi640 & ~w5162;
assign w8615 = ~pi496 & w5162;
assign w8616 = ~w8614 & ~w8615;
assign w8617 = pi641 & ~w5162;
assign w8618 = ~pi475 & w5162;
assign w8619 = ~w8617 & ~w8618;
assign w8620 = pi642 & ~w5162;
assign w8621 = ~pi350 & w5162;
assign w8622 = ~w8620 & ~w8621;
assign w8623 = pi643 & ~w5162;
assign w8624 = ~pi501 & w5162;
assign w8625 = ~w8623 & ~w8624;
assign w8626 = pi644 & ~w5162;
assign w8627 = ~pi449 & w5162;
assign w8628 = ~w8626 & ~w8627;
assign w8629 = pi645 & ~w5162;
assign w8630 = ~pi486 & w5162;
assign w8631 = ~w8629 & ~w8630;
assign w8632 = pi646 & ~w5162;
assign w8633 = ~pi532 & w5162;
assign w8634 = ~w8632 & ~w8633;
assign w8635 = pi647 & ~w5162;
assign w8636 = ~pi454 & w5162;
assign w8637 = ~w8635 & ~w8636;
assign w8638 = pi648 & ~w5162;
assign w8639 = ~pi508 & w5162;
assign w8640 = ~w8638 & ~w8639;
assign w8641 = pi649 & ~w5162;
assign w8642 = ~pi515 & w5162;
assign w8643 = ~w8641 & ~w8642;
assign w8644 = pi650 & ~w5162;
assign w8645 = ~pi471 & w5162;
assign w8646 = ~w8644 & ~w8645;
assign w8647 = pi651 & ~w5162;
assign w8648 = ~pi440 & w5162;
assign w8649 = ~w8647 & ~w8648;
assign w8650 = pi652 & ~w5162;
assign w8651 = ~pi473 & w5162;
assign w8652 = ~w8650 & ~w8651;
assign w8653 = pi653 & ~w5162;
assign w8654 = ~pi442 & w5162;
assign w8655 = ~w8653 & ~w8654;
assign w8656 = pi654 & ~w5162;
assign w8657 = ~pi429 & w5162;
assign w8658 = ~w8656 & ~w8657;
assign w8659 = pi655 & ~w5162;
assign w8660 = ~pi455 & w5162;
assign w8661 = ~w8659 & ~w8660;
assign w8662 = pi656 & ~w5162;
assign w8663 = ~pi424 & w5162;
assign w8664 = ~w8662 & ~w8663;
assign w8665 = pi657 & ~w5162;
assign w8666 = ~pi441 & w5162;
assign w8667 = ~w8665 & ~w8666;
assign w8668 = pi658 & ~w5162;
assign w8669 = ~pi494 & w5162;
assign w8670 = ~w8668 & ~w8669;
assign w8671 = pi659 & ~w5162;
assign w8672 = ~pi481 & w5162;
assign w8673 = ~w8671 & ~w8672;
assign w8674 = pi660 & ~w5162;
assign w8675 = ~pi516 & w5162;
assign w8676 = ~w8674 & ~w8675;
assign w8677 = pi661 & ~w5162;
assign w8678 = ~pi542 & w5162;
assign w8679 = ~w8677 & ~w8678;
assign w8680 = pi662 & ~w5162;
assign w8681 = ~pi526 & w5162;
assign w8682 = ~w8680 & ~w8681;
assign w8683 = pi663 & ~w5162;
assign w8684 = ~pi444 & w5162;
assign w8685 = ~w8683 & ~w8684;
assign w8686 = pi664 & ~w5162;
assign w8687 = ~pi347 & w5162;
assign w8688 = ~w8686 & ~w8687;
assign w8689 = ~w102 & ~w424;
assign w8690 = pi668 & pi000;
assign w8691 = ~w26 & pi813;
assign w8692 = w26 & pi000;
assign w8693 = w29 & ~w2;
assign w8694 = w48 & ~w46;
assign w8695 = w45 & pi190;
assign w8696 = pi006 & ~pi007;
assign w8697 = w66 & pi164;
assign w8698 = w45 & ~w42;
assign w8699 = w66 & pi190;
assign w8700 = ~w102 & ~w100;
assign w8701 = w105 & pi673;
assign w8702 = w66 & ~w42;
assign w8703 = w45 & ~w82;
assign w8704 = w66 & pi195;
assign w8705 = w45 & pi164;
assign w8706 = w149 & pi165;
assign w8707 = w66 & pi132;
assign w8708 = w66 & pi192;
assign w8709 = w45 & pi110;
assign w8710 = w66 & pi165;
assign w8711 = w45 & pi132;
assign w8712 = w149 & pi110;
assign w8713 = w200 & ~w109;
assign w8714 = ~w109 & ~w203;
assign w8715 = w26 & pi133;
assign w8716 = ~w26 & ~pi909;
assign w8717 = w26 & pi045;
assign w8718 = ~w26 & pi877;
assign w8719 = ~w26 & ~pi845;
assign w8720 = w26 & ~pi012;
assign w8721 = pi668 & ~pi000;
assign w8722 = w29 & ~w227;
assign w8723 = w95 & ~w109;
assign w8724 = w149 & pi192;
assign w8725 = w45 & pi165;
assign w8726 = w26 & pi134;
assign w8727 = ~w26 & ~pi910;
assign w8728 = ~w26 & ~pi878;
assign w8729 = w26 & ~pi044;
assign w8730 = pi668 & ~pi001;
assign w8731 = w26 & pi013;
assign w8732 = ~w26 & pi846;
assign w8733 = ~w26 & ~pi814;
assign w8734 = w26 & ~pi001;
assign w8735 = ~w1 & ~w268;
assign w8736 = w26 & pi048;
assign w8737 = ~w26 & pi879;
assign w8738 = ~w26 & ~pi847;
assign w8739 = w26 & ~pi014;
assign w8740 = ~w200 & w109;
assign w8741 = ~w26 & ~pi911;
assign w8742 = w26 & ~pi167;
assign w8743 = ~w308 & ~w311;
assign w8744 = w308 & w311;
assign w8745 = w26 & ~pi002;
assign w8746 = ~w26 & ~pi815;
assign w8747 = ~w291 & w1;
assign w8748 = pi668 & ~pi002;
assign w8749 = w319 & ~w325;
assign w8750 = ~w324 & w326;
assign w8751 = w26 & pi049;
assign w8752 = ~w26 & pi880;
assign w8753 = ~w26 & ~pi848;
assign w8754 = w26 & ~pi015;
assign w8755 = ~w26 & ~pi912;
assign w8756 = w26 & ~pi166;
assign w8757 = ~w352 & ~w355;
assign w8758 = w352 & w355;
assign w8759 = ~w338 & w1;
assign w8760 = pi668 & pi003;
assign w8761 = w26 & ~pi003;
assign w8762 = ~w26 & ~pi816;
assign w8763 = w364 & ~w362;
assign w8764 = ~w361 & w367;
assign w8765 = pi668 & pi004;
assign w8766 = ~w26 & pi817;
assign w8767 = w26 & pi004;
assign w8768 = w376 & ~w374;
assign w8769 = w26 & pi155;
assign w8770 = ~w26 & ~pi913;
assign w8771 = w26 & pi057;
assign w8772 = ~w26 & pi881;
assign w8773 = ~w26 & ~pi849;
assign w8774 = w26 & ~pi016;
assign w8775 = pi668 & ~pi004;
assign w8776 = w376 & ~w414;
assign w8777 = ~w3 & ~w23;
assign w8778 = w26 & pi199;
assign w8779 = ~w26 & pi832;
assign w8780 = ~pi668 & pi824;
assign w8781 = pi668 & pi816;
assign w8782 = pi668 & pi808;
assign w8783 = ~w26 & ~w430;
assign w8784 = pi668 & pi209;
assign w8785 = ~pi668 & pi221;
assign w8786 = w26 & ~w436;
assign w8787 = ~w431 & ~w437;
assign w8788 = ~pi673 & ~pi280;
assign w8789 = pi673 & ~pi601;
assign w8790 = w536 & w540;
assign w8791 = ~pi673 & ~pi398;
assign w8792 = pi673 & ~pi640;
assign w8793 = w105 & ~w546;
assign w8794 = ~pi568 & pi642;
assign w8795 = ~pi568 & pi300;
assign w8796 = w26 & pi196;
assign w8797 = ~w26 & pi830;
assign w8798 = ~pi668 & pi222;
assign w8799 = pi668 & pi001;
assign w8800 = pi668 & pi207;
assign w8801 = w26 & w629;
assign w8802 = pi668 & pi814;
assign w8803 = pi668 & pi806;
assign w8804 = ~pi668 & pi822;
assign w8805 = ~w26 & w635;
assign w8806 = ~pi568 & pi324;
assign w8807 = ~pi568 & pi653;
assign w8808 = w25 & pi827;
assign w8809 = ~w25 & pi202;
assign w8810 = pi668 & pi803;
assign w8811 = pi668 & pi811;
assign w8812 = ~pi668 & pi819;
assign w8813 = ~w26 & w723;
assign w8814 = ~pi668 & pi216;
assign w8815 = pi668 & pi011;
assign w8816 = pi668 & pi211;
assign w8817 = w26 & w729;
assign w8818 = ~pi568 & pi660;
assign w8819 = ~pi568 & pi281;
assign w8820 = w26 & pi201;
assign w8821 = ~w26 & pi833;
assign w8822 = pi668 & pi213;
assign w8823 = ~pi668 & pi212;
assign w8824 = w26 & w817;
assign w8825 = pi668 & pi817;
assign w8826 = pi668 & pi809;
assign w8827 = ~pi668 & pi825;
assign w8828 = ~w26 & w823;
assign w8829 = w826 & ~w109;
assign w8830 = pi673 & ~pi594;
assign w8831 = ~pi673 & ~pi269;
assign w8832 = w536 & w859;
assign w8833 = w26 & pi010;
assign w8834 = ~w26 & pi812;
assign w8835 = w25 & pi828;
assign w8836 = ~w25 & pi203;
assign w8837 = ~pi668 & pi219;
assign w8838 = pi668 & pi205;
assign w8839 = w26 & w915;
assign w8840 = ~pi668 & pi820;
assign w8841 = pi668 & pi804;
assign w8842 = ~w26 & w919;
assign w8843 = ~w638 & w109;
assign w8844 = w26 & pi198;
assign w8845 = ~w26 & pi831;
assign w8846 = pi668 & pi807;
assign w8847 = pi668 & pi815;
assign w8848 = ~pi668 & pi823;
assign w8849 = ~w26 & ~w937;
assign w8850 = pi668 & pi208;
assign w8851 = pi668 & pi002;
assign w8852 = ~pi668 & pi220;
assign w8853 = w26 & ~w943;
assign w8854 = ~w938 & ~w944;
assign w8855 = ~pi673 & ~pi277;
assign w8856 = pi673 & ~pi615;
assign w8857 = w536 & w1010;
assign w8858 = w926 & w1016;
assign w8859 = ~w926 & ~w639;
assign w8860 = w109 & ~w1024;
assign w8861 = ~pi568 & pi647;
assign w8862 = ~pi568 & pi322;
assign w8863 = w26 & pi200;
assign w8864 = ~w26 & pi826;
assign w8865 = ~pi668 & pi217;
assign w8866 = pi668 & pi009;
assign w8867 = pi668 & pi210;
assign w8868 = w26 & w1106;
assign w8869 = pi668 & pi802;
assign w8870 = pi668 & pi810;
assign w8871 = ~pi668 & pi818;
assign w8872 = ~w26 & w1112;
assign w8873 = w26 & pi197;
assign w8874 = ~w26 & pi829;
assign w8875 = pi668 & pi805;
assign w8876 = pi668 & pi813;
assign w8877 = ~pi668 & pi821;
assign w8878 = ~w26 & ~w1129;
assign w8879 = pi668 & pi206;
assign w8880 = ~pi668 & pi218;
assign w8881 = w26 & ~w1135;
assign w8882 = ~w1130 & ~w1136;
assign w8883 = pi673 & ~pi624;
assign w8884 = ~pi673 & ~pi272;
assign w8885 = w536 & w1186;
assign w8886 = ~w1138 & ~w109;
assign w8887 = ~w1120 & ~w1209;
assign w8888 = ~w731 & ~w109;
assign w8889 = ~w1115 & w109;
assign w8890 = w1115 & w109;
assign w8891 = w638 & ~w109;
assign w8892 = w1138 & w109;
assign w8893 = ~w1138 & w109;
assign w8894 = ~w1115 & ~w109;
assign w8895 = w926 & w1272;
assign w8896 = ~w926 & w1014;
assign w8897 = w1213 & ~w1250;
assign w8898 = ~w1235 & ~w1321;
assign w8899 = ~w1251 & ~w1330;
assign w8900 = w1275 & ~w1276;
assign w8901 = ~w109 & ~w303;
assign w8902 = w26 & pi017;
assign w8903 = ~w26 & pi842;
assign w8904 = w26 & pi056;
assign w8905 = ~w26 & pi874;
assign w8906 = w26 & pi136;
assign w8907 = ~w26 & ~pi906;
assign w8908 = w26 & ~pi009;
assign w8909 = ~w26 & ~pi810;
assign w8910 = w1374 & w1;
assign w8911 = w1379 & ~w1385;
assign w8912 = ~w1384 & w1386;
assign w8913 = ~w1392 & ~w171;
assign w8914 = w26 & pi188;
assign w8915 = ~w26 & ~pi908;
assign w8916 = w26 & pi046;
assign w8917 = ~w26 & ~pi876;
assign w8918 = ~w26 & ~pi844;
assign w8919 = w26 & ~pi042;
assign w8920 = ~w1390 & w1412;
assign w8921 = pi668 & ~pi010;
assign w8922 = ~w1 & ~w1416;
assign w8923 = pi668 & ~pi011;
assign w8924 = ~w26 & pi811;
assign w8925 = w26 & pi011;
assign w8926 = w1427 & ~w1425;
assign w8927 = w26 & pi176;
assign w8928 = ~w26 & ~pi907;
assign w8929 = w26 & pi043;
assign w8930 = ~w26 & pi843;
assign w8931 = w26 & pi047;
assign w8932 = ~w26 & ~pi875;
assign w8933 = w109 & ~w1445;
assign w8934 = ~w1444 & ~w1445;
assign w8935 = ~w1444 & w8933;
assign w8936 = w1451 & ~w1429;
assign w8937 = w1427 & ~w1454;
assign w8938 = ~pi568 & pi018;
assign w8939 = pi568 & pi022;
assign w8940 = ~w1469 & w1467;
assign w8941 = ~w1464 & ~pi018;
assign w8942 = ~w308 & w1472;
assign w8943 = ~w535 & pi018;
assign w8944 = ~w535 & ~w8941;
assign w8945 = ~pi568 & pi019;
assign w8946 = pi568 & pi023;
assign w8947 = ~w1464 & ~pi019;
assign w8948 = ~w352 & w1472;
assign w8949 = ~w535 & pi019;
assign w8950 = ~w535 & ~w8947;
assign w8951 = ~pi568 & pi020;
assign w8952 = pi568 & pi024;
assign w8953 = ~w1469 & ~w1467;
assign w8954 = ~w1487 & ~pi020;
assign w8955 = ~w308 & w1489;
assign w8956 = ~w535 & pi020;
assign w8957 = ~w535 & ~w8954;
assign w8958 = ~pi568 & pi021;
assign w8959 = pi568 & pi025;
assign w8960 = ~w1487 & ~pi021;
assign w8961 = ~w352 & w1489;
assign w8962 = ~w535 & pi021;
assign w8963 = ~w535 & ~w8960;
assign w8964 = ~pi568 & pi022;
assign w8965 = pi568 & pi018;
assign w8966 = ~w1487 & ~pi022;
assign w8967 = ~w308 & w1504;
assign w8968 = ~w535 & pi022;
assign w8969 = ~w535 & ~w8966;
assign w8970 = ~pi568 & pi023;
assign w8971 = pi568 & pi019;
assign w8972 = ~w1487 & ~pi023;
assign w8973 = ~w352 & w1504;
assign w8974 = ~w535 & pi023;
assign w8975 = ~w535 & ~w8972;
assign w8976 = ~pi568 & pi024;
assign w8977 = pi568 & pi020;
assign w8978 = ~w1464 & ~pi024;
assign w8979 = ~w308 & w1519;
assign w8980 = ~w535 & pi024;
assign w8981 = ~w535 & ~w8978;
assign w8982 = ~pi568 & pi025;
assign w8983 = pi568 & pi021;
assign w8984 = ~w1464 & ~pi025;
assign w8985 = ~w352 & w1519;
assign w8986 = ~w535 & pi025;
assign w8987 = ~w535 & ~w8984;
assign w8988 = ~pi568 & pi026;
assign w8989 = pi568 & ~w1533;
assign w8990 = pi673 & w1534;
assign w8991 = ~w1537 & ~pi026;
assign w8992 = ~w352 & w1538;
assign w8993 = ~w1532 & ~w1534;
assign w8994 = ~w1532 & ~w8990;
assign w8995 = ~pi568 & pi027;
assign w8996 = pi568 & ~w1546;
assign w8997 = pi673 & w1547;
assign w8998 = ~w308 & w1538;
assign w8999 = pi027 & ~w535;
assign w9000 = ~w1545 & ~w1547;
assign w9001 = ~w1545 & ~w8997;
assign w9002 = ~pi568 & pi028;
assign w9003 = ~pi566 & ~pi568;
assign w9004 = ~w1560 & ~pi028;
assign w9005 = ~w352 & w1561;
assign w9006 = ~pi568 & pi029;
assign w9007 = ~w1560 & ~pi029;
assign w9008 = ~w308 & w1561;
assign w9009 = ~w9008 & w1574;
assign w9010 = ~pi568 & pi030;
assign w9011 = pi566 & ~pi568;
assign w9012 = ~pi563 & w1585;
assign w9013 = ~w9012 & ~pi030;
assign w9014 = ~w308 & w1586;
assign w9015 = ~w9014 & w1588;
assign w9016 = ~pi568 & pi031;
assign w9017 = ~w9012 & ~pi031;
assign w9018 = ~w352 & w1586;
assign w9019 = ~pi568 & pi032;
assign w9020 = ~w308 & w1604;
assign w9021 = pi032 & ~w535;
assign w9022 = ~w308 & pi673;
assign w9023 = pi568 & ~w1608;
assign w9024 = ~w9022 & w1609;
assign w9025 = ~pi568 & pi033;
assign w9026 = ~w352 & w1604;
assign w9027 = pi033 & ~w535;
assign w9028 = ~w352 & pi673;
assign w9029 = pi568 & ~w1616;
assign w9030 = ~w1615 & ~w1613;
assign w9031 = ~pi568 & pi034;
assign w9032 = ~pi563 & w1560;
assign w9033 = ~w308 & w1627;
assign w9034 = pi034 & ~w535;
assign w9035 = ~pi568 & pi035;
assign w9036 = ~w352 & w1627;
assign w9037 = pi035 & ~w535;
assign w9038 = ~pi568 & pi036;
assign w9039 = ~pi568 & pi037;
assign w9040 = ~pi568 & pi038;
assign w9041 = ~w1537 & ~pi038;
assign w9042 = ~w352 & w1660;
assign w9043 = ~pi568 & pi039;
assign w9044 = ~w1537 & ~pi039;
assign w9045 = ~w308 & w1660;
assign w9046 = ~w9045 & w1673;
assign w9047 = ~pi568 & pi040;
assign w9048 = ~w1682 & ~pi040;
assign w9049 = ~w308 & w1683;
assign w9050 = ~w9049 & w1685;
assign w9051 = ~pi568 & pi041;
assign w9052 = ~w1682 & ~pi041;
assign w9053 = ~w352 & w1683;
assign w9054 = pi668 & ~pi046;
assign w9055 = ~w1 & ~w1707;
assign w9056 = w1 & w1403;
assign w9057 = w1712 & ~w1445;
assign w9058 = w1712 & w8933;
assign w9059 = w1714 & w1445;
assign w9060 = w1714 & ~w8933;
assign w9061 = pi668 & pi047;
assign w9062 = ~w1 & ~w1718;
assign w9063 = w308 & w1728;
assign w9064 = ~w1464 & pi050;
assign w9065 = w352 & w1728;
assign w9066 = ~w1464 & pi051;
assign w9067 = ~w441 & w1487;
assign w9068 = w308 & w1735;
assign w9069 = ~w441 & w1464;
assign w9070 = w352 & w1739;
assign w9071 = w352 & w1735;
assign w9072 = w308 & w1739;
assign w9073 = ~pi568 & pi058;
assign w9074 = pi568 & pi059;
assign w9075 = ~w1464 & ~pi058;
assign w9076 = ~w535 & pi058;
assign w9077 = ~w535 & ~w9075;
assign w9078 = ~pi568 & pi059;
assign w9079 = pi568 & pi058;
assign w9080 = ~w1487 & ~pi059;
assign w9081 = ~w535 & pi059;
assign w9082 = ~w535 & ~w9080;
assign w9083 = ~pi568 & pi060;
assign w9084 = pi568 & pi061;
assign w9085 = ~w1464 & ~pi060;
assign w9086 = ~w535 & pi060;
assign w9087 = ~w535 & ~w9085;
assign w9088 = ~pi568 & pi061;
assign w9089 = pi568 & pi060;
assign w9090 = ~w1487 & ~pi061;
assign w9091 = ~w535 & pi061;
assign w9092 = ~w535 & ~w9090;
assign w9093 = ~pi568 & pi062;
assign w9094 = ~pi568 & pi063;
assign w9095 = ~w1560 & ~pi063;
assign w9096 = ~w1561 & w1798;
assign w9097 = ~pi568 & pi064;
assign w9098 = ~w9012 & ~pi064;
assign w9099 = ~w1586 & w1808;
assign w9100 = ~pi568 & pi065;
assign w9101 = ~w1537 & ~pi065;
assign w9102 = ~w1660 & w1818;
assign w9103 = ~pi568 & pi066;
assign w9104 = ~w1682 & ~pi066;
assign w9105 = ~w1683 & w1828;
assign w9106 = ~w1537 & ~pi067;
assign w9107 = ~w1538 & w1833;
assign w9108 = pi568 & ~w1836;
assign w9109 = pi673 & w1837;
assign w9110 = ~pi568 & pi068;
assign w9111 = pi068 & ~w535;
assign w9112 = w308 & w1851;
assign w9113 = ~w1487 & pi069;
assign w9114 = w352 & w1851;
assign w9115 = ~w1487 & pi070;
assign w9116 = w308 & w427;
assign w9117 = ~pi668 & ~pi071;
assign w9118 = w352 & w427;
assign w9119 = ~pi668 & ~pi072;
assign w9120 = ~pi568 & pi073;
assign w9121 = pi568 & pi080;
assign w9122 = ~w1464 & ~pi073;
assign w9123 = ~w535 & pi073;
assign w9124 = ~w535 & ~w9122;
assign w9125 = ~pi568 & pi074;
assign w9126 = pi568 & pi079;
assign w9127 = ~w1464 & ~pi074;
assign w9128 = ~w535 & pi074;
assign w9129 = ~w535 & ~w9127;
assign w9130 = ~pi568 & pi075;
assign w9131 = pi568 & pi081;
assign w9132 = ~w1464 & ~pi075;
assign w9133 = w348 & ~w384;
assign w9134 = ~w348 & w384;
assign w9135 = ~w535 & pi075;
assign w9136 = ~w535 & ~w9132;
assign w9137 = ~pi568 & pi076;
assign w9138 = pi568 & pi082;
assign w9139 = ~w1487 & ~pi076;
assign w9140 = ~w535 & pi076;
assign w9141 = ~w535 & ~w9139;
assign w9142 = ~pi568 & pi077;
assign w9143 = pi568 & pi083;
assign w9144 = ~w1487 & ~pi077;
assign w9145 = ~w535 & pi077;
assign w9146 = ~w535 & ~w9144;
assign w9147 = ~pi568 & pi078;
assign w9148 = pi568 & pi084;
assign w9149 = ~w1487 & ~pi078;
assign w9150 = ~w535 & pi078;
assign w9151 = ~w535 & ~w9149;
assign w9152 = ~pi568 & pi079;
assign w9153 = pi568 & pi074;
assign w9154 = ~w1487 & ~pi079;
assign w9155 = ~w535 & pi079;
assign w9156 = ~w535 & ~w9154;
assign w9157 = ~pi568 & pi080;
assign w9158 = pi568 & pi073;
assign w9159 = ~w1487 & ~pi080;
assign w9160 = ~w535 & pi080;
assign w9161 = ~w535 & ~w9159;
assign w9162 = ~pi568 & pi081;
assign w9163 = pi568 & pi075;
assign w9164 = ~w1487 & ~pi081;
assign w9165 = ~w535 & pi081;
assign w9166 = ~w535 & ~w9164;
assign w9167 = ~pi568 & pi082;
assign w9168 = pi568 & pi076;
assign w9169 = ~w1464 & ~pi082;
assign w9170 = ~w535 & pi082;
assign w9171 = ~w535 & ~w9169;
assign w9172 = ~pi568 & pi083;
assign w9173 = pi568 & pi077;
assign w9174 = ~w1464 & ~pi083;
assign w9175 = ~w535 & pi083;
assign w9176 = ~w535 & ~w9174;
assign w9177 = ~pi568 & pi084;
assign w9178 = pi568 & pi078;
assign w9179 = ~w1464 & ~pi084;
assign w9180 = ~w535 & pi084;
assign w9181 = ~w535 & ~w9179;
assign w9182 = ~w1537 & ~pi085;
assign w9183 = ~w1538 & w1952;
assign w9184 = pi568 & ~w1955;
assign w9185 = pi673 & w1956;
assign w9186 = ~pi568 & pi086;
assign w9187 = ~w1560 & ~pi086;
assign w9188 = ~w1561 & w1966;
assign w9189 = ~pi568 & pi087;
assign w9190 = ~w1560 & ~pi087;
assign w9191 = ~w1561 & w1976;
assign w9192 = ~pi568 & pi088;
assign w9193 = ~w1560 & ~pi088;
assign w9194 = ~w1561 & w1986;
assign w9195 = ~pi568 & pi089;
assign w9196 = ~w9012 & ~pi089;
assign w9197 = ~w1586 & w1996;
assign w9198 = ~pi568 & pi090;
assign w9199 = ~w9012 & ~pi090;
assign w9200 = ~w1586 & w2006;
assign w9201 = ~pi568 & pi091;
assign w9202 = ~w9012 & ~pi091;
assign w9203 = ~w1586 & w2016;
assign w9204 = ~pi568 & pi092;
assign w9205 = pi568 & ~w2021;
assign w9206 = ~pi673 & w2022;
assign w9207 = pi092 & ~w535;
assign w9208 = ~w2020 & ~w2022;
assign w9209 = ~w2020 & ~w9206;
assign w9210 = ~pi568 & pi093;
assign w9211 = ~pi568 & pi094;
assign w9212 = pi094 & ~w535;
assign w9213 = ~pi568 & pi095;
assign w9214 = pi095 & ~w535;
assign w9215 = ~pi568 & pi096;
assign w9216 = pi096 & ~w535;
assign w9217 = ~pi568 & pi097;
assign w9218 = pi097 & ~w535;
assign w9219 = pi568 & ~w2068;
assign w9220 = ~pi673 & w2069;
assign w9221 = ~pi568 & pi098;
assign w9222 = ~w1537 & ~pi098;
assign w9223 = ~w1660 & w2079;
assign w9224 = ~pi568 & pi099;
assign w9225 = ~w1537 & ~pi099;
assign w9226 = ~w1660 & w2089;
assign w9227 = ~pi568 & pi100;
assign w9228 = ~pi568 & pi101;
assign w9229 = ~pi568 & pi102;
assign w9230 = ~w1537 & ~pi102;
assign w9231 = ~w1660 & w2111;
assign w9232 = ~pi568 & pi103;
assign w9233 = ~w1682 & ~pi103;
assign w9234 = ~w1683 & w2121;
assign w9235 = ~pi568 & pi104;
assign w9236 = ~w1682 & ~pi104;
assign w9237 = ~w1683 & w2131;
assign w9238 = ~pi568 & pi105;
assign w9239 = ~w1682 & ~pi105;
assign w9240 = ~w1683 & w2141;
assign w9241 = ~w1464 & pi106;
assign w9242 = ~w1487 & pi108;
assign w9243 = w352 & w102;
assign w9244 = ~pi668 & ~pi111;
assign w9245 = ~pi568 & pi112;
assign w9246 = ~w1537 & ~pi112;
assign w9247 = ~w1538 & w2164;
assign w9248 = pi568 & ~w2166;
assign w9249 = pi673 & w2167;
assign w9250 = w352 & w424;
assign w9251 = w308 & w424;
assign w9252 = pi668 & ~pi114;
assign w9253 = ~pi568 & pi115;
assign w9254 = pi115 & ~w535;
assign w9255 = pi568 & ~w2181;
assign w9256 = ~pi673 & w2182;
assign w9257 = pi568 & ~w2186;
assign w9258 = ~pi673 & w2187;
assign w9259 = pi116 & ~w535;
assign w9260 = ~w2188 & ~w2187;
assign w9261 = ~w2188 & ~w9258;
assign w9262 = w308 & w102;
assign w9263 = ~pi568 & pi118;
assign w9264 = ~w1537 & ~pi118;
assign w9265 = ~w1538 & w2199;
assign w9266 = pi568 & ~w2201;
assign w9267 = pi673 & w2202;
assign w9268 = ~w1464 & pi119;
assign w9269 = ~w1464 & pi120;
assign w9270 = ~w1464 & pi121;
assign w9271 = ~w1487 & pi125;
assign w9272 = ~w1487 & pi126;
assign w9273 = ~w1487 & pi127;
assign w9274 = ~pi668 & pi131;
assign w9275 = pi668 & pi133;
assign w9276 = pi668 & pi134;
assign w9277 = ~pi668 & pi135;
assign w9278 = pi668 & ~pi136;
assign w9279 = ~pi668 & pi137;
assign w9280 = ~pi668 & pi138;
assign w9281 = ~w1464 & ~pi139;
assign w9282 = ~w535 & pi139;
assign w9283 = ~w535 & ~w9281;
assign w9284 = ~pi568 & pi139;
assign w9285 = pi568 & pi142;
assign w9286 = ~w1487 & ~pi140;
assign w9287 = ~w535 & pi140;
assign w9288 = ~w535 & ~w9286;
assign w9289 = ~pi568 & pi140;
assign w9290 = pi568 & pi141;
assign w9291 = ~w1464 & ~pi141;
assign w9292 = ~w535 & pi141;
assign w9293 = ~w535 & ~w9291;
assign w9294 = ~pi568 & pi141;
assign w9295 = pi568 & pi140;
assign w9296 = ~w1487 & ~pi142;
assign w9297 = ~w535 & pi142;
assign w9298 = ~w535 & ~w9296;
assign w9299 = ~pi568 & pi142;
assign w9300 = pi568 & pi139;
assign w9301 = ~w1560 & ~pi143;
assign w9302 = ~w1561 & w2292;
assign w9303 = ~pi668 & pi144;
assign w9304 = pi668 & pi145;
assign w9305 = pi668 & pi146;
assign w9306 = ~w9012 & ~pi147;
assign w9307 = ~w1586 & w2311;
assign w9308 = ~pi568 & pi148;
assign w9309 = pi149 & ~w535;
assign w9310 = ~pi568 & pi149;
assign w9311 = ~w1537 & ~pi150;
assign w9312 = ~w1660 & w2337;
assign w9313 = ~w1682 & ~pi151;
assign w9314 = ~w1683 & w2347;
assign w9315 = ~w1537 & ~pi152;
assign w9316 = ~w1538 & w2357;
assign w9317 = ~w164 & ~pi673;
assign w9318 = pi568 & ~w2360;
assign w9319 = ~w2364 & ~w2359;
assign w9320 = pi668 & pi153;
assign w9321 = ~pi668 & pi154;
assign w9322 = pi668 & pi155;
assign w9323 = ~pi668 & pi156;
assign w9324 = ~pi668 & pi157;
assign w9325 = pi568 & pi673;
assign w9326 = ~pi568 & pi158;
assign w9327 = pi568 & w2386;
assign w9328 = ~w2385 & ~w2387;
assign w9329 = pi668 & pi159;
assign w9330 = ~w1464 & ~pi160;
assign w9331 = ~w1487 & ~pi162;
assign w9332 = ~pi568 & pi168;
assign w9333 = pi568 & pi169;
assign w9334 = ~w1464 & ~pi168;
assign w9335 = w1472 & ~w1445;
assign w9336 = w1472 & w8933;
assign w9337 = ~w535 & pi168;
assign w9338 = ~w535 & ~w9334;
assign w9339 = ~pi568 & pi169;
assign w9340 = pi568 & pi168;
assign w9341 = ~w1487 & ~pi169;
assign w9342 = w1504 & ~w1445;
assign w9343 = w1504 & w8933;
assign w9344 = ~w535 & pi169;
assign w9345 = ~w535 & ~w9341;
assign w9346 = ~pi568 & pi170;
assign w9347 = pi568 & pi171;
assign w9348 = ~w1464 & ~pi170;
assign w9349 = w1519 & ~w1445;
assign w9350 = w1519 & w8933;
assign w9351 = ~w535 & pi170;
assign w9352 = ~w535 & ~w9348;
assign w9353 = ~pi568 & pi171;
assign w9354 = pi568 & pi170;
assign w9355 = ~w1487 & ~pi171;
assign w9356 = w1489 & ~w1445;
assign w9357 = w1489 & w8933;
assign w9358 = ~w535 & pi171;
assign w9359 = ~w535 & ~w9355;
assign w9360 = ~pi568 & pi172;
assign w9361 = ~w9012 & ~pi172;
assign w9362 = w1586 & ~w1445;
assign w9363 = w1586 & w8933;
assign w9364 = w2442 & ~w9362;
assign w9365 = w2442 & ~w9363;
assign w9366 = ~pi568 & pi173;
assign w9367 = ~pi568 & pi174;
assign w9368 = ~w1537 & ~pi174;
assign w9369 = w1660 & ~w1445;
assign w9370 = w1660 & w8933;
assign w9371 = w2458 & ~w9369;
assign w9372 = w2458 & ~w9370;
assign w9373 = ~pi568 & pi175;
assign w9374 = pi568 & ~w2463;
assign w9375 = pi673 & w2464;
assign w9376 = w1538 & ~w1445;
assign w9377 = w1538 & w8933;
assign w9378 = pi175 & ~w535;
assign w9379 = ~w2462 & ~w2464;
assign w9380 = ~w2462 & ~w9375;
assign w9381 = pi668 & pi176;
assign w9382 = ~pi668 & pi177;
assign w9383 = ~pi568 & pi179;
assign w9384 = ~w1682 & ~pi179;
assign w9385 = w1683 & ~w1445;
assign w9386 = w1683 & w8933;
assign w9387 = w2481 & ~w9385;
assign w9388 = w2481 & ~w9386;
assign w9389 = ~pi568 & pi180;
assign w9390 = w1627 & ~w1445;
assign w9391 = w1627 & w8933;
assign w9392 = pi180 & ~w535;
assign w9393 = ~pi568 & pi181;
assign w9394 = ~w1560 & ~pi181;
assign w9395 = w1561 & ~w1445;
assign w9396 = w1561 & w8933;
assign w9397 = w2501 & ~w9395;
assign w9398 = w2501 & ~w9396;
assign w9399 = ~pi568 & pi182;
assign w9400 = pi673 & ~w1445;
assign w9401 = pi673 & w8933;
assign w9402 = pi568 & ~w2506;
assign w9403 = w2507 & ~w9400;
assign w9404 = w2507 & ~w9401;
assign w9405 = w1604 & ~w1445;
assign w9406 = w1604 & w8933;
assign w9407 = pi182 & ~w535;
assign w9408 = w1851 & w1445;
assign w9409 = w1851 & ~w8933;
assign w9410 = ~w1487 & ~pi183;
assign w9411 = w1739 & w1445;
assign w9412 = w1739 & ~w8933;
assign w9413 = w1735 & w1445;
assign w9414 = w1735 & ~w8933;
assign w9415 = ~pi668 & pi186;
assign w9416 = w1728 & w1445;
assign w9417 = w1728 & ~w8933;
assign w9418 = ~w1464 & ~pi187;
assign w9419 = w1 & ~w1397;
assign w9420 = pi668 & pi188;
assign w9421 = ~w2530 & ~w2531;
assign w9422 = pi668 & pi189;
assign w9423 = w427 & w1445;
assign w9424 = w427 & ~w8933;
assign w9425 = ~pi668 & ~pi191;
assign w9426 = w102 & w1445;
assign w9427 = w102 & ~w8933;
assign w9428 = ~pi668 & ~pi193;
assign w9429 = w424 & w1445;
assign w9430 = w424 & ~w8933;
assign w9431 = pi668 & ~pi194;
assign w9432 = pi668 & pi196;
assign w9433 = pi550 & pi552;
assign w9434 = ~pi665 & ~w2552;
assign w9435 = pi551 & ~w2552;
assign w9436 = pi551 & w9434;
assign w9437 = ~pi550 & ~pi552;
assign w9438 = w2562 & ~w2552;
assign w9439 = w2562 & w9434;
assign w9440 = pi665 & ~w2568;
assign w9441 = ~pi665 & ~pi390;
assign w9442 = w2550 & ~pi559;
assign w9443 = ~pi665 & ~pi559;
assign w9444 = w2578 & ~pi559;
assign w9445 = w2578 & w9443;
assign w9446 = ~w2580 & w2564;
assign w9447 = ~w26 & ~pi926;
assign w9448 = w26 & ~pi288;
assign w9449 = w26 & pi228;
assign w9450 = ~w26 & ~pi894;
assign w9451 = w26 & pi204;
assign w9452 = ~w26 & ~pi862;
assign w9453 = w623 & w1;
assign w9454 = w26 & pi238;
assign w9455 = ~w26 & pi893;
assign w9456 = ~w26 & ~pi925;
assign w9457 = w26 & ~pi333;
assign w9458 = w26 & pi215;
assign w9459 = ~w26 & ~pi861;
assign w9460 = pi668 & pi197;
assign w9461 = pi668 & ~pi198;
assign w9462 = w26 & pi332;
assign w9463 = ~w26 & pi927;
assign w9464 = w2582 & w2649;
assign w9465 = ~w2582 & ~w2649;
assign w9466 = w26 & pi239;
assign w9467 = ~w26 & ~pi895;
assign w9468 = w26 & pi214;
assign w9469 = ~w26 & ~pi863;
assign w9470 = w931 & w1;
assign w9471 = pi668 & pi199;
assign w9472 = ~w2574 & ~w2564;
assign w9473 = ~w26 & ~pi928;
assign w9474 = w26 & ~pi394;
assign w9475 = ~w26 & ~pi896;
assign w9476 = w26 & ~pi249;
assign w9477 = w26 & pi226;
assign w9478 = ~w26 & ~pi864;
assign w9479 = w1 & w422;
assign w9480 = ~w1 & w2695;
assign w9481 = ~w9479 & ~w2669;
assign w9482 = pi668 & pi200;
assign w9483 = w2580 & w2564;
assign w9484 = ~w26 & ~pi922;
assign w9485 = w26 & ~pi387;
assign w9486 = ~w26 & ~pi890;
assign w9487 = w26 & ~pi248;
assign w9488 = w26 & pi227;
assign w9489 = ~w26 & ~pi858;
assign w9490 = w1100 & w1;
assign w9491 = pi668 & pi201;
assign w9492 = ~w26 & ~pi929;
assign w9493 = w26 & ~pi389;
assign w9494 = ~w26 & ~pi897;
assign w9495 = w26 & ~pi250;
assign w9496 = w26 & pi225;
assign w9497 = ~w26 & ~pi865;
assign w9498 = w1 & w811;
assign w9499 = ~w1 & w2750;
assign w9500 = ~w9498 & ~w2726;
assign w9501 = pi668 & ~pi202;
assign w9502 = w26 & pi251;
assign w9503 = ~w26 & pi891;
assign w9504 = w2583 & pi193;
assign w9505 = ~w2583 & ~pi193;
assign w9506 = ~w26 & ~pi923;
assign w9507 = w26 & ~pi388;
assign w9508 = w26 & pi223;
assign w9509 = ~w26 & ~pi859;
assign w9510 = ~w1 & ~w2754;
assign w9511 = ~w1 & w2778;
assign w9512 = pi668 & ~pi203;
assign w9513 = w2671 & w2564;
assign w9514 = w26 & ~pi396;
assign w9515 = w2785 & pi186;
assign w9516 = ~w2785 & ~pi186;
assign w9517 = w26 & pi247;
assign w9518 = ~w26 & ~pi892;
assign w9519 = w26 & pi224;
assign w9520 = ~w26 & ~pi860;
assign w9521 = ~w1 & ~w2782;
assign w9522 = w1 & ~w911;
assign w9523 = pi668 & pi204;
assign w9524 = pi668 & ~pi205;
assign w9525 = ~w26 & ~pi900;
assign w9526 = w26 & ~pi414;
assign w9527 = ~w26 & ~pi868;
assign w9528 = w26 & ~pi292;
assign w9529 = w26 & pi231;
assign w9530 = ~w26 & ~pi836;
assign w9531 = w26 & pi205;
assign w9532 = ~w26 & pi804;
assign w9533 = w2833 & w1;
assign w9534 = pi668 & ~pi206;
assign w9535 = ~w26 & ~pi901;
assign w9536 = w26 & ~pi437;
assign w9537 = ~w26 & ~pi869;
assign w9538 = w26 & ~pi291;
assign w9539 = w26 & pi232;
assign w9540 = ~w26 & ~pi837;
assign w9541 = w26 & pi206;
assign w9542 = ~w26 & pi805;
assign w9543 = w2859 & w1;
assign w9544 = pi668 & ~pi207;
assign w9545 = ~w26 & ~pi902;
assign w9546 = w26 & ~pi415;
assign one = 1;
assign po000 = pi564;// level 0
assign po001 = pi266;// level 0
assign po002 = pi303;// level 0
assign po003 = pi312;// level 0
assign po004 = pi270;// level 0
assign po005 = pi326;// level 0
assign po006 = pi297;// level 0
assign po007 = pi256;// level 0
assign po008 = pi308;// level 0
assign po009 = pi264;// level 0
assign po010 = pi323;// level 0
assign po011 = pi282;// level 0
assign po012 = pi319;// level 0
assign po013 = pi327;// level 0
assign po014 = pi283;// level 0
assign po015 = pi329;// level 0
assign po016 = pi331;// level 0
assign po017 = pi400;// level 0
assign po018 = pi386;// level 0
assign po019 = pi407;// level 0
assign po020 = pi404;// level 0
assign po021 = pi355;// level 0
assign po022 = pi358;// level 0
assign po023 = pi360;// level 0
assign po024 = pi363;// level 0
assign po025 = pi306;// level 0
assign po026 = pi258;// level 0
assign po027 = pi262;// level 0
assign po028 = pi340;// level 0
assign po029 = pi309;// level 0
assign po030 = pi263;// level 0
assign po031 = pi311;// level 0
assign po032 = pi313;// level 0
assign po033 = pi374;// level 0
assign po034 = pi343;// level 0
assign po035 = pi317;// level 0
assign po036 = pi346;// level 0
assign po037 = pi378;// level 0
assign po038 = pi380;// level 0
assign po039 = pi381;// level 0
assign po040 = pi382;// level 0
assign po041 = pi299;// level 0
assign po042 = pi271;// level 0
assign po043 = pi273;// level 0
assign po044 = pi274;// level 0
assign po045 = pi275;// level 0
assign po046 = pi325;// level 0
assign po047 = pi278;// level 0
assign po048 = pi279;// level 0
assign po049 = pi408;// level 0
assign po050 = pi383;// level 0
assign po051 = pi406;// level 0
assign po052 = pi405;// level 0
assign po053 = pi384;// level 0
assign po054 = pi402;// level 0
assign po055 = pi398;// level 0
assign po056 = pi385;// level 0
assign po057 = pi330;// level 0
assign po058 = pi286;// level 0
assign po059 = pi285;// level 0
assign po060 = pi287;// level 0
assign po061 = pi253;// level 0
assign po062 = pi301;// level 0
assign po063 = pi302;// level 0
assign po064 = pi255;// level 0
assign po065 = pi353;// level 0
assign po066 = pi354;// level 0
assign po067 = pi356;// level 0
assign po068 = pi357;// level 0
assign po069 = pi401;// level 0
assign po070 = pi359;// level 0
assign po071 = pi361;// level 0
assign po072 = pi399;// level 0
assign po073 = pi307;// level 0
assign po074 = pi304;// level 0
assign po075 = pi305;// level 0
assign po076 = pi341;// level 0
assign po077 = pi257;// level 0
assign po078 = pi259;// level 0
assign po079 = pi260;// level 0
assign po080 = pi261;// level 0
assign po081 = pi366;// level 0
assign po082 = pi367;// level 0
assign po083 = pi395;// level 0
assign po084 = pi368;// level 0
assign po085 = pi371;// level 0
assign po086 = pi369;// level 0
assign po087 = pi370;// level 0
assign po088 = pi372;// level 0
assign po089 = pi373;// level 0
assign po090 = pi392;// level 0
assign po091 = pi314;// level 0
assign po092 = pi315;// level 0
assign po093 = pi316;// level 0
assign po094 = pi318;// level 0
assign po095 = pi320;// level 0
assign po096 = pi321;// level 0
assign po097 = pi376;// level 0
assign po098 = pi377;// level 0
assign po099 = pi345;// level 0
assign po100 = pi379;// level 0
assign po101 = pi342;// level 0
assign po102 = pi351;// level 0
assign po103 = pi362;// level 0
assign po104 = pi344;// level 0
assign po105 = pi310;// level 0
assign po106 = pi265;// level 0
assign po107 = pi267;// level 0
assign po108 = pi268;// level 0
assign po109 = pi276;// level 0
assign po110 = pi328;// level 0
assign po111 = pi284;// level 0
assign po112 = pi254;// level 0
assign po113 = pi352;// level 0
assign po114 = pi403;// level 0
assign po115 = pi397;// level 0
assign po116 = pi364;// level 0
assign po117 = pi365;// level 0
assign po118 = pi393;// level 0
assign po119 = pi391;// level 0
assign po120 = pi375;// level 0
assign po121 = pi322;// level 0
assign po122 = pi324;// level 0
assign po123 = pi269;// level 0
assign po124 = pi272;// level 0
assign po125 = pi300;// level 0
assign po126 = pi277;// level 0
assign po127 = pi280;// level 0
assign po128 = pi281;// level 0
assign po129 = pi671;// level 0
assign po130 = one;// level 0
assign po131 = pi670;// level 0
assign po132 = ~w230;// level 23
assign po133 = w282;// level 24
assign po134 = ~w329;// level 23
assign po135 = w373;// level 23
assign po136 = ~w417;// level 25
assign po137 = ~w1299;// level 25
assign po138 = ~w1319;// level 25
assign po139 = w1337;// level 24
assign po140 = w1352;// level 24
assign po141 = w1389;// level 24
assign po142 = ~w1424;// level 23
assign po143 = w1457;// level 23
assign po144 = ~w225;// level 21
assign po145 = ~w1;// level 2
assign po146 = pi012;// level 0
assign po147 = w1460;// level 24
assign po148 = pi013;// level 0
assign po149 = w317;// level 21
assign po150 = pi014;// level 0
assign po151 = ~w371;// level 21
assign po152 = pi015;// level 0
assign po153 = ~w412;// level 23
assign po154 = pi016;// level 0
assign po155 = ~w1377;// level 22
assign po156 = pi017;// level 0
assign po157 = ~w1477;// level 20
assign po158 = ~w1484;// level 20
assign po159 = ~w1494;// level 20
assign po160 = ~w1501;// level 20
assign po161 = ~w1509;// level 20
assign po162 = ~w1516;// level 20
assign po163 = ~w1524;// level 20
assign po164 = ~w1531;// level 20
assign po165 = ~w1544;// level 20
assign po166 = ~w1552;// level 20
assign po167 = ~w1567;// level 20
assign po168 = ~w1577;// level 19
assign po169 = ~w1591;// level 19
assign po170 = ~w1602;// level 20
assign po171 = ~w1612;// level 21
assign po172 = ~w1621;// level 20
assign po173 = ~w1632;// level 20
assign po174 = ~w1642;// level 20
assign po175 = ~w1648;// level 5
assign po176 = ~w1654;// level 5
assign po177 = ~w1666;// level 20
assign po178 = ~w1676;// level 19
assign po179 = ~w1688;// level 19
assign po180 = ~w1699;// level 20
assign po181 = ~w1702;// level 22
assign po182 = pi042;// level 0
assign po183 = w1452;// level 21
assign po184 = pi043;// level 0
assign po185 = ~w267;// level 22
assign po186 = pi044;// level 0
assign po187 = ~w1705;// level 21
assign po188 = pi045;// level 0
assign po189 = w1711;// level 23
assign po190 = w1721;// level 22
assign po191 = ~w1724;// level 21
assign po192 = pi048;// level 0
assign po193 = ~w1727;// level 21
assign po194 = pi049;// level 0
assign po195 = ~w1731;// level 19
assign po196 = ~w1734;// level 19
assign po197 = ~w1738;// level 19
assign po198 = ~w1742;// level 19
assign po199 = ~w1745;// level 19
assign po200 = ~w1748;// level 19
assign po201 = ~w1754;// level 24
assign po202 = pi056;// level 0
assign po203 = w1757;// level 23
assign po204 = pi057;// level 0
assign po205 = ~w1764;// level 23
assign po206 = ~w1771;// level 23
assign po207 = ~w1778;// level 23
assign po208 = ~w1785;// level 23
assign po209 = w1791;// level 5
assign po210 = ~w1801;// level 22
assign po211 = ~w1811;// level 22
assign po212 = ~w1821;// level 22
assign po213 = ~w1831;// level 22
assign po214 = ~w1840;// level 23
assign po215 = ~w1850;// level 23
assign po216 = ~w1854;// level 19
assign po217 = ~w1857;// level 19
assign po218 = ~w1860;// level 19
assign po219 = ~w1863;// level 19
assign po220 = ~w1870;// level 20
assign po221 = ~w1877;// level 21
assign po222 = ~w1887;// level 23
assign po223 = ~w1894;// level 20
assign po224 = ~w1901;// level 21
assign po225 = ~w1908;// level 23
assign po226 = ~w1915;// level 21
assign po227 = ~w1922;// level 20
assign po228 = ~w1929;// level 23
assign po229 = ~w1936;// level 20
assign po230 = ~w1943;// level 21
assign po231 = ~w1950;// level 23
assign po232 = ~w1959;// level 23
assign po233 = ~w1969;// level 19
assign po234 = ~w1979;// level 20
assign po235 = ~w1989;// level 22
assign po236 = ~w1999;// level 20
assign po237 = ~w2009;// level 19
assign po238 = ~w2019;// level 22
assign po239 = ~w2027;// level 23
assign po240 = ~w2033;// level 5
assign po241 = ~w2043;// level 20
assign po242 = ~w2053;// level 21
assign po243 = ~w2063;// level 23
assign po244 = ~w2072;// level 22
assign po245 = ~w2082;// level 20
assign po246 = ~w2092;// level 19
assign po247 = ~w2098;// level 5
assign po248 = ~w2104;// level 5
assign po249 = ~w2114;// level 22
assign po250 = ~w2124;// level 20
assign po251 = ~w2134;// level 19
assign po252 = ~w2144;// level 22
assign po253 = ~w2147;// level 22
assign po254 = ~w2150;// level 22
assign po255 = ~w2153;// level 22
assign po256 = ~w2156;// level 22
assign po257 = ~w2158;// level 21
assign po258 = ~w2161;// level 19
assign po259 = ~w2170;// level 21
assign po260 = ~w2173;// level 19
assign po261 = ~w2176;// level 19
assign po262 = ~w2185;// level 21
assign po263 = ~w2193;// level 23
assign po264 = ~w2196;// level 19
assign po265 = ~w2205;// level 20
assign po266 = ~w2208;// level 19
assign po267 = ~w2211;// level 20
assign po268 = ~w2214;// level 22
assign po269 = ~w2217;// level 19
assign po270 = ~w2220;// level 20
assign po271 = ~w2223;// level 22
assign po272 = ~w2226;// level 19
assign po273 = ~w2229;// level 20
assign po274 = ~w2232;// level 22
assign po275 = ~w2235;// level 22
assign po276 = ~w2238;// level 19
assign po277 = ~w2241;// level 20
assign po278 = w2244;// level 22
assign po279 = w1275;// level 15
assign po280 = w2247;// level 21
assign po281 = w2250;// level 22
assign po282 = w2253;// level 20
assign po283 = ~w2256;// level 24
assign po284 = w2259;// level 22
assign po285 = w2262;// level 19
assign po286 = ~w2269;// level 23
assign po287 = ~w2276;// level 23
assign po288 = ~w2283;// level 23
assign po289 = ~w2290;// level 23
assign po290 = ~w2300;// level 22
assign po291 = w2303;// level 22
assign po292 = w2306;// level 19
assign po293 = w2309;// level 20
assign po294 = ~w2319;// level 22
assign po295 = ~w2325;// level 5
assign po296 = ~w2335;// level 23
assign po297 = ~w2345;// level 22
assign po298 = ~w2355;// level 22
assign po299 = ~w2366;// level 22
assign po300 = w2369;// level 22
assign po301 = w2372;// level 20
assign po302 = w2375;// level 23
assign po303 = w2378;// level 19
assign po304 = w2381;// level 22
assign po305 = ~w2389;// level 22
assign po306 = w2392;// level 22
assign po307 = w2395;// level 22
assign po308 = w2398;// level 22
assign po309 = w2401;// level 22
assign po310 = w2404;// level 22
assign po311 = w1219;// level 19
assign po312 = w2407;// level 21
assign po313 = w358;// level 19
assign po314 = pi166;// level 0
assign po315 = w314;// level 19
assign po316 = pi167;// level 0
assign po317 = ~w2414;// level 21
assign po318 = ~w2421;// level 21
assign po319 = ~w2428;// level 21
assign po320 = ~w2435;// level 21
assign po321 = ~w2445;// level 20
assign po322 = w2451;// level 5
assign po323 = ~w2461;// level 20
assign po324 = ~w2469;// level 21
assign po325 = w2471;// level 21
assign po326 = w2474;// level 22
assign po327 = ~w1265;// level 19
assign po328 = ~w2484;// level 20
assign po329 = ~w2494;// level 21
assign po330 = ~w2504;// level 20
assign po331 = ~w2513;// level 21
assign po332 = ~w2516;// level 20
assign po333 = ~w2519;// level 20
assign po334 = ~w2522;// level 20
assign po335 = w2525;// level 22
assign po336 = ~w2528;// level 20
assign po337 = w2533;// level 22
assign po338 = w2536;// level 22
assign po339 = w1339;// level 19
assign po340 = ~w2539;// level 20
assign po341 = ~w2541;// level 19
assign po342 = ~w2544;// level 20
assign po343 = ~w2547;// level 20
assign po344 = ~w1022;// level 17
assign po345 = ~w2610;// level 20
assign po346 = ~w2641;// level 23
assign po347 = w2668;// level 19
assign po348 = ~w2698;// level 20
assign po349 = ~w2725;// level 20
assign po350 = ~w2753;// level 20
assign po351 = ~w2781;// level 20
assign po352 = ~w2808;// level 21
assign po353 = w2811;// level 19
assign po354 = w2837;// level 16
assign po355 = w2863;// level 16
assign po356 = w2890;// level 17
assign po357 = ~w2918;// level 17
assign po358 = ~w2945;// level 18
assign po359 = w2972;// level 18
assign po360 = w2999;// level 18
assign po361 = w3026;// level 18
assign po362 = ~w3053;// level 18
assign po363 = w3056;// level 18
assign po364 = w3059;// level 21
assign po365 = w3086;// level 18
assign po366 = w3113;// level 18
assign po367 = w3140;// level 18
assign po368 = w3167;// level 18
assign po369 = w3194;// level 18
assign po370 = w3221;// level 18
assign po371 = w3248;// level 18
assign po372 = w3250;// level 20
assign po373 = w3252;// level 20
assign po374 = ~w3254;// level 20
assign po375 = ~w3256;// level 20
assign po376 = w3259;// level 19
assign po377 = w3262;// level 17
assign po378 = w3265;// level 16
assign po379 = w3268;// level 16
assign po380 = w3271;// level 15
assign po381 = w3274;// level 15
assign po382 = w3277;// level 15
assign po383 = w3280;// level 16
assign po384 = w3283;// level 16
assign po385 = w3286;// level 16
assign po386 = w3288;// level 16
assign po387 = ~w3291;// level 19
assign po388 = w3294;// level 16
assign po389 = w3297;// level 16
assign po390 = w3300;// level 16
assign po391 = w3303;// level 16
assign po392 = w3306;// level 16
assign po393 = w3309;// level 16
assign po394 = w3312;// level 16
assign po395 = w3315;// level 16
assign po396 = w3318;// level 18
assign po397 = ~w3321;// level 17
assign po398 = ~w3324;// level 18
assign po399 = ~w3327;// level 18
assign po400 = ~w3330;// level 18
assign po401 = ~w3333;// level 14
assign po402 = ~w3375;// level 16
assign po403 = ~w3398;// level 16
assign po404 = ~w3421;// level 16
assign po405 = ~w3444;// level 16
assign po406 = ~w3467;// level 16
assign po407 = ~w3490;// level 16
assign po408 = ~w3513;// level 16
assign po409 = ~w3536;// level 16
assign po410 = ~w3559;// level 16
assign po411 = ~w3582;// level 16
assign po412 = ~w3605;// level 16
assign po413 = ~w3628;// level 16
assign po414 = ~w3651;// level 16
assign po415 = ~w3674;// level 16
assign po416 = ~w3697;// level 16
assign po417 = ~w3720;// level 16
assign po418 = ~w3743;// level 16
assign po419 = ~w3766;// level 16
assign po420 = ~w3789;// level 16
assign po421 = ~w3812;// level 16
assign po422 = ~w3835;// level 16
assign po423 = ~w3858;// level 16
assign po424 = ~w3881;// level 16
assign po425 = ~w3904;// level 16
assign po426 = ~w3927;// level 16
assign po427 = ~w3950;// level 16
assign po428 = ~w3973;// level 16
assign po429 = ~w3996;// level 16
assign po430 = ~w4019;// level 16
assign po431 = ~w4042;// level 16
assign po432 = ~w4065;// level 16
assign po433 = ~w4088;// level 16
assign po434 = ~w4111;// level 16
assign po435 = ~w4134;// level 16
assign po436 = ~w4157;// level 16
assign po437 = ~w4160;// level 15
assign po438 = ~w4163;// level 14
assign po439 = ~w4166;// level 14
assign po440 = ~w4169;// level 13
assign po441 = ~w4172;// level 13
assign po442 = ~w4175;// level 13
assign po443 = ~w4178;// level 14
assign po444 = ~w4181;// level 14
assign po445 = ~w4184;// level 14
assign po446 = ~w4207;// level 16
assign po447 = ~w4210;// level 14
assign po448 = ~w4233;// level 16
assign po449 = ~w4256;// level 16
assign po450 = ~w4279;// level 16
assign po451 = ~w4302;// level 16
assign po452 = ~w4325;// level 16
assign po453 = ~w4348;// level 16
assign po454 = ~w4371;// level 16
assign po455 = ~w4394;// level 16
assign po456 = ~w4417;// level 16
assign po457 = ~w4440;// level 16
assign po458 = ~w4463;// level 16
assign po459 = ~w4486;// level 16
assign po460 = ~w4509;// level 16
assign po461 = ~w4532;// level 16
assign po462 = ~w4555;// level 16
assign po463 = ~w4578;// level 16
assign po464 = ~w4601;// level 16
assign po465 = ~w4624;// level 16
assign po466 = ~w4647;// level 16
assign po467 = ~w4670;// level 16
assign po468 = ~w4693;// level 16
assign po469 = ~w4716;// level 16
assign po470 = ~w4739;// level 16
assign po471 = ~w4762;// level 16
assign po472 = ~w4785;// level 16
assign po473 = ~w4808;// level 16
assign po474 = ~w4831;// level 16
assign po475 = ~w4854;// level 16
assign po476 = ~w4877;// level 16
assign po477 = ~w4900;// level 16
assign po478 = ~w4923;// level 16
assign po479 = ~w4946;// level 16
assign po480 = ~w4969;// level 16
assign po481 = ~w4972;// level 14
assign po482 = ~w4975;// level 17
assign po483 = ~w4978;// level 14
assign po484 = ~w4981;// level 14
assign po485 = ~w4984;// level 14
assign po486 = ~w4987;// level 14
assign po487 = ~w4990;// level 14
assign po488 = ~w4993;// level 14
assign po489 = ~w5016;// level 16
assign po490 = ~w5039;// level 16
assign po491 = ~w5062;// level 16
assign po492 = ~w5085;// level 16
assign po493 = ~w5108;// level 16
assign po494 = ~w5131;// level 16
assign po495 = ~w5154;// level 16
assign po496 = w5614;// level 25
assign po497 = w5760;// level 25
assign po498 = w5799;// level 25
assign po499 = w5818;// level 25
assign po500 = ~w5841;// level 16
assign po501 = ~w5864;// level 16
assign po502 = ~w5893;// level 16
assign po503 = ~w5921;// level 16
assign po504 = ~w5949;// level 16
assign po505 = ~w5977;// level 16
assign po506 = ~w6005;// level 16
assign po507 = ~w6033;// level 16
assign po508 = ~w6061;// level 16
assign po509 = ~w6089;// level 16
assign po510 = ~w6117;// level 16
assign po511 = ~w6145;// level 16
assign po512 = ~w6173;// level 16
assign po513 = ~w6201;// level 16
assign po514 = ~w6229;// level 16
assign po515 = ~w6257;// level 16
assign po516 = ~w6285;// level 16
assign po517 = ~w6313;// level 16
assign po518 = ~w6341;// level 16
assign po519 = ~w6369;// level 16
assign po520 = ~w6397;// level 16
assign po521 = ~w6425;// level 16
assign po522 = ~w6448;// level 16
assign po523 = ~w6476;// level 16
assign po524 = ~w6504;// level 16
assign po525 = ~w6532;// level 16
assign po526 = ~w6560;// level 18
assign po527 = ~w6588;// level 16
assign po528 = ~w6616;// level 16
assign po529 = ~w6644;// level 16
assign po530 = ~w6672;// level 16
assign po531 = ~w6700;// level 16
assign po532 = ~w6728;// level 16
assign po533 = ~w6756;// level 16
assign po534 = ~w6784;// level 16
assign po535 = ~w6812;// level 16
assign po536 = ~w6815;// level 15
assign po537 = ~w6818;// level 16
assign po538 = ~w6821;// level 16
assign po539 = w6822;// level 9
assign po540 = ~w6850;// level 16
assign po541 = ~w6873;// level 16
assign po542 = ~w6901;// level 16
assign po543 = ~w6904;// level 16
assign po544 = ~w6932;// level 16
assign po545 = ~w6935;// level 16
assign po546 = ~w6963;// level 16
assign po547 = ~w6991;// level 16
assign po548 = ~w7019;// level 16
assign po549 = ~w7047;// level 16
assign po550 = ~w7075;// level 16
assign po551 = ~w7103;// level 16
assign po552 = ~w7131;// level 16
assign po553 = ~w7159;// level 16
assign po554 = ~w7187;// level 16
assign po555 = ~w7215;// level 16
assign po556 = ~w7243;// level 16
assign po557 = ~w7271;// level 16
assign po558 = ~w7274;// level 12
assign po559 = w7392;// level 25
assign po560 = w7424;// level 25
assign po561 = w7446;// level 25
assign po562 = ~w7449;// level 12
assign po563 = ~w7452;// level 11
assign po564 = ~w7455;// level 11
assign po565 = ~w7458;// level 12
assign po566 = ~w7461;// level 12
assign po567 = ~w7464;// level 12
assign po568 = ~w7467;// level 12
assign po569 = w7487;// level 25
assign po570 = ~w7490;// level 12
assign po571 = w7496;// level 25
assign po572 = w7502;// level 25
assign po573 = w7508;// level 25
assign po574 = w7514;// level 25
assign po575 = w7520;// level 25
assign po576 = w7526;// level 25
assign po577 = w7532;// level 25
assign po578 = w7538;// level 25
assign po579 = ~w7541;// level 12
assign po580 = ~w7544;// level 12
assign po581 = ~w7547;// level 12
assign po582 = ~w7550;// level 12
assign po583 = ~w7553;// level 12
assign po584 = w7554;// level 6
assign po585 = ~w7557;// level 12
assign po586 = ~w7560;// level 11
assign po587 = w7582;// level 25
assign po588 = w7604;// level 23
assign po589 = w7620;// level 25
assign po590 = w7642;// level 25
assign po591 = w7657;// level 25
assign po592 = w7666;// level 25
assign po593 = w7676;// level 25
assign po594 = w7686;// level 25
assign po595 = w7696;// level 25
assign po596 = w7706;// level 25
assign po597 = w7716;// level 25
assign po598 = w7726;// level 25
assign po599 = w7739;// level 25
assign po600 = ~w7748;// level 25
assign po601 = w7758;// level 25
assign po602 = w7768;// level 25
assign po603 = w7778;// level 22
assign po604 = w7803;// level 25
assign po605 = w7828;// level 25
assign po606 = w7853;// level 23
assign po607 = w7862;// level 21
assign po608 = w7872;// level 21
assign po609 = w7881;// level 21
assign po610 = w7897;// level 25
assign po611 = ~w7906;// level 25
assign po612 = ~w7915;// level 23
assign po613 = w7930;// level 25
assign po614 = ~w7939;// level 25
assign po615 = ~w7946;// level 25
assign po616 = ~w7953;// level 25
assign po617 = w7959;// level 25
assign po618 = ~w7965;// level 25
assign po619 = w7975;// level 25
assign po620 = ~w7978;// level 25
assign po621 = w7981;// level 23
assign po622 = w7991;// level 25
assign po623 = w8001;// level 25
assign po624 = w8004;// level 25
assign po625 = w8007;// level 25
assign po626 = w8010;// level 25
assign po627 = w8020;// level 25
assign po628 = ~w8023;// level 25
assign po629 = w8026;// level 23
assign po630 = w8036;// level 25
assign po631 = w8046;// level 25
assign po632 = w8049;// level 25
assign po633 = w8052;// level 25
assign po634 = w8055;// level 25
assign po635 = w8058;// level 25
assign po636 = w8061;// level 25
assign po637 = ~w8064;// level 25
assign po638 = w8067;// level 25
assign po639 = ~w8070;// level 25
assign po640 = w8073;// level 25
assign po641 = w8076;// level 25
assign po642 = w8086;// level 25
assign po643 = ~w8089;// level 23
assign po644 = ~w8092;// level 25
assign po645 = w8095;// level 23
assign po646 = ~w8098;// level 23
assign po647 = ~w8101;// level 25
assign po648 = w8104;// level 23
assign po649 = w8107;// level 25
assign po650 = w8110;// level 21
assign po651 = w8113;// level 21
assign po652 = w8116;// level 22
assign po653 = w8119;// level 21
assign po654 = w8122;// level 22
assign po655 = w8125;// level 21
assign po656 = w8128;// level 21
assign po657 = w8131;// level 21
assign po658 = ~w8145;// level 25
assign po659 = ~w8151;// level 25
assign po660 = w8161;// level 25
assign po661 = w8164;// level 25
assign po662 = w8167;// level 25
assign po663 = w8186;// level 21
assign po664 = w8202;// level 23
assign po665 = w8217;// level 23
assign po666 = w8226;// level 21
assign po667 = w8234;// level 25
assign po668 = ~w8237;// level 25
assign po669 = w8247;// level 25
assign po670 = w8250;// level 25
assign po671 = ~w8253;// level 25
assign po672 = w8261;// level 25
assign po673 = ~w8264;// level 25
assign po674 = ~w8267;// level 23
assign po675 = w8270;// level 23
assign po676 = ~w8273;// level 21
assign po677 = w8276;// level 21
assign po678 = w8279;// level 21
assign po679 = ~w8282;// level 25
assign po680 = ~w8285;// level 25
assign po681 = w8288;// level 23
assign po682 = ~w8291;// level 23
assign po683 = ~w8294;// level 25
assign po684 = ~w8297;// level 21
assign po685 = w8300;// level 23
assign po686 = w8303;// level 21
assign po687 = ~w8306;// level 23
assign po688 = ~w8309;// level 25
assign po689 = ~w8312;// level 21
assign po690 = ~w8315;// level 22
assign po691 = w8318;// level 23
assign po692 = ~w8321;// level 25
assign po693 = ~w8324;// level 25
assign po694 = w8327;// level 21
assign po695 = w8330;// level 21
assign po696 = ~w8333;// level 21
assign po697 = ~w8336;// level 23
assign po698 = ~w8339;// level 23
assign po699 = ~w8341;// level 6
assign po700 = ~w8343;// level 8
assign po701 = ~w8345;// level 6
assign po702 = ~w8346;// level 7
assign po703 = w427;// level 2
assign po704 = ~w8361;// level 11
assign po705 = ~w8373;// level 11
assign po706 = w8378;// level 11
assign po707 = ~w8386;// level 12
assign po708 = w8390;// level 10
assign po709 = ~w8391;// level 8
assign po710 = ~w8392;// level 2
assign po711 = w8393;// level 6
assign po712 = ~w8394;// level 7
assign po713 = w8351;// level 5
assign po714 = ~w8397;// level 4
assign po715 = w8398;// level 3
assign po716 = ~w1468;// level 2
assign po717 = ~w8400;// level 7
assign po718 = ~w8403;// level 3
assign po719 = ~w8406;// level 3
assign po720 = ~w8409;// level 3
assign po721 = ~w8412;// level 3
assign po722 = ~w8415;// level 3
assign po723 = ~w8418;// level 3
assign po724 = ~w8421;// level 3
assign po725 = ~w8424;// level 3
assign po726 = ~w8427;// level 3
assign po727 = ~w8430;// level 3
assign po728 = ~w8433;// level 3
assign po729 = ~w8436;// level 3
assign po730 = ~w8439;// level 3
assign po731 = ~w8442;// level 3
assign po732 = ~w8445;// level 3
assign po733 = ~w8448;// level 3
assign po734 = ~w8451;// level 3
assign po735 = ~w8454;// level 3
assign po736 = ~w8457;// level 3
assign po737 = ~w8460;// level 3
assign po738 = ~w8463;// level 3
assign po739 = ~w8466;// level 3
assign po740 = ~w8469;// level 3
assign po741 = ~w8472;// level 3
assign po742 = ~w8475;// level 3
assign po743 = ~w8478;// level 3
assign po744 = ~w8481;// level 3
assign po745 = ~w8484;// level 3
assign po746 = ~w8487;// level 3
assign po747 = ~w8490;// level 3
assign po748 = ~w8493;// level 3
assign po749 = ~w8496;// level 3
assign po750 = ~w8499;// level 3
assign po751 = ~w8502;// level 3
assign po752 = ~w8505;// level 3
assign po753 = ~w8508;// level 3
assign po754 = ~w8511;// level 3
assign po755 = ~w8514;// level 3
assign po756 = ~w8517;// level 3
assign po757 = ~w8520;// level 3
assign po758 = ~w8523;// level 3
assign po759 = ~w8526;// level 3
assign po760 = ~w8529;// level 3
assign po761 = ~w8532;// level 3
assign po762 = ~w8535;// level 3
assign po763 = ~w8538;// level 3
assign po764 = ~w8541;// level 3
assign po765 = ~w8544;// level 3
assign po766 = ~w8547;// level 3
assign po767 = ~w8550;// level 3
assign po768 = ~w8553;// level 3
assign po769 = ~w8556;// level 3
assign po770 = ~w8559;// level 3
assign po771 = ~w8562;// level 3
assign po772 = ~w8565;// level 3
assign po773 = ~w8568;// level 3
assign po774 = ~w8571;// level 3
assign po775 = ~w8574;// level 3
assign po776 = ~w8577;// level 3
assign po777 = ~w8580;// level 3
assign po778 = ~w8583;// level 3
assign po779 = ~w8586;// level 3
assign po780 = ~w8589;// level 3
assign po781 = ~w8592;// level 3
assign po782 = ~w8595;// level 3
assign po783 = ~w8598;// level 3
assign po784 = ~w8601;// level 3
assign po785 = ~w8604;// level 3
assign po786 = ~w8607;// level 3
assign po787 = ~w8610;// level 3
assign po788 = ~w8613;// level 3
assign po789 = ~w8616;// level 3
assign po790 = ~w8619;// level 3
assign po791 = ~w8622;// level 3
assign po792 = ~w8625;// level 3
assign po793 = ~w8628;// level 3
assign po794 = ~w8631;// level 3
assign po795 = ~w8634;// level 3
assign po796 = ~w8637;// level 3
assign po797 = ~w8640;// level 3
assign po798 = ~w8643;// level 3
assign po799 = ~w8646;// level 3
assign po800 = ~w8649;// level 3
assign po801 = ~w8652;// level 3
assign po802 = ~w8655;// level 3
assign po803 = ~w8658;// level 3
assign po804 = ~w8661;// level 3
assign po805 = ~w8664;// level 3
assign po806 = ~w8667;// level 3
assign po807 = ~w8670;// level 3
assign po808 = ~w8673;// level 3
assign po809 = ~w8676;// level 3
assign po810 = ~w8679;// level 3
assign po811 = ~w8682;// level 3
assign po812 = ~w8685;// level 3
assign po813 = ~w8688;// level 3
assign po814 = w1;// level 2
assign po815 = w5162;// level 1
assign po816 = w8347;// level 1
assign po817 = ~w8689;// level 3
assign po818 = w1462;// level 3
endmodule
