module pci_bridge32 ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205,
    pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214,
    pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223,
    pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232,
    pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241,
    pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250,
    pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259,
    pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268,
    pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277,
    pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286,
    pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295,
    pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304,
    pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313,
    pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322,
    pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331,
    pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340,
    pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349,
    pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358,
    pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367,
    pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376,
    pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385,
    pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394,
    pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403,
    pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412,
    pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421,
    pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430,
    pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439,
    pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448,
    pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457,
    pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466,
    pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475,
    pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484,
    pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493,
    pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502,
    pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511,
    pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520,
    pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529,
    pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538,
    pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547,
    pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556,
    pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565,
    pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574,
    pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583,
    pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592,
    pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601,
    pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610,
    pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619,
    pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628,
    pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637,
    pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646,
    pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655,
    pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664,
    pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673,
    pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682,
    pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691,
    pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700,
    pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709,
    pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718,
    pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727,
    pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736,
    pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745,
    pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754,
    pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763,
    pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772,
    pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781,
    pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790,
    pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799,
    pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808,
    pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817,
    pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826,
    pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835,
    pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844,
    pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853,
    pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862,
    pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871,
    pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880,
    pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889,
    pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898,
    pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907,
    pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916,
    pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925,
    pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934,
    pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943,
    pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952,
    pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961,
    pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970,
    pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979,
    pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988,
    pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997,
    pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006,
    pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015,
    pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024,
    pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033,
    pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042,
    pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051,
    pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060,
    pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069,
    pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078,
    pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087,
    pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096,
    pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105,
    pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114,
    pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123,
    pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132,
    pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141,
    pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150,
    pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159,
    pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168,
    pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177,
    pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186,
    pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195,
    pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204,
    pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213,
    pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222,
    pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231,
    pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240,
    pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249,
    pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258,
    pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267,
    pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276,
    pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285,
    pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294,
    pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303,
    pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312,
    pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321,
    pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330,
    pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339,
    pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348,
    pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357,
    pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366,
    pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375,
    pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384,
    pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393,
    pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402,
    pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411,
    pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420,
    pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429,
    pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438,
    pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447,
    pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456,
    pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465,
    pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474,
    pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483,
    pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492,
    pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501,
    pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510,
    pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519,
    pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528,
    pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537,
    pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546,
    pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555,
    pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564,
    pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573,
    pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582,
    pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591,
    pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600,
    pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609,
    pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618,
    pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627,
    pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636,
    pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645,
    pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654,
    pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663,
    pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672,
    pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681,
    pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690,
    pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699,
    pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708,
    pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717,
    pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726,
    pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735,
    pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744,
    pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753,
    pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762,
    pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771,
    pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780,
    pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789,
    pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798,
    pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807,
    pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816,
    pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825,
    pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834,
    pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843,
    pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852,
    pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861,
    pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870,
    pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879,
    pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888,
    pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897,
    pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906,
    pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915,
    pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924,
    pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933,
    pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942,
    pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951,
    pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960,
    pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969,
    pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978,
    pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987,
    pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996,
    pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005,
    pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014,
    pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023,
    pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032,
    pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041,
    pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050,
    pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059,
    pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068,
    pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077,
    pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086,
    pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095,
    pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104,
    pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113,
    pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122,
    pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131,
    pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140,
    pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149,
    pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158,
    pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167,
    pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176,
    pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185,
    pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194,
    pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203,
    pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212,
    pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221,
    pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230,
    pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239,
    pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248,
    pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257,
    pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266,
    pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275,
    pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284,
    pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293,
    pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302,
    pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311,
    pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320,
    pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329,
    pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338,
    pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347,
    pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356,
    pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365,
    pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374,
    pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383,
    pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392,
    pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401,
    pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410,
    pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419,
    pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428,
    pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437,
    pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446,
    pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455,
    pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464,
    pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473,
    pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482,
    pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491,
    pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500,
    pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509,
    pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511,
    po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520,
    po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529,
    po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538,
    po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547,
    po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556,
    po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565,
    po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574,
    po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583,
    po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592,
    po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601,
    po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610,
    po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619,
    po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628,
    po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637,
    po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646,
    po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655,
    po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664,
    po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673,
    po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682,
    po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691,
    po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700,
    po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709,
    po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718,
    po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727,
    po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736,
    po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745,
    po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754,
    po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763,
    po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772,
    po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781,
    po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790,
    po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799,
    po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808,
    po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817,
    po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826,
    po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835,
    po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844,
    po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853,
    po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862,
    po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871,
    po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880,
    po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889,
    po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898,
    po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907,
    po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916,
    po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925,
    po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934,
    po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943,
    po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952,
    po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961,
    po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970,
    po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979,
    po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988,
    po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997,
    po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006,
    po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015,
    po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024,
    po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033,
    po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042,
    po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051,
    po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060,
    po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069,
    po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078,
    po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087,
    po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096,
    po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105,
    po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114,
    po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123,
    po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132,
    po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141,
    po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150,
    po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159,
    po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168,
    po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177,
    po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186,
    po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195,
    po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204,
    po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213,
    po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222,
    po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231,
    po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240,
    po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249,
    po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258,
    po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267,
    po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276,
    po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285,
    po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294,
    po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303,
    po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312,
    po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321,
    po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330,
    po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339,
    po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348,
    po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357,
    po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366,
    po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375,
    po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384,
    po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393,
    po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402,
    po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411,
    po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420,
    po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429,
    po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438,
    po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447,
    po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456,
    po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465,
    po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474,
    po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483,
    po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492,
    po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501,
    po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510,
    po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519,
    po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528,
    po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537,
    po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546,
    po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555,
    po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564,
    po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573,
    po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582,
    po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591,
    po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600,
    po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609,
    po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618,
    po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627,
    po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636,
    po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645,
    po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654,
    po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663,
    po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672,
    po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681,
    po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690,
    po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699,
    po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708,
    po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717,
    po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726,
    po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735,
    po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744,
    po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753,
    po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762,
    po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771,
    po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780,
    po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789,
    po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798,
    po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807,
    po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816,
    po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825,
    po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834,
    po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843,
    po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852,
    po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861,
    po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870,
    po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879,
    po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888,
    po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897,
    po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906,
    po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915,
    po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924,
    po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933,
    po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942,
    po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951,
    po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960,
    po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969,
    po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978,
    po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987,
    po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996,
    po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005,
    po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014,
    po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023,
    po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032,
    po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041,
    po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050,
    po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059,
    po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068,
    po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077,
    po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086,
    po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095,
    po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104,
    po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113,
    po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122,
    po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131,
    po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140,
    po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149,
    po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158,
    po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167,
    po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176,
    po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185,
    po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194,
    po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203,
    po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212,
    po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221,
    po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230,
    po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239,
    po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248,
    po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257,
    po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266,
    po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275,
    po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284,
    po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293,
    po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302,
    po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311,
    po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320,
    po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329,
    po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338,
    po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347,
    po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356,
    po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365,
    po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374,
    po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383,
    po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392,
    po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401,
    po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410,
    po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419,
    po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428,
    po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437,
    po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446,
    po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455,
    po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464,
    po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473,
    po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482,
    po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491,
    po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500,
    po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509,
    po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518,
    po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204,
    pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213,
    pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222,
    pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231,
    pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240,
    pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249,
    pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258,
    pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267,
    pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276,
    pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285,
    pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294,
    pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303,
    pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312,
    pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321,
    pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330,
    pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339,
    pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348,
    pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357,
    pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366,
    pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375,
    pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384,
    pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393,
    pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402,
    pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411,
    pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420,
    pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429,
    pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438,
    pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447,
    pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456,
    pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465,
    pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474,
    pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483,
    pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492,
    pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501,
    pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510,
    pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519,
    pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528,
    pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537,
    pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546,
    pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555,
    pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564,
    pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573,
    pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582,
    pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591,
    pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600,
    pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609,
    pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618,
    pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627,
    pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636,
    pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645,
    pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654,
    pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663,
    pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672,
    pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681,
    pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690,
    pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699,
    pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708,
    pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717,
    pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726,
    pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735,
    pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744,
    pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753,
    pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762,
    pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771,
    pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780,
    pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789,
    pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798,
    pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807,
    pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816,
    pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825,
    pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834,
    pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843,
    pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852,
    pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861,
    pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870,
    pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879,
    pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888,
    pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897,
    pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906,
    pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915,
    pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924,
    pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933,
    pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942,
    pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951,
    pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960,
    pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969,
    pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978,
    pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987,
    pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996,
    pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005,
    pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014,
    pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023,
    pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032,
    pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041,
    pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050,
    pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059,
    pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068,
    pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077,
    pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086,
    pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095,
    pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104,
    pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113,
    pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122,
    pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131,
    pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140,
    pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149,
    pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158,
    pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167,
    pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176,
    pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185,
    pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194,
    pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203,
    pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212,
    pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221,
    pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230,
    pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239,
    pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248,
    pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257,
    pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266,
    pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275,
    pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284,
    pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293,
    pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302,
    pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311,
    pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320,
    pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329,
    pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338,
    pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347,
    pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356,
    pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365,
    pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374,
    pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383,
    pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392,
    pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401,
    pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410,
    pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419,
    pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428,
    pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437,
    pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446,
    pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455,
    pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464,
    pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473,
    pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482,
    pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491,
    pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500,
    pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509,
    pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518,
    pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527,
    pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536,
    pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545,
    pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554,
    pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563,
    pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572,
    pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581,
    pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590,
    pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599,
    pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608,
    pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617,
    pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626,
    pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635,
    pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644,
    pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653,
    pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662,
    pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671,
    pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680,
    pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689,
    pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698,
    pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707,
    pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716,
    pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725,
    pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734,
    pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743,
    pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752,
    pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761,
    pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770,
    pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779,
    pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788,
    pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797,
    pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806,
    pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815,
    pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824,
    pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833,
    pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842,
    pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851,
    pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860,
    pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869,
    pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878,
    pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887,
    pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896,
    pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905,
    pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914,
    pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923,
    pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932,
    pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941,
    pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950,
    pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959,
    pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968,
    pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977,
    pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986,
    pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995,
    pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004,
    pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013,
    pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022,
    pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031,
    pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040,
    pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049,
    pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058,
    pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067,
    pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076,
    pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085,
    pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094,
    pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103,
    pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112,
    pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121,
    pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130,
    pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139,
    pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148,
    pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157,
    pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166,
    pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175,
    pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184,
    pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193,
    pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202,
    pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211,
    pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220,
    pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229,
    pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238,
    pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247,
    pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256,
    pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265,
    pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274,
    pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283,
    pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292,
    pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301,
    pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310,
    pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319,
    pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328,
    pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337,
    pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346,
    pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355,
    pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364,
    pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373,
    pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382,
    pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391,
    pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400,
    pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409,
    pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418,
    pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427,
    pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436,
    pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445,
    pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454,
    pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463,
    pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472,
    pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481,
    pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490,
    pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499,
    pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508,
    pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517,
    pi3518;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510,
    po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519,
    po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528,
    po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537,
    po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546,
    po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555,
    po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564,
    po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573,
    po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582,
    po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591,
    po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600,
    po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609,
    po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618,
    po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627,
    po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636,
    po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645,
    po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654,
    po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663,
    po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672,
    po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681,
    po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690,
    po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699,
    po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708,
    po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717,
    po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726,
    po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735,
    po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744,
    po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753,
    po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762,
    po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771,
    po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780,
    po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789,
    po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798,
    po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807,
    po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816,
    po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825,
    po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834,
    po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843,
    po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852,
    po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861,
    po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870,
    po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879,
    po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888,
    po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897,
    po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906,
    po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915,
    po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924,
    po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933,
    po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942,
    po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951,
    po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960,
    po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969,
    po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978,
    po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987,
    po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996,
    po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005,
    po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014,
    po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023,
    po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032,
    po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041,
    po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050,
    po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059,
    po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068,
    po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077,
    po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086,
    po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095,
    po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104,
    po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113,
    po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122,
    po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131,
    po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140,
    po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149,
    po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158,
    po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167,
    po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176,
    po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185,
    po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194,
    po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203,
    po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212,
    po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221,
    po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230,
    po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239,
    po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248,
    po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257,
    po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266,
    po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275,
    po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284,
    po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293,
    po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302,
    po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311,
    po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320,
    po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329,
    po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338,
    po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347,
    po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356,
    po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365,
    po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374,
    po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383,
    po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392,
    po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401,
    po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410,
    po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419,
    po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428,
    po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437,
    po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446,
    po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455,
    po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464,
    po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473,
    po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482,
    po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491,
    po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500,
    po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509,
    po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518,
    po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527,
    po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536,
    po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545,
    po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554,
    po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563,
    po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572,
    po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581,
    po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590,
    po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599,
    po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608,
    po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617,
    po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626,
    po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635,
    po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644,
    po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653,
    po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662,
    po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671,
    po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680,
    po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689,
    po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698,
    po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707,
    po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716,
    po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725,
    po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734,
    po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743,
    po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752,
    po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761,
    po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770,
    po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779,
    po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788,
    po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797,
    po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806,
    po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815,
    po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824,
    po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833,
    po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842,
    po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851,
    po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860,
    po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869,
    po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878,
    po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887,
    po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896,
    po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905,
    po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914,
    po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923,
    po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932,
    po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941,
    po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950,
    po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959,
    po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968,
    po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977,
    po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986,
    po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995,
    po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004,
    po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013,
    po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022,
    po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031,
    po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040,
    po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049,
    po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058,
    po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067,
    po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076,
    po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085,
    po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094,
    po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103,
    po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112,
    po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121,
    po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130,
    po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139,
    po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148,
    po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157,
    po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166,
    po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175,
    po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184,
    po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193,
    po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202,
    po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211,
    po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220,
    po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229,
    po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238,
    po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247,
    po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256,
    po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265,
    po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274,
    po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283,
    po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292,
    po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301,
    po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310,
    po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319,
    po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328,
    po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337,
    po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346,
    po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355,
    po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364,
    po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373,
    po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382,
    po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391,
    po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400,
    po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409,
    po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418,
    po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427,
    po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436,
    po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445,
    po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454,
    po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463,
    po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472,
    po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481,
    po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490,
    po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499,
    po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508,
    po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517,
    po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526,
    po3527;
  wire n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
    n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
    n7110, n7111, n7112, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
    n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
    n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7234,
    n7235, n7236, n7237, n7238, n7239, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7260, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7275, n7276, n7277,
    n7278, n7279, n7280, n7281, n7282, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7302, n7303, n7304, n7305, n7306, n7308, n7309, n7310, n7311,
    n7312, n7314, n7315, n7316, n7317, n7318, n7320, n7321, n7322, n7323,
    n7324, n7326, n7327, n7328, n7329, n7330, n7332, n7333, n7334, n7335,
    n7336, n7338, n7339, n7340, n7341, n7342, n7344, n7345, n7346, n7347,
    n7348, n7350, n7351, n7352, n7353, n7354, n7356, n7357, n7358, n7359,
    n7360, n7362, n7363, n7364, n7365, n7366, n7368, n7369, n7370, n7371,
    n7372, n7374, n7375, n7376, n7377, n7378, n7380, n7381, n7382, n7383,
    n7384, n7386, n7387, n7388, n7389, n7390, n7392, n7393, n7394, n7395,
    n7396, n7398, n7399, n7400, n7401, n7402, n7404, n7405, n7406, n7407,
    n7408, n7410, n7411, n7412, n7413, n7414, n7416, n7417, n7418, n7419,
    n7420, n7422, n7423, n7424, n7425, n7426, n7428, n7429, n7430, n7431,
    n7432, n7434, n7435, n7436, n7437, n7438, n7440, n7441, n7442, n7443,
    n7444, n7446, n7447, n7448, n7449, n7450, n7452, n7453, n7454, n7455,
    n7456, n7458, n7459, n7460, n7461, n7462, n7464, n7465, n7466, n7467,
    n7468, n7470, n7471, n7472, n7473, n7474, n7476, n7477, n7478, n7479,
    n7480, n7482, n7483, n7484, n7485, n7486, n7488, n7489, n7490, n7491,
    n7492, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
    n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
    n7554, n7555, n7556, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
    n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
    n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
    n7712, n7713, n7714, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
    n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
    n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
    n7766, n7767, n7768, n7769, n7771, n7772, n7773, n7774, n7775, n7776,
    n7777, n7778, n7779, n7780, n7781, n7783, n7784, n7785, n7786, n7787,
    n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
    n7842, n7843, n7844, n7845, n7846, n7847, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7885,
    n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
    n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
    n7962, n7963, n7964, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7975, n7976, n7977, n7978, n7979, n7981, n7982, n7983, n7985,
    n7986, n7988, n7989, n7991, n7992, n7994, n7995, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
    n8102, n8103, n8104, n8105, n8106, n8107, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
    n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
    n8173, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
    n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8251, n8252, n8253, n8254, n8255,
    n8256, n8258, n8259, n8260, n8262, n8263, n8264, n8265, n8266, n8267,
    n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
    n8309, n8310, n8311, n8313, n8314, n8316, n8317, n8319, n8320, n8321,
    n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
    n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347, n8349, n8350, n8351, n8352,
    n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
    n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8394, n8395,
    n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422, n8424, n8425, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
    n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
    n8492, n8493, n8494, n8495, n8496, n8497, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
    n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
    n8524, n8525, n8526, n8527, n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8544, n8545,
    n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572, n8574, n8575, n8576, n8577,
    n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
    n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
    n8642, n8643, n8644, n8645, n8646, n8647, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
    n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
    n8674, n8675, n8676, n8677, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
    n8706, n8707, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
    n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8754, n8755, n8756, n8757, n8758, n8759,
    n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
    n8792, n8793, n8794, n8795, n8796, n8797, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
    n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
    n8856, n8857, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
    n8867, n8868, n8869, n8870, n8871, n8872, n8874, n8875, n8876, n8877,
    n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
    n8889, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
    n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
    n8952, n8953, n8954, n8955, n8956, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
    n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
    n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
    n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
    n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9371, n9372, n9373, n9374, n9375, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
    n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
    n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
    n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9528, n9530,
    n9531, n9532, n9533, n9534, n9536, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9574,
    n9575, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
    n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9595, n9596,
    n9598, n9599, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
    n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9645, n9646, n9647, n9648, n9649,
    n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
    n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
    n9680, n9681, n9682, n9683, n9684, n9685, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
    n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
    n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
    n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
    n9772, n9773, n9774, n9775, n9776, n9777, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
    n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9823,
    n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
    n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
    n9864, n9865, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
    n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
    n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
    n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
    n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
    n9946, n9947, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
    n9977, n9978, n9979, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
    n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
    n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
    n10007, n10008, n10009, n10010, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
    n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
    n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
    n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
    n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
    n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
    n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
    n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
    n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
    n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
    n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10242, n10243, n10244, n10245, n10246, n10247,
    n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
    n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10284,
    n10286, n10288, n10290, n10292, n10294, n10296, n10298, n10300, n10302,
    n10304, n10306, n10308, n10310, n10312, n10314, n10315, n10316, n10317,
    n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
    n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
    n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10353, n10354,
    n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
    n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
    n10391, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
    n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
    n10428, n10429, n10430, n10431, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
    n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
    n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
    n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10553, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
    n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10633, n10635, n10637, n10639, n10641, n10643, n10645, n10647,
    n10649, n10651, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
    n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
    n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
    n10714, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10760,
    n10762, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10804, n10806, n10807, n10808, n10809,
    n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10856,
    n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
    n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
    n10921, n10922, n10923, n10925, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
    n10968, n10969, n10970, n10971, n10973, n10975, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10986, n10987, n10988, n10989,
    n10990, n10992, n10993, n10994, n10995, n10996, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
    n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11022, n11023, n11025, n11026, n11028, n11029, n11031,
    n11032, n11034, n11035, n11037, n11038, n11040, n11041, n11043, n11044,
    n11046, n11047, n11049, n11050, n11053, n11054, n11055, n11056, n11057,
    n11060, n11061, n11063, n11064, n11066, n11067, n11069, n11070, n11072,
    n11073, n11075, n11076, n11078, n11079, n11081, n11082, n11084, n11085,
    n11087, n11088, n11090, n11091, n11093, n11094, n11096, n11097, n11099,
    n11100, n11102, n11103, n11105, n11106, n11108, n11109, n11111, n11112,
    n11114, n11115, n11117, n11118, n11120, n11121, n11123, n11124, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
    n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
    n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
    n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
    n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
    n11200, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11215, n11216, n11217, n11218, n11219,
    n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234, n11236, n11237, n11238,
    n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
    n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
    n11257, n11258, n11259, n11261, n11262, n11263, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310, n11312, n11313, n11314,
    n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
    n11324, n11325, n11326, n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11347, n11348, n11349, n11350, n11351, n11352,
    n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
    n11362, n11363, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
    n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
    n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
    n11390, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
    n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
    n11419, n11420, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
    n11429, n11430, n11431, n11432, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444, n11446, n11447, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
    n11469, n11470, n11471, n11472, n11473, n11474, n11476, n11478, n11479,
    n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11490,
    n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
    n11500, n11501, n11502, n11503, n11505, n11506, n11507, n11508, n11509,
    n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
    n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11551, n11552, n11554, n11555, n11557, n11558, n11559,
    n11560, n11561, n11563, n11564, n11565, n11566, n11567, n11569, n11570,
    n11571, n11572, n11573, n11575, n11576, n11577, n11578, n11579, n11581,
    n11582, n11583, n11584, n11585, n11587, n11588, n11589, n11590, n11591,
    n11593, n11594, n11595, n11596, n11597, n11599, n11600, n11601, n11602,
    n11603, n11605, n11606, n11607, n11608, n11609, n11611, n11612, n11613,
    n11614, n11615, n11617, n11618, n11619, n11620, n11621, n11623, n11624,
    n11625, n11626, n11627, n11629, n11630, n11631, n11632, n11633, n11635,
    n11636, n11637, n11638, n11639, n11641, n11642, n11643, n11644, n11645,
    n11647, n11648, n11649, n11650, n11651, n11653, n11654, n11655, n11656,
    n11657, n11659, n11660, n11661, n11662, n11663, n11665, n11666, n11667,
    n11668, n11669, n11671, n11672, n11673, n11674, n11675, n11677, n11678,
    n11679, n11680, n11681, n11683, n11684, n11685, n11686, n11687, n11689,
    n11690, n11691, n11692, n11693, n11695, n11696, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705, n11707, n11708, n11709,
    n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11719,
    n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11744, n11745, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754, n11756, n11757, n11758,
    n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11780, n11781, n11782, n11783, n11784, n11786, n11787, n11788,
    n11789, n11790, n11792, n11793, n11794, n11795, n11796, n11798, n11799,
    n11800, n11801, n11802, n11804, n11805, n11807, n11808, n11810, n11811,
    n11812, n11813, n11814, n11816, n11817, n11818, n11819, n11820, n11821,
    n11823, n11824, n11826, n11827, n11829, n11830, n11832, n11833, n11835,
    n11836, n11838, n11839, n11841, n11842, n11844, n11845, n11847, n11848,
    n11849, n11850, n11851, n11853, n11854, n11855, n11856, n11857, n11859,
    n11860, n11862, n11863, n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11877, n11878, n11879, n11880,
    n11881, n11883, n11884, n11885, n11886, n11887, n11889, n11890, n11891,
    n11892, n11893, n11895, n11896, n11897, n11898, n11899, n11901, n11902,
    n11903, n11904, n11905, n11907, n11908, n11909, n11910, n11911, n11913,
    n11914, n11916, n11917, n11918, n11919, n11920, n11922, n11923, n11924,
    n11925, n11926, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
    n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
    n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
    n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
    n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
    n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
    n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
    n12046, n12047, n12048, n12050, n12051, n12052, n12053, n12054, n12055,
    n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
    n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
    n12074, n12075, n12076, n12077, n12078, n12079, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
    n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
    n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
    n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
    n12139, n12140, n12141, n12143, n12144, n12145, n12146, n12147, n12148,
    n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
    n12167, n12168, n12169, n12170, n12171, n12172, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
    n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
    n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
    n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
    n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
    n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
    n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
    n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
    n12325, n12326, n12327, n12329, n12330, n12331, n12332, n12333, n12335,
    n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
    n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12394, n12395, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
    n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
    n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12552, n12553, n12554, n12555, n12556, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12568, n12569,
    n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
    n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
    n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
    n12625, n12626, n12627, n12628, n12630, n12631, n12632, n12633, n12634,
    n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
    n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
    n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
    n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
    n12690, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
    n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
    n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12721, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
    n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12754, n12755,
    n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
    n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
    n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
    n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
    n12811, n12812, n12813, n12814, n12816, n12817, n12818, n12819, n12820,
    n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
    n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
    n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
    n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
    n12876, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
    n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
    n12904, n12905, n12906, n12907, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
    n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
    n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12940, n12941,
    n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
    n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
    n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
    n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13002, n13003, n13004, n13005, n13006,
    n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
    n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
    n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
    n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
    n13062, n13064, n13065, n13067, n13068, n13070, n13071, n13073, n13074,
    n13076, n13077, n13079, n13080, n13082, n13083, n13085, n13086, n13088,
    n13089, n13091, n13092, n13094, n13095, n13097, n13098, n13100, n13101,
    n13103, n13104, n13106, n13107, n13109, n13110, n13112, n13113, n13115,
    n13116, n13118, n13119, n13121, n13122, n13124, n13125, n13127, n13128,
    n13130, n13131, n13133, n13134, n13136, n13137, n13139, n13140, n13142,
    n13143, n13145, n13146, n13148, n13149, n13151, n13152, n13154, n13155,
    n13157, n13158, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13175, n13176,
    n13178, n13179, n13180, n13182, n13183, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
    n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
    n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13239, n13240, n13241, n13242, n13243,
    n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
    n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
    n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13270, n13271,
    n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
    n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
    n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
    n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
    n13327, n13328, n13329, n13330, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
    n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
    n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
    n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
    n13392, n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
    n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
    n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
    n13420, n13421, n13422, n13423, n13425, n13426, n13427, n13428, n13429,
    n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
    n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
    n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13456, n13457,
    n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
    n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
    n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
    n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
    n13513, n13514, n13515, n13516, n13518, n13519, n13520, n13521, n13522,
    n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
    n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
    n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
    n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
    n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
    n13606, n13607, n13608, n13609, n13611, n13612, n13613, n13614, n13615,
    n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
    n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
    n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13642, n13643,
    n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
    n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
    n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
    n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
    n13699, n13700, n13701, n13702, n13704, n13705, n13706, n13707, n13708,
    n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
    n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
    n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
    n13764, n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
    n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
    n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
    n13792, n13793, n13794, n13795, n13797, n13798, n13799, n13800, n13801,
    n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
    n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
    n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
    n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
    n13885, n13886, n13887, n13888, n13890, n13891, n13892, n13893, n13894,
    n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
    n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
    n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
    n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
    n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
    n13978, n13979, n13980, n13981, n13983, n13984, n13985, n13986, n13987,
    n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
    n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14014, n14015,
    n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
    n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
    n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
    n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
    n14071, n14072, n14073, n14074, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
    n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
    n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
    n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
    n14136, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
    n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
    n14164, n14165, n14166, n14167, n14169, n14170, n14171, n14172, n14173,
    n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
    n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14200, n14201,
    n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
    n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
    n14257, n14258, n14259, n14260, n14262, n14263, n14264, n14265, n14266,
    n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
    n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
    n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
    n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
    n14322, n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
    n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
    n14350, n14351, n14352, n14353, n14355, n14356, n14357, n14358, n14359,
    n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
    n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
    n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
    n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
    n14396, n14397, n14398, n14399, n14401, n14402, n14403, n14404, n14405,
    n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
    n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
    n14425, n14426, n14427, n14428, n14429, n14431, n14432, n14433, n14434,
    n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
    n14454, n14455, n14456, n14457, n14458, n14459, n14461, n14462, n14463,
    n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
    n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
    n14502, n14503, n14504, n14506, n14507, n14508, n14509, n14510, n14511,
    n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
    n14531, n14532, n14533, n14534, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
    n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
    n14579, n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594, n14596, n14597, n14598,
    n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
    n14608, n14609, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14626, n14627,
    n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14641, n14642, n14643, n14644, n14645, n14646,
    n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14656,
    n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14671, n14672, n14673, n14674, n14675,
    n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
    n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14701, n14702, n14703, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
    n14724, n14725, n14726, n14727, n14728, n14729, n14731, n14732, n14733,
    n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
    n14743, n14744, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
    n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
    n14772, n14773, n14774, n14776, n14777, n14778, n14779, n14780, n14781,
    n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14791,
    n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
    n14801, n14802, n14803, n14804, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
    n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
    n14830, n14831, n14832, n14833, n14834, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
    n14849, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14866, n14867, n14868,
    n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
    n14878, n14879, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14918, n14919, n14920, n14921, n14923, n14924, n14925,
    n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
    n14935, n14936, n14937, n14938, n14940, n14941, n14942, n14943, n14944,
    n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
    n14964, n14965, n14966, n14967, n14968, n14970, n14971, n14972, n14973,
    n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
    n14993, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
    n15022, n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15040, n15041,
    n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15055, n15056, n15057, n15058, n15059, n15060,
    n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15070,
    n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15084, n15085, n15086, n15087, n15088, n15089,
    n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15099,
    n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
    n15109, n15110, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
    n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
    n15148, n15149, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
    n15167, n15168, n15169, n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192, n15194, n15195, n15196,
    n15197, n15198, n15199, n15200, n15201, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15212, n15213, n15214, n15215, n15216,
    n15217, n15218, n15219, n15221, n15222, n15223, n15224, n15225, n15226,
    n15227, n15228, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242, n15244, n15245, n15246,
    n15247, n15248, n15249, n15250, n15251, n15253, n15254, n15255, n15256,
    n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15275, n15276,
    n15277, n15278, n15279, n15280, n15281, n15282, n15284, n15285, n15286,
    n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302, n15304, n15305, n15306,
    n15307, n15308, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
    n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15330, n15331, n15332, n15333, n15334, n15335,
    n15336, n15337, n15338, n15339, n15340, n15342, n15343, n15344, n15345,
    n15346, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
    n15365, n15366, n15367, n15368, n15369, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15383, n15384,
    n15385, n15386, n15387, n15388, n15389, n15390, n15392, n15393, n15394,
    n15395, n15396, n15397, n15399, n15400, n15401, n15402, n15403, n15404,
    n15406, n15407, n15408, n15409, n15410, n15411, n15413, n15414, n15415,
    n15416, n15417, n15418, n15420, n15421, n15422, n15423, n15424, n15426,
    n15427, n15428, n15429, n15430, n15431, n15433, n15434, n15435, n15436,
    n15437, n15438, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
    n15458, n15459, n15460, n15461, n15462, n15464, n15465, n15466, n15467,
    n15468, n15469, n15470, n15471, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15482, n15483, n15484, n15485, n15486, n15487,
    n15488, n15489, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
    n15498, n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
    n15509, n15510, n15511, n15512, n15513, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15524, n15525, n15526, n15527, n15528,
    n15529, n15530, n15531, n15533, n15534, n15535, n15536, n15537, n15538,
    n15539, n15540, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
    n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15569,
    n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15578, n15579,
    n15580, n15581, n15582, n15583, n15584, n15585, n15587, n15588, n15589,
    n15590, n15591, n15592, n15593, n15594, n15596, n15597, n15598, n15599,
    n15600, n15601, n15602, n15603, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
    n15630, n15632, n15633, n15634, n15635, n15636, n15638, n15639, n15640,
    n15641, n15642, n15644, n15645, n15646, n15647, n15648, n15650, n15651,
    n15652, n15653, n15654, n15656, n15657, n15658, n15659, n15660, n15662,
    n15663, n15664, n15665, n15666, n15668, n15669, n15670, n15671, n15672,
    n15674, n15675, n15676, n15677, n15678, n15680, n15681, n15682, n15683,
    n15684, n15686, n15687, n15688, n15689, n15690, n15692, n15693, n15694,
    n15695, n15696, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
    n15716, n15717, n15718, n15719, n15720, n15722, n15723, n15724, n15725,
    n15726, n15728, n15729, n15730, n15731, n15732, n15734, n15735, n15736,
    n15737, n15738, n15740, n15741, n15742, n15743, n15744, n15746, n15747,
    n15748, n15749, n15750, n15752, n15753, n15754, n15755, n15756, n15758,
    n15759, n15760, n15761, n15762, n15764, n15765, n15766, n15767, n15768,
    n15770, n15771, n15772, n15773, n15774, n15776, n15777, n15778, n15779,
    n15780, n15782, n15783, n15784, n15785, n15786, n15788, n15789, n15790,
    n15791, n15792, n15794, n15795, n15796, n15797, n15798, n15800, n15801,
    n15802, n15803, n15804, n15806, n15807, n15808, n15809, n15810, n15812,
    n15813, n15814, n15815, n15816, n15818, n15819, n15820, n15821, n15822,
    n15824, n15825, n15826, n15827, n15828, n15830, n15831, n15832, n15833,
    n15834, n15836, n15837, n15838, n15839, n15840, n15842, n15843, n15844,
    n15845, n15846, n15848, n15849, n15850, n15851, n15852, n15854, n15855,
    n15856, n15857, n15858, n15860, n15861, n15862, n15863, n15864, n15866,
    n15867, n15868, n15869, n15870, n15872, n15873, n15874, n15875, n15876,
    n15878, n15879, n15880, n15881, n15882, n15884, n15885, n15886, n15887,
    n15888, n15890, n15891, n15892, n15893, n15894, n15896, n15897, n15898,
    n15899, n15900, n15902, n15903, n15904, n15905, n15906, n15908, n15909,
    n15910, n15911, n15912, n15914, n15915, n15916, n15917, n15918, n15920,
    n15921, n15922, n15923, n15924, n15926, n15927, n15928, n15929, n15930,
    n15932, n15933, n15934, n15935, n15936, n15938, n15939, n15940, n15941,
    n15942, n15944, n15945, n15946, n15947, n15948, n15950, n15951, n15952,
    n15953, n15954, n15956, n15957, n15958, n15959, n15960, n15962, n15963,
    n15964, n15965, n15966, n15968, n15969, n15970, n15971, n15972, n15974,
    n15975, n15976, n15977, n15978, n15980, n15981, n15982, n15983, n15984,
    n15986, n15987, n15988, n15989, n15990, n15992, n15993, n15994, n15995,
    n15996, n15998, n15999, n16000, n16001, n16002, n16004, n16005, n16006,
    n16007, n16008, n16010, n16011, n16012, n16013, n16014, n16016, n16017,
    n16018, n16019, n16020, n16022, n16023, n16024, n16025, n16026, n16028,
    n16029, n16030, n16031, n16032, n16034, n16035, n16036, n16037, n16038,
    n16040, n16041, n16042, n16043, n16044, n16046, n16047, n16048, n16049,
    n16050, n16052, n16053, n16054, n16055, n16056, n16058, n16059, n16060,
    n16061, n16062, n16064, n16065, n16066, n16067, n16068, n16070, n16071,
    n16072, n16073, n16074, n16076, n16077, n16078, n16079, n16080, n16082,
    n16083, n16084, n16085, n16086, n16088, n16089, n16090, n16091, n16092,
    n16094, n16095, n16096, n16097, n16098, n16100, n16101, n16102, n16103,
    n16104, n16106, n16107, n16108, n16109, n16110, n16112, n16113, n16114,
    n16115, n16116, n16118, n16119, n16120, n16121, n16122, n16124, n16125,
    n16126, n16127, n16128, n16130, n16131, n16132, n16133, n16134, n16136,
    n16137, n16138, n16139, n16140, n16141, n16143, n16144, n16145, n16146,
    n16147, n16149, n16150, n16151, n16152, n16153, n16155, n16156, n16157,
    n16158, n16159, n16161, n16162, n16163, n16164, n16165, n16167, n16168,
    n16169, n16170, n16171, n16173, n16174, n16175, n16176, n16177, n16179,
    n16180, n16181, n16182, n16183, n16185, n16186, n16187, n16188, n16189,
    n16191, n16192, n16193, n16194, n16195, n16197, n16198, n16199, n16200,
    n16201, n16203, n16204, n16205, n16206, n16207, n16209, n16210, n16211,
    n16212, n16213, n16215, n16216, n16217, n16218, n16219, n16221, n16222,
    n16223, n16224, n16225, n16227, n16228, n16229, n16230, n16231, n16233,
    n16234, n16235, n16236, n16237, n16239, n16240, n16241, n16242, n16243,
    n16245, n16246, n16247, n16248, n16249, n16251, n16252, n16253, n16254,
    n16255, n16257, n16258, n16259, n16260, n16261, n16263, n16264, n16265,
    n16266, n16267, n16269, n16270, n16271, n16272, n16273, n16275, n16276,
    n16277, n16278, n16279, n16281, n16282, n16283, n16284, n16285, n16287,
    n16288, n16289, n16290, n16291, n16293, n16294, n16295, n16296, n16297,
    n16299, n16300, n16301, n16302, n16303, n16305, n16306, n16307, n16308,
    n16309, n16311, n16312, n16313, n16314, n16315, n16317, n16318, n16319,
    n16320, n16321, n16323, n16324, n16325, n16326, n16327, n16329, n16330,
    n16331, n16332, n16333, n16335, n16336, n16337, n16338, n16339, n16341,
    n16342, n16343, n16344, n16345, n16347, n16348, n16349, n16350, n16351,
    n16353, n16354, n16355, n16356, n16357, n16359, n16360, n16361, n16362,
    n16363, n16365, n16366, n16367, n16368, n16369, n16371, n16372, n16373,
    n16374, n16375, n16377, n16378, n16379, n16380, n16381, n16383, n16384,
    n16385, n16386, n16387, n16389, n16390, n16391, n16392, n16393, n16395,
    n16396, n16397, n16398, n16399, n16401, n16402, n16403, n16404, n16405,
    n16407, n16408, n16409, n16410, n16411, n16413, n16414, n16415, n16416,
    n16417, n16419, n16420, n16421, n16422, n16423, n16425, n16426, n16427,
    n16428, n16429, n16431, n16432, n16433, n16434, n16435, n16437, n16438,
    n16439, n16440, n16441, n16443, n16444, n16445, n16446, n16447, n16449,
    n16450, n16451, n16452, n16453, n16455, n16456, n16457, n16458, n16459,
    n16461, n16462, n16463, n16464, n16465, n16467, n16468, n16469, n16470,
    n16471, n16473, n16474, n16475, n16476, n16477, n16479, n16480, n16481,
    n16482, n16483, n16485, n16486, n16487, n16488, n16489, n16491, n16492,
    n16493, n16494, n16495, n16497, n16498, n16499, n16500, n16501, n16503,
    n16504, n16505, n16506, n16507, n16509, n16510, n16511, n16512, n16513,
    n16515, n16516, n16517, n16518, n16519, n16521, n16522, n16523, n16524,
    n16525, n16527, n16528, n16529, n16530, n16531, n16533, n16534, n16535,
    n16536, n16537, n16539, n16540, n16541, n16542, n16543, n16545, n16546,
    n16547, n16548, n16549, n16551, n16552, n16553, n16554, n16555, n16557,
    n16558, n16559, n16560, n16561, n16563, n16564, n16565, n16566, n16567,
    n16569, n16570, n16571, n16572, n16573, n16575, n16576, n16577, n16578,
    n16579, n16581, n16582, n16583, n16584, n16585, n16587, n16588, n16589,
    n16590, n16591, n16593, n16594, n16595, n16596, n16597, n16599, n16600,
    n16601, n16602, n16603, n16605, n16606, n16607, n16608, n16609, n16611,
    n16612, n16613, n16614, n16615, n16617, n16618, n16619, n16620, n16621,
    n16623, n16624, n16625, n16626, n16627, n16629, n16630, n16631, n16632,
    n16633, n16635, n16636, n16637, n16638, n16639, n16640, n16642, n16643,
    n16644, n16645, n16646, n16648, n16649, n16650, n16651, n16652, n16654,
    n16655, n16656, n16657, n16658, n16660, n16661, n16662, n16663, n16664,
    n16666, n16667, n16668, n16669, n16670, n16672, n16673, n16674, n16675,
    n16676, n16678, n16679, n16680, n16681, n16682, n16684, n16685, n16686,
    n16687, n16688, n16690, n16691, n16692, n16693, n16694, n16696, n16697,
    n16698, n16699, n16700, n16702, n16703, n16704, n16705, n16706, n16708,
    n16709, n16710, n16711, n16712, n16714, n16715, n16716, n16717, n16718,
    n16720, n16721, n16722, n16723, n16724, n16726, n16727, n16728, n16729,
    n16730, n16732, n16733, n16734, n16735, n16736, n16738, n16739, n16740,
    n16741, n16742, n16744, n16745, n16746, n16747, n16748, n16750, n16751,
    n16752, n16753, n16754, n16756, n16757, n16758, n16759, n16760, n16762,
    n16763, n16764, n16765, n16766, n16768, n16769, n16770, n16771, n16772,
    n16774, n16775, n16776, n16777, n16778, n16780, n16781, n16782, n16783,
    n16784, n16786, n16787, n16788, n16789, n16790, n16792, n16793, n16794,
    n16795, n16796, n16798, n16799, n16800, n16801, n16802, n16804, n16805,
    n16806, n16807, n16808, n16810, n16811, n16812, n16813, n16814, n16816,
    n16817, n16818, n16819, n16820, n16822, n16823, n16824, n16825, n16826,
    n16828, n16829, n16830, n16831, n16832, n16834, n16835, n16836, n16837,
    n16838, n16840, n16841, n16842, n16843, n16844, n16846, n16847, n16848,
    n16849, n16850, n16852, n16853, n16854, n16855, n16856, n16858, n16859,
    n16860, n16861, n16862, n16864, n16865, n16866, n16867, n16868, n16870,
    n16871, n16872, n16873, n16874, n16875, n16877, n16878, n16879, n16880,
    n16881, n16883, n16884, n16885, n16886, n16887, n16889, n16890, n16891,
    n16892, n16893, n16895, n16896, n16897, n16898, n16899, n16901, n16902,
    n16903, n16904, n16905, n16907, n16908, n16909, n16910, n16911, n16913,
    n16914, n16915, n16916, n16917, n16919, n16920, n16921, n16922, n16923,
    n16925, n16926, n16927, n16928, n16929, n16931, n16932, n16933, n16934,
    n16935, n16937, n16938, n16939, n16940, n16941, n16943, n16944, n16945,
    n16946, n16947, n16949, n16950, n16951, n16952, n16953, n16955, n16956,
    n16957, n16958, n16959, n16961, n16962, n16963, n16964, n16965, n16967,
    n16968, n16969, n16970, n16971, n16973, n16974, n16975, n16976, n16977,
    n16979, n16980, n16981, n16982, n16983, n16985, n16986, n16987, n16988,
    n16989, n16991, n16992, n16993, n16994, n16995, n16997, n16998, n16999,
    n17000, n17001, n17003, n17004, n17005, n17006, n17007, n17009, n17010,
    n17011, n17012, n17013, n17015, n17016, n17017, n17018, n17019, n17020,
    n17022, n17023, n17024, n17025, n17026, n17028, n17029, n17030, n17031,
    n17032, n17034, n17035, n17036, n17037, n17038, n17040, n17041, n17042,
    n17043, n17044, n17046, n17047, n17048, n17049, n17050, n17052, n17053,
    n17054, n17055, n17056, n17058, n17059, n17060, n17061, n17062, n17064,
    n17065, n17066, n17067, n17068, n17070, n17071, n17072, n17073, n17074,
    n17076, n17077, n17078, n17079, n17080, n17082, n17083, n17084, n17085,
    n17086, n17088, n17089, n17090, n17091, n17092, n17094, n17095, n17096,
    n17097, n17098, n17100, n17101, n17102, n17103, n17104, n17106, n17107,
    n17108, n17109, n17110, n17112, n17113, n17114, n17115, n17116, n17118,
    n17119, n17120, n17121, n17122, n17124, n17125, n17126, n17127, n17128,
    n17130, n17131, n17132, n17133, n17134, n17136, n17137, n17138, n17139,
    n17140, n17142, n17143, n17144, n17145, n17146, n17148, n17149, n17150,
    n17151, n17152, n17154, n17155, n17156, n17157, n17158, n17159, n17161,
    n17162, n17163, n17164, n17165, n17167, n17168, n17169, n17170, n17171,
    n17173, n17174, n17175, n17176, n17177, n17179, n17180, n17181, n17182,
    n17183, n17185, n17186, n17187, n17188, n17189, n17191, n17192, n17193,
    n17194, n17195, n17197, n17198, n17199, n17200, n17201, n17203, n17204,
    n17205, n17206, n17207, n17209, n17210, n17211, n17212, n17213, n17215,
    n17216, n17217, n17218, n17219, n17221, n17222, n17223, n17224, n17225,
    n17227, n17228, n17229, n17230, n17231, n17233, n17234, n17235, n17236,
    n17237, n17239, n17240, n17241, n17242, n17243, n17245, n17246, n17247,
    n17248, n17249, n17251, n17252, n17253, n17254, n17255, n17257, n17258,
    n17259, n17260, n17261, n17263, n17264, n17265, n17266, n17267, n17269,
    n17270, n17271, n17272, n17273, n17275, n17276, n17277, n17278, n17279,
    n17281, n17282, n17283, n17284, n17285, n17287, n17288, n17289, n17290,
    n17291, n17293, n17294, n17295, n17296, n17297, n17299, n17300, n17301,
    n17302, n17303, n17305, n17306, n17307, n17308, n17309, n17311, n17312,
    n17313, n17314, n17315, n17317, n17318, n17319, n17320, n17321, n17323,
    n17324, n17325, n17326, n17327, n17329, n17330, n17331, n17332, n17333,
    n17335, n17336, n17337, n17338, n17339, n17341, n17342, n17343, n17344,
    n17345, n17347, n17348, n17349, n17350, n17351, n17353, n17354, n17355,
    n17356, n17357, n17359, n17360, n17361, n17362, n17363, n17365, n17366,
    n17367, n17368, n17369, n17371, n17372, n17373, n17374, n17375, n17377,
    n17378, n17379, n17380, n17381, n17383, n17384, n17385, n17386, n17387,
    n17389, n17390, n17391, n17392, n17393, n17395, n17396, n17397, n17398,
    n17399, n17401, n17402, n17403, n17404, n17405, n17407, n17408, n17409,
    n17410, n17411, n17413, n17414, n17415, n17416, n17417, n17419, n17420,
    n17421, n17422, n17423, n17425, n17426, n17427, n17428, n17429, n17431,
    n17432, n17433, n17434, n17435, n17437, n17438, n17439, n17440, n17441,
    n17442, n17444, n17445, n17446, n17447, n17448, n17450, n17451, n17452,
    n17453, n17454, n17456, n17457, n17458, n17459, n17460, n17463, n17464,
    n17465, n17466, n17467, n17469, n17470, n17471, n17472, n17473, n17475,
    n17476, n17477, n17478, n17479, n17481, n17482, n17483, n17484, n17485,
    n17487, n17488, n17489, n17490, n17491, n17493, n17494, n17495, n17496,
    n17497, n17499, n17500, n17501, n17502, n17503, n17505, n17506, n17507,
    n17508, n17509, n17511, n17512, n17513, n17514, n17515, n17517, n17518,
    n17519, n17520, n17521, n17523, n17524, n17525, n17526, n17527, n17529,
    n17530, n17531, n17532, n17533, n17535, n17536, n17537, n17538, n17539,
    n17541, n17542, n17543, n17544, n17545, n17547, n17548, n17549, n17550,
    n17551, n17553, n17554, n17555, n17556, n17557, n17559, n17560, n17561,
    n17562, n17563, n17565, n17566, n17567, n17568, n17569, n17571, n17573,
    n17574, n17575, n17576, n17577, n17579, n17580, n17581, n17582, n17583,
    n17585, n17586, n17587, n17588, n17589, n17591, n17592, n17593, n17594,
    n17595, n17597, n17598, n17599, n17600, n17601, n17603, n17604, n17605,
    n17606, n17607, n17609, n17610, n17611, n17612, n17613, n17615, n17616,
    n17617, n17618, n17619, n17621, n17622, n17623, n17624, n17625, n17627,
    n17628, n17629, n17630, n17631, n17633, n17634, n17635, n17636, n17637,
    n17639, n17640, n17641, n17642, n17643, n17645, n17646, n17647, n17648,
    n17649, n17651, n17652, n17653, n17654, n17655, n17657, n17658, n17659,
    n17660, n17661, n17663, n17664, n17665, n17666, n17667, n17669, n17670,
    n17671, n17672, n17673, n17675, n17676, n17677, n17678, n17679, n17681,
    n17682, n17683, n17684, n17685, n17687, n17688, n17689, n17690, n17691,
    n17693, n17694, n17695, n17696, n17697, n17699, n17700, n17701, n17702,
    n17703, n17705, n17706, n17707, n17708, n17709, n17711, n17712, n17713,
    n17714, n17715, n17717, n17718, n17719, n17720, n17721, n17723, n17724,
    n17725, n17726, n17727, n17729, n17730, n17731, n17732, n17733, n17735,
    n17736, n17737, n17738, n17739, n17741, n17742, n17743, n17744, n17745,
    n17747, n17748, n17749, n17750, n17751, n17753, n17754, n17755, n17756,
    n17757, n17759, n17760, n17761, n17762, n17763, n17765, n17766, n17767,
    n17768, n17769, n17771, n17772, n17773, n17774, n17775, n17777, n17778,
    n17779, n17780, n17781, n17783, n17784, n17785, n17786, n17787, n17789,
    n17790, n17791, n17792, n17793, n17795, n17796, n17797, n17798, n17799,
    n17801, n17802, n17803, n17804, n17805, n17807, n17808, n17809, n17810,
    n17811, n17813, n17814, n17815, n17816, n17817, n17819, n17820, n17821,
    n17822, n17823, n17825, n17826, n17827, n17828, n17829, n17831, n17832,
    n17833, n17834, n17835, n17837, n17838, n17839, n17840, n17841, n17843,
    n17844, n17845, n17846, n17847, n17848, n17849, n17851, n17852, n17853,
    n17854, n17855, n17856, n17858, n17859, n17860, n17861, n17862, n17864,
    n17865, n17866, n17867, n17868, n17870, n17871, n17872, n17873, n17874,
    n17876, n17877, n17878, n17879, n17880, n17882, n17883, n17884, n17885,
    n17886, n17888, n17889, n17890, n17891, n17892, n17894, n17895, n17896,
    n17897, n17898, n17900, n17901, n17902, n17903, n17904, n17906, n17907,
    n17908, n17909, n17910, n17912, n17913, n17914, n17915, n17916, n17918,
    n17919, n17920, n17921, n17922, n17924, n17925, n17926, n17927, n17928,
    n17930, n17931, n17932, n17933, n17934, n17936, n17937, n17938, n17939,
    n17940, n17942, n17943, n17944, n17945, n17946, n17948, n17949, n17950,
    n17951, n17952, n17954, n17955, n17956, n17957, n17958, n17960, n17961,
    n17962, n17963, n17964, n17966, n17967, n17968, n17969, n17970, n17972,
    n17973, n17974, n17975, n17976, n17978, n17979, n17980, n17981, n17982,
    n17984, n17985, n17986, n17987, n17988, n17990, n17991, n17992, n17993,
    n17994, n17996, n17997, n17999, n18000, n18001, n18002, n18003, n18004,
    n18006, n18007, n18008, n18009, n18010, n18012, n18013, n18014, n18015,
    n18016, n18018, n18019, n18020, n18021, n18022, n18024, n18025, n18026,
    n18027, n18028, n18030, n18031, n18032, n18033, n18034, n18036, n18037,
    n18038, n18039, n18040, n18042, n18043, n18044, n18045, n18046, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054, n18056, n18057, n18058,
    n18059, n18060, n18061, n18062, n18063, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18074, n18075, n18076, n18077, n18078,
    n18079, n18080, n18081, n18083, n18084, n18085, n18086, n18087, n18088,
    n18089, n18090, n18092, n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
    n18110, n18112, n18113, n18114, n18115, n18116, n18118, n18119, n18120,
    n18121, n18122, n18124, n18125, n18126, n18127, n18128, n18130, n18131,
    n18132, n18133, n18134, n18136, n18137, n18138, n18139, n18140, n18142,
    n18143, n18144, n18145, n18146, n18148, n18149, n18150, n18151, n18152,
    n18154, n18155, n18156, n18157, n18158, n18160, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18169, n18170, n18171, n18172, n18173,
    n18175, n18176, n18177, n18178, n18179, n18181, n18182, n18183, n18184,
    n18185, n18187, n18188, n18189, n18190, n18191, n18193, n18194, n18195,
    n18196, n18197, n18199, n18200, n18201, n18202, n18203, n18205, n18206,
    n18207, n18208, n18209, n18211, n18212, n18213, n18214, n18215, n18216,
    n18217, n18218, n18220, n18221, n18222, n18223, n18224, n18226, n18227,
    n18228, n18229, n18230, n18232, n18233, n18234, n18235, n18236, n18238,
    n18239, n18240, n18241, n18242, n18244, n18245, n18246, n18247, n18248,
    n18250, n18251, n18252, n18253, n18254, n18256, n18257, n18258, n18259,
    n18260, n18262, n18263, n18264, n18265, n18266, n18268, n18269, n18270,
    n18271, n18272, n18274, n18275, n18276, n18277, n18278, n18280, n18281,
    n18282, n18283, n18284, n18286, n18287, n18288, n18289, n18290, n18292,
    n18293, n18294, n18295, n18296, n18298, n18299, n18300, n18301, n18302,
    n18304, n18305, n18306, n18307, n18308, n18310, n18311, n18312, n18313,
    n18314, n18316, n18317, n18318, n18319, n18320, n18322, n18323, n18324,
    n18325, n18326, n18328, n18329, n18330, n18331, n18332, n18334, n18335,
    n18336, n18337, n18338, n18340, n18341, n18342, n18343, n18344, n18346,
    n18347, n18348, n18349, n18350, n18352, n18353, n18354, n18355, n18356,
    n18358, n18359, n18360, n18361, n18362, n18364, n18365, n18366, n18367,
    n18368, n18370, n18371, n18372, n18373, n18374, n18376, n18377, n18378,
    n18379, n18380, n18382, n18383, n18384, n18385, n18386, n18388, n18389,
    n18390, n18391, n18392, n18394, n18395, n18396, n18397, n18398, n18400,
    n18401, n18402, n18403, n18404, n18406, n18407, n18408, n18409, n18410,
    n18412, n18413, n18414, n18415, n18416, n18418, n18419, n18420, n18421,
    n18422, n18424, n18425, n18426, n18427, n18428, n18430, n18431, n18432,
    n18433, n18434, n18436, n18437, n18438, n18439, n18440, n18442, n18443,
    n18444, n18445, n18446, n18448, n18449, n18450, n18451, n18452, n18454,
    n18455, n18456, n18457, n18458, n18460, n18461, n18462, n18463, n18464,
    n18466, n18467, n18468, n18469, n18470, n18472, n18473, n18474, n18475,
    n18476, n18478, n18479, n18480, n18481, n18482, n18484, n18485, n18486,
    n18487, n18488, n18490, n18491, n18492, n18493, n18494, n18496, n18497,
    n18498, n18499, n18500, n18502, n18503, n18504, n18505, n18506, n18508,
    n18509, n18510, n18511, n18512, n18514, n18515, n18516, n18517, n18518,
    n18520, n18521, n18522, n18523, n18524, n18526, n18527, n18528, n18529,
    n18530, n18532, n18533, n18534, n18535, n18536, n18538, n18539, n18540,
    n18541, n18542, n18544, n18545, n18546, n18547, n18548, n18550, n18551,
    n18552, n18553, n18554, n18556, n18557, n18558, n18559, n18560, n18562,
    n18563, n18564, n18565, n18566, n18568, n18569, n18570, n18571, n18572,
    n18574, n18575, n18576, n18577, n18578, n18580, n18581, n18582, n18583,
    n18584, n18586, n18587, n18588, n18589, n18590, n18592, n18593, n18594,
    n18595, n18596, n18598, n18599, n18600, n18601, n18602, n18604, n18605,
    n18606, n18607, n18608, n18610, n18611, n18612, n18613, n18614, n18616,
    n18617, n18618, n18619, n18620, n18622, n18623, n18624, n18625, n18626,
    n18628, n18629, n18630, n18631, n18632, n18634, n18635, n18636, n18637,
    n18638, n18640, n18641, n18642, n18643, n18644, n18646, n18647, n18648,
    n18649, n18650, n18652, n18653, n18654, n18655, n18656, n18658, n18659,
    n18660, n18661, n18662, n18664, n18665, n18666, n18667, n18668, n18670,
    n18671, n18672, n18673, n18674, n18676, n18677, n18678, n18679, n18680,
    n18682, n18683, n18684, n18685, n18686, n18688, n18689, n18690, n18691,
    n18692, n18694, n18695, n18696, n18697, n18698, n18700, n18701, n18702,
    n18703, n18704, n18706, n18707, n18708, n18709, n18710, n18712, n18713,
    n18714, n18715, n18716, n18718, n18719, n18720, n18721, n18722, n18724,
    n18725, n18726, n18727, n18728, n18730, n18731, n18732, n18733, n18734,
    n18736, n18737, n18738, n18739, n18740, n18742, n18743, n18744, n18745,
    n18746, n18748, n18749, n18750, n18751, n18752, n18754, n18755, n18756,
    n18757, n18758, n18760, n18761, n18762, n18763, n18764, n18766, n18767,
    n18768, n18769, n18770, n18772, n18773, n18774, n18775, n18776, n18778,
    n18779, n18780, n18781, n18782, n18784, n18785, n18786, n18787, n18788,
    n18790, n18791, n18792, n18793, n18794, n18796, n18797, n18798, n18799,
    n18800, n18802, n18803, n18804, n18805, n18806, n18808, n18809, n18810,
    n18811, n18812, n18814, n18815, n18816, n18817, n18818, n18820, n18821,
    n18822, n18823, n18824, n18826, n18827, n18828, n18829, n18830, n18832,
    n18833, n18834, n18835, n18836, n18838, n18839, n18840, n18841, n18842,
    n18844, n18845, n18846, n18847, n18848, n18850, n18851, n18852, n18853,
    n18854, n18856, n18857, n18858, n18859, n18860, n18862, n18863, n18864,
    n18865, n18866, n18868, n18869, n18870, n18871, n18872, n18874, n18875,
    n18876, n18877, n18878, n18880, n18881, n18882, n18883, n18884, n18886,
    n18887, n18888, n18889, n18890, n18892, n18893, n18894, n18895, n18896,
    n18898, n18899, n18900, n18901, n18902, n18904, n18905, n18906, n18907,
    n18908, n18910, n18911, n18912, n18913, n18914, n18916, n18917, n18918,
    n18919, n18920, n18922, n18923, n18924, n18925, n18926, n18928, n18929,
    n18930, n18931, n18932, n18934, n18935, n18936, n18937, n18938, n18940,
    n18941, n18942, n18944, n18945, n18946, n18947, n18949, n18950, n18952,
    n18953, n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18965, n18966, n18968, n18969, n18971, n18972, n18974, n18975,
    n18977, n18978, n18980, n18981, n18983, n18984, n18986, n18987, n18989,
    n18990, n18992, n18993, n18995, n18996, n18998, n18999, n19001, n19002,
    n19004, n19005, n19007, n19008, n19010, n19011, n19013, n19014, n19016,
    n19017, n19019, n19020, n19022, n19023, n19024, n19025, n19026, n19028,
    n19030, n19031, n19033, n19034, n19036, n19037, n19039, n19040, n19042,
    n19043, n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19061, n19062,
    n19064, n19065, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
    n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19083,
    n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19092, n19093,
    n19094, n19095, n19096, n19097, n19098, n19099, n19101, n19102, n19103,
    n19104, n19105, n19107, n19108, n19109, n19111, n19112, n19113, n19114,
    n19115, n19116, n19118, n19119, n19121, n19122, n19124, n19125, n19127,
    n19128, n19130, n19131, n19132, n19133, n19134, n19136, n19137, n19138,
    n19139, n19140, n19142, n19143, n19144, n19145, n19146, n19148, n19149,
    n19151, n19152, n19153, n19154, n19155, n19156, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19179, n19180,
    n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19194, n19195, n19196, n19197, n19198, n19200,
    n19201, n19203, n19204, n19205, n19206, n19207, n19208, n19210, n19211,
    n19213, n19214, n19216, n19217, n19219, n19220, n19222, n19223, n19225,
    n19226, n19227, n19228, n19229, n19231, n19232, n19233, n19234, n19235,
    n19237, n19238, n19239, n19240, n19241, n19243, n19244, n19246, n19247,
    n19249, n19250, n19252, n19254, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19263, n19264, n19265, n19266, n19268, n19269, n19270,
    n19271, n19272, n19274, n19275, n19276, n19277, n19278, n19280, n19281,
    n19282, n19283, n19284, n19286, n19287, n19288, n19289, n19290, n19292,
    n19293, n19294, n19295, n19296, n19298, n19299, n19300, n19301, n19302,
    n19304, n19305, n19306, n19307, n19308, n19310, n19311, n19312, n19313,
    n19314, n19316, n19317, n19318, n19319, n19320, n19322, n19323, n19324,
    n19325, n19326, n19328, n19329, n19330, n19331, n19332, n19334, n19335,
    n19337, n19338, n19340, n19341, n19343, n19344, n19345, n19346, n19347,
    n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
    n19357, n19359, n19360, n19362, n19363, n19365, n19366, n19367, n19368,
    n19369, n19371, n19372, n19373, n19374, n19375, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19384, n19386, n19387, n19388, n19389,
    n19390, n19391, n19392, n19393, n19395, n19396, n19397, n19398, n19399,
    n19400, n19402, n19403, n19404, n19405, n19406, n19408, n19409, n19411,
    n19412, n19413, n19414, n19415, n19417, n19418, n19419, n19420, n19421,
    n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431,
    n19432, n19433, n19435, n19436, n19437, n19438, n19439, n19441, n19442,
    n19444, n19445, n19446, n19447, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
    n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19478, n19479, n19480, n19481,
    n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19491,
    n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
    n19502, n19504, n19505, n19506, n19507, n19508, n19509, n19511, n19512,
    n19513, n19514, n19515, n19516, n19517, n19519, n19520, n19521, n19522,
    n19523, n19524, n19525, n19526, n19527, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19537, n19538, n19539, n19540, n19541, n19542,
    n19544, n19545, n19546, n19547, n19548, n19549, n19551, n19552, n19553,
    n19554, n19555, n19557, n19558, n19560, n19561, n19563, n19564, n19566,
    n19567, n19569, n19570, n19572, n19573, n19575, n19576, n19577, n19578,
    n19579, n19581, n19582, n19583, n19584, n19585, n19587, n19588, n19590,
    n19591, n19593, n19594, n19595, n19596, n19597, n19599, n19600, n19602,
    n19603, n19604, n19605, n19606, n19607, n19608, n19610, n19611, n19612,
    n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19621, n19623,
    n19624, n19625, n19626, n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19636, n19637, n19639, n19640, n19642, n19643, n19645, n19646,
    n19648, n19650, n19651, n19653, n19654, n19655, n19656, n19657, n19659,
    n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
    n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19677, n19678,
    n19679, n19681, n19682, n19683, n19685, n19686, n19688, n19689, n19691,
    n19692, n19694, n19695, n19697, n19698, n19700, n19701, n19703, n19704,
    n19706, n19707, n19709, n19710, n19712, n19713, n19715, n19716, n19718,
    n19719, n19721, n19722, n19724, n19725, n19727, n19728, n19730, n19731,
    n19733, n19734, n19736, n19737, n19739, n19740, n19742, n19743, n19745,
    n19746, n19748, n19749, n19751, n19752, n19755, n19756, n19757, n19758,
    n19759, n19760, n19761, n19762, n19763, n19764, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19774, n19775, n19776, n19777, n19778,
    n19779, n19781, n19782, n19784, n19785, n19787, n19788, n19789, n19790,
    n19791, n19792, n19794, n19795, n19796, n19797, n19798, n19799, n19801,
    n19802, n19803, n19805, n19806, n19808, n19809, n19811, n19812, n19814,
    n19815, n19816, n19817, n19818, n19821, n19822, n19823, n19824, n19825,
    n19826, n19827, n19829, n19830, n19832, n19833, n19834, n19836, n19837,
    n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19847, n19848,
    n19850, n19851, n19852, n19853, n19854, n19855, n19857, n19858, n19859,
    n19860, n19861, n19862, n19864, n19865, n19867, n19868, n19870, n19871,
    n19873, n19874, n19876, n19877, n19879, n19880, n19882, n19883, n19885,
    n19886, n19888, n19889, n19891, n19892, n19894, n19895, n19897, n19898,
    n19899, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
    n19909, n19911, n19912, n19914, n19915, n19916, n19917, n19918, n19919,
    n19920, n19921, n19922, n19923, n19924, n19926, n19927, n19928, n19929,
    n19930, n19931, n19932, n19934, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
    n19950, n19951, n19952, n19954, n19955, n19956, n19957, n19958, n19959,
    n19960, n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968,
    n19969, n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
    n19978, n19979, n19980, n19981, n19983, n19984, n19985, n19986, n19987,
    n19988, n19989, n19990, n19991, n19992, n19994, n19995, n19996, n19998,
    n19999, n20000, n20001, n20002, n20003, n20005, n20006, n20007, n20008,
    n20009, n20010, n20011, n20012, n20013, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20025, n20026, n20028, n20029,
    n20030, n20031, n20032, n20033, n20034, n20036, n20037, n20038, n20040,
    n20041, n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
    n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
    n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
    n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
    n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
    n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103,
    n20104, n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112,
    n20113, n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
    n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
    n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
    n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20172, n20173, n20174, n20175, n20176,
    n20177, n20178, n20179, n20180, n20182, n20183, n20184, n20185, n20186,
    n20187, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
    n20197, n20199, n20200, n20201, n20202, n20203, n20205, n20206, n20208,
    n20209, n20210, n20212, n20213, n20215, n20216, n20218, n20219, n20221,
    n20222, n20224, n20225, n20227, n20228, n20230, n20231, n20232, n20233,
    n20235, n20236, n20238, n20239, n20241, n20242, n20243, n20244, n20246,
    n20247, n20248, n20249, n20251, n20252, n20253, n20254, n20256, n20257,
    n20258, n20260, n20261, n20262, n20263, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
    n20278, n20279, n20281, n20282, n20283, n20284, n20286, n20287, n20288,
    n20289, n20291, n20292, n20293, n20294, n20296, n20297, n20299, n20300,
    n20301, n20302, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
    n20312, n20313, n20314, n20316, n20319, n20320, n20321, n20323, n20324,
    n20325, n20327, n20328, n20330, n20331, n20332, n20333, n20334, n20335,
    n20337, n20338, n20339, n20340, n20341, n20342, n20344, n20345, n20346,
    n20347, n20348, n20350, n20351, n20353, n20354, n20355, n20356, n20357,
    n20359, n20360, n20361, n20362, n20363, n20365, n20366, n20367, n20368,
    n20369, n20371, n20372, n20373, n20374, n20375, n20377, n20378, n20379,
    n20380, n20381, n20383, n20384, n20385, n20386, n20387, n20389, n20390,
    n20391, n20392, n20393, n20395, n20396, n20397, n20398, n20399, n20401,
    n20402, n20403, n20404, n20405, n20407, n20408, n20409, n20410, n20411,
    n20413, n20414, n20415, n20416, n20417, n20419, n20420, n20421, n20422,
    n20423, n20424, n20426, n20427, n20429, n20430, n20432, n20433, n20434,
    n20435, n20436, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
    n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20455,
    n20456, n20457, n20458, n20459, n20460, n20462, n20463, n20464, n20465,
    n20466, n20467, n20469, n20470, n20471, n20472, n20473, n20475, n20476,
    n20477, n20478, n20479, n20481, n20482, n20483, n20484, n20486, n20487,
    n20488, n20489, n20491, n20492, n20494, n20495, n20497, n20498, n20500,
    n20501, n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20511,
    n20512, n20513, n20514, n20515, n20517, n20518, n20519, n20520, n20521,
    n20523, n20524, n20525, n20526, n20527, n20529, n20530, n20531, n20532,
    n20533, n20535, n20536, n20537, n20538, n20539, n20541, n20542, n20543,
    n20544, n20545, n20547, n20548, n20549, n20550, n20551, n20553, n20554,
    n20555, n20556, n20557, n20559, n20560, n20561, n20562, n20563, n20565,
    n20566, n20567, n20568, n20569, n20571, n20572, n20573, n20574, n20575,
    n20577, n20578, n20579, n20580, n20581, n20583, n20584, n20585, n20586,
    n20587, n20589, n20590, n20591, n20592, n20593, n20595, n20596, n20597,
    n20598, n20599, n20601, n20602, n20603, n20604, n20605, n20607, n20608,
    n20609, n20610, n20611, n20613, n20614, n20615, n20616, n20617, n20619,
    n20620, n20621, n20622, n20623, n20624, n20626, n20627, n20628, n20629,
    n20630, n20632, n20633, n20634, n20635, n20636, n20638, n20639, n20640,
    n20641, n20642, n20644, n20645, n20646, n20647, n20648, n20650, n20651,
    n20652, n20653, n20654, n20656, n20657, n20658, n20659, n20660, n20662,
    n20663, n20664, n20665, n20666, n20668, n20669, n20670, n20671, n20672,
    n20674, n20675, n20676, n20677, n20678, n20680, n20681, n20682, n20683,
    n20684, n20686, n20687, n20688, n20689, n20690, n20692, n20693, n20694,
    n20695, n20696, n20698, n20699, n20700, n20701, n20702, n20704, n20705,
    n20706, n20707, n20708, n20710, n20711, n20712, n20713, n20714, n20716,
    n20717, n20718, n20719, n20720, n20722, n20723, n20724, n20725, n20726,
    n20728, n20729, n20730, n20731, n20732, n20734, n20735, n20736, n20737,
    n20738, n20740, n20741, n20742, n20743, n20744, n20746, n20747, n20748,
    n20749, n20750, n20752, n20753, n20754, n20755, n20756, n20757, n20759,
    n20760, n20761, n20762, n20763, n20765, n20766, n20767, n20768, n20769,
    n20771, n20772, n20773, n20774, n20775, n20777, n20778, n20779, n20780,
    n20781, n20783, n20784, n20785, n20786, n20787, n20789, n20790, n20791,
    n20792, n20793, n20795, n20796, n20797, n20798, n20799, n20801, n20802,
    n20803, n20804, n20805, n20807, n20808, n20809, n20810, n20811, n20813,
    n20814, n20815, n20816, n20817, n20819, n20820, n20821, n20822, n20823,
    n20825, n20826, n20827, n20828, n20829, n20831, n20832, n20833, n20834,
    n20835, n20837, n20838, n20839, n20840, n20841, n20843, n20844, n20845,
    n20846, n20847, n20849, n20850, n20851, n20852, n20853, n20855, n20856,
    n20857, n20858, n20859, n20861, n20862, n20863, n20864, n20865, n20867,
    n20868, n20869, n20870, n20871, n20873, n20874, n20875, n20876, n20877,
    n20879, n20880, n20881, n20882, n20883, n20885, n20886, n20887, n20888,
    n20889, n20891, n20892, n20893, n20894, n20895, n20897, n20898, n20899,
    n20900, n20901, n20903, n20904, n20905, n20906, n20907, n20909, n20910,
    n20911, n20912, n20913, n20915, n20916, n20917, n20918, n20919, n20921,
    n20922, n20923, n20924, n20925, n20927, n20928, n20929, n20930, n20931,
    n20933, n20934, n20935, n20936, n20937, n20939, n20940, n20941, n20942,
    n20943, n20945, n20946, n20947, n20948, n20949, n20951, n20952, n20953,
    n20954, n20955, n20957, n20958, n20959, n20960, n20961, n20963, n20964,
    n20965, n20966, n20967, n20969, n20970, n20971, n20972, n20973, n20975,
    n20976, n20977, n20978, n20979, n20981, n20982, n20983, n20984, n20985,
    n20987, n20988, n20989, n20990, n20991, n20993, n20994, n20995, n20996,
    n20997, n20999, n21000, n21001, n21002, n21003, n21005, n21006, n21007,
    n21008, n21009, n21011, n21012, n21013, n21014, n21015, n21016, n21018,
    n21019, n21020, n21021, n21022, n21024, n21025, n21026, n21027, n21028,
    n21030, n21031, n21032, n21033, n21034, n21036, n21037, n21038, n21039,
    n21040, n21042, n21043, n21044, n21045, n21046, n21048, n21049, n21050,
    n21051, n21052, n21054, n21055, n21056, n21057, n21058, n21060, n21061,
    n21062, n21063, n21064, n21066, n21067, n21068, n21069, n21070, n21072,
    n21073, n21074, n21075, n21076, n21078, n21079, n21080, n21081, n21082,
    n21084, n21085, n21086, n21087, n21088, n21090, n21091, n21092, n21093,
    n21094, n21096, n21097, n21098, n21099, n21100, n21102, n21103, n21104,
    n21105, n21106, n21108, n21109, n21110, n21111, n21112, n21114, n21115,
    n21116, n21117, n21118, n21120, n21121, n21122, n21123, n21124, n21126,
    n21127, n21128, n21129, n21130, n21132, n21133, n21134, n21135, n21136,
    n21138, n21139, n21140, n21141, n21142, n21144, n21145, n21146, n21147,
    n21148, n21150, n21151, n21152, n21153, n21154, n21156, n21157, n21158,
    n21159, n21160, n21162, n21163, n21164, n21165, n21166, n21168, n21169,
    n21170, n21171, n21172, n21174, n21175, n21176, n21177, n21178, n21180,
    n21181, n21182, n21183, n21184, n21186, n21187, n21188, n21189, n21190,
    n21192, n21193, n21194, n21195, n21196, n21198, n21199, n21200, n21201,
    n21202, n21204, n21205, n21206, n21207, n21208, n21210, n21211, n21212,
    n21213, n21214, n21216, n21217, n21218, n21219, n21220, n21222, n21223,
    n21224, n21225, n21226, n21228, n21229, n21230, n21231, n21232, n21234,
    n21235, n21236, n21237, n21238, n21240, n21241, n21242, n21243, n21244,
    n21246, n21247, n21248, n21249, n21250, n21252, n21253, n21254, n21255,
    n21256, n21258, n21259, n21260, n21261, n21262, n21264, n21265, n21266,
    n21267, n21268, n21270, n21271, n21272, n21273, n21274, n21276, n21277,
    n21278, n21279, n21280, n21282, n21283, n21284, n21285, n21286, n21288,
    n21289, n21290, n21291, n21292, n21294, n21295, n21296, n21297, n21298,
    n21300, n21301, n21302, n21303, n21304, n21306, n21307, n21308, n21309,
    n21310, n21312, n21313, n21314, n21315, n21316, n21318, n21319, n21320,
    n21321, n21322, n21324, n21325, n21326, n21327, n21328, n21330, n21331,
    n21332, n21333, n21334, n21336, n21337, n21338, n21339, n21340, n21342,
    n21343, n21344, n21345, n21346, n21348, n21349, n21350, n21351, n21352,
    n21354, n21355, n21356, n21357, n21358, n21360, n21361, n21362, n21363,
    n21364, n21366, n21367, n21368, n21369, n21370, n21371, n21373, n21374,
    n21375, n21376, n21377, n21379, n21380, n21381, n21382, n21383, n21385,
    n21386, n21387, n21388, n21389, n21391, n21392, n21393, n21394, n21395,
    n21397, n21398, n21399, n21400, n21401, n21403, n21404, n21405, n21406,
    n21407, n21409, n21410, n21411, n21412, n21413, n21415, n21416, n21417,
    n21418, n21419, n21421, n21422, n21423, n21424, n21425, n21427, n21428,
    n21429, n21430, n21431, n21433, n21434, n21435, n21436, n21437, n21439,
    n21440, n21441, n21442, n21443, n21445, n21446, n21447, n21448, n21449,
    n21451, n21452, n21453, n21454, n21455, n21457, n21458, n21459, n21460,
    n21461, n21463, n21464, n21465, n21466, n21467, n21469, n21470, n21471,
    n21472, n21473, n21475, n21476, n21477, n21478, n21479, n21481, n21482,
    n21483, n21484, n21485, n21487, n21488, n21489, n21490, n21491, n21493,
    n21494, n21495, n21496, n21497, n21499, n21500, n21501, n21502, n21503,
    n21505, n21506, n21507, n21508, n21509, n21511, n21512, n21513, n21514,
    n21515, n21517, n21518, n21519, n21520, n21521, n21523, n21524, n21525,
    n21526, n21527, n21529, n21530, n21531, n21532, n21533, n21535, n21536,
    n21537, n21538, n21539, n21541, n21542, n21543, n21544, n21545, n21547,
    n21548, n21549, n21550, n21551, n21553, n21554, n21555, n21556, n21557,
    n21559, n21560, n21561, n21562, n21563, n21565, n21566, n21567, n21568,
    n21569, n21571, n21572, n21573, n21574, n21575, n21577, n21578, n21579,
    n21580, n21581, n21582, n21584, n21585, n21586, n21587, n21588, n21590,
    n21591, n21592, n21593, n21594, n21596, n21597, n21598, n21599, n21600,
    n21602, n21603, n21604, n21605, n21606, n21608, n21609, n21610, n21611,
    n21612, n21614, n21615, n21616, n21617, n21618, n21620, n21621, n21622,
    n21623, n21624, n21626, n21627, n21628, n21629, n21630, n21632, n21633,
    n21634, n21635, n21636, n21638, n21639, n21640, n21641, n21642, n21644,
    n21645, n21646, n21647, n21648, n21650, n21651, n21652, n21653, n21654,
    n21656, n21657, n21658, n21659, n21660, n21662, n21663, n21664, n21665,
    n21666, n21668, n21669, n21670, n21671, n21672, n21674, n21675, n21676,
    n21677, n21678, n21680, n21681, n21682, n21683, n21684, n21686, n21687,
    n21688, n21689, n21690, n21692, n21693, n21694, n21695, n21696, n21698,
    n21699, n21700, n21701, n21702, n21704, n21705, n21706, n21707, n21708,
    n21710, n21711, n21712, n21713, n21714, n21716, n21717, n21718, n21719,
    n21720, n21722, n21723, n21724, n21725, n21726, n21728, n21729, n21730,
    n21731, n21732, n21734, n21735, n21736, n21737, n21738, n21740, n21741,
    n21742, n21743, n21744, n21746, n21747, n21748, n21749, n21750, n21752,
    n21753, n21754, n21755, n21756, n21758, n21759, n21760, n21761, n21762,
    n21764, n21765, n21766, n21767, n21768, n21770, n21771, n21772, n21773,
    n21774, n21776, n21777, n21778, n21779, n21780, n21782, n21783, n21784,
    n21785, n21786, n21788, n21789, n21790, n21791, n21792, n21794, n21795,
    n21796, n21797, n21798, n21800, n21801, n21802, n21803, n21804, n21806,
    n21807, n21808, n21809, n21810, n21812, n21813, n21814, n21815, n21816,
    n21818, n21819, n21820, n21821, n21822, n21824, n21825, n21826, n21827,
    n21828, n21830, n21831, n21832, n21833, n21834, n21836, n21837, n21838,
    n21839, n21840, n21842, n21843, n21844, n21845, n21846, n21848, n21849,
    n21850, n21851, n21852, n21854, n21855, n21856, n21857, n21858, n21860,
    n21861, n21862, n21863, n21864, n21866, n21867, n21868, n21869, n21870,
    n21872, n21873, n21874, n21875, n21876, n21878, n21879, n21880, n21881,
    n21882, n21884, n21885, n21886, n21887, n21888, n21890, n21891, n21892,
    n21893, n21894, n21896, n21897, n21898, n21899, n21900, n21902, n21903,
    n21904, n21905, n21906, n21908, n21909, n21910, n21911, n21912, n21914,
    n21915, n21916, n21917, n21918, n21920, n21921, n21922, n21923, n21924,
    n21926, n21927, n21928, n21929, n21930, n21932, n21933, n21934, n21935,
    n21936, n21938, n21939, n21940, n21941, n21942, n21944, n21945, n21946,
    n21947, n21948, n21950, n21951, n21952, n21953, n21954, n21956, n21957,
    n21958, n21959, n21960, n21962, n21963, n21964, n21965, n21966, n21968,
    n21969, n21970, n21971, n21972, n21974, n21975, n21976, n21977, n21978,
    n21980, n21981, n21982, n21983, n21984, n21986, n21987, n21988, n21989,
    n21990, n21992, n21993, n21994, n21995, n21996, n21998, n21999, n22000,
    n22001, n22002, n22004, n22005, n22006, n22007, n22008, n22010, n22011,
    n22012, n22013, n22014, n22016, n22017, n22019, n22020, n22022, n22023,
    n22025, n22026, n22028, n22029, n22031, n22032, n22034, n22035, n22036,
    n22037, n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
    n22047, n22048, n22050, n22051, n22052, n22053, n22054, n22056, n22057,
    n22059, n22060, n22062, n22063, n22065, n22066, n22068, n22069, n22071,
    n22072, n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
    n22083, n22084, n22085, n22087, n22088, n22089, n22090, n22091, n22092,
    n22093, n22095, n22096, n22097, n22098, n22099, n22101, n22102, n22103,
    n22104, n22105, n22106, n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22118, n22119, n22120, n22121, n22122,
    n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132,
    n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
    n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
    n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159,
    n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168,
    n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
    n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
    n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
    n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204,
    n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
    n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
    n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231,
    n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240,
    n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
    n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
    n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
    n22268, n22270, n22271, n22272, n22273, n22274, n22276, n22277, n22278,
    n22279, n22280, n22281, n22282, n22283, n22284, n22286, n22287, n22288,
    n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22301, n22302, n22303, n22304, n22305, n22306, n22307, n22308,
    n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22318, n22319,
    n22320, n22321, n22322, n22323, n22325, n22326, n22327, n22328, n22329,
    n22330, n22331, n22333, n22334, n22335, n22336, n22338, n22339, n22341,
    n22342, n22343, n22345, n22346, n22347, n22348, n22349, n22350, n22351,
    n22353, n22354, n22355, n22356, n22357, n22359, n22360, n22361, n22363,
    n22364, n22365, n22366, n22367, n22369, n22370, n22372, n22373, n22374,
    n22376, n22377, n22378, n22380, n22381, n22383, n22384, n22385, n22387,
    n22388, n22389, n22391, n22392, n22393, n22395, n22396, n22397, n22399,
    n22400, n22402, n22403, n22405, n22406, n22408, n22409, n22411, n22412,
    n22413, n22414, n22416, n22417, n22419, n22420, n22421, n22423, n22424,
    n22425, n22427, n22428, n22429, n22431, n22432, n22433, n22435, n22436,
    n22438, n22439, n22440, n22442, n22443, n22444, n22445, n22447, n22448,
    n22450, n22451, n22453, n22454, n22456, n22457, n22459, n22460, n22461,
    n22462, n22463, n22464, n22465, n22466, n22467, n22469, n22470, n22471,
    n22472, n22473, n22474, n22475, n22476, n22477, n22479, n22480, n22482,
    n22483, n22485, n22486, n22488, n22489, n22491, n22492, n22494, n22495,
    n22497, n22498, n22500, n22501, n22503, n22504, n22506, n22507, n22509,
    n22510, n22512, n22513, n22515, n22516, n22518, n22519, n22521, n22522,
    n22524, n22525, n22527, n22528, n22530, n22531, n22533, n22534, n22536,
    n22537, n22539, n22540, n22541, n22542, n22543, n22544, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22554, n22555, n22556, n22557,
    n22558, n22559, n22561, n22562, n22563, n22564, n22565, n22566, n22568,
    n22569, n22570, n22571, n22572, n22573, n22574, n22575, n22577, n22578,
    n22580, n22581, n22582, n22584, n22585, n22587, n22588, n22589, n22591,
    n22592, n22593, n22595, n22596, n22597, n22598, n22599, n22600, n22602,
    n22603, n22604, n22606, n22607, n22608, n22610, n22611, n22612, n22613,
    n22614, n22615, n22617, n22618, n22620, n22621, n22622, n22623, n22624,
    n22625, n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22642, n22643,
    n22644, n22645, n22646, n22648, n22649, n22650, n22652, n22653, n22655,
    n22656, n22658, n22659, n22661, n22662, n22664, n22665, n22666, n22668,
    n22669, n22671, n22672, n22674, n22675, n22677, n22678, n22680, n22681,
    n22683, n22684, n22686, n22687, n22689, n22690, n22692, n22693, n22695,
    n22696, n22698, n22699, n22701, n22702, n22704, n22705, n22707, n22708,
    n22710, n22711, n22713, n22714, n22716, n22717, n22719, n22720, n22722,
    n22723, n22725, n22726, n22728, n22729, n22731, n22732, n22734, n22735,
    n22737, n22738, n22740, n22741, n22743, n22744, n22746, n22747, n22748,
    n22749, n22750, n22752, n22753, n22755, n22756, n22758, n22759, n22761,
    n22762, n22764, n22765, n22767, n22768, n22770, n22771, n22773, n22774,
    n22776, n22777, n22778, n22779, n22780, n22782, n22783, n22785, n22786,
    n22788, n22789, n22791, n22792, n22794, n22795, n22798, n22799, n22800,
    n22801, n22802, n22804, n22805, n22806, n22808, n22809, n22810, n22812,
    n22813, n22814, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
    n22823, n22825, n22826, n22828, n22829, n22831, n22832, n22834, n22835,
    n22837, n22838, n22840, n22841, n22843, n22844, n22846, n22847, n22849,
    n22850, n22852, n22853, n22855, n22856, n22857, n22858, n22860, n22861,
    n22862, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
    n22872, n22873, n22874, n22875, n22877, n22878, n22879, n22880, n22881,
    n22882, n22883, n22885, n22886, n22887, n22888, n22889, n22890, n22892,
    n22893, n22894, n22895, n22896, n22897, n22899, n22900, n22901, n22902,
    n22903, n22904, n22906, n22907, n22908, n22909, n22910, n22911, n22912,
    n22913, n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22923,
    n22924, n22925, n22926, n22927, n22928, n22930, n22931, n22932, n22933,
    n22934, n22935, n22937, n22938, n22939, n22940, n22941, n22942, n22944,
    n22945, n22946, n22947, n22948, n22949, n22951, n22952, n22953, n22954,
    n22955, n22956, n22958, n22959, n22960, n22961, n22962, n22963, n22965,
    n22966, n22967, n22968, n22969, n22970, n22972, n22973, n22974, n22975,
    n22976, n22977, n22979, n22980, n22981, n22982, n22983, n22984, n22986,
    n22987, n22989, n22990, n22992, n22993, n22995, n22996, n22998, n22999,
    n23001, n23002, n23004, n23005, n23007, n23008, n23010, n23011, n23013,
    n23014, n23016, n23017, n23019, n23020, n23021, n23022, n23023, n23025,
    n23026, n23027, n23028, n23029, n23031, n23032, n23033, n23035, n23036,
    n23037, n23038, n23039, n23041, n23042, n23043, n23044, n23045, n23047,
    n23048, n23049, n23050, n23051, n23053, n23054, n23055, n23056, n23057,
    n23059, n23060, n23061, n23062, n23063, n23065, n23066, n23067, n23068,
    n23069, n23071, n23072, n23073, n23074, n23075, n23077, n23078, n23079,
    n23080, n23081, n23083, n23084, n23085, n23086, n23087, n23089, n23090,
    n23091, n23092, n23093, n23095, n23096, n23097, n23098, n23099, n23101,
    n23102, n23103, n23104, n23105, n23107, n23108, n23109, n23110, n23111,
    n23113, n23114, n23115, n23116, n23117, n23119, n23120, n23121, n23122,
    n23123, n23125, n23126, n23127, n23128, n23129, n23131, n23132, n23133,
    n23134, n23135, n23137, n23138, n23139, n23140, n23141, n23143, n23145,
    n23146, n23148, n23149, n23150, n23151, n23152, n23154, n23155, n23156,
    n23157, n23158, n23160, n23161, n23162, n23163, n23164, n23166, n23167,
    n23168, n23169, n23170, n23172, n23173, n23174, n23175, n23176, n23178,
    n23179, n23180, n23181, n23182, n23184, n23185, n23186, n23187, n23188,
    n23190, n23191, n23192, n23193, n23194, n23196, n23197, n23198, n23199,
    n23200, n23202, n23203, n23204, n23205, n23206, n23208, n23209, n23210,
    n23211, n23212, n23214, n23215, n23216, n23217, n23218, n23220, n23221,
    n23222, n23223, n23224, n23226, n23227, n23228, n23229, n23230, n23232,
    n23233, n23234, n23235, n23236, n23238, n23239, n23240, n23241, n23242,
    n23244, n23245, n23246, n23247, n23248, n23250, n23251, n23252, n23253,
    n23254, n23256, n23257, n23258, n23259, n23260, n23262, n23263, n23264,
    n23265, n23266, n23268, n23269, n23270, n23271, n23272, n23274, n23275,
    n23276, n23277, n23278, n23280, n23281, n23282, n23283, n23284, n23286,
    n23287, n23288, n23289, n23290, n23292, n23293, n23294, n23295, n23296,
    n23298, n23299, n23300, n23301, n23302, n23304, n23305, n23306, n23307,
    n23308, n23309, n23311, n23312, n23313, n23314, n23315, n23316, n23318,
    n23319, n23320, n23321, n23322, n23323, n23325, n23326, n23327, n23328,
    n23329, n23330, n23332, n23333, n23334, n23335, n23336, n23337, n23339,
    n23340, n23341, n23342, n23343, n23344, n23346, n23347, n23348, n23349,
    n23350, n23351, n23353, n23354, n23355, n23356, n23357, n23358, n23360,
    n23361, n23362, n23363, n23364, n23366, n23367, n23368, n23369, n23370,
    n23371, n23373, n23374, n23375, n23376, n23377, n23379, n23380, n23381,
    n23382, n23383, n23384, n23386, n23387, n23388, n23389, n23390, n23391,
    n23393, n23394, n23395, n23396, n23397, n23398, n23400, n23401, n23402,
    n23403, n23404, n23406, n23407, n23408, n23409, n23410, n23411, n23413,
    n23414, n23415, n23416, n23417, n23418, n23420, n23421, n23422, n23423,
    n23424, n23427, n23428, n23429, n23430, n23431, n23432, n23434, n23435,
    n23436, n23437, n23438, n23440, n23441, n23442, n23443, n23444, n23446,
    n23447, n23448, n23449, n23450, n23451, n23453, n23454, n23455, n23456,
    n23457, n23459, n23460, n23461, n23462, n23463, n23464, n23466, n23467,
    n23468, n23469, n23470, n23472, n23473, n23474, n23475, n23476, n23477,
    n23479, n23480, n23481, n23482, n23483, n23484, n23486, n23487, n23488,
    n23489, n23490, n23492, n23493, n23494, n23495, n23496, n23498, n23499,
    n23500, n23501, n23502, n23504, n23505, n23506, n23507, n23508, n23510,
    n23511, n23512, n23513, n23514, n23515, n23517, n23518, n23519, n23520,
    n23521, n23522, n23524, n23525, n23526, n23527, n23528, n23530, n23531,
    n23532, n23533, n23534, n23536, n23537, n23538, n23539, n23540, n23541,
    n23543, n23544, n23545, n23546, n23547, n23549, n23550, n23551, n23552,
    n23553, n23554, n23556, n23557, n23558, n23559, n23560, n23561, n23563,
    n23564, n23565, n23566, n23567, n23569, n23570, n23571, n23572, n23573,
    n23574, n23576, n23577, n23578, n23579, n23580, n23582, n23583, n23584,
    n23585, n23586, n23588, n23589, n23590, n23591, n23592, n23594, n23595,
    n23596, n23597, n23598, n23600, n23601, n23602, n23603, n23604, n23606,
    n23607, n23608, n23609, n23610, n23612, n23613, n23614, n23615, n23616,
    n23618, n23619, n23620, n23621, n23622, n23624, n23625, n23626, n23627,
    n23628, n23629, n23631, n23632, n23633, n23634, n23635, n23637, n23638,
    n23639, n23640, n23641, n23642, n23644, n23645, n23646, n23647, n23648,
    n23649, n23651, n23652, n23653, n23654, n23655, n23657, n23658, n23659,
    n23660, n23661, n23663, n23664, n23665, n23666, n23667, n23668, n23670,
    n23671, n23672, n23673, n23674, n23676, n23677, n23678, n23679, n23680,
    n23682, n23683, n23684, n23685, n23686, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699, n23700,
    n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
    n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23722, n23723,
    n23725, n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
    n23734, n23735, n23736, n23738, n23739, n23740, n23741, n23742, n23743,
    n23744, n23745, n23747, n23748, n23749, n23750, n23751, n23753, n23754,
    n23755, n23756, n23757, n23759, n23760, n23761, n23762, n23763, n23765,
    n23766, n23767, n23768, n23769, n23771, n23772, n23773, n23774, n23775,
    n23777, n23778, n23779, n23780, n23781, n23783, n23784, n23785, n23786,
    n23787, n23789, n23790, n23792, n23793, n23795, n23796, n23798, n23799,
    n23801, n23802, n23803, n23804, n23805, n23807, n23808, n23809, n23810,
    n23811, n23813, n23814, n23815, n23816, n23817, n23819, n23820, n23821,
    n23822, n23823, n23825, n23826, n23827, n23828, n23829, n23831, n23832,
    n23833, n23834, n23835, n23837, n23838, n23839, n23840, n23841, n23843,
    n23844, n23845, n23846, n23847, n23849, n23850, n23851, n23852, n23853,
    n23855, n23856, n23857, n23858, n23859, n23861, n23862, n23863, n23864,
    n23865, n23866, n23868, n23869, n23870, n23871, n23872, n23874, n23875,
    n23876, n23877, n23878, n23880, n23881, n23882, n23883, n23884, n23886,
    n23887, n23888, n23889, n23890, n23892, n23893, n23894, n23895, n23896,
    n23898, n23899, n23900, n23901, n23902, n23904, n23905, n23906, n23907,
    n23908, n23910, n23911, n23912, n23913, n23914, n23916, n23917, n23918,
    n23919, n23920, n23922, n23923, n23924, n23925, n23926, n23928, n23929,
    n23930, n23931, n23932, n23934, n23935, n23936, n23937, n23938, n23940,
    n23941, n23942, n23943, n23944, n23946, n23947, n23948, n23949, n23950,
    n23952, n23953, n23954, n23955, n23956, n23957, n23959, n23960, n23961,
    n23962, n23963, n23965, n23966, n23967, n23968, n23969, n23971, n23972,
    n23973, n23974, n23975, n23977, n23978, n23979, n23980, n23981, n23983,
    n23984, n23985, n23986, n23987, n23989, n23990, n23991, n23992, n23993,
    n23995, n23996, n23997, n23998, n23999, n24001, n24002, n24003, n24004,
    n24005, n24006, n24008, n24009, n24010, n24011, n24012, n24014, n24015,
    n24016, n24017, n24018, n24020, n24021, n24022, n24023, n24024, n24026,
    n24027, n24028, n24029, n24030, n24032, n24033, n24034, n24035, n24036,
    n24038, n24039, n24040, n24041, n24042, n24044, n24045, n24046, n24047,
    n24048, n24050, n24051, n24052, n24053, n24054, n24056, n24057, n24058,
    n24059, n24060, n24062, n24063, n24064, n24065, n24066, n24068, n24069,
    n24070, n24071, n24072, n24074, n24075, n24076, n24077, n24078, n24080,
    n24081, n24082, n24083, n24084, n24086, n24087, n24088, n24089, n24090,
    n24092, n24093, n24094, n24095, n24096, n24098, n24099, n24100, n24101,
    n24102, n24104, n24105, n24106, n24107, n24108, n24110, n24111, n24112,
    n24113, n24114, n24116, n24117, n24118, n24119, n24120, n24122, n24123,
    n24124, n24125, n24126, n24128, n24129, n24130, n24131, n24132, n24134,
    n24135, n24136, n24137, n24138, n24140, n24141, n24142, n24143, n24144,
    n24146, n24147, n24148, n24149, n24150, n24152, n24153, n24154, n24155,
    n24156, n24158, n24159, n24160, n24161, n24162, n24164, n24165, n24166,
    n24167, n24168, n24170, n24171, n24172, n24173, n24174, n24176, n24177,
    n24178, n24179, n24180, n24182, n24183, n24184, n24185, n24186, n24188,
    n24189, n24190, n24191, n24192, n24194, n24195, n24196, n24197, n24198,
    n24200, n24201, n24202, n24203, n24204, n24206, n24207, n24208, n24209,
    n24210, n24212, n24213, n24214, n24215, n24216, n24218, n24219, n24220,
    n24221, n24222, n24224, n24225, n24226, n24227, n24228, n24230, n24231,
    n24232, n24233, n24234, n24236, n24237, n24238, n24239, n24240, n24242,
    n24243, n24244, n24245, n24246, n24248, n24249, n24250, n24251, n24252,
    n24254, n24255, n24256, n24257, n24258, n24260, n24261, n24262, n24263,
    n24264, n24266, n24267, n24268, n24269, n24270, n24272, n24273, n24274,
    n24275, n24276, n24278, n24279, n24280, n24281, n24282, n24284, n24285,
    n24286, n24287, n24288, n24290, n24291, n24292, n24293, n24294, n24296,
    n24297, n24298, n24299, n24300, n24302, n24303, n24304, n24305, n24306,
    n24308, n24309, n24310, n24311, n24312, n24314, n24315, n24316, n24317,
    n24318, n24320, n24321, n24322, n24323, n24324, n24326, n24327, n24328,
    n24329, n24330, n24332, n24333, n24334, n24335, n24336, n24338, n24339,
    n24340, n24341, n24342, n24344, n24345, n24346, n24347, n24348, n24350,
    n24351, n24352, n24353, n24354, n24356, n24357, n24358, n24359, n24360,
    n24362, n24363, n24364, n24365, n24366, n24368, n24369, n24370, n24371,
    n24372, n24374, n24375, n24376, n24377, n24378, n24380, n24381, n24382,
    n24383, n24384, n24386, n24387, n24388, n24389, n24390, n24392, n24393,
    n24394, n24395, n24396, n24398, n24399, n24400, n24401, n24402, n24404,
    n24405, n24406, n24407, n24408, n24410, n24411, n24412, n24413, n24414,
    n24416, n24417, n24418, n24419, n24420, n24422, n24423, n24424, n24425,
    n24426, n24428, n24429, n24430, n24431, n24432, n24434, n24435, n24436,
    n24437, n24438, n24440, n24441, n24442, n24443, n24444, n24446, n24447,
    n24448, n24449, n24450, n24452, n24453, n24454, n24455, n24456, n24458,
    n24459, n24460, n24461, n24462, n24464, n24465, n24466, n24467, n24468,
    n24470, n24471, n24472, n24473, n24474, n24476, n24477, n24478, n24479,
    n24480, n24482, n24483, n24484, n24485, n24486, n24488, n24489, n24490,
    n24491, n24492, n24494, n24495, n24496, n24497, n24498, n24500, n24501,
    n24502, n24503, n24504, n24506, n24507, n24508, n24509, n24510, n24512,
    n24513, n24514, n24515, n24516, n24518, n24519, n24520, n24521, n24522,
    n24524, n24525, n24526, n24527, n24528, n24530, n24531, n24532, n24533,
    n24534, n24536, n24537, n24538, n24539, n24540, n24542, n24543, n24544,
    n24545, n24546, n24548, n24549, n24550, n24551, n24552, n24554, n24555,
    n24556, n24557, n24558, n24560, n24561, n24562, n24563, n24564, n24566,
    n24567, n24568, n24569, n24570, n24572, n24573, n24574, n24575, n24576,
    n24578, n24579, n24580, n24581, n24582, n24584, n24585, n24586, n24587,
    n24588, n24590, n24591, n24592, n24593, n24594, n24596, n24597, n24598,
    n24599, n24600, n24602, n24603, n24604, n24605, n24606, n24608, n24609,
    n24610, n24611, n24612, n24614, n24615, n24616, n24617, n24618, n24620,
    n24621, n24622, n24623, n24624, n24626, n24627, n24628, n24629, n24630,
    n24632, n24633, n24634, n24635, n24636, n24638, n24639, n24640, n24641,
    n24642, n24644, n24645, n24646, n24647, n24648, n24650, n24651, n24652,
    n24653, n24654, n24656, n24657, n24658, n24659, n24660, n24662, n24663,
    n24664, n24665, n24666, n24668, n24669, n24670, n24671, n24672, n24674,
    n24675, n24676, n24677, n24678, n24680, n24681, n24682, n24683, n24684,
    n24686, n24687, n24688, n24689, n24690, n24692, n24693, n24694, n24695,
    n24696, n24698, n24699, n24700, n24701, n24702, n24704, n24705, n24706,
    n24707, n24708, n24710, n24711, n24712, n24713, n24714, n24716, n24717,
    n24718, n24719, n24720, n24722, n24723, n24724, n24725, n24726, n24728,
    n24729, n24730, n24731, n24732, n24734, n24735, n24736, n24737, n24738,
    n24740, n24741, n24742, n24743, n24744, n24746, n24747, n24748, n24749,
    n24750, n24752, n24753, n24754, n24755, n24756, n24758, n24759, n24760,
    n24761, n24762, n24764, n24765, n24766, n24767, n24768, n24770, n24771,
    n24772, n24773, n24774, n24776, n24777, n24778, n24779, n24780, n24782,
    n24783, n24784, n24785, n24786, n24788, n24789, n24790, n24791, n24792,
    n24794, n24795, n24796, n24797, n24798, n24800, n24801, n24802, n24803,
    n24804, n24806, n24807, n24808, n24809, n24810, n24812, n24813, n24814,
    n24815, n24816, n24818, n24819, n24820, n24821, n24822, n24824, n24825,
    n24826, n24827, n24828, n24830, n24831, n24832, n24833, n24834, n24836,
    n24837, n24838, n24839, n24840, n24842, n24843, n24844, n24845, n24846,
    n24848, n24849, n24850, n24851, n24852, n24854, n24855, n24856, n24857,
    n24858, n24860, n24861, n24862, n24863, n24864, n24866, n24867, n24868,
    n24869, n24870, n24872, n24873, n24874, n24875, n24876, n24878, n24879,
    n24880, n24881, n24882, n24884, n24885, n24886, n24887, n24888, n24890,
    n24891, n24892, n24893, n24894, n24896, n24897, n24898, n24899, n24900,
    n24902, n24903, n24904, n24905, n24906, n24908, n24909, n24910, n24911,
    n24912, n24914, n24915, n24916, n24917, n24918, n24920, n24921, n24922,
    n24923, n24924, n24926, n24927, n24928, n24929, n24930, n24932, n24933,
    n24934, n24935, n24936, n24938, n24939, n24940, n24941, n24942, n24944,
    n24945, n24946, n24947, n24948, n24950, n24951, n24952, n24953, n24954,
    n24956, n24957, n24958, n24959, n24960, n24962, n24963, n24964, n24965,
    n24966, n24968, n24969, n24970, n24971, n24972, n24974, n24975, n24976,
    n24977, n24978, n24980, n24981, n24982, n24983, n24984, n24986, n24987,
    n24988, n24989, n24990, n24992, n24993, n24994, n24995, n24996, n24998,
    n24999, n25000, n25001, n25002, n25004, n25005, n25006, n25007, n25008,
    n25010, n25011, n25012, n25013, n25014, n25016, n25017, n25018, n25019,
    n25020, n25022, n25023, n25024, n25025, n25026, n25028, n25029, n25030,
    n25031, n25032, n25034, n25035, n25036, n25037, n25038, n25040, n25041,
    n25042, n25043, n25044, n25046, n25047, n25048, n25049, n25050, n25052,
    n25053, n25054, n25055, n25056, n25058, n25059, n25060, n25061, n25062,
    n25064, n25065, n25066, n25067, n25068, n25070, n25071, n25072, n25073,
    n25074, n25076, n25077, n25078, n25079, n25080, n25082, n25083, n25084,
    n25085, n25086, n25088, n25089, n25090, n25091, n25092, n25094, n25095,
    n25096, n25097, n25098, n25100, n25101, n25102, n25103, n25104, n25106,
    n25107, n25108, n25109, n25110, n25112, n25113, n25114, n25115, n25116,
    n25118, n25119, n25120, n25121, n25122, n25124, n25125, n25126, n25127,
    n25128, n25130, n25131, n25132, n25133, n25134, n25136, n25137, n25138,
    n25139, n25140, n25142, n25143, n25144, n25145, n25146, n25148, n25149,
    n25150, n25151, n25152, n25154, n25155, n25156, n25157, n25158, n25160,
    n25161, n25162, n25163, n25164, n25166, n25167, n25168, n25169, n25170,
    n25172, n25173, n25174, n25175, n25176, n25178, n25179, n25180, n25181,
    n25182, n25184, n25185, n25186, n25187, n25188, n25190, n25191, n25192,
    n25193, n25194, n25196, n25197, n25198, n25199, n25200, n25202, n25203,
    n25204, n25205, n25206, n25208, n25209, n25210, n25211, n25212, n25214,
    n25215, n25216, n25217, n25218, n25220, n25221, n25222, n25223, n25224,
    n25226, n25227, n25228, n25229, n25230, n25232, n25233, n25234, n25235,
    n25236, n25238, n25239, n25240, n25241, n25242, n25244, n25245, n25246,
    n25247, n25248, n25250, n25251, n25252, n25253, n25254, n25256, n25257,
    n25258, n25259, n25260, n25262, n25263, n25264, n25265, n25266, n25268,
    n25269, n25270, n25271, n25272, n25274, n25275, n25276, n25277, n25278,
    n25280, n25281, n25282, n25283, n25284, n25286, n25287, n25288, n25289,
    n25290, n25292, n25293, n25294, n25295, n25296, n25298, n25299, n25300,
    n25301, n25302, n25304, n25305, n25306, n25307, n25308, n25310, n25311,
    n25312, n25313, n25314, n25316, n25317, n25318, n25319, n25320, n25322,
    n25323, n25324, n25325, n25326, n25328, n25329, n25330, n25331, n25332,
    n25334, n25335, n25336, n25337, n25338, n25340, n25341, n25342, n25343,
    n25344, n25346, n25347, n25348, n25349, n25350, n25352, n25353, n25354,
    n25355, n25356, n25358, n25359, n25360, n25361, n25362, n25364, n25365,
    n25366, n25367, n25368, n25370, n25371, n25372, n25373, n25374, n25376,
    n25377, n25378, n25379, n25380, n25382, n25383, n25384, n25385, n25386,
    n25388, n25389, n25390, n25391, n25392, n25394, n25395, n25396, n25397,
    n25398, n25399, n25400, n25401, n25403, n25404, n25405, n25406, n25407,
    n25409, n25410, n25411, n25412, n25413, n25415, n25416, n25417, n25418,
    n25419, n25421, n25422, n25423, n25424, n25425, n25427, n25428, n25429,
    n25430, n25431, n25433, n25434, n25435, n25436, n25437, n25439, n25440,
    n25441, n25442, n25443, n25445, n25446, n25447, n25448, n25449, n25451,
    n25452, n25453, n25454, n25455, n25457, n25458, n25459, n25460, n25461,
    n25463, n25464, n25465, n25466, n25467, n25469, n25470, n25471, n25472,
    n25473, n25475, n25476, n25477, n25478, n25479, n25481, n25482, n25483,
    n25484, n25485, n25487, n25488, n25489, n25490, n25491, n25493, n25494,
    n25495, n25496, n25497, n25499, n25500, n25501, n25502, n25503, n25505,
    n25506, n25507, n25508, n25509, n25511, n25512, n25513, n25514, n25515,
    n25517, n25518, n25519, n25520, n25521, n25523, n25524, n25525, n25526,
    n25527, n25529, n25530, n25531, n25532, n25533, n25535, n25536, n25537,
    n25538, n25539, n25541, n25542, n25543, n25544, n25545, n25547, n25548,
    n25549, n25550, n25551, n25553, n25554, n25555, n25556, n25557, n25559,
    n25560, n25561, n25562, n25563, n25565, n25566, n25567, n25568, n25569,
    n25571, n25572, n25573, n25574, n25575, n25577, n25578, n25579, n25580,
    n25581, n25583, n25584, n25585, n25586, n25587, n25589, n25590, n25591,
    n25592, n25593, n25595, n25596, n25598, n25599, n25600, n25601, n25602,
    n25604, n25605, n25606, n25607, n25608, n25610, n25611, n25612, n25613,
    n25614, n25616, n25617, n25618, n25619, n25620, n25622, n25623, n25624,
    n25625, n25626, n25628, n25629, n25630, n25631, n25632, n25634, n25635,
    n25636, n25637, n25638, n25640, n25641, n25642, n25643, n25644, n25646,
    n25647, n25648, n25649, n25650, n25652, n25653, n25654, n25655, n25656,
    n25658, n25659, n25660, n25661, n25662, n25664, n25665, n25666, n25667,
    n25668, n25670, n25671, n25672, n25673, n25674, n25676, n25677, n25678,
    n25679, n25680, n25682, n25683, n25684, n25685, n25686, n25688, n25689,
    n25690, n25691, n25692, n25694, n25695, n25696, n25697, n25698, n25700,
    n25701, n25702, n25703, n25704, n25706, n25707, n25708, n25709, n25710,
    n25712, n25713, n25714, n25715, n25716, n25718, n25719, n25720, n25721,
    n25722, n25724, n25725, n25726, n25727, n25728, n25730, n25731, n25732,
    n25733, n25734, n25736, n25737, n25738, n25739, n25740, n25742, n25743,
    n25744, n25745, n25746, n25748, n25749, n25750, n25751, n25752, n25754,
    n25755, n25756, n25757, n25758, n25760, n25761, n25762, n25763, n25764,
    n25766, n25767, n25768, n25769, n25770, n25772, n25773, n25774, n25775,
    n25776, n25778, n25779, n25780, n25781, n25782, n25784, n25785, n25786,
    n25787, n25788, n25790, n25791, n25792, n25793, n25794, n25796, n25797,
    n25798, n25799, n25800, n25802, n25803, n25804, n25805, n25806, n25808,
    n25809, n25810, n25811, n25812, n25814, n25815, n25816, n25817, n25818,
    n25820, n25821, n25822, n25823, n25824, n25826, n25827, n25828, n25829,
    n25830, n25832, n25833, n25834, n25835, n25836, n25838, n25839, n25840,
    n25841, n25842, n25844, n25845, n25846, n25847, n25848, n25850, n25851,
    n25852, n25853, n25854, n25856, n25857, n25858, n25859, n25860, n25862,
    n25863, n25864, n25865, n25866, n25868, n25869, n25870, n25871, n25872,
    n25874, n25875, n25876, n25877, n25878, n25880, n25881, n25882, n25883,
    n25884, n25886, n25887, n25888, n25889, n25890, n25892, n25893, n25894,
    n25895, n25896, n25898, n25899, n25900, n25901, n25902, n25904, n25905,
    n25906, n25907, n25908, n25910, n25911, n25912, n25913, n25914, n25916,
    n25917, n25918, n25919, n25920, n25922, n25923, n25924, n25925, n25926,
    n25928, n25929, n25930, n25931, n25932, n25934, n25935, n25936, n25937,
    n25938, n25940, n25941, n25942, n25943, n25944, n25946, n25947, n25948,
    n25949, n25950, n25952, n25953, n25954, n25955, n25956, n25958, n25959,
    n25960, n25961, n25962, n25964, n25965, n25966, n25967, n25968, n25970,
    n25971, n25972, n25973, n25974, n25976, n25977, n25978, n25979, n25980,
    n25982, n25983, n25984, n25985, n25986, n25988, n25989, n25990, n25991,
    n25992, n25994, n25995, n25996, n25997, n25998, n26000, n26001, n26002,
    n26003, n26004, n26006, n26007, n26008, n26009, n26010, n26012, n26013,
    n26014, n26015, n26016, n26018, n26019, n26020, n26021, n26022, n26024,
    n26025, n26026, n26027, n26028, n26030, n26031, n26032, n26033, n26034,
    n26036, n26037, n26038, n26039, n26040, n26042, n26043, n26044, n26045,
    n26046, n26048, n26049, n26050, n26051, n26052, n26054, n26055, n26056,
    n26057, n26058, n26060, n26061, n26062, n26063, n26064, n26066, n26067,
    n26068, n26069, n26070, n26072, n26073, n26074, n26075, n26076, n26078,
    n26079, n26080, n26081, n26082, n26084, n26085, n26086, n26087, n26088,
    n26090, n26091, n26092, n26093, n26094, n26096, n26097, n26098, n26099,
    n26100, n26102, n26103, n26104, n26105, n26106, n26108, n26109, n26110,
    n26111, n26112, n26114, n26115, n26116, n26117, n26118, n26120, n26121,
    n26122, n26123, n26124, n26126, n26127, n26128, n26129, n26130, n26132,
    n26133, n26134, n26135, n26136, n26138, n26139, n26140, n26141, n26142,
    n26144, n26145, n26146, n26147, n26148, n26150, n26151, n26152, n26153,
    n26154, n26156, n26157, n26158, n26159, n26160, n26162, n26163, n26164,
    n26165, n26166, n26168, n26169, n26170, n26171, n26172, n26174, n26175,
    n26176, n26177, n26178, n26180, n26181, n26182, n26183, n26184, n26186,
    n26187, n26188, n26190, n26191, n26192, n26193, n26194, n26196, n26197,
    n26198, n26199, n26200, n26202, n26203, n26204, n26205, n26206, n26208,
    n26209, n26210, n26211, n26212, n26214, n26215, n26216, n26217, n26218,
    n26220, n26221, n26222, n26223, n26224, n26226, n26227, n26228, n26229,
    n26230, n26232, n26233, n26234, n26235, n26236, n26238, n26239, n26240,
    n26241, n26242, n26244, n26245, n26246, n26247, n26248, n26250, n26251,
    n26252, n26253, n26254, n26256, n26257, n26258, n26259, n26260, n26262,
    n26263, n26264, n26265, n26266, n26268, n26269, n26270, n26271, n26272,
    n26274, n26275, n26276, n26277, n26278, n26280, n26281, n26282, n26283,
    n26284, n26286, n26287, n26288, n26289, n26290, n26292, n26293, n26294,
    n26295, n26296, n26298, n26299, n26300, n26301, n26302, n26304, n26305,
    n26306, n26307, n26308, n26310, n26311, n26312, n26313, n26314, n26316,
    n26317, n26318, n26319, n26320, n26322, n26323, n26324, n26325, n26326,
    n26328, n26329, n26330, n26331, n26332, n26334, n26335, n26336, n26337,
    n26338, n26340, n26341, n26342, n26343, n26344, n26346, n26347, n26348,
    n26349, n26350, n26352, n26353, n26354, n26355, n26356, n26358, n26359,
    n26360, n26361, n26362, n26364, n26365, n26366, n26367, n26368, n26370,
    n26371, n26372, n26373, n26374, n26376, n26377, n26378, n26379, n26380,
    n26382, n26383, n26384, n26385, n26386, n26388, n26389, n26390, n26391,
    n26392, n26394, n26395, n26396, n26397, n26398, n26400, n26401, n26402,
    n26403, n26404, n26406, n26407, n26408, n26409, n26410, n26412, n26413,
    n26414, n26415, n26416, n26418, n26419, n26420, n26421, n26422, n26424,
    n26425, n26426, n26427, n26428, n26430, n26431, n26432, n26433, n26434,
    n26436, n26437, n26438, n26439, n26440, n26442, n26443, n26444, n26445,
    n26446, n26448, n26449, n26450, n26451, n26452, n26454, n26455, n26456,
    n26457, n26458, n26460, n26461, n26462, n26463, n26464, n26466, n26467,
    n26468, n26469, n26470, n26472, n26473, n26474, n26475, n26476, n26478,
    n26479, n26480, n26481, n26482, n26484, n26485, n26486, n26487, n26488,
    n26490, n26491, n26492, n26493, n26494, n26496, n26497, n26498, n26499,
    n26500, n26502, n26503, n26504, n26505, n26506, n26508, n26509, n26510,
    n26511, n26512, n26514, n26515, n26516, n26517, n26518, n26520, n26521,
    n26522, n26523, n26524, n26526, n26527, n26528, n26529, n26530, n26532,
    n26533, n26534, n26535, n26536, n26538, n26539, n26540, n26541, n26542,
    n26544, n26545, n26546, n26547, n26548, n26550, n26551, n26552, n26553,
    n26554, n26556, n26557, n26558, n26559, n26560, n26562, n26563, n26564,
    n26565, n26566, n26568, n26569, n26570, n26571, n26572, n26574, n26575,
    n26576, n26577, n26578, n26580, n26581, n26582, n26583, n26584, n26586,
    n26587, n26588, n26589, n26590, n26592, n26593, n26594, n26595, n26596,
    n26598, n26599, n26600, n26601, n26602, n26604, n26605, n26606, n26607,
    n26608, n26610, n26611, n26612, n26613, n26614, n26616, n26617, n26618,
    n26619, n26620, n26622, n26623, n26624, n26625, n26626, n26628, n26629,
    n26630, n26631, n26632, n26634, n26635, n26636, n26637, n26638, n26639,
    n26640, n26641, n26642, n26643, n26644, n26646, n26647, n26648, n26649,
    n26650, n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26660,
    n26661, n26662, n26663, n26664, n26666, n26667, n26668, n26669, n26670,
    n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678, n26679,
    n26680, n26681, n26683, n26684, n26685, n26686, n26687, n26689, n26690,
    n26691, n26692, n26693, n26695, n26696, n26697, n26698, n26699, n26701,
    n26702, n26703, n26704, n26705, n26707, n26708, n26709, n26710, n26711,
    n26713, n26714, n26715, n26716, n26717, n26719, n26720, n26721, n26722,
    n26723, n26725, n26726, n26727, n26728, n26729, n26731, n26732, n26733,
    n26734, n26735, n26737, n26738, n26739, n26740, n26741, n26743, n26744,
    n26745, n26746, n26747, n26749, n26750, n26751, n26752, n26753, n26755,
    n26756, n26757, n26758, n26759, n26761, n26762, n26764, n26765, n26767,
    n26768, n26769, n26770, n26771, n26773, n26774, n26776, n26777, n26779,
    n26780, n26781, n26782, n26783, n26785, n26786, n26788, n26789, n26790,
    n26791, n26793, n26794, n26795, n26796, n26797, n26799, n26800, n26802,
    n26803, n26805, n26806, n26807, n26808, n26809, n26811, n26812, n26813,
    n26814, n26815, n26817, n26818, n26819, n26820, n26821, n26823, n26824,
    n26825, n26826, n26827, n26829, n26830, n26831, n26832, n26833, n26835,
    n26836, n26837, n26838, n26839, n26841, n26842, n26844, n26845, n26846,
    n26847, n26848, n26850, n26851, n26852, n26853, n26854, n26856, n26857,
    n26859, n26860, n26861, n26862, n26863, n26865, n26866, n26868, n26869,
    n26871, n26872, n26874, n26875, n26876, n26877, n26878, n26880, n26881,
    n26883, n26884, n26886, n26887, n26888, n26889, n26890, n26892, n26893,
    n26895, n26896, n26897, n26898, n26899, n26901, n26902, n26903, n26904,
    n26905, n26907, n26908, n26909, n26910, n26911, n26913, n26914, n26915,
    n26916, n26917, n26919, n26920, n26921, n26922, n26923, n26925, n26926,
    n26927, n26928, n26929, n26931, n26932, n26933, n26934, n26935, n26937,
    n26938, n26939, n26940, n26941, n26943, n26944, n26945, n26946, n26947,
    n26949, n26950, n26952, n26953, n26954, n26955, n26957, n26958, n26960,
    n26962, n26963, n26965, n26966, n26968, n26969, n26971, n26972, n26973,
    n26974, n26975, n26976, n26978, n26979, n26980, n26981, n26982, n26983,
    n26984, n26985, n26987, n26988, n26990, n26991, n26993, n26994, n26996,
    n26997, n26999, n27000, n27002, n27003, n27005, n27006, n27008, n27009,
    n27011, n27012, n27014, n27015, n27017, n27018, n27020, n27021, n27023,
    n27024, n27026, n27027, n27029, n27030, n27032, n27033, n27035, n27036,
    n27038, n27039, n27041, n27042, n27044, n27045, n27047, n27048, n27050,
    n27051, n27053, n27054, n27056, n27057, n27059, n27060, n27062, n27063,
    n27065, n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
    n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
    n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
    n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099, n27100,
    n27101, n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
    n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117, n27118,
    n27119, n27120, n27121, n27122, n27123, n27124, n27125, n27126, n27127,
    n27128, n27129, n27130, n27131, n27132, n27133, n27134, n27135, n27136,
    n27137, n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
    n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
    n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
    n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171, n27172,
    n27173, n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
    n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189, n27190,
    n27191, n27192, n27193, n27194, n27195, n27196, n27197, n27198, n27199,
    n27200, n27201, n27202, n27203, n27204, n27205, n27206, n27207, n27208,
    n27209, n27211, n27212, n27214, n27215, n27217, n27218, n27220, n27221,
    n27223, n27224, n27226, n27227, n27229, n27230, n27232, n27233, n27235,
    n27236, n27238, n27239, n27241, n27242, n27244, n27245, n27247, n27248,
    n27250, n27251, n27253, n27254, n27256, n27257, n27259, n27260, n27262,
    n27263, n27265, n27266, n27268, n27269, n27271, n27272, n27274, n27275,
    n27277, n27278, n27280, n27281, n27283, n27284, n27286, n27287, n27289,
    n27290, n27292, n27293, n27295, n27296, n27298, n27299, n27301, n27302,
    n27304, n27305, n27307, n27308, n27310, n27311, n27313, n27314, n27316,
    n27317, n27319, n27320, n27322, n27323, n27325, n27326, n27328, n27329,
    n27330, n27331, n27332, n27333, n27335, n27337, n27338, n27339, n27340,
    n27341, n27343, n27344, n27345, n27346, n27347, n27349, n27350, n27351,
    n27352, n27353, n27355, n27356, n27357, n27358, n27359, n27361, n27362,
    n27363, n27364, n27365, n27367, n27368, n27369, n27370, n27371, n27373,
    n27374, n27375, n27376, n27377, n27379, n27380, n27381, n27382, n27383,
    n27385, n27386, n27387, n27388, n27389, n27391, n27392, n27393, n27394,
    n27395, n27397, n27398, n27399, n27400, n27401, n27403, n27404, n27405,
    n27406, n27407, n27409, n27410, n27411, n27412, n27413, n27415, n27416,
    n27417, n27418, n27419, n27421, n27422, n27423, n27424, n27425, n27427,
    n27428, n27429, n27430, n27431, n27433, n27434, n27435, n27436, n27437,
    n27439, n27440, n27441, n27442, n27443, n27445, n27446, n27447, n27448,
    n27449, n27451, n27452, n27453, n27454, n27455, n27457, n27458, n27459,
    n27460, n27461, n27463, n27464, n27465, n27466, n27467, n27469, n27470,
    n27471, n27472, n27473, n27475, n27476, n27477, n27478, n27479, n27481,
    n27482, n27483, n27484, n27485, n27487, n27488, n27489, n27490, n27491,
    n27493, n27494, n27495, n27496, n27497, n27499, n27500, n27501, n27502,
    n27503, n27505, n27506, n27507, n27508, n27509, n27511, n27512, n27513,
    n27514, n27515, n27517, n27518, n27519, n27520, n27521, n27523, n27524,
    n27525, n27526, n27527, n27529, n27530, n27531, n27532, n27533, n27535,
    n27536, n27537, n27538, n27539, n27541, n27542, n27543, n27544, n27545,
    n27547, n27548, n27549, n27550, n27551, n27553, n27554, n27555, n27556,
    n27557, n27559, n27560, n27561, n27562, n27563, n27565, n27566, n27567,
    n27568, n27569, n27571, n27572, n27573, n27574, n27575, n27577, n27578,
    n27579, n27580, n27581, n27583, n27584, n27585, n27586, n27587, n27589,
    n27590, n27591, n27592, n27593, n27595, n27596, n27597, n27598, n27599,
    n27601, n27602, n27603, n27604, n27605, n27607, n27608, n27609, n27610,
    n27611, n27613, n27614, n27615, n27616, n27617, n27619, n27620, n27621,
    n27622, n27623, n27625, n27626, n27627, n27628, n27629, n27631, n27632,
    n27633, n27634, n27635, n27637, n27638, n27639, n27640, n27641, n27643,
    n27644, n27645, n27646, n27647, n27649, n27650, n27651, n27652, n27653,
    n27655, n27656, n27657, n27658, n27659, n27661, n27662, n27663, n27664,
    n27665, n27667, n27668, n27669, n27670, n27671, n27673, n27674, n27675,
    n27676, n27677, n27679, n27680, n27681, n27682, n27683, n27685, n27686,
    n27687, n27688, n27689, n27691, n27692, n27693, n27694, n27695, n27697,
    n27698, n27699, n27700, n27701, n27703, n27704, n27705, n27706, n27707,
    n27709, n27710, n27711, n27712, n27713, n27715, n27716, n27717, n27718,
    n27719, n27721, n27722, n27723, n27724, n27725, n27727, n27728, n27729,
    n27730, n27731, n27733, n27734, n27735, n27736, n27737, n27739, n27740,
    n27741, n27742, n27743, n27745, n27746, n27747, n27748, n27749, n27751,
    n27752, n27753, n27754, n27755, n27757, n27758, n27759, n27760, n27761,
    n27763, n27764, n27765, n27766, n27767, n27769, n27770, n27771, n27772,
    n27773, n27775, n27776, n27777, n27778, n27779, n27781, n27782, n27783,
    n27784, n27785, n27787, n27788, n27789, n27790, n27791, n27793, n27794,
    n27795, n27796, n27797, n27799, n27800, n27801, n27802, n27803, n27805,
    n27806, n27807, n27808, n27809, n27811, n27812, n27813, n27814, n27815,
    n27817, n27818, n27819, n27820, n27821, n27823, n27824, n27825, n27826,
    n27827, n27829, n27830, n27831, n27832, n27833, n27835, n27836, n27837,
    n27838, n27839, n27841, n27842, n27843, n27844, n27845, n27847, n27848,
    n27849, n27850, n27851, n27853, n27854, n27855, n27856, n27857, n27859,
    n27860, n27861, n27862, n27863, n27865, n27866, n27867, n27868, n27869,
    n27871, n27872, n27873, n27874, n27875, n27877, n27878, n27879, n27880,
    n27881, n27883, n27884, n27885, n27886, n27887, n27889, n27890, n27891,
    n27892, n27893, n27895, n27896, n27897, n27898, n27899, n27901, n27902,
    n27903, n27904, n27905, n27907, n27908, n27909, n27910, n27911, n27913,
    n27914, n27915, n27916, n27917, n27919, n27920, n27921, n27922, n27923,
    n27925, n27926, n27927, n27928, n27929, n27931, n27932, n27933, n27934,
    n27935, n27937, n27938, n27939, n27940, n27941, n27943, n27944, n27945,
    n27946, n27947, n27949, n27950, n27951, n27952, n27953, n27955, n27956,
    n27957, n27958, n27959, n27961, n27962, n27963, n27964, n27965, n27967,
    n27968, n27969, n27970, n27971, n27973, n27974, n27975, n27976, n27977,
    n27979, n27980, n27981, n27982, n27983, n27985, n27986, n27987, n27988,
    n27989, n27991, n27992, n27993, n27994, n27995, n27997, n27998, n28000,
    n28001, n28002, n28003, n28004, n28006, n28007, n28008, n28009, n28010,
    n28012, n28013, n28014, n28015, n28016, n28018, n28019, n28020, n28021,
    n28022, n28024, n28025, n28026, n28027, n28028, n28030, n28031, n28032,
    n28033, n28034, n28036, n28037, n28038, n28039, n28040, n28042, n28043,
    n28044, n28045, n28046, n28048, n28049, n28050, n28051, n28052, n28054,
    n28055, n28056, n28057, n28058, n28060, n28061, n28062, n28063, n28064,
    n28066, n28067, n28068, n28069, n28070, n28072, n28073, n28074, n28075,
    n28076, n28078, n28079, n28080, n28081, n28082, n28084, n28085, n28086,
    n28087, n28088, n28090, n28091, n28092, n28093, n28094, n28096, n28097,
    n28098, n28099, n28100, n28102, n28103, n28104, n28105, n28106, n28108,
    n28109, n28110, n28111, n28112, n28114, n28115, n28116, n28117, n28118,
    n28120, n28121, n28122, n28123, n28124, n28126, n28127, n28128, n28129,
    n28130, n28132, n28133, n28134, n28135, n28136, n28138, n28139, n28140,
    n28141, n28142, n28144, n28145, n28146, n28147, n28148, n28150, n28151,
    n28152, n28153, n28154, n28156, n28157, n28158, n28159, n28160, n28162,
    n28163, n28165, n28166, n28167, n28168, n28169, n28171, n28172, n28173,
    n28174, n28175, n28177, n28178, n28180, n28181, n28183, n28184, n28186,
    n28187, n28188, n28189, n28190, n28192, n28193, n28194, n28195, n28196,
    n28198, n28199, n28200, n28201, n28202, n28204, n28205, n28206, n28207,
    n28208, n28210, n28211, n28212, n28213, n28214, n28216, n28217, n28218,
    n28219, n28220, n28222, n28223, n28224, n28225, n28226, n28228, n28229,
    n28230, n28231, n28232, n28234, n28235, n28236, n28237, n28238, n28240,
    n28241, n28242, n28243, n28244, n28246, n28247, n28249, n28250, n28251,
    n28252, n28253, n28255, n28256, n28257, n28258, n28259, n28261, n28262,
    n28264, n28265, n28266, n28267, n28268, n28270, n28271, n28272, n28273,
    n28274, n28276, n28277, n28278, n28280, n28281, n28282, n28283, n28284,
    n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28293, n28294,
    n28296, n28298, n28299, n28300, n28301, n28302, n28304, n28305, n28307,
    n28308, n28310, n28311, n28313, n28314, n28315, n28316, n28317, n28319,
    n28320, n28321, n28322, n28323, n28325, n28326, n28328, n28329, n28331,
    n28332, n28334, n28335, n28336, n28337, n28338, n28340, n28341, n28342,
    n28343, n28344, n28346, n28347, n28348, n28349, n28350, n28352, n28353,
    n28354, n28355, n28356, n28358, n28359, n28360, n28361, n28362, n28364,
    n28365, n28366, n28367, n28368, n28370, n28371, n28372, n28373, n28374,
    n28376, n28377, n28378, n28379, n28380, n28382, n28383, n28384, n28385,
    n28386, n28388, n28389, n28390, n28391, n28392, n28394, n28395, n28396,
    n28397, n28398, n28400, n28401, n28403, n28404, n28405, n28406, n28407,
    n28409, n28410, n28411, n28412, n28413, n28415, n28416, n28417, n28418,
    n28419, n28421, n28422, n28423, n28424, n28425, n28427, n28428, n28429,
    n28430, n28431, n28433, n28434, n28435, n28436, n28437, n28439, n28440,
    n28441, n28442, n28443, n28445, n28446, n28448, n28449, n28450, n28451,
    n28452, n28454, n28455, n28456, n28457, n28458, n28460, n28461, n28462,
    n28463, n28464, n28466, n28467, n28468, n28469, n28470, n28472, n28473,
    n28474, n28475, n28476, n28478, n28479, n28480, n28481, n28482, n28484,
    n28485, n28486, n28487, n28488, n28490, n28491, n28493, n28494, n28495,
    n28496, n28497, n28499, n28500, n28501, n28502, n28503, n28505, n28506,
    n28507, n28508, n28509, n28511, n28512, n28513, n28514, n28515, n28517,
    n28518, n28519, n28520, n28521, n28523, n28524, n28525, n28526, n28527,
    n28529, n28530, n28531, n28532, n28533, n28535, n28536, n28537, n28538,
    n28539, n28541, n28542, n28543, n28544, n28545, n28547, n28548, n28549,
    n28550, n28551, n28553, n28554, n28555, n28556, n28557, n28559, n28560,
    n28561, n28562, n28563, n28565, n28566, n28567, n28568, n28569, n28571,
    n28572, n28573, n28574, n28575, n28577, n28578, n28579, n28580, n28581,
    n28583, n28584, n28585, n28586, n28587, n28589, n28590, n28591, n28592,
    n28593, n28595, n28596, n28597, n28598, n28599, n28601, n28602, n28603,
    n28604, n28605, n28607, n28608, n28609, n28610, n28611, n28613, n28614,
    n28615, n28616, n28617, n28619, n28620, n28621, n28622, n28623, n28625,
    n28626, n28628, n28629, n28631, n28632, n28633, n28634, n28635, n28637,
    n28638, n28639, n28640, n28641, n28643, n28644, n28645, n28646, n28647,
    n28649, n28650, n28651, n28652, n28653, n28655, n28656, n28657, n28658,
    n28659, n28661, n28662, n28663, n28664, n28665, n28667, n28668, n28669,
    n28670, n28671, n28673, n28674, n28675, n28676, n28677, n28679, n28680,
    n28681, n28682, n28683, n28685, n28686, n28687, n28688, n28689, n28691,
    n28692, n28693, n28694, n28695, n28697, n28698, n28699, n28700, n28701,
    n28703, n28704, n28705, n28706, n28707, n28709, n28710, n28711, n28712,
    n28713, n28715, n28716, n28718, n28719, n28720, n28721, n28722, n28724,
    n28725, n28726, n28727, n28728, n28730, n28731, n28732, n28733, n28734,
    n28736, n28737, n28739, n28740, n28741, n28742, n28743, n28745, n28746,
    n28748, n28749, n28751, n28752, n28754, n28755, n28757, n28758, n28759,
    n28760, n28761, n28763, n28764, n28766, n28767, n28769, n28770, n28772,
    n28773, n28775, n28776, n28778, n28779, n28781, n28782, n28784, n28785,
    n28787, n28788, n28790, n28791, n28793, n28794, n28795, n28796, n28797,
    n28799, n28800, n28802, n28803, n28804, n28805, n28806, n28808, n28809,
    n28811, n28812, n28814, n28815, n28816, n28817, n28818, n28820, n28821,
    n28823, n28824, n28826, n28827, n28829, n28830, n28832, n28833, n28835,
    n28836, n28838, n28839, n28841, n28842, n28844, n28845, n28847, n28848,
    n28850, n28851, n28853, n28854, n28856, n28857, n28859, n28860, n28861,
    n28862, n28864, n28865, n28866, n28867, n28868, n28870, n28871, n28872,
    n28873, n28874, n28876, n28877, n28878, n28879, n28880, n28882, n28883,
    n28884, n28885, n28886, n28888, n28889, n28890, n28891, n28892, n28894,
    n28895, n28896, n28897, n28898, n28900, n28901, n28902, n28903, n28904,
    n28906, n28907, n28908, n28909, n28910, n28912, n28913, n28914, n28915,
    n28916, n28918, n28919, n28921, n28922, n28924, n28925, n28926, n28927,
    n28928, n28930, n28931, n28932, n28933, n28934, n28936, n28937, n28939,
    n28940, n28942, n28943, n28944, n28945, n28946, n28948, n28949, n28950,
    n28951, n28952, n28954, n28955, n28956, n28957, n28958, n28960, n28961,
    n28962, n28963, n28964, n28966, n28967, n28969, n28970, n28972, n28973,
    n28974, n28975, n28976, n28978, n28979, n28980, n28981, n28982, n28984,
    n28985, n28986, n28987, n28988, n28990, n28991, n28992, n28993, n28994,
    n28996, n28997, n28998, n28999, n29000, n29002, n29003, n29005, n29006,
    n29007, n29008, n29009, n29011, n29012, n29013, n29014, n29015, n29017,
    n29018, n29020, n29021, n29022, n29023, n29024, n29026, n29027, n29029,
    n29030, n29032, n29033, n29034, n29036, n29037, n29038, n29039, n29040,
    n29041, n29042, n29043, n29044, n29046, n29047, n29049, n29050, n29051,
    n29052, n29053, n29055, n29056, n29057, n29059, n29060, n29061, n29063,
    n29064, n29065, n29066, n29067, n29069, n29071, n29072, n29074, n29075,
    n29077, n29078, n29080, n29081, n29083, n29084, n29085, n29086, n29087,
    n29089, n29090, n29092, n29094, n29095, n29098, n29099, n29100, n29101,
    n29102, n29104, n29105, n29106, n29107, n29108, n29110, n29111, n29112,
    n29113, n29114, n29116, n29117, n29118, n29119, n29120, n29122, n29123,
    n29124, n29125, n29126, n29128, n29129, n29130, n29131, n29132, n29134,
    n29135, n29136, n29137, n29138, n29140, n29141, n29142, n29143, n29144,
    n29146, n29147, n29149, n29150, n29152, n29153, n29155, n29157, n29158,
    n29160, n29161, n29162, n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29170, n29171, n29172, n29174, n29175, n29177, n29178, n29180,
    n29181, n29183, n29184, n29185, n29187, n29188, n29190, n29191, n29193,
    n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
    n29203, n29204, n29205, n29206, n29207, n29208, n29210, n29211, n29212,
    n29213, n29214, n29215, n29216, n29217, n29218, n29219, n29220, n29223,
    n29224, n29225, n29226, n29227, n29229, n29230, n29232, n29233, n29234,
    n29235, n29236, n29238, n29239, n29241, n29242, n29243, n29244, n29245,
    n29246, n29248, n29249, n29251, n29252, n29254, n29255, n29257, n29258,
    n29259, n29261, n29262, n29264, n29265, n29267, n29268, n29270, n29271,
    n29272, n29273, n29275, n29276, n29277, n29279, n29281, n29282, n29284,
    n29285, n29287, n29288, n29293, n29295, n29296, n29298, n29299, n29300,
    n29301, n29302, n29303, n29305, n29306, n29308, n29309, n29310, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
    n29322, n29323, n29325, n29327, n29328, n29330, n29331, n29332, n29334,
    n29335, n29336, n29338, n29339, n29341, n29342, n29344, n29345, n29347,
    n29348, n29350, n29351, n29352, n29354, n29356, n29357, n29359, n29360,
    n29361, n29363, n29364, n29366, n29368, n29370, n29371, n29373, n29375,
    n29376, n29378, n29379, n29381, n29382, n29384, n29385, n29387, n29388,
    n29389, n29391, n29392, n29394, n29396, n29397, n29400, n29402, n29403,
    n29405, n29406, n29408, n29409, n29411, n29412, n29414, n29415, n29417,
    n29418, n29420, n29421, n29423, n29424, n29426, n29427, n29429, n29430,
    n29432, n29433, n29435, n29436, n29438, n29439, n29441, n29442, n29444,
    n29445, n29447, n29448, n29450, n29451, n29453, n29454, n29456, n29457,
    n29459, n29460, n29462, n29463, n29465, n29466, n29468, n29469, n29471,
    n29473, n29474, n29476, n29477, n29479, n29480, n29482, n29483, n29485,
    n29486, n29488, n29489, n29491, n29492, n29494, n29495, n29497, n29499,
    n29500, n29502, n29503, n29505, n29506, n29508, n29509, n29511, n29512,
    n29514, n29515, n29517, n29518, n29520, n29521, n29523, n29524, n29526,
    n29527, n29529, n29530, n29532, n29533, n29535, n29536, n29538, n29539,
    n29541, n29542, n29544, n29545, n29547, n29548, n29550, n29551, n29553,
    n29554, n29556, n29557, n29559, n29560, n29562, n29563, n29565, n29566,
    n29568, n29569, n29571, n29572, n29574, n29575, n29577, n29578, n29580,
    n29581, n29583, n29584, n29586, n29587, n29589, n29590, n29592, n29593,
    n29595, n29596, n29598, n29599, n29601, n29602, n29604, n29605, n29607,
    n29608, n29610, n29611, n29613, n29614, n29616, n29617, n29619, n29620,
    n29622, n29623, n29625, n29626, n29628, n29629, n29631, n29633, n29634,
    n29636, n29637, n29639, n29640, n29642, n29643, n29645, n29646, n29648,
    n29649, n29651, n29652, n29654, n29655, n29657, n29658, n29660, n29661,
    n29663, n29664, n29666, n29667, n29669, n29670, n29672, n29673, n29675,
    n29676, n29678, n29679, n29681, n29682, n29684, n29685, n29687, n29688,
    n29691, n29693, n29694, n29696, n29698, n29699, n29701, n29703, n29705,
    n29707, n29708, n29710, n29711, n29713, n29714, n29716, n29717, n29719,
    n29720, n29722, n29723, n29725, n29726, n29728, n29729, n29731, n29733,
    n29734, n29737, n29738, n29739, n29741, n29742, n29744, n29745, n29747,
    n29748, n29750, n29751, n29753, n29754, n29756, n29757, n29759, n29760,
    n29763, n29766, n29767, n29769, n29770, n29772, n29773, n29774, n29776,
    n29777, n29779, n29780, n29782, n29783, n29785, n29786, n29788, n29789,
    n29791, n29792, n29794, n29795, n29797, n29798, n29800, n29801, n29803,
    n29804, n29806, n29807, n29809, n29810, n29812, n29813, n29815, n29816,
    n29819, n29820, n29822, n29823, n29825, n29826, n29828, n29829, n29831,
    n29832, n29834, n29835, n29837, n29838, n29840, n29841, n29843, n29844,
    n29846, n29847, n29849, n29850;
  assign po0000 = pi1677 | ~pi3368;
  assign n7050 = ~pi0315 & ~pi3235;
  assign n7051 = pi0315 & pi3235;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = ~pi0314 & ~pi3229;
  assign n7054 = pi0314 & pi3229;
  assign n7055 = ~n7053 & ~n7054;
  assign n7056 = ~n7052 & ~n7055;
  assign n7057 = ~pi0313 & pi3225;
  assign n7058 = pi0313 & ~pi3225;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = n7056 & n7059;
  assign n7061 = ~pi0085 & ~n7060;
  assign n7062 = ~pi1687 & pi1778;
  assign n7063 = ~pi0452 & n7062;
  assign n7064 = n7061 & n7063;
  assign n7065 = pi0452 & ~pi1778;
  assign n7066 = ~pi1687 & n7065;
  assign n7067 = ~pi3364 & ~pi3366;
  assign n7068 = pi3365 & n7067;
  assign n7069 = pi1233 & pi1258;
  assign n7070 = pi1234 & n7069;
  assign n7071 = pi1237 & pi1257;
  assign n7072 = ~pi1228 & pi1236;
  assign n7073 = pi1238 & n7072;
  assign n7074 = n7071 & n7073;
  assign n7075 = n7070 & n7074;
  assign n7076 = n7068 & n7075;
  assign n7077 = ~pi3365 & pi3366;
  assign n7078 = ~pi3364 & n7077;
  assign n7079 = n7061 & n7078;
  assign n7080 = ~n7076 & ~n7079;
  assign n7081 = n7066 & ~n7080;
  assign n7082 = ~pi3365 & ~pi3366;
  assign n7083 = pi3364 & n7082;
  assign n7084 = ~n7068 & ~n7078;
  assign n7085 = ~n7083 & n7084;
  assign n7086 = pi3102 & pi3112;
  assign n7087 = ~pi3007 & ~pi3111;
  assign n7088 = pi1813 & n7087;
  assign n7089 = pi3034 & n7088;
  assign n7090 = n7086 & n7089;
  assign n7091 = pi3034 & ~pi3111;
  assign n7092 = pi3007 & n7091;
  assign n7093 = pi3112 & n7092;
  assign n7094 = n7086 & n7091;
  assign n7095 = ~n7093 & ~n7094;
  assign n7096 = pi1813 & n7093;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = ~n7090 & n7097;
  assign n7099 = n7083 & n7098;
  assign n7100 = ~n7085 & ~n7099;
  assign n7101 = pi0452 & n7062;
  assign n7102 = ~n7100 & n7101;
  assign n7103 = ~n7081 & ~n7102;
  assign n7104 = ~pi1332 & pi1686;
  assign n7105 = ~n7057 & n7104;
  assign n7106 = ~n7058 & n7105;
  assign n7107 = ~n7052 & n7106;
  assign n7108 = ~n7055 & n7107;
  assign n7109 = ~pi0452 & ~pi1778;
  assign n7110 = ~pi1687 & n7109;
  assign n7111 = n7108 & n7110;
  assign n7112 = n7103 & ~n7111;
  assign po1955 = n7064 | ~n7112;
  assign n7114 = ~pi0222 & n7068;
  assign n7115 = ~n7078 & ~n7114;
  assign n7116 = n7083 & ~n7098;
  assign n7117 = n7115 & ~n7116;
  assign n7118 = ~n7076 & n7117;
  assign n7119 = n7101 & ~n7118;
  assign n7120 = ~n7061 & n7083;
  assign n7121 = n7066 & n7120;
  assign n7122 = ~n7061 & n7078;
  assign n7123 = n7066 & n7122;
  assign n7124 = pi1687 & n7109;
  assign n7125 = pi1686 & n7124;
  assign n7126 = ~n7123 & ~n7125;
  assign n7127 = ~n7121 & n7126;
  assign po1864 = n7119 | ~n7127;
  assign n7129 = ~po1955 & ~po1864;
  assign n7130 = ~n7108 & n7110;
  assign n7131 = pi1332 & n7130;
  assign n7132 = ~n7078 & ~n7085;
  assign n7133 = ~n7083 & n7132;
  assign n7134 = ~n7114 & n7133;
  assign n7135 = n7101 & ~n7134;
  assign n7136 = ~n7111 & ~n7135;
  assign n7137 = ~pi2967 & n7108;
  assign n7138 = ~n7055 & ~n7057;
  assign n7139 = ~n7058 & n7104;
  assign n7140 = n7138 & n7139;
  assign n7141 = ~n7052 & n7140;
  assign n7142 = ~pi2967 & pi3254;
  assign n7143 = ~n7141 & n7142;
  assign n7144 = pi1332 & n7143;
  assign n7145 = pi0085 & n7144;
  assign n7146 = ~n7137 & ~n7145;
  assign po1399 = n7110 & ~n7146;
  assign n7148 = ~pi0083 & pi0084;
  assign n7149 = ~n7060 & n7148;
  assign n7150 = ~po1399 & n7149;
  assign n7151 = pi3034 & n7110;
  assign n7152 = n7108 & n7151;
  assign n7153 = pi3125 & ~pi3242;
  assign n7154 = pi3188 & ~n7087;
  assign n7155 = pi3243 & ~pi3247;
  assign n7156 = ~pi3244 & n7155;
  assign n7157 = ~pi3245 & n7156;
  assign n7158 = n7154 & n7157;
  assign n7159 = pi3125 & n7158;
  assign n7160 = ~n7153 & ~n7159;
  assign n7161 = pi3125 & ~n7158;
  assign n7162 = n7160 & ~n7161;
  assign n7163 = n7152 & ~n7162;
  assign n7164 = ~n7146 & n7163;
  assign n7165 = ~pi0975 & ~n7164;
  assign n7166 = ~n7150 & n7165;
  assign n7167 = pi0076 & n7061;
  assign n7168 = ~n7166 & n7167;
  assign n7169 = n7083 & ~n7168;
  assign n7170 = n7066 & n7169;
  assign n7171 = ~n7085 & ~n7122;
  assign n7172 = n7066 & ~n7171;
  assign n7173 = ~n7170 & ~n7172;
  assign n7174 = n7136 & n7173;
  assign po0652 = n7131 | ~n7174;
  assign n7176 = n7129 & po0652;
  assign n7177 = po1955 & ~po1864;
  assign n7178 = po0652 & n7177;
  assign n7179 = ~n7176 & n7178;
  assign n7180 = pi0339 & pi2967;
  assign n7181 = pi0340 & pi3364;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = ~pi1219 & n7182;
  assign n7184 = pi1725 & ~pi1796;
  assign n7185 = ~n7166 & ~n7184;
  assign n7186 = ~n7183 & ~n7185;
  assign n7187 = n7179 & n7186;
  assign n7188 = pi0339 & ~pi3254;
  assign n7189 = n7183 & ~n7188;
  assign n7190 = n7068 & n7070;
  assign n7191 = ~pi0085 & n7190;
  assign n7192 = n7074 & n7191;
  assign n7193 = ~n7060 & n7192;
  assign n7194 = ~n7060 & n7078;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = pi0076 & n7195;
  assign n7197 = ~n7166 & n7196;
  assign n7198 = n7061 & n7083;
  assign n7199 = n7195 & ~n7198;
  assign n7200 = n7066 & ~n7199;
  assign n7201 = ~n7197 & n7200;
  assign n7202 = ~pi2967 & ~n7141;
  assign n7203 = pi1332 & n7202;
  assign n7204 = n7110 & n7203;
  assign n7205 = ~pi1219 & ~n7204;
  assign n7206 = ~n7064 & n7205;
  assign n7207 = ~n7201 & n7206;
  assign n7208 = ~n7166 & n7207;
  assign n7209 = pi0113 & n7208;
  assign n7210 = ~n7189 & ~n7209;
  assign n7211 = pi0322 & pi3229;
  assign n7212 = ~pi0322 & ~pi3229;
  assign n7213 = ~n7211 & ~n7212;
  assign n7214 = pi0321 & pi3225;
  assign n7215 = ~pi0321 & ~pi3225;
  assign n7216 = ~n7214 & ~n7215;
  assign n7217 = n7213 & n7216;
  assign n7218 = pi0323 & pi3235;
  assign n7219 = ~pi0323 & ~pi3235;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = n7217 & n7220;
  assign n7222 = pi0113 & ~n7221;
  assign n7223 = ~pi0083 & n7222;
  assign n7224 = ~n7166 & n7223;
  assign n7225 = n7210 & ~n7224;
  assign n7226 = pi0000 & n7189;
  assign n7227 = ~n7225 & ~n7226;
  assign n7228 = n7176 & ~n7178;
  assign n7229 = ~n7227 & n7228;
  assign n7230 = pi0000 & n7179;
  assign n7231 = n7183 & n7230;
  assign n7232 = ~n7229 & ~n7231;
  assign po0205 = n7187 | ~n7232;
  assign n7234 = pi0001 & n7189;
  assign n7235 = ~n7225 & ~n7234;
  assign n7236 = n7228 & ~n7235;
  assign n7237 = pi0001 & n7179;
  assign n7238 = n7183 & n7237;
  assign n7239 = ~n7236 & ~n7238;
  assign po0206 = n7187 | ~n7239;
  assign n7241 = ~pi2995 & ~pi3001;
  assign n7242 = ~pi2982 & ~pi2996;
  assign n7243 = ~pi2981 & ~pi2997;
  assign n7244 = n7242 & n7243;
  assign n7245 = n7241 & n7244;
  assign n7246 = pi2920 & ~pi2966;
  assign n7247 = n7245 & n7246;
  assign n7248 = ~pi3018 & pi3138;
  assign n7249 = n7247 & n7248;
  assign n7250 = ~pi1335 & ~pi2984;
  assign n7251 = ~pi3129 & ~n7250;
  assign n7252 = ~pi3120 & pi3207;
  assign n7253 = n7251 & n7252;
  assign n7254 = pi2969 & n7253;
  assign n7255 = n7249 & n7254;
  assign n7256 = pi0002 & ~n7255;
  assign n7257 = pi1379 & pi3160;
  assign n7258 = pi0071 & n7257;
  assign n7259 = ~pi0202 & ~n7258;
  assign n7260 = ~pi3144 & ~n7259;
  assign po0208 = n7256 | n7260;
  assign n7262 = pi2971 & n7178;
  assign n7263 = ~n7176 & ~n7178;
  assign n7264 = pi0003 & n7263;
  assign n7265 = ~n7262 & ~n7264;
  assign n7266 = ~n7166 & n7178;
  assign n7267 = ~po1399 & ~n7207;
  assign n7268 = ~pi1219 & ~n7267;
  assign n7269 = ~pi0109 & ~n7268;
  assign n7270 = pi0003 & n7268;
  assign n7271 = ~n7269 & ~n7270;
  assign n7272 = n7176 & ~n7271;
  assign n7273 = ~n7266 & ~n7272;
  assign po0209 = ~n7265 | ~n7273;
  assign n7275 = pi3016 & n7178;
  assign n7276 = pi0004 & n7263;
  assign n7277 = ~n7275 & ~n7276;
  assign n7278 = ~pi0110 & ~n7268;
  assign n7279 = pi0004 & n7268;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = n7176 & ~n7280;
  assign n7282 = ~n7266 & ~n7281;
  assign po0210 = ~n7277 | ~n7282;
  assign n7284 = pi3064 & n7178;
  assign n7285 = pi0005 & n7263;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 = ~pi0111 & ~n7268;
  assign n7288 = pi0005 & n7268;
  assign n7289 = ~n7287 & ~n7288;
  assign n7290 = n7176 & ~n7289;
  assign n7291 = ~n7266 & ~n7290;
  assign po0211 = ~n7286 | ~n7291;
  assign n7293 = pi3070 & n7178;
  assign n7294 = pi0006 & n7263;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = ~pi0112 & ~n7268;
  assign n7297 = pi0006 & n7268;
  assign n7298 = ~n7296 & ~n7297;
  assign n7299 = n7176 & ~n7298;
  assign n7300 = ~n7266 & ~n7299;
  assign po0212 = ~n7295 | ~n7300;
  assign n7302 = pi0007 & ~n7176;
  assign n7303 = pi0089 & ~n7268;
  assign n7304 = pi0007 & n7268;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = n7176 & ~n7305;
  assign po0213 = n7302 | n7306;
  assign n7308 = pi0008 & ~n7176;
  assign n7309 = pi0086 & ~n7268;
  assign n7310 = pi0008 & n7268;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = n7176 & ~n7311;
  assign po0214 = n7308 | n7312;
  assign n7314 = pi0009 & ~n7176;
  assign n7315 = pi0087 & ~n7268;
  assign n7316 = pi0009 & n7268;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = n7176 & ~n7317;
  assign po0215 = n7314 | n7318;
  assign n7320 = pi0010 & ~n7176;
  assign n7321 = pi0088 & ~n7268;
  assign n7322 = pi0010 & n7268;
  assign n7323 = ~n7321 & ~n7322;
  assign n7324 = n7176 & ~n7323;
  assign po0216 = n7320 | n7324;
  assign n7326 = pi0011 & ~n7176;
  assign n7327 = pi0090 & ~n7268;
  assign n7328 = pi0011 & n7268;
  assign n7329 = ~n7327 & ~n7328;
  assign n7330 = n7176 & ~n7329;
  assign po0217 = n7326 | n7330;
  assign n7332 = pi0012 & ~n7176;
  assign n7333 = pi0091 & ~n7268;
  assign n7334 = pi0012 & n7268;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = n7176 & ~n7335;
  assign po0218 = n7332 | n7336;
  assign n7338 = pi0013 & ~n7176;
  assign n7339 = pi0093 & ~n7268;
  assign n7340 = pi0013 & n7268;
  assign n7341 = ~n7339 & ~n7340;
  assign n7342 = n7176 & ~n7341;
  assign po0219 = n7338 | n7342;
  assign n7344 = pi0014 & ~n7176;
  assign n7345 = pi0094 & ~n7268;
  assign n7346 = pi0014 & n7268;
  assign n7347 = ~n7345 & ~n7346;
  assign n7348 = n7176 & ~n7347;
  assign po0220 = n7344 | n7348;
  assign n7350 = pi0015 & ~n7176;
  assign n7351 = pi0095 & ~n7268;
  assign n7352 = pi0015 & n7268;
  assign n7353 = ~n7351 & ~n7352;
  assign n7354 = n7176 & ~n7353;
  assign po0221 = n7350 | n7354;
  assign n7356 = pi0016 & ~n7176;
  assign n7357 = pi0096 & ~n7268;
  assign n7358 = pi0016 & n7268;
  assign n7359 = ~n7357 & ~n7358;
  assign n7360 = n7176 & ~n7359;
  assign po0222 = n7356 | n7360;
  assign n7362 = pi0017 & ~n7176;
  assign n7363 = pi0097 & ~n7268;
  assign n7364 = pi0017 & n7268;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = n7176 & ~n7365;
  assign po0223 = n7362 | n7366;
  assign n7368 = pi0018 & ~n7176;
  assign n7369 = pi0018 & n7268;
  assign n7370 = pi0098 & ~n7268;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = n7176 & ~n7371;
  assign po0224 = n7368 | n7372;
  assign n7374 = pi0019 & ~n7176;
  assign n7375 = pi0099 & ~n7268;
  assign n7376 = pi0019 & n7268;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = n7176 & ~n7377;
  assign po0225 = n7374 | n7378;
  assign n7380 = pi0020 & ~n7176;
  assign n7381 = pi0100 & ~n7268;
  assign n7382 = pi0020 & n7268;
  assign n7383 = ~n7381 & ~n7382;
  assign n7384 = n7176 & ~n7383;
  assign po0226 = n7380 | n7384;
  assign n7386 = pi0021 & ~n7176;
  assign n7387 = pi0101 & ~n7268;
  assign n7388 = pi0021 & n7268;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = n7176 & ~n7389;
  assign po0227 = n7386 | n7390;
  assign n7392 = pi0022 & ~n7176;
  assign n7393 = pi0102 & ~n7268;
  assign n7394 = pi0022 & n7268;
  assign n7395 = ~n7393 & ~n7394;
  assign n7396 = n7176 & ~n7395;
  assign po0228 = n7392 | n7396;
  assign n7398 = pi0023 & ~n7176;
  assign n7399 = pi0103 & ~n7268;
  assign n7400 = pi0023 & n7268;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = n7176 & ~n7401;
  assign po0229 = n7398 | n7402;
  assign n7404 = pi0024 & ~n7176;
  assign n7405 = pi0104 & ~n7268;
  assign n7406 = pi0024 & n7268;
  assign n7407 = ~n7405 & ~n7406;
  assign n7408 = n7176 & ~n7407;
  assign po0230 = n7404 | n7408;
  assign n7410 = pi0025 & ~n7176;
  assign n7411 = pi0105 & ~n7268;
  assign n7412 = pi0025 & n7268;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = n7176 & ~n7413;
  assign po0231 = n7410 | n7414;
  assign n7416 = pi0026 & ~n7176;
  assign n7417 = pi0106 & ~n7268;
  assign n7418 = pi0026 & n7268;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = n7176 & ~n7419;
  assign po0232 = n7416 | n7420;
  assign n7422 = pi0027 & ~n7176;
  assign n7423 = pi0108 & ~n7268;
  assign n7424 = pi0027 & n7268;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = n7176 & ~n7425;
  assign po0233 = n7422 | n7426;
  assign n7428 = pi0028 & ~n7176;
  assign n7429 = pi0114 & ~n7268;
  assign n7430 = pi0028 & n7268;
  assign n7431 = ~n7429 & ~n7430;
  assign n7432 = n7176 & ~n7431;
  assign po0234 = n7428 | n7432;
  assign n7434 = pi0029 & ~n7176;
  assign n7435 = pi0115 & ~n7268;
  assign n7436 = pi0029 & n7268;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = n7176 & ~n7437;
  assign po0235 = n7434 | n7438;
  assign n7440 = pi0030 & ~n7176;
  assign n7441 = pi0116 & ~n7268;
  assign n7442 = pi0030 & n7268;
  assign n7443 = ~n7441 & ~n7442;
  assign n7444 = n7176 & ~n7443;
  assign po0236 = n7440 | n7444;
  assign n7446 = pi0031 & ~n7176;
  assign n7447 = pi0117 & ~n7268;
  assign n7448 = pi0031 & n7268;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = n7176 & ~n7449;
  assign po0237 = n7446 | n7450;
  assign n7452 = pi0032 & ~n7176;
  assign n7453 = pi0118 & ~n7268;
  assign n7454 = pi0032 & n7268;
  assign n7455 = ~n7453 & ~n7454;
  assign n7456 = n7176 & ~n7455;
  assign po0238 = n7452 | n7456;
  assign n7458 = pi0033 & ~n7176;
  assign n7459 = pi0119 & ~n7268;
  assign n7460 = pi0033 & n7268;
  assign n7461 = ~n7459 & ~n7460;
  assign n7462 = n7176 & ~n7461;
  assign po0239 = n7458 | n7462;
  assign n7464 = pi0034 & ~n7176;
  assign n7465 = pi0107 & ~n7268;
  assign n7466 = pi0034 & n7268;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = n7176 & ~n7467;
  assign po0240 = n7464 | n7468;
  assign n7470 = pi0035 & ~n7176;
  assign n7471 = pi0092 & ~n7268;
  assign n7472 = pi0035 & n7268;
  assign n7473 = ~n7471 & ~n7472;
  assign n7474 = n7176 & ~n7473;
  assign po0241 = n7470 | n7474;
  assign n7476 = pi0036 & ~n7176;
  assign n7477 = pi0123 & ~n7268;
  assign n7478 = pi0036 & n7268;
  assign n7479 = ~n7477 & ~n7478;
  assign n7480 = n7176 & ~n7479;
  assign po0242 = n7476 | n7480;
  assign n7482 = pi0037 & ~n7176;
  assign n7483 = pi0124 & ~n7268;
  assign n7484 = pi0037 & n7268;
  assign n7485 = ~n7483 & ~n7484;
  assign n7486 = n7176 & ~n7485;
  assign po0243 = n7482 | n7486;
  assign n7488 = pi0038 & ~n7176;
  assign n7489 = pi0122 & ~n7268;
  assign n7490 = pi0038 & n7268;
  assign n7491 = ~n7489 & ~n7490;
  assign n7492 = n7176 & ~n7491;
  assign po0244 = n7488 | n7492;
  assign n7494 = n7083 & ~n7101;
  assign n7495 = n7066 & n7494;
  assign n7496 = n7083 & n7101;
  assign n7497 = ~n7066 & n7496;
  assign n7498 = ~n7495 & ~n7497;
  assign n7499 = pi0039 & n7498;
  assign n7500 = pi0061 & pi0062;
  assign n7501 = pi0059 & n7500;
  assign n7502 = pi0060 & n7501;
  assign n7503 = pi0051 & pi0064;
  assign n7504 = pi0063 & pi0068;
  assign n7505 = n7503 & n7504;
  assign n7506 = pi0052 & pi0053;
  assign n7507 = pi0055 & pi0056;
  assign n7508 = n7506 & n7507;
  assign n7509 = n7505 & n7508;
  assign n7510 = n7502 & n7509;
  assign n7511 = pi0054 & pi0067;
  assign n7512 = pi0050 & pi0066;
  assign n7513 = n7511 & n7512;
  assign n7514 = n7510 & n7513;
  assign n7515 = pi0065 & n7514;
  assign n7516 = pi0039 & ~n7515;
  assign n7517 = ~pi0039 & n7515;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = ~n7498 & ~n7518;
  assign n7520 = ~n7499 & ~n7519;
  assign n7521 = ~po1399 & ~n7520;
  assign n7522 = pi3072 & n7108;
  assign n7523 = pi0094 & ~n7108;
  assign n7524 = ~n7522 & ~n7523;
  assign n7525 = po1399 & ~n7524;
  assign po0245 = n7521 | n7525;
  assign n7527 = pi0040 & n7498;
  assign n7528 = pi0055 & pi0067;
  assign n7529 = pi0050 & pi0054;
  assign n7530 = n7528 & n7529;
  assign n7531 = pi0039 & pi0066;
  assign n7532 = pi0042 & pi0044;
  assign n7533 = n7531 & n7532;
  assign n7534 = n7530 & n7533;
  assign n7535 = pi0059 & pi0065;
  assign n7536 = pi0060 & n7535;
  assign n7537 = pi0061 & n7536;
  assign n7538 = pi0063 & pi0064;
  assign n7539 = pi0062 & pi0068;
  assign n7540 = n7538 & n7539;
  assign n7541 = pi0051 & pi0052;
  assign n7542 = pi0053 & pi0056;
  assign n7543 = n7541 & n7542;
  assign n7544 = n7540 & n7543;
  assign n7545 = n7537 & n7544;
  assign n7546 = n7534 & n7545;
  assign n7547 = pi0040 & ~n7546;
  assign n7548 = ~pi0040 & n7546;
  assign n7549 = ~n7547 & ~n7548;
  assign n7550 = ~n7498 & ~n7549;
  assign n7551 = ~n7527 & ~n7550;
  assign n7552 = ~po1399 & ~n7551;
  assign n7553 = pi3005 & n7108;
  assign n7554 = pi0098 & ~n7108;
  assign n7555 = ~n7553 & ~n7554;
  assign n7556 = po1399 & ~n7555;
  assign po0246 = n7552 | n7556;
  assign n7558 = pi0041 & n7498;
  assign n7559 = n7529 & n7531;
  assign n7560 = pi0060 & pi0061;
  assign n7561 = n7539 & n7560;
  assign n7562 = n7535 & n7561;
  assign n7563 = n7538 & n7541;
  assign n7564 = n7528 & n7542;
  assign n7565 = n7563 & n7564;
  assign n7566 = pi0040 & pi0057;
  assign n7567 = n7532 & n7566;
  assign n7568 = n7565 & n7567;
  assign n7569 = n7562 & n7568;
  assign n7570 = n7559 & n7569;
  assign n7571 = pi0041 & ~n7570;
  assign n7572 = ~pi0041 & n7570;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = ~n7498 & ~n7573;
  assign n7575 = ~n7558 & ~n7574;
  assign n7576 = ~po1399 & ~n7575;
  assign n7577 = pi3030 & n7108;
  assign n7578 = pi0100 & ~n7108;
  assign n7579 = ~n7577 & ~n7578;
  assign n7580 = po1399 & ~n7579;
  assign po0247 = n7576 | n7580;
  assign n7582 = pi0042 & n7498;
  assign n7583 = n7561 & n7565;
  assign n7584 = n7535 & n7583;
  assign n7585 = n7559 & n7584;
  assign n7586 = pi0042 & ~n7585;
  assign n7587 = ~pi0042 & n7585;
  assign n7588 = ~n7586 & ~n7587;
  assign n7589 = ~n7498 & ~n7588;
  assign n7590 = ~n7582 & ~n7589;
  assign n7591 = ~po1399 & ~n7590;
  assign n7592 = pi3033 & n7108;
  assign n7593 = pi0096 & ~n7108;
  assign n7594 = ~n7592 & ~n7593;
  assign n7595 = po1399 & ~n7594;
  assign po0248 = n7591 | n7595;
  assign n7597 = pi0043 & n7498;
  assign n7598 = pi0039 & pi0042;
  assign n7599 = pi0040 & pi0044;
  assign n7600 = n7598 & n7599;
  assign n7601 = pi0041 & pi0057;
  assign n7602 = pi0046 & pi0058;
  assign n7603 = n7601 & n7602;
  assign n7604 = pi0065 & n7502;
  assign n7605 = n7505 & n7604;
  assign n7606 = n7508 & n7605;
  assign n7607 = n7513 & n7606;
  assign n7608 = n7603 & n7607;
  assign n7609 = n7600 & n7608;
  assign n7610 = pi0043 & ~n7609;
  assign n7611 = ~pi0043 & n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n7498 & ~n7612;
  assign n7614 = ~n7597 & ~n7613;
  assign n7615 = ~po1399 & ~n7614;
  assign n7616 = pi3044 & n7108;
  assign n7617 = pi0103 & ~n7108;
  assign n7618 = ~n7616 & ~n7617;
  assign n7619 = po1399 & ~n7618;
  assign po0249 = n7615 | n7619;
  assign n7621 = pi0044 & n7498;
  assign n7622 = n7503 & n7506;
  assign n7623 = n7507 & n7511;
  assign n7624 = n7622 & n7623;
  assign n7625 = n7512 & n7598;
  assign n7626 = n7624 & n7625;
  assign n7627 = n7500 & n7504;
  assign n7628 = n7536 & n7627;
  assign n7629 = n7626 & n7628;
  assign n7630 = pi0044 & ~n7629;
  assign n7631 = ~pi0044 & n7629;
  assign n7632 = ~n7630 & ~n7631;
  assign n7633 = ~n7498 & ~n7632;
  assign n7634 = ~n7621 & ~n7633;
  assign n7635 = ~po1399 & ~n7634;
  assign n7636 = pi3006 & n7108;
  assign n7637 = pi0097 & ~n7108;
  assign n7638 = ~n7636 & ~n7637;
  assign n7639 = po1399 & ~n7638;
  assign po0250 = n7635 | n7639;
  assign n7641 = pi0045 & n7498;
  assign n7642 = pi0041 & pi0046;
  assign n7643 = n7566 & n7642;
  assign n7644 = n7537 & n7540;
  assign n7645 = n7543 & n7644;
  assign n7646 = n7534 & n7645;
  assign n7647 = n7643 & n7646;
  assign n7648 = pi0043 & pi0058;
  assign n7649 = pi0047 & n7648;
  assign n7650 = pi0049 & n7649;
  assign n7651 = n7647 & n7650;
  assign n7652 = pi0045 & ~n7651;
  assign n7653 = ~pi0045 & n7651;
  assign n7654 = ~n7652 & ~n7653;
  assign n7655 = ~n7498 & ~n7654;
  assign n7656 = ~n7641 & ~n7655;
  assign n7657 = ~po1399 & ~n7656;
  assign n7658 = pi3074 & n7108;
  assign n7659 = pi0107 & ~n7108;
  assign n7660 = ~n7658 & ~n7659;
  assign n7661 = po1399 & ~n7660;
  assign po0251 = n7657 | n7661;
  assign n7663 = pi0046 & n7498;
  assign n7664 = n7599 & n7601;
  assign n7665 = n7624 & n7664;
  assign n7666 = n7628 & n7665;
  assign n7667 = n7625 & n7666;
  assign n7668 = pi0046 & ~n7667;
  assign n7669 = ~pi0046 & n7667;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~n7498 & ~n7670;
  assign n7672 = ~n7663 & ~n7671;
  assign n7673 = ~po1399 & ~n7672;
  assign n7674 = pi3029 & n7108;
  assign n7675 = pi0101 & ~n7108;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = po1399 & ~n7676;
  assign po0252 = n7673 | n7677;
  assign n7679 = pi0047 & n7498;
  assign n7680 = n7562 & n7563;
  assign n7681 = n7567 & n7680;
  assign n7682 = n7564 & n7681;
  assign n7683 = n7559 & n7642;
  assign n7684 = n7648 & n7683;
  assign n7685 = n7682 & n7684;
  assign n7686 = pi0047 & ~n7685;
  assign n7687 = ~pi0047 & n7685;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n7498 & ~n7688;
  assign n7690 = ~n7679 & ~n7689;
  assign n7691 = ~po1399 & ~n7690;
  assign n7692 = pi3032 & n7108;
  assign n7693 = pi0104 & ~n7108;
  assign n7694 = ~n7692 & ~n7693;
  assign n7695 = po1399 & ~n7694;
  assign po0253 = n7691 | n7695;
  assign n7697 = pi0048 & n7498;
  assign n7698 = n7513 & n7600;
  assign n7699 = n7606 & n7698;
  assign n7700 = n7603 & n7699;
  assign n7701 = pi0043 & pi0047;
  assign n7702 = pi0049 & n7701;
  assign n7703 = pi0045 & n7702;
  assign n7704 = n7700 & n7703;
  assign n7705 = pi0048 & ~n7704;
  assign n7706 = ~pi0048 & n7704;
  assign n7707 = ~n7705 & ~n7706;
  assign n7708 = ~n7498 & ~n7707;
  assign n7709 = ~n7697 & ~n7708;
  assign n7710 = ~po1399 & ~n7709;
  assign n7711 = pi3051 & n7108;
  assign n7712 = pi0108 & ~n7108;
  assign n7713 = ~n7711 & ~n7712;
  assign n7714 = po1399 & ~n7713;
  assign po0254 = n7710 | n7714;
  assign n7716 = pi0049 & n7498;
  assign n7717 = n7622 & n7628;
  assign n7718 = n7664 & n7717;
  assign n7719 = n7623 & n7718;
  assign n7720 = n7602 & n7625;
  assign n7721 = n7701 & n7720;
  assign n7722 = n7719 & n7721;
  assign n7723 = pi0049 & ~n7722;
  assign n7724 = ~pi0049 & n7722;
  assign n7725 = ~n7723 & ~n7724;
  assign n7726 = ~n7498 & ~n7725;
  assign n7727 = ~n7716 & ~n7726;
  assign n7728 = ~po1399 & ~n7727;
  assign n7729 = pi3113 & n7108;
  assign n7730 = pi0105 & ~n7108;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = po1399 & ~n7731;
  assign po0255 = n7728 | n7732;
  assign n7734 = pi0050 & n7498;
  assign n7735 = n7624 & n7628;
  assign n7736 = pi0050 & ~n7735;
  assign n7737 = ~pi0050 & n7735;
  assign n7738 = ~n7736 & ~n7737;
  assign n7739 = ~n7498 & ~n7738;
  assign n7740 = ~n7734 & ~n7739;
  assign n7741 = ~po1399 & ~n7740;
  assign n7742 = pi3116 & n7108;
  assign n7743 = pi0093 & ~n7108;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = po1399 & ~n7744;
  assign po0256 = n7741 | n7745;
  assign n7747 = pi0051 & n7498;
  assign n7748 = pi0051 & ~n7644;
  assign n7749 = ~pi0051 & n7644;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = ~n7498 & ~n7750;
  assign n7752 = ~n7747 & ~n7751;
  assign n7753 = ~po1399 & ~n7752;
  assign n7754 = pi3081 & n7108;
  assign n7755 = pi0086 & ~n7108;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = po1399 & ~n7756;
  assign po0257 = n7753 | n7757;
  assign n7759 = pi0052 & n7498;
  assign n7760 = pi0052 & ~n7605;
  assign n7761 = ~pi0052 & n7605;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = ~n7498 & ~n7762;
  assign n7764 = ~n7759 & ~n7763;
  assign n7765 = ~po1399 & ~n7764;
  assign n7766 = pi3069 & n7108;
  assign n7767 = pi0087 & ~n7108;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = po1399 & ~n7768;
  assign po0258 = n7765 | n7769;
  assign n7771 = pi0053 & n7498;
  assign n7772 = pi0053 & ~n7680;
  assign n7773 = ~pi0053 & n7680;
  assign n7774 = ~n7772 & ~n7773;
  assign n7775 = ~n7498 & ~n7774;
  assign n7776 = ~n7771 & ~n7775;
  assign n7777 = ~po1399 & ~n7776;
  assign n7778 = pi3080 & n7108;
  assign n7779 = pi0088 & ~n7108;
  assign n7780 = ~n7778 & ~n7779;
  assign n7781 = po1399 & ~n7780;
  assign po0259 = n7777 | n7781;
  assign n7783 = pi0054 & n7498;
  assign n7784 = n7564 & n7680;
  assign n7785 = pi0054 & ~n7784;
  assign n7786 = ~pi0054 & n7784;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = ~n7498 & ~n7787;
  assign n7789 = ~n7783 & ~n7788;
  assign n7790 = ~po1399 & ~n7789;
  assign n7791 = pi3013 & n7108;
  assign n7792 = pi0091 & ~n7108;
  assign n7793 = ~n7791 & ~n7792;
  assign n7794 = po1399 & ~n7793;
  assign po0260 = n7790 | n7794;
  assign n7796 = pi0055 & n7498;
  assign n7797 = pi0055 & ~n7645;
  assign n7798 = ~pi0055 & n7645;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = ~n7498 & ~n7799;
  assign n7801 = ~n7796 & ~n7800;
  assign n7802 = ~po1399 & ~n7801;
  assign n7803 = pi3067 & n7108;
  assign n7804 = pi0092 & ~n7108;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = po1399 & ~n7805;
  assign po0261 = n7802 | n7806;
  assign n7808 = pi0056 & n7498;
  assign n7809 = pi0056 & ~n7717;
  assign n7810 = ~pi0056 & n7717;
  assign n7811 = ~n7809 & ~n7810;
  assign n7812 = ~n7498 & ~n7811;
  assign n7813 = ~n7808 & ~n7812;
  assign n7814 = ~po1399 & ~n7813;
  assign n7815 = pi3078 & n7108;
  assign n7816 = pi0090 & ~n7108;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = po1399 & ~n7817;
  assign po0262 = n7814 | n7818;
  assign n7820 = pi0057 & n7498;
  assign n7821 = n7604 & n7698;
  assign n7822 = n7509 & n7821;
  assign n7823 = pi0057 & ~n7822;
  assign n7824 = ~pi0057 & n7822;
  assign n7825 = ~n7823 & ~n7824;
  assign n7826 = ~n7498 & ~n7825;
  assign n7827 = ~n7820 & ~n7826;
  assign n7828 = ~po1399 & ~n7827;
  assign n7829 = pi3031 & n7108;
  assign n7830 = pi0099 & ~n7108;
  assign n7831 = ~n7829 & ~n7830;
  assign n7832 = po1399 & ~n7831;
  assign po0263 = n7828 | n7832;
  assign n7834 = pi0058 & n7498;
  assign n7835 = n7530 & n7645;
  assign n7836 = n7533 & n7643;
  assign n7837 = n7835 & n7836;
  assign n7838 = pi0058 & ~n7837;
  assign n7839 = ~pi0058 & n7837;
  assign n7840 = ~n7838 & ~n7839;
  assign n7841 = ~n7498 & ~n7840;
  assign n7842 = ~n7834 & ~n7841;
  assign n7843 = ~po1399 & ~n7842;
  assign n7844 = pi3028 & n7108;
  assign n7845 = pi0102 & ~n7108;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = po1399 & ~n7846;
  assign po0264 = n7843 | n7847;
  assign n7849 = pi0059 & n7498;
  assign n7850 = ~pi0059 & pi0065;
  assign n7851 = pi0059 & ~pi0065;
  assign n7852 = ~n7850 & ~n7851;
  assign n7853 = ~n7498 & ~n7852;
  assign n7854 = ~n7849 & ~n7853;
  assign n7855 = ~po1399 & ~n7854;
  assign n7856 = pi3076 & n7108;
  assign n7857 = pi0114 & ~n7108;
  assign n7858 = ~n7856 & ~n7857;
  assign n7859 = po1399 & ~n7858;
  assign po0265 = n7855 | n7859;
  assign n7861 = pi0060 & n7498;
  assign n7862 = pi0060 & ~n7535;
  assign n7863 = ~pi0060 & n7535;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = ~n7498 & ~n7864;
  assign n7866 = ~n7861 & ~n7865;
  assign n7867 = ~po1399 & ~n7866;
  assign n7868 = pi3035 & n7108;
  assign n7869 = pi0115 & ~n7108;
  assign n7870 = ~n7868 & ~n7869;
  assign n7871 = po1399 & ~n7870;
  assign po0266 = n7867 | n7871;
  assign n7873 = pi0061 & n7498;
  assign n7874 = pi0061 & ~n7536;
  assign n7875 = ~pi0061 & n7536;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = ~n7498 & ~n7876;
  assign n7878 = ~n7873 & ~n7877;
  assign n7879 = ~po1399 & ~n7878;
  assign n7880 = pi3105 & n7108;
  assign n7881 = pi0116 & ~n7108;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = po1399 & ~n7882;
  assign po0267 = n7879 | n7883;
  assign n7885 = pi0062 & n7498;
  assign n7886 = pi0062 & ~n7537;
  assign n7887 = ~pi0062 & n7537;
  assign n7888 = ~n7886 & ~n7887;
  assign n7889 = ~n7498 & ~n7888;
  assign n7890 = ~n7885 & ~n7889;
  assign n7891 = ~po1399 & ~n7890;
  assign n7892 = pi3068 & n7108;
  assign n7893 = pi0117 & ~n7108;
  assign n7894 = ~n7892 & ~n7893;
  assign n7895 = po1399 & ~n7894;
  assign po0268 = n7891 | n7895;
  assign n7897 = pi0063 & n7498;
  assign n7898 = pi0063 & ~n7562;
  assign n7899 = ~pi0063 & n7562;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = ~n7498 & ~n7900;
  assign n7902 = ~n7897 & ~n7901;
  assign n7903 = ~po1399 & ~n7902;
  assign n7904 = pi3075 & n7108;
  assign n7905 = pi0118 & ~n7108;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = po1399 & ~n7906;
  assign po0269 = n7903 | n7907;
  assign n7909 = pi0064 & n7498;
  assign n7910 = pi0064 & ~n7628;
  assign n7911 = ~pi0064 & n7628;
  assign n7912 = ~n7910 & ~n7911;
  assign n7913 = ~n7498 & ~n7912;
  assign n7914 = ~n7909 & ~n7913;
  assign n7915 = ~po1399 & ~n7914;
  assign n7916 = pi3046 & n7108;
  assign n7917 = pi0119 & ~n7108;
  assign n7918 = ~n7916 & ~n7917;
  assign n7919 = po1399 & ~n7918;
  assign po0270 = n7915 | n7919;
  assign n7921 = pi0065 & n7498;
  assign n7922 = ~pi0065 & ~n7498;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = ~po1399 & ~n7923;
  assign n7925 = pi3026 & n7108;
  assign n7926 = pi0106 & ~n7108;
  assign n7927 = ~n7925 & ~n7926;
  assign n7928 = po1399 & ~n7927;
  assign po0271 = n7924 | n7928;
  assign n7930 = pi0066 & n7498;
  assign n7931 = pi0066 & ~n7835;
  assign n7932 = ~pi0066 & n7835;
  assign n7933 = ~n7931 & ~n7932;
  assign n7934 = ~n7498 & ~n7933;
  assign n7935 = ~n7930 & ~n7934;
  assign n7936 = ~po1399 & ~n7935;
  assign n7937 = pi3114 & n7108;
  assign n7938 = pi0123 & ~n7108;
  assign n7939 = ~n7937 & ~n7938;
  assign n7940 = po1399 & ~n7939;
  assign po0272 = n7936 | n7940;
  assign n7942 = pi0067 & n7498;
  assign n7943 = pi0067 & ~n7606;
  assign n7944 = ~pi0067 & n7606;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = ~n7498 & ~n7945;
  assign n7947 = ~n7942 & ~n7946;
  assign n7948 = ~po1399 & ~n7947;
  assign n7949 = pi3073 & n7108;
  assign n7950 = pi0122 & ~n7108;
  assign n7951 = ~n7949 & ~n7950;
  assign n7952 = po1399 & ~n7951;
  assign po0273 = n7948 | n7952;
  assign n7954 = pi0068 & n7498;
  assign n7955 = pi0068 & ~n7604;
  assign n7956 = ~pi0068 & n7604;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = ~n7498 & ~n7957;
  assign n7959 = ~n7954 & ~n7958;
  assign n7960 = ~po1399 & ~n7959;
  assign n7961 = pi3037 & n7108;
  assign n7962 = pi0124 & ~n7108;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = po1399 & ~n7963;
  assign po0274 = n7960 | n7964;
  assign n7966 = pi0069 & ~po1399;
  assign n7967 = ~pi3112 & pi3115;
  assign n7968 = ~pi3102 & po1399;
  assign n7969 = n7108 & n7968;
  assign n7970 = n7967 & n7969;
  assign n7971 = ~n7108 & po1399;
  assign n7972 = pi0089 & n7971;
  assign n7973 = ~n7970 & ~n7972;
  assign po0275 = n7966 | ~n7973;
  assign n7975 = pi0070 & ~po1399;
  assign n7976 = pi3066 & ~pi3112;
  assign n7977 = n7969 & n7976;
  assign n7978 = pi0095 & n7971;
  assign n7979 = ~n7977 & ~n7978;
  assign po0276 = n7975 | ~n7979;
  assign n7981 = ~pi0129 & ~pi3377;
  assign n7982 = pi0129 & pi0223;
  assign n7983 = ~n7981 & ~n7982;
  assign po0277 = ~pi0380 & ~n7983;
  assign n7985 = ~pi0072 & ~po1399;
  assign n7986 = pi0109 & po1399;
  assign po0278 = n7985 | n7986;
  assign n7988 = ~pi0073 & ~po1399;
  assign n7989 = pi0110 & po1399;
  assign po0279 = n7988 | n7989;
  assign n7991 = ~pi0074 & ~po1399;
  assign n7992 = pi0111 & po1399;
  assign po0280 = n7991 | n7992;
  assign n7994 = ~pi0075 & ~po1399;
  assign n7995 = pi0112 & po1399;
  assign po0281 = n7994 | n7995;
  assign n7997 = pi0310 & pi3218;
  assign n7998 = ~pi0310 & ~pi3218;
  assign n7999 = ~n7997 & ~n7998;
  assign n8000 = pi0266 & pi3217;
  assign n8001 = ~pi0266 & ~pi3217;
  assign n8002 = ~n8000 & ~n8001;
  assign n8003 = n7999 & n8002;
  assign n8004 = pi0076 & n7082;
  assign n8005 = ~pi3364 & n8004;
  assign n8006 = pi0113 & ~n8005;
  assign po0282 = ~n8003 & ~n8006;
  assign n8008 = ~pi1973 & ~pi3117;
  assign n8009 = pi3130 & n8008;
  assign n8010 = pi2972 & pi3020;
  assign n8011 = pi3109 & n8010;
  assign n8012 = pi3057 & n8011;
  assign n8013 = pi2980 & n8012;
  assign n8014 = pi2993 & ~pi3024;
  assign n8015 = ~pi3025 & n8014;
  assign n8016 = ~n8013 & n8015;
  assign n8017 = ~n8009 & n8016;
  assign n8018 = ~pi2980 & ~pi3109;
  assign n8019 = pi3018 & pi3057;
  assign n8020 = n8010 & n8019;
  assign n8021 = pi2972 & ~n8020;
  assign n8022 = n8018 & ~n8021;
  assign n8023 = n8017 & ~n8022;
  assign n8024 = pi2980 & ~pi3109;
  assign n8025 = ~pi2980 & pi3109;
  assign n8026 = ~n8024 & ~n8025;
  assign n8027 = ~pi3020 & pi3057;
  assign n8028 = pi2972 & n8027;
  assign n8029 = ~n8020 & ~n8028;
  assign n8030 = ~pi3109 & n8029;
  assign n8031 = pi2972 & ~pi3057;
  assign n8032 = pi3109 & ~n8031;
  assign n8033 = ~n8020 & n8032;
  assign n8034 = ~n8030 & ~n8033;
  assign n8035 = ~n8026 & n8034;
  assign n8036 = n8023 & ~n8035;
  assign n8037 = pi2984 & ~n8036;
  assign n8038 = ~pi2969 & ~pi2984;
  assign n8039 = ~n8036 & n8038;
  assign n8040 = pi1335 & ~pi2553;
  assign n8041 = n8039 & n8040;
  assign n8042 = ~n8037 & ~n8041;
  assign n8043 = ~pi1160 & ~pi1161;
  assign n8044 = pi1159 & n8043;
  assign n8045 = ~pi1159 & pi1160;
  assign n8046 = ~pi1161 & n8045;
  assign n8047 = ~pi1214 & ~pi3193;
  assign n8048 = pi1215 & pi3220;
  assign n8049 = ~n8047 & ~n8048;
  assign n8050 = ~pi1215 & ~pi3220;
  assign n8051 = pi1222 & pi3204;
  assign n8052 = ~n8050 & ~n8051;
  assign n8053 = ~pi1222 & ~pi3204;
  assign n8054 = pi1214 & pi3193;
  assign n8055 = ~n8053 & ~n8054;
  assign n8056 = n8052 & n8055;
  assign n8057 = n8049 & n8056;
  assign n8058 = pi0476 & ~n8057;
  assign n8059 = n7252 & ~n8057;
  assign n8060 = n8058 & n8059;
  assign n8061 = pi0360 & ~n8059;
  assign n8062 = ~n8060 & ~n8061;
  assign n8063 = n7250 & ~n8062;
  assign n8064 = pi1261 & pi2553;
  assign n8065 = n8039 & n8064;
  assign n8066 = ~n8063 & n8065;
  assign n8067 = pi1331 & pi2969;
  assign n8068 = ~pi2984 & n8067;
  assign n8069 = ~n8036 & n8068;
  assign n8070 = ~n8066 & ~n8069;
  assign n8071 = n8046 & n8070;
  assign n8072 = ~n8044 & n8071;
  assign n8073 = n8042 & n8072;
  assign n8074 = ~pi1159 & ~pi1160;
  assign n8075 = pi1161 & n8074;
  assign n8076 = ~pi1973 & pi3370;
  assign n8077 = pi1232 & pi1973;
  assign n8078 = ~n8076 & ~n8077;
  assign n8079 = pi2969 & ~pi3117;
  assign n8080 = ~pi2914 & ~pi3205;
  assign n8081 = pi2914 & pi3205;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = ~pi2921 & ~pi3199;
  assign n8084 = pi2921 & pi3199;
  assign n8085 = ~n8083 & ~n8084;
  assign n8086 = ~n8082 & ~n8085;
  assign n8087 = pi2940 & ~pi3208;
  assign n8088 = ~pi2940 & pi3208;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = n8086 & n8089;
  assign n8091 = pi2937 & pi2969;
  assign po3257 = pi0077 & n8075;
  assign n8093 = ~pi3129 & n7252;
  assign n8094 = ~po3257 & n8093;
  assign n8095 = ~pi2984 & n8094;
  assign n8096 = ~pi2984 & n8046;
  assign n8097 = ~n8036 & n8096;
  assign n8098 = ~n8095 & ~n8097;
  assign n8099 = n8091 & ~n8098;
  assign n8100 = ~pi1335 & n8099;
  assign n8101 = pi2969 & ~pi2984;
  assign n8102 = pi3083 & ~po3257;
  assign n8103 = pi3207 & ~n8102;
  assign n8104 = pi2937 & ~pi3120;
  assign n8105 = ~pi1335 & n8104;
  assign n8106 = n8103 & n8105;
  assign n8107 = n8101 & n8106;
  assign po1484 = n8100 | n8107;
  assign n8109 = ~pi2951 & ~pi3199;
  assign n8110 = pi2951 & pi3199;
  assign n8111 = ~n8109 & ~n8110;
  assign n8112 = pi2916 & ~pi3205;
  assign n8113 = ~pi2916 & pi3205;
  assign n8114 = ~n8112 & ~n8113;
  assign n8115 = ~n8111 & n8114;
  assign n8116 = pi2942 & ~pi3208;
  assign n8117 = ~pi2942 & pi3208;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = n8115 & n8118;
  assign n8120 = po1484 & n8119;
  assign n8121 = ~pi2956 & ~pi3205;
  assign n8122 = pi2956 & pi3205;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = ~pi2954 & ~pi3199;
  assign n8125 = pi2954 & pi3199;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = ~n8123 & ~n8126;
  assign n8128 = pi2934 & ~pi3208;
  assign n8129 = ~pi2934 & pi3208;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = n8127 & n8130;
  assign n8132 = ~pi2935 & ~pi3205;
  assign n8133 = pi2935 & pi3205;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = ~pi2945 & ~pi3199;
  assign n8136 = pi2945 & pi3199;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = ~n8134 & ~n8137;
  assign n8139 = ~pi2936 & pi3208;
  assign n8140 = pi2936 & ~pi3208;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = n8138 & n8141;
  assign n8143 = ~n8131 & ~n8142;
  assign n8144 = ~n8120 & n8143;
  assign n8145 = ~n8090 & n8144;
  assign n8146 = ~pi0484 & n8145;
  assign n8147 = ~pi3024 & ~pi3025;
  assign n8148 = n8018 & ~n8147;
  assign n8149 = n8146 & n8148;
  assign n8150 = n8079 & ~n8149;
  assign n8151 = pi1271 & pi3025;
  assign n8152 = ~pi3024 & ~n8151;
  assign n8153 = n8018 & ~n8152;
  assign n8154 = ~n8057 & n8153;
  assign n8155 = ~n8147 & n8154;
  assign n8156 = ~pi2969 & ~pi3117;
  assign n8157 = ~n8155 & n8156;
  assign n8158 = ~n7250 & n8075;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = ~n8150 & n8159;
  assign n8161 = ~n8063 & n8160;
  assign n8162 = ~pi2969 & n8161;
  assign n8163 = ~n8036 & n8162;
  assign n8164 = n8078 & ~n8163;
  assign n8165 = n8075 & n8164;
  assign n8166 = pi2969 & n8160;
  assign n8167 = n8165 & ~n8166;
  assign n8168 = ~pi3227 & pi3371;
  assign n8169 = pi3121 & pi3227;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = n8167 & n8170;
  assign n8172 = ~pi0077 & ~n8171;
  assign n8173 = ~n8044 & ~n8172;
  assign po0283 = n8073 | n8173;
  assign n8175 = pi0483 & ~pi2960;
  assign n8176 = pi3514 & pi3516;
  assign n8177 = pi3515 & n8176;
  assign n8178 = pi3362 & ~n8177;
  assign n8179 = pi2465 & n8178;
  assign n8180 = ~pi0988 & ~pi1312;
  assign n8181 = ~pi1210 & n8180;
  assign n8182 = ~n8179 & ~n8181;
  assign n8183 = n8175 & ~n8182;
  assign n8184 = pi0483 & pi2960;
  assign n8185 = pi0509 & n8184;
  assign n8186 = ~n8183 & ~n8185;
  assign n8187 = n8175 & ~n8186;
  assign n8188 = n8184 & ~n8186;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = ~pi1798 & ~pi1806;
  assign n8191 = ~pi1967 & n8190;
  assign n8192 = ~pi1923 & ~pi1968;
  assign n8193 = n8191 & n8192;
  assign n8194 = ~n8189 & ~n8193;
  assign n8195 = ~pi0358 & ~pi0359;
  assign n8196 = pi0079 & pi1811;
  assign n8197 = ~pi0082 & n8196;
  assign n8198 = ~pi1969 & n8197;
  assign n8199 = ~n8188 & n8198;
  assign n8200 = pi0483 & pi2465;
  assign n8201 = pi1762 & n8200;
  assign n8202 = n8199 & ~n8201;
  assign n8203 = pi1682 & pi1684;
  assign n8204 = n8187 & ~n8203;
  assign n8205 = ~pi1678 & n8188;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = n8202 & n8206;
  assign n8208 = ~n8195 & n8207;
  assign n8209 = n8194 & n8208;
  assign n8210 = pi1178 & ~pi3219;
  assign n8211 = ~pi1178 & pi3219;
  assign n8212 = ~n8210 & ~n8211;
  assign n8213 = pi1165 & ~pi3216;
  assign n8214 = ~pi1165 & pi3216;
  assign n8215 = ~n8213 & ~n8214;
  assign n8216 = ~n8212 & ~n8215;
  assign n8217 = pi1163 & ~pi3180;
  assign n8218 = ~pi1163 & pi3180;
  assign n8219 = ~n8217 & ~n8218;
  assign n8220 = pi1164 & ~pi3222;
  assign n8221 = ~pi1164 & pi3222;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = ~n8219 & ~n8222;
  assign n8224 = n8216 & n8223;
  assign n8225 = n8195 & ~n8224;
  assign n8226 = n8187 & ~n8225;
  assign n8227 = n8200 & ~n8226;
  assign n8228 = pi0082 & ~pi1811;
  assign n8229 = pi0079 & n8228;
  assign n8230 = ~n8227 & n8229;
  assign n8231 = ~n8209 & ~n8230;
  assign n8232 = pi1318 & n8231;
  assign n8233 = pi0078 & n8232;
  assign po0284 = ~pi3187 & ~n8233;
  assign n8235 = ~pi0079 & ~pi1811;
  assign n8236 = pi3149 & ~n8189;
  assign n8237 = ~pi0082 & n8236;
  assign n8238 = n8235 & n8237;
  assign n8239 = n8227 & n8229;
  assign n8240 = pi1969 & n8187;
  assign n8241 = ~n8188 & n8240;
  assign n8242 = n8195 & n8206;
  assign n8243 = ~pi1969 & ~n8188;
  assign n8244 = n8194 & n8243;
  assign n8245 = ~n8201 & n8244;
  assign n8246 = n8242 & n8245;
  assign n8247 = ~n8241 & ~n8246;
  assign n8248 = n8197 & ~n8247;
  assign n8249 = ~n8239 & ~n8248;
  assign po0285 = n8238 | ~n8249;
  assign n8251 = ~pi0080 & n7183;
  assign n8252 = n7179 & ~n8251;
  assign n8253 = ~pi0080 & n7189;
  assign n8254 = n7228 & ~n8253;
  assign n8255 = ~n7179 & ~n7228;
  assign n8256 = ~n8254 & ~n8255;
  assign po0286 = n8252 | ~n8256;
  assign n8258 = pi0078 & pi3230;
  assign n8259 = ~pi0078 & pi0081;
  assign n8260 = ~n8258 & ~n8259;
  assign po0287 = n8232 & ~n8260;
  assign n8262 = ~pi1170 & ~pi3192;
  assign n8263 = pi1170 & pi3192;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = ~pi1169 & ~pi3198;
  assign n8266 = pi1169 & pi3198;
  assign n8267 = ~n8265 & ~n8266;
  assign n8268 = ~pi1168 & ~pi3194;
  assign n8269 = pi1168 & pi3194;
  assign n8270 = ~n8268 & ~n8269;
  assign n8271 = ~pi1171 & ~pi3209;
  assign n8272 = pi1171 & pi3209;
  assign n8273 = ~n8271 & ~n8272;
  assign n8274 = ~n8270 & ~n8273;
  assign n8275 = ~n8267 & n8274;
  assign n8276 = ~n8264 & n8275;
  assign n8277 = n8188 & n8276;
  assign n8278 = n8200 & ~n8277;
  assign n8279 = ~pi1175 & ~pi3209;
  assign n8280 = pi1175 & pi3209;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 = ~pi1172 & ~pi3192;
  assign n8283 = pi1172 & pi3192;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = ~n8281 & ~n8284;
  assign n8286 = ~pi1166 & ~pi3198;
  assign n8287 = pi1166 & pi3198;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = ~pi1153 & ~pi3194;
  assign n8290 = pi1153 & pi3194;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = ~n8288 & ~n8291;
  assign n8293 = n8285 & n8292;
  assign n8294 = n8188 & n8293;
  assign n8295 = n8278 & ~n8294;
  assign n8296 = pi0082 & n8235;
  assign n8297 = n8295 & n8296;
  assign n8298 = n8188 & n8206;
  assign n8299 = ~n8242 & ~n8298;
  assign n8300 = ~pi1969 & ~n8201;
  assign n8301 = n8197 & n8300;
  assign n8302 = n8194 & n8301;
  assign n8303 = ~n8299 & n8302;
  assign n8304 = pi1969 & ~n8189;
  assign n8305 = n8197 & n8304;
  assign n8306 = ~n8239 & ~n8305;
  assign n8307 = ~n8303 & n8306;
  assign po0288 = n8297 | ~n8307;
  assign n8309 = ~n7060 & ~n7207;
  assign n8310 = ~pi0312 & n8309;
  assign n8311 = ~pi0338 & ~n8309;
  assign po0539 = n8310 | n8311;
  assign n8313 = ~pi0267 & n8309;
  assign n8314 = ~pi0335 & ~n8309;
  assign po0536 = n8313 | n8314;
  assign n8316 = ~pi0311 & n8309;
  assign n8317 = ~pi0337 & ~n8309;
  assign po0538 = n8316 | n8317;
  assign n8319 = po0536 & ~po0538;
  assign n8320 = ~po0539 & n8319;
  assign n8321 = ~pi1890 & n8320;
  assign n8322 = ~po0539 & ~po0536;
  assign n8323 = ~po0538 & n8322;
  assign n8324 = ~pi1904 & n8323;
  assign n8325 = ~n8321 & ~n8324;
  assign n8326 = po0539 & po0538;
  assign n8327 = ~po0536 & n8326;
  assign n8328 = ~pi2163 & n8327;
  assign n8329 = po0536 & po0538;
  assign n8330 = po0539 & n8329;
  assign n8331 = ~pi2157 & n8330;
  assign n8332 = ~n8328 & ~n8331;
  assign n8333 = n8325 & n8332;
  assign n8334 = ~po0536 & po0538;
  assign n8335 = ~po0539 & n8334;
  assign n8336 = ~pi1883 & n8335;
  assign n8337 = ~po0539 & n8329;
  assign n8338 = ~pi1901 & n8337;
  assign n8339 = ~n8336 & ~n8338;
  assign n8340 = po0539 & ~po0536;
  assign n8341 = ~po0538 & n8340;
  assign n8342 = ~pi2164 & n8341;
  assign n8343 = po0539 & po0536;
  assign n8344 = ~po0538 & n8343;
  assign n8345 = ~pi2158 & n8344;
  assign n8346 = ~n8342 & ~n8345;
  assign n8347 = n8339 & n8346;
  assign po0289 = ~n8333 | ~n8347;
  assign n8349 = ~pi2691 & n8323;
  assign n8350 = ~pi2692 & n8320;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = ~pi2690 & n8341;
  assign n8353 = ~pi2689 & n8344;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = n8351 & n8354;
  assign n8356 = ~pi2836 & n8337;
  assign n8357 = ~pi2824 & n8335;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = ~pi2905 & n8327;
  assign n8360 = ~pi2857 & n8330;
  assign n8361 = ~n8359 & ~n8360;
  assign n8362 = n8358 & n8361;
  assign po0290 = ~n8355 | ~n8362;
  assign n8364 = ~pi2926 & n8337;
  assign n8365 = ~pi2929 & n8335;
  assign n8366 = ~n8364 & ~n8365;
  assign n8367 = ~pi2932 & n8327;
  assign n8368 = ~pi2928 & n8330;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = n8366 & n8369;
  assign n8371 = ~pi2933 & n8341;
  assign n8372 = ~pi2931 & n8344;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~pi2930 & n8323;
  assign n8375 = ~pi2927 & n8320;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = n8373 & n8376;
  assign po0291 = ~n8370 | ~n8377;
  assign n8379 = ~pi2844 & n8337;
  assign n8380 = ~pi2673 & n8335;
  assign n8381 = ~n8379 & ~n8380;
  assign n8382 = ~pi2638 & n8327;
  assign n8383 = ~pi2829 & n8330;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~pi2741 & n8323;
  assign n8386 = ~pi2802 & n8320;
  assign n8387 = ~n8385 & ~n8386;
  assign n8388 = n8384 & n8387;
  assign n8389 = ~pi2784 & n8341;
  assign n8390 = ~pi2620 & n8344;
  assign n8391 = ~n8389 & ~n8390;
  assign n8392 = n8388 & n8391;
  assign po0292 = ~n8381 | ~n8392;
  assign n8394 = ~pi2680 & n8337;
  assign n8395 = ~pi2745 & n8335;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = ~pi2606 & n8341;
  assign n8398 = ~pi2723 & n8344;
  assign n8399 = ~n8397 & ~n8398;
  assign n8400 = ~pi2597 & n8327;
  assign n8401 = ~pi2860 & n8330;
  assign n8402 = ~n8400 & ~n8401;
  assign n8403 = n8399 & n8402;
  assign n8404 = ~pi2654 & n8323;
  assign n8405 = ~pi2808 & n8320;
  assign n8406 = ~n8404 & ~n8405;
  assign n8407 = n8403 & n8406;
  assign po0293 = ~n8396 | ~n8407;
  assign n8409 = ~pi2701 & n8330;
  assign n8410 = ~pi2596 & n8327;
  assign n8411 = ~n8409 & ~n8410;
  assign n8412 = ~pi2839 & n8337;
  assign n8413 = ~pi2646 & n8335;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = ~pi2739 & n8323;
  assign n8416 = ~pi2809 & n8320;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = n8414 & n8417;
  assign n8419 = ~pi2621 & n8344;
  assign n8420 = ~pi2515 & n8341;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = n8418 & n8421;
  assign po0294 = ~n8411 | ~n8422;
  assign n8424 = ~pi2292 & n8327;
  assign n8425 = ~pi1975 & n8330;
  assign n8426 = ~n8424 & ~n8425;
  assign n8427 = ~pi2289 & n8341;
  assign n8428 = ~pi1974 & n8344;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~pi1980 & n8337;
  assign n8431 = ~pi1979 & n8335;
  assign n8432 = ~n8430 & ~n8431;
  assign n8433 = n8429 & n8432;
  assign n8434 = ~pi1976 & n8323;
  assign n8435 = ~pi1977 & n8320;
  assign n8436 = ~n8434 & ~n8435;
  assign n8437 = n8433 & n8436;
  assign po0295 = ~n8426 | ~n8437;
  assign n8439 = ~pi2695 & n8327;
  assign n8440 = ~pi2881 & n8330;
  assign n8441 = ~n8439 & ~n8440;
  assign n8442 = ~pi2763 & n8337;
  assign n8443 = ~pi2693 & n8335;
  assign n8444 = ~n8442 & ~n8443;
  assign n8445 = ~pi2655 & n8323;
  assign n8446 = ~pi2811 & n8320;
  assign n8447 = ~n8445 & ~n8446;
  assign n8448 = n8444 & n8447;
  assign n8449 = ~pi2724 & n8344;
  assign n8450 = ~pi2607 & n8341;
  assign n8451 = ~n8449 & ~n8450;
  assign n8452 = n8448 & n8451;
  assign po0296 = ~n8441 | ~n8452;
  assign n8454 = ~pi2898 & n8330;
  assign n8455 = ~pi2627 & n8327;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = ~pi2826 & n8337;
  assign n8458 = ~pi2514 & n8335;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = ~pi2490 & n8323;
  assign n8461 = ~pi2665 & n8320;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = n8459 & n8462;
  assign n8464 = ~pi2650 & n8344;
  assign n8465 = ~pi2748 & n8341;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = n8463 & n8466;
  assign po0297 = ~n8456 | ~n8467;
  assign n8469 = ~pi2653 & n8327;
  assign n8470 = ~pi2637 & n8330;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = ~pi2837 & n8337;
  assign n8473 = ~pi2674 & n8335;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = ~pi2726 & n8341;
  assign n8476 = ~pi2702 & n8344;
  assign n8477 = ~n8475 & ~n8476;
  assign n8478 = n8474 & n8477;
  assign n8479 = ~pi2492 & n8323;
  assign n8480 = ~pi2806 & n8320;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = n8478 & n8481;
  assign po0298 = ~n8471 | ~n8482;
  assign n8484 = ~pi2609 & n8341;
  assign n8485 = ~pi2622 & n8344;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = ~pi2900 & n8335;
  assign n8488 = ~pi2815 & n8337;
  assign n8489 = ~n8487 & ~n8488;
  assign n8490 = n8486 & n8489;
  assign n8491 = ~pi2595 & n8327;
  assign n8492 = ~pi2639 & n8330;
  assign n8493 = ~n8491 & ~n8492;
  assign n8494 = ~pi2657 & n8323;
  assign n8495 = ~pi2793 & n8320;
  assign n8496 = ~n8494 & ~n8495;
  assign n8497 = n8493 & n8496;
  assign po0299 = ~n8490 | ~n8497;
  assign n8499 = ~pi2800 & n8320;
  assign n8500 = ~pi2896 & n8330;
  assign n8501 = ~pi2658 & n8323;
  assign n8502 = ~pi2628 & n8327;
  assign n8503 = ~n8501 & ~n8502;
  assign n8504 = ~n8500 & n8503;
  assign n8505 = ~n8499 & n8504;
  assign n8506 = ~pi2697 & n8344;
  assign n8507 = ~pi2727 & n8341;
  assign n8508 = ~pi2676 & n8335;
  assign n8509 = ~pi2813 & n8337;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = ~n8507 & n8510;
  assign n8512 = ~n8506 & n8511;
  assign po0300 = ~n8505 | ~n8512;
  assign n8514 = ~pi2434 & n8337;
  assign n8515 = ~pi2432 & n8335;
  assign n8516 = ~n8514 & ~n8515;
  assign n8517 = ~pi2295 & n8341;
  assign n8518 = ~pi2284 & n8344;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = ~pi2467 & n8327;
  assign n8521 = ~pi2293 & n8330;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = n8519 & n8522;
  assign n8524 = ~pi2436 & n8323;
  assign n8525 = ~pi1978 & n8320;
  assign n8526 = ~n8524 & ~n8525;
  assign n8527 = n8523 & n8526;
  assign po0301 = ~n8516 | ~n8527;
  assign n8529 = ~pi2598 & n8327;
  assign n8530 = ~pi2640 & n8330;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = ~pi2835 & n8337;
  assign n8533 = ~pi2764 & n8335;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = ~pi2481 & n8323;
  assign n8536 = ~pi2666 & n8320;
  assign n8537 = ~n8535 & ~n8536;
  assign n8538 = n8534 & n8537;
  assign n8539 = ~pi2699 & n8344;
  assign n8540 = ~pi2610 & n8341;
  assign n8541 = ~n8539 & ~n8540;
  assign n8542 = n8538 & n8541;
  assign po0302 = ~n8531 | ~n8542;
  assign n8544 = ~pi2497 & n8323;
  assign n8545 = ~pi2799 & n8320;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = ~pi2681 & n8337;
  assign n8548 = ~pi2513 & n8335;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = ~pi2512 & n8327;
  assign n8551 = ~pi2882 & n8330;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = n8549 & n8552;
  assign n8554 = ~pi2652 & n8344;
  assign n8555 = ~pi2644 & n8341;
  assign n8556 = ~n8554 & ~n8555;
  assign n8557 = n8553 & n8556;
  assign po0303 = ~n8546 | ~n8557;
  assign n8559 = ~pi2493 & n8341;
  assign n8560 = ~pi2623 & n8344;
  assign n8561 = ~n8559 & ~n8560;
  assign n8562 = ~pi2756 & n8337;
  assign n8563 = ~pi2510 & n8335;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = ~pi2716 & n8323;
  assign n8566 = ~pi2667 & n8320;
  assign n8567 = ~n8565 & ~n8566;
  assign n8568 = n8564 & n8567;
  assign n8569 = ~pi2629 & n8327;
  assign n8570 = ~pi2641 & n8330;
  assign n8571 = ~n8569 & ~n8570;
  assign n8572 = n8568 & n8571;
  assign po0304 = ~n8561 | ~n8572;
  assign n8574 = ~pi2509 & n8323;
  assign n8575 = ~pi2782 & n8320;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = ~pi2771 & n8337;
  assign n8578 = ~pi2677 & n8335;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = ~pi2611 & n8341;
  assign n8581 = ~pi2651 & n8344;
  assign n8582 = ~n8580 & ~n8581;
  assign n8583 = n8579 & n8582;
  assign n8584 = ~pi2715 & n8327;
  assign n8585 = ~pi2643 & n8330;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = n8583 & n8586;
  assign po0305 = ~n8576 | ~n8587;
  assign n8589 = ~pi2498 & n8323;
  assign n8590 = ~pi2791 & n8320;
  assign n8591 = ~n8589 & ~n8590;
  assign n8592 = ~pi2775 & n8335;
  assign n8593 = ~pi2682 & n8337;
  assign n8594 = ~n8592 & ~n8593;
  assign n8595 = ~pi2600 & n8327;
  assign n8596 = ~pi2880 & n8330;
  assign n8597 = ~n8595 & ~n8596;
  assign n8598 = n8594 & n8597;
  assign n8599 = ~pi2642 & n8341;
  assign n8600 = ~pi2624 & n8344;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = n8598 & n8601;
  assign po0306 = ~n8591 | ~n8602;
  assign n8604 = ~pi2645 & n8330;
  assign n8605 = ~pi2696 & n8327;
  assign n8606 = ~n8604 & ~n8605;
  assign n8607 = ~pi2814 & n8337;
  assign n8608 = ~pi2876 & n8335;
  assign n8609 = ~n8607 & ~n8608;
  assign n8610 = ~pi2612 & n8341;
  assign n8611 = ~pi2781 & n8344;
  assign n8612 = ~n8610 & ~n8611;
  assign n8613 = n8609 & n8612;
  assign n8614 = ~pi2484 & n8323;
  assign n8615 = ~pi2788 & n8320;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = n8613 & n8616;
  assign po0307 = ~n8606 | ~n8617;
  assign n8619 = ~pi2776 & n8323;
  assign n8620 = ~pi2773 & n8320;
  assign n8621 = ~n8619 & ~n8620;
  assign n8622 = ~pi2630 & n8341;
  assign n8623 = ~pi2780 & n8344;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = ~pi2517 & n8327;
  assign n8626 = ~pi2827 & n8330;
  assign n8627 = ~n8625 & ~n8626;
  assign n8628 = ~pi2688 & n8337;
  assign n8629 = ~pi2883 & n8335;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 = n8627 & n8630;
  assign n8632 = n8624 & n8631;
  assign po0308 = ~n8621 | ~n8632;
  assign n8634 = ~pi2683 & n8337;
  assign n8635 = ~pi2890 & n8335;
  assign n8636 = ~n8634 & ~n8635;
  assign n8637 = ~pi2734 & n8341;
  assign n8638 = ~pi2707 & n8344;
  assign n8639 = ~n8637 & ~n8638;
  assign n8640 = ~pi2500 & n8327;
  assign n8641 = ~pi2828 & n8330;
  assign n8642 = ~n8640 & ~n8641;
  assign n8643 = ~pi2659 & n8323;
  assign n8644 = ~pi2668 & n8320;
  assign n8645 = ~n8643 & ~n8644;
  assign n8646 = n8642 & n8645;
  assign n8647 = n8639 & n8646;
  assign po0309 = ~n8636 | ~n8647;
  assign n8649 = ~pi2899 & n8323;
  assign n8650 = ~pi2746 & n8320;
  assign n8651 = ~n8649 & ~n8650;
  assign n8652 = ~pi2700 & n8327;
  assign n8653 = ~pi2892 & n8330;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = ~pi2822 & n8337;
  assign n8656 = ~pi2678 & n8335;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = n8654 & n8657;
  assign n8659 = ~pi2613 & n8341;
  assign n8660 = ~pi2825 & n8344;
  assign n8661 = ~n8659 & ~n8660;
  assign n8662 = n8658 & n8661;
  assign po0310 = ~n8651 | ~n8662;
  assign n8664 = ~pi2507 & n8327;
  assign n8665 = ~pi2778 & n8330;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = ~pi2744 & n8337;
  assign n8668 = ~pi2893 & n8335;
  assign n8669 = ~n8667 & ~n8668;
  assign n8670 = ~pi2686 & n8323;
  assign n8671 = ~pi2669 & n8320;
  assign n8672 = ~n8670 & ~n8671;
  assign n8673 = n8669 & n8672;
  assign n8674 = ~pi2735 & n8341;
  assign n8675 = ~pi2605 & n8344;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = n8673 & n8676;
  assign po0311 = ~n8666 | ~n8677;
  assign n8679 = ~pi2731 & n8341;
  assign n8680 = ~pi2879 & n8344;
  assign n8681 = ~n8679 & ~n8680;
  assign n8682 = ~pi2684 & n8337;
  assign n8683 = ~pi2902 & n8335;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = ~pi2660 & n8323;
  assign n8686 = ~pi2769 & n8320;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = n8684 & n8687;
  assign n8689 = ~pi2631 & n8327;
  assign n8690 = ~pi2786 & n8330;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = n8688 & n8691;
  assign po0312 = ~n8681 | ~n8692;
  assign n8694 = ~pi2891 & n8323;
  assign n8695 = ~pi2770 & n8320;
  assign n8696 = ~n8694 & ~n8695;
  assign n8697 = ~pi2615 & n8341;
  assign n8698 = ~pi2886 & n8344;
  assign n8699 = ~n8697 & ~n8698;
  assign n8700 = ~pi2816 & n8337;
  assign n8701 = ~pi2887 & n8335;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = n8699 & n8702;
  assign n8704 = ~pi2495 & n8327;
  assign n8705 = ~pi2721 & n8330;
  assign n8706 = ~n8704 & ~n8705;
  assign n8707 = n8703 & n8706;
  assign po0313 = ~n8696 | ~n8707;
  assign n8709 = ~pi2732 & n8341;
  assign n8710 = ~pi2625 & n8344;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = ~pi2794 & n8337;
  assign n8713 = ~pi2754 & n8335;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = ~pi2878 & n8327;
  assign n8716 = ~pi2785 & n8330;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = n8714 & n8717;
  assign n8719 = ~pi2777 & n8323;
  assign n8720 = ~pi2751 & n8320;
  assign n8721 = ~n8719 & ~n8720;
  assign n8722 = n8718 & n8721;
  assign po0314 = ~n8711 | ~n8722;
  assign n8724 = ~pi1881 & n8323;
  assign n8725 = ~pi1882 & n8320;
  assign n8726 = ~n8724 & ~n8725;
  assign n8727 = ~pi1884 & n8337;
  assign n8728 = ~pi1903 & n8335;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = ~pi1880 & n8341;
  assign n8731 = ~pi1879 & n8344;
  assign n8732 = ~n8730 & ~n8731;
  assign n8733 = n8729 & n8732;
  assign n8734 = ~pi1857 & n8327;
  assign n8735 = ~pi1856 & n8330;
  assign n8736 = ~n8734 & ~n8735;
  assign n8737 = n8733 & n8736;
  assign po0315 = ~n8726 | ~n8737;
  assign n8739 = ~pi2633 & n8327;
  assign n8740 = ~pi2730 & n8330;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = ~pi2801 & n8337;
  assign n8743 = ~pi2877 & n8335;
  assign n8744 = ~n8742 & ~n8743;
  assign n8745 = ~pi2796 & n8323;
  assign n8746 = ~pi2670 & n8320;
  assign n8747 = ~n8745 & ~n8746;
  assign n8748 = n8744 & n8747;
  assign n8749 = ~pi2603 & n8344;
  assign n8750 = ~pi2706 & n8341;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = n8748 & n8751;
  assign po0316 = ~n8741 | ~n8752;
  assign n8754 = ~pi2616 & n8341;
  assign n8755 = ~pi2602 & n8344;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = ~pi2807 & n8337;
  assign n8758 = ~pi2810 & n8335;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = ~pi2820 & n8323;
  assign n8761 = ~pi2759 & n8320;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = n8759 & n8762;
  assign n8764 = ~pi2632 & n8327;
  assign n8765 = ~pi2647 & n8330;
  assign n8766 = ~n8764 & ~n8765;
  assign n8767 = n8763 & n8766;
  assign po0317 = ~n8756 | ~n8767;
  assign n8769 = ~pi2687 & n8337;
  assign n8770 = ~pi2821 & n8335;
  assign n8771 = ~n8769 & ~n8770;
  assign n8772 = ~pi2709 & n8327;
  assign n8773 = ~pi2897 & n8330;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = ~pi2617 & n8341;
  assign n8776 = ~pi2516 & n8344;
  assign n8777 = ~n8775 & ~n8776;
  assign n8778 = n8774 & n8777;
  assign n8779 = ~pi2823 & n8323;
  assign n8780 = ~pi2753 & n8320;
  assign n8781 = ~n8779 & ~n8780;
  assign n8782 = n8778 & n8781;
  assign po0318 = ~n8771 | ~n8782;
  assign n8784 = ~pi1688 & n8341;
  assign n8785 = ~pi1749 & n8344;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = ~pi1689 & n8327;
  assign n8788 = ~pi1748 & n8330;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = ~pi1690 & n8323;
  assign n8791 = ~pi1747 & n8320;
  assign n8792 = ~n8790 & ~n8791;
  assign n8793 = n8789 & n8792;
  assign n8794 = ~pi1691 & n8337;
  assign n8795 = ~pi1746 & n8335;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = n8793 & n8796;
  assign po0319 = ~n8786 | ~n8797;
  assign n8799 = ~pi2729 & n8341;
  assign n8800 = ~pi2713 & n8344;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~pi2875 & n8335;
  assign n8803 = ~pi2804 & n8337;
  assign n8804 = ~n8802 & ~n8803;
  assign n8805 = n8801 & n8804;
  assign n8806 = ~pi2601 & n8327;
  assign n8807 = ~pi2903 & n8330;
  assign n8808 = ~n8806 & ~n8807;
  assign n8809 = ~pi2661 & n8323;
  assign n8810 = ~pi2740 & n8320;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = n8808 & n8811;
  assign po0320 = ~n8805 | ~n8812;
  assign n8814 = ~pi2662 & n8323;
  assign n8815 = ~pi2743 & n8320;
  assign n8816 = ~n8814 & ~n8815;
  assign n8817 = ~pi2750 & n8335;
  assign n8818 = ~pi2772 & n8337;
  assign n8819 = ~n8817 & ~n8818;
  assign n8820 = ~pi2494 & n8327;
  assign n8821 = ~pi2491 & n8330;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = n8819 & n8822;
  assign n8824 = ~pi2728 & n8341;
  assign n8825 = ~pi2717 & n8344;
  assign n8826 = ~n8824 & ~n8825;
  assign n8827 = n8823 & n8826;
  assign po0321 = ~n8816 | ~n8827;
  assign n8829 = ~pi2783 & n8337;
  assign n8830 = ~pi2855 & n8335;
  assign n8831 = ~n8829 & ~n8830;
  assign n8832 = ~pi2618 & n8341;
  assign n8833 = ~pi2710 & n8344;
  assign n8834 = ~n8832 & ~n8833;
  assign n8835 = ~pi2634 & n8327;
  assign n8836 = ~pi2648 & n8330;
  assign n8837 = ~n8835 & ~n8836;
  assign n8838 = n8834 & n8837;
  assign n8839 = ~pi2817 & n8323;
  assign n8840 = ~pi2747 & n8320;
  assign n8841 = ~n8839 & ~n8840;
  assign n8842 = n8838 & n8841;
  assign po0322 = ~n8831 | ~n8842;
  assign n8844 = ~pi2790 & n8337;
  assign n8845 = ~pi2768 & n8335;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = ~pi2719 & n8327;
  assign n8848 = ~pi2708 & n8330;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~pi2712 & n8341;
  assign n8851 = ~pi2711 & n8344;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = n8849 & n8852;
  assign n8854 = ~pi2663 & n8323;
  assign n8855 = ~pi2671 & n8320;
  assign n8856 = ~n8854 & ~n8855;
  assign n8857 = n8853 & n8856;
  assign po0323 = ~n8846 | ~n8857;
  assign n8859 = ~pi2792 & n8337;
  assign n8860 = ~pi2679 & n8335;
  assign n8861 = ~n8859 & ~n8860;
  assign n8862 = ~pi2831 & n8341;
  assign n8863 = ~pi2626 & n8344;
  assign n8864 = ~n8862 & ~n8863;
  assign n8865 = ~pi2722 & n8327;
  assign n8866 = ~pi2714 & n8330;
  assign n8867 = ~n8865 & ~n8866;
  assign n8868 = n8864 & n8867;
  assign n8869 = ~pi2812 & n8323;
  assign n8870 = ~pi2672 & n8320;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = n8868 & n8871;
  assign po0324 = ~n8861 | ~n8872;
  assign n8874 = ~pi2718 & n8341;
  assign n8875 = ~pi2725 & n8344;
  assign n8876 = ~n8874 & ~n8875;
  assign n8877 = ~pi2675 & n8335;
  assign n8878 = ~pi2789 & n8337;
  assign n8879 = ~n8877 & ~n8878;
  assign n8880 = n8876 & n8879;
  assign n8881 = ~pi2636 & n8327;
  assign n8882 = ~pi2703 & n8330;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = ~pi2797 & n8323;
  assign n8885 = ~pi2487 & n8320;
  assign n8886 = ~n8884 & ~n8885;
  assign n8887 = n8883 & n8886;
  assign po0325 = ~n8880 | ~n8887;
  assign n8889 = ~pi1335 & ~pi2969;
  assign po3302 = ~pi0077 & n8075;
  assign n8891 = ~pi2984 & po3302;
  assign n8892 = n8078 & n8891;
  assign n8893 = n8889 & n8892;
  assign n8894 = n8161 & n8893;
  assign n8895 = pi1261 & n8096;
  assign n8896 = pi2553 & ~pi2969;
  assign n8897 = ~n8036 & ~n8063;
  assign n8898 = n8896 & n8897;
  assign n8899 = n8895 & n8898;
  assign n8900 = ~pi2553 & ~pi2969;
  assign n8901 = n8097 & n8900;
  assign n8902 = pi1335 & n8901;
  assign n8903 = ~pi1335 & pi2969;
  assign n8904 = n8078 & n8160;
  assign n8905 = n8891 & n8904;
  assign n8906 = n8903 & n8905;
  assign n8907 = n8037 & n8046;
  assign n8908 = n8067 & n8097;
  assign n8909 = ~n8907 & ~n8908;
  assign n8910 = ~n8906 & n8909;
  assign n8911 = ~n8902 & n8910;
  assign n8912 = ~n8899 & n8911;
  assign n8913 = ~pi1335 & ~n8147;
  assign n8914 = ~pi2969 & n8063;
  assign n8915 = ~pi2969 & n8153;
  assign n8916 = pi2969 & n8018;
  assign n8917 = ~n8915 & ~n8916;
  assign n8918 = ~n8914 & ~n8917;
  assign n8919 = n8913 & n8918;
  assign n8920 = n8078 & n8919;
  assign n8921 = pi3120 & n8920;
  assign n8922 = n8891 & n8921;
  assign n8923 = n8912 & ~n8922;
  assign n8924 = ~n8894 & n8923;
  assign n8925 = pi0120 & n8078;
  assign n8926 = ~n8170 & n8925;
  assign po0326 = n8924 & ~n8926;
  assign n8928 = ~pi2656 & n8323;
  assign n8929 = ~pi2805 & n8320;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = ~pi2604 & n8330;
  assign n8932 = ~pi2698 & n8327;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = ~pi2803 & n8337;
  assign n8935 = ~pi2504 & n8335;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~pi2720 & n8344;
  assign n8938 = ~pi2608 & n8341;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = n8936 & n8939;
  assign n8941 = n8933 & n8940;
  assign po0327 = ~n8930 | ~n8941;
  assign n8943 = ~pi2685 & n8323;
  assign n8944 = ~pi2798 & n8320;
  assign n8945 = ~n8943 & ~n8944;
  assign n8946 = ~pi2704 & n8330;
  assign n8947 = ~pi2511 & n8327;
  assign n8948 = ~n8946 & ~n8947;
  assign n8949 = ~pi2832 & n8337;
  assign n8950 = ~pi2833 & n8335;
  assign n8951 = ~n8949 & ~n8950;
  assign n8952 = ~pi2694 & n8344;
  assign n8953 = ~pi2614 & n8341;
  assign n8954 = ~n8952 & ~n8953;
  assign n8955 = n8951 & n8954;
  assign n8956 = n8948 & n8955;
  assign po0328 = ~n8945 | ~n8956;
  assign n8958 = ~pi2664 & n8323;
  assign n8959 = ~pi2742 & n8320;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = ~pi2649 & n8330;
  assign n8962 = ~pi2635 & n8327;
  assign n8963 = ~n8961 & ~n8962;
  assign n8964 = ~pi2774 & n8337;
  assign n8965 = ~pi2830 & n8335;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = ~pi2599 & n8344;
  assign n8968 = ~pi2619 & n8341;
  assign n8969 = ~n8967 & ~n8968;
  assign n8970 = n8966 & n8969;
  assign n8971 = n8963 & n8970;
  assign po0329 = ~n8960 | ~n8971;
  assign n8973 = n8038 & n8046;
  assign n8974 = pi2553 & n8973;
  assign n8975 = ~pi1261 & n8974;
  assign n8976 = n8063 & n8895;
  assign n8977 = n8896 & n8976;
  assign n8978 = pi0126 & po3257;
  assign n8979 = n8078 & n8978;
  assign n8980 = pi2969 & n8096;
  assign n8981 = ~pi1331 & n8980;
  assign n8982 = n8036 & n8046;
  assign n8983 = ~n8981 & ~n8982;
  assign n8984 = ~pi2553 & n8889;
  assign n8985 = n8096 & n8984;
  assign n8986 = n8983 & ~n8985;
  assign n8987 = ~n8979 & n8986;
  assign n8988 = ~n8977 & n8987;
  assign n8989 = ~n8975 & n8988;
  assign n8990 = ~pi2969 & po3302;
  assign n8991 = n8063 & n8990;
  assign n8992 = ~n8160 & po3302;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = n8078 & n8170;
  assign n8995 = ~n8993 & n8994;
  assign po0330 = n8989 & ~n8995;
  assign n8997 = ~pi3136 & ~pi3163;
  assign n8998 = pi3161 & n8027;
  assign n8999 = pi3018 & n8998;
  assign n9000 = n8997 & n8999;
  assign n9001 = n8009 & n9000;
  assign n9002 = pi1722 & pi3133;
  assign n9003 = ~pi1722 & ~pi3133;
  assign n9004 = ~n9002 & ~n9003;
  assign n9005 = ~pi1713 & ~pi3134;
  assign n9006 = pi1713 & pi3134;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = ~pi1718 & ~pi3171;
  assign n9009 = pi1718 & pi3171;
  assign n9010 = ~n9008 & ~n9009;
  assign n9011 = ~n9007 & ~n9010;
  assign n9012 = ~pi1716 & ~pi3164;
  assign n9013 = pi1716 & pi3164;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~pi1711 & ~pi3132;
  assign n9016 = pi1711 & pi3132;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = ~n9014 & ~n9017;
  assign n9019 = ~pi1707 & ~pi3147;
  assign n9020 = pi1707 & pi3147;
  assign n9021 = ~n9019 & ~n9020;
  assign n9022 = ~pi1668 & ~pi3141;
  assign n9023 = pi1668 & pi3141;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = ~n9021 & ~n9024;
  assign n9026 = ~pi1717 & ~pi3153;
  assign n9027 = pi1717 & pi3153;
  assign n9028 = ~n9026 & ~n9027;
  assign n9029 = ~pi1710 & ~pi3143;
  assign n9030 = pi1710 & pi3143;
  assign n9031 = ~n9029 & ~n9030;
  assign n9032 = ~n9028 & ~n9031;
  assign n9033 = n9025 & n9032;
  assign n9034 = n9018 & n9033;
  assign n9035 = n9011 & n9034;
  assign n9036 = ~pi1719 & ~pi3151;
  assign n9037 = pi1719 & pi3151;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = ~pi1752 & ~pi3157;
  assign n9040 = pi1752 & pi3157;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = ~n9038 & ~n9041;
  assign n9043 = ~pi1753 & ~pi3138;
  assign n9044 = pi1753 & pi3138;
  assign n9045 = ~n9043 & ~n9044;
  assign n9046 = ~pi1720 & ~pi3172;
  assign n9047 = pi1720 & pi3172;
  assign n9048 = ~n9046 & ~n9047;
  assign n9049 = ~n9045 & ~n9048;
  assign n9050 = ~pi1715 & ~pi3154;
  assign n9051 = pi1715 & pi3154;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = ~pi1755 & ~pi3165;
  assign n9054 = pi1755 & pi3165;
  assign n9055 = ~n9053 & ~n9054;
  assign n9056 = ~n9052 & ~n9055;
  assign n9057 = ~pi1754 & ~pi3162;
  assign n9058 = pi1754 & pi3162;
  assign n9059 = ~n9057 & ~n9058;
  assign n9060 = ~pi1714 & ~pi3155;
  assign n9061 = pi1714 & pi3155;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~n9059 & ~n9062;
  assign n9064 = n9056 & n9063;
  assign n9065 = n9049 & n9064;
  assign n9066 = n9042 & n9065;
  assign n9067 = pi1723 & ~pi3150;
  assign n9068 = ~pi1723 & pi3150;
  assign n9069 = ~n9067 & ~n9068;
  assign n9070 = ~pi1721 & ~pi3135;
  assign n9071 = pi1721 & pi3135;
  assign n9072 = ~n9070 & ~n9071;
  assign n9073 = n9069 & ~n9072;
  assign n9074 = n9066 & n9073;
  assign n9075 = n9035 & n9074;
  assign n9076 = ~pi1751 & ~pi3158;
  assign n9077 = pi1751 & pi3158;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = n9075 & ~n9078;
  assign n9080 = ~pi3018 & ~pi3057;
  assign n9081 = n9079 & ~n9080;
  assign n9082 = ~n9004 & n9081;
  assign n9083 = pi3020 & n9082;
  assign n9084 = pi3020 & ~pi3057;
  assign n9085 = pi3018 & n9084;
  assign n9086 = pi2972 & n9085;
  assign n9087 = n9083 & ~n9086;
  assign n9088 = pi3160 & n9087;
  assign n9089 = pi1361 & n9088;
  assign n9090 = pi1768 & pi1790;
  assign n9091 = pi1790 & pi3151;
  assign n9092 = n9090 & n9091;
  assign n9093 = ~n9090 & ~n9091;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = pi1770 & pi1810;
  assign n9096 = pi1810 & pi3172;
  assign n9097 = n9095 & n9096;
  assign n9098 = ~n9095 & ~n9096;
  assign n9099 = ~n9097 & ~n9098;
  assign n9100 = pi1793 & pi1797;
  assign n9101 = pi1793 & pi3158;
  assign n9102 = n9100 & ~n9101;
  assign n9103 = ~n9100 & n9101;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = pi1794 & pi3133;
  assign n9106 = pi1772 & pi1794;
  assign n9107 = n9105 & ~n9106;
  assign n9108 = ~n9105 & n9106;
  assign n9109 = ~n9107 & ~n9108;
  assign n9110 = n9104 & n9109;
  assign n9111 = pi1771 & pi1792;
  assign n9112 = pi1792 & pi3150;
  assign n9113 = n9111 & ~n9112;
  assign n9114 = ~n9111 & n9112;
  assign n9115 = ~n9113 & ~n9114;
  assign n9116 = pi1795 & pi1802;
  assign n9117 = pi1795 & pi3135;
  assign n9118 = n9116 & ~n9117;
  assign n9119 = ~n9116 & n9117;
  assign n9120 = ~n9118 & ~n9119;
  assign n9121 = n9115 & n9120;
  assign n9122 = pi1775 & pi1783;
  assign n9123 = pi1783 & pi3143;
  assign n9124 = n9122 & n9123;
  assign n9125 = ~n9122 & ~n9123;
  assign n9126 = ~n9124 & ~n9125;
  assign n9127 = pi1774 & pi1781;
  assign n9128 = pi1781 & pi3141;
  assign n9129 = n9127 & n9128;
  assign n9130 = ~n9127 & ~n9128;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = pi1757 & pi1760;
  assign n9133 = pi1757 & pi3153;
  assign n9134 = n9132 & n9133;
  assign n9135 = ~n9132 & ~n9133;
  assign n9136 = ~n9134 & ~n9135;
  assign n9137 = pi1776 & pi1787;
  assign n9138 = pi1787 & pi3147;
  assign n9139 = n9137 & n9138;
  assign n9140 = ~n9137 & ~n9138;
  assign n9141 = ~n9139 & ~n9140;
  assign n9142 = ~n9136 & ~n9141;
  assign n9143 = ~n9131 & n9142;
  assign n9144 = ~n9126 & n9143;
  assign n9145 = pi1785 & pi1804;
  assign n9146 = pi1785 & pi3132;
  assign n9147 = n9145 & n9146;
  assign n9148 = ~n9145 & ~n9146;
  assign n9149 = ~n9147 & ~n9148;
  assign n9150 = pi1756 & pi1777;
  assign n9151 = pi1756 & pi3134;
  assign n9152 = n9150 & n9151;
  assign n9153 = ~n9150 & ~n9151;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = pi1764 & pi1791;
  assign n9156 = pi1791 & pi3171;
  assign n9157 = n9155 & n9156;
  assign n9158 = ~n9155 & ~n9156;
  assign n9159 = ~n9157 & ~n9158;
  assign n9160 = pi1763 & pi1784;
  assign n9161 = pi1784 & pi3164;
  assign n9162 = n9160 & n9161;
  assign n9163 = ~n9160 & ~n9161;
  assign n9164 = ~n9162 & ~n9163;
  assign n9165 = ~n9159 & ~n9164;
  assign n9166 = ~n9154 & n9165;
  assign n9167 = ~n9149 & n9166;
  assign n9168 = n9144 & n9167;
  assign n9169 = pi1767 & pi1789;
  assign n9170 = pi1789 & pi3154;
  assign n9171 = n9169 & n9170;
  assign n9172 = ~n9169 & ~n9170;
  assign n9173 = ~n9171 & ~n9172;
  assign n9174 = pi1765 & pi1786;
  assign n9175 = pi1786 & pi3155;
  assign n9176 = n9174 & n9175;
  assign n9177 = ~n9174 & ~n9175;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = pi1766 & pi1779;
  assign n9180 = pi1779 & pi3162;
  assign n9181 = n9179 & n9180;
  assign n9182 = ~n9179 & ~n9180;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = pi1788 & pi1801;
  assign n9185 = pi1788 & pi3165;
  assign n9186 = n9184 & n9185;
  assign n9187 = ~n9184 & ~n9185;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = ~n9183 & ~n9188;
  assign n9190 = ~n9178 & n9189;
  assign n9191 = ~n9173 & n9190;
  assign n9192 = pi1800 & pi1809;
  assign n9193 = pi1809 & pi3146;
  assign n9194 = n9192 & n9193;
  assign n9195 = ~n9192 & ~n9193;
  assign n9196 = ~n9194 & ~n9195;
  assign n9197 = pi1799 & pi1808;
  assign n9198 = pi1808 & pi3170;
  assign n9199 = n9197 & n9198;
  assign n9200 = ~n9197 & ~n9198;
  assign n9201 = ~n9199 & ~n9200;
  assign n9202 = pi1759 & pi1782;
  assign n9203 = pi1782 & pi3168;
  assign n9204 = n9202 & n9203;
  assign n9205 = ~n9202 & ~n9203;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = pi1773 & pi1780;
  assign n9208 = pi1780 & pi3139;
  assign n9209 = n9207 & n9208;
  assign n9210 = ~n9207 & ~n9208;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = ~n9206 & ~n9211;
  assign n9213 = ~n9201 & n9212;
  assign n9214 = ~n9196 & n9213;
  assign n9215 = n9191 & n9214;
  assign n9216 = n9168 & n9215;
  assign n9217 = n9121 & n9216;
  assign n9218 = n9110 & n9217;
  assign n9219 = pi1758 & pi1803;
  assign n9220 = pi1758 & pi3138;
  assign n9221 = n9219 & ~n9220;
  assign n9222 = ~n9219 & n9220;
  assign n9223 = ~n9221 & ~n9222;
  assign n9224 = n9218 & n9223;
  assign n9225 = pi1769 & pi1807;
  assign n9226 = pi1807 & pi3157;
  assign n9227 = n9225 & n9226;
  assign n9228 = ~n9225 & ~n9226;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = n9224 & ~n9229;
  assign n9231 = ~n9099 & n9230;
  assign n9232 = ~n9094 & n9231;
  assign n9233 = pi1360 & ~n9086;
  assign n9234 = pi3160 & n9233;
  assign n9235 = pi1793 & n9234;
  assign n9236 = ~pi3018 & n8027;
  assign n9237 = n9235 & n9236;
  assign n9238 = n9232 & n9237;
  assign n9239 = ~n9089 & ~n9238;
  assign n9240 = n8009 & ~n9000;
  assign n9241 = ~n9239 & n9240;
  assign n9242 = ~n9001 & ~n9241;
  assign n9243 = n8063 & n8064;
  assign n9244 = n8038 & n9243;
  assign n9245 = ~n8036 & n8046;
  assign n9246 = ~n9244 & n9245;
  assign n9247 = n9242 & ~n9246;
  assign n9248 = n8063 & ~n8170;
  assign n9249 = n8990 & n9248;
  assign n9250 = n8078 & n9249;
  assign n9251 = pi0128 & po3257;
  assign n9252 = pi2969 & po3302;
  assign n9253 = ~n8063 & n8990;
  assign n9254 = ~n9252 & ~n9253;
  assign n9255 = ~n9251 & n9254;
  assign n9256 = n8078 & ~n9255;
  assign n9257 = ~n9250 & ~n9256;
  assign po0331 = n9247 & n9257;
  assign n9259 = ~pi0411 & ~pi1346;
  assign n9260 = pi0411 & pi3376;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = ~pi3138 & pi3151;
  assign n9263 = pi3138 & ~pi3151;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = ~pi3157 & pi3172;
  assign n9266 = pi3157 & ~pi3172;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = ~n9264 & n9267;
  assign n9269 = n9264 & ~n9267;
  assign n9270 = ~n9268 & ~n9269;
  assign n9271 = pi3154 & ~pi3165;
  assign n9272 = ~pi3154 & pi3165;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = ~pi3155 & pi3162;
  assign n9275 = pi3155 & ~pi3162;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = ~n9273 & n9276;
  assign n9278 = n9273 & ~n9276;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = ~n9270 & n9279;
  assign n9281 = n9270 & ~n9279;
  assign n9282 = ~n9280 & ~n9281;
  assign n9283 = pi3132 & ~pi3134;
  assign n9284 = ~pi3132 & pi3134;
  assign n9285 = ~n9283 & ~n9284;
  assign n9286 = ~pi3164 & pi3171;
  assign n9287 = pi3164 & ~pi3171;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = ~n9285 & n9288;
  assign n9290 = n9285 & ~n9288;
  assign n9291 = ~n9289 & ~n9290;
  assign n9292 = ~pi3141 & pi3143;
  assign n9293 = pi3141 & ~pi3143;
  assign n9294 = ~n9292 & ~n9293;
  assign n9295 = ~pi3147 & pi3153;
  assign n9296 = pi3147 & ~pi3153;
  assign n9297 = ~n9295 & ~n9296;
  assign n9298 = ~n9294 & n9297;
  assign n9299 = n9294 & ~n9297;
  assign n9300 = ~n9298 & ~n9299;
  assign n9301 = ~n9291 & n9300;
  assign n9302 = n9291 & ~n9300;
  assign n9303 = ~n9301 & ~n9302;
  assign n9304 = ~n9282 & n9303;
  assign n9305 = n9282 & ~n9303;
  assign n9306 = ~n9304 & ~n9305;
  assign n9307 = pi3131 & ~pi3159;
  assign n9308 = ~pi3131 & pi3159;
  assign n9309 = ~n9307 & ~n9308;
  assign n9310 = ~pi3145 & pi3169;
  assign n9311 = pi3145 & ~pi3169;
  assign n9312 = ~n9310 & ~n9311;
  assign n9313 = ~n9309 & n9312;
  assign n9314 = n9309 & ~n9312;
  assign n9315 = ~n9313 & ~n9314;
  assign n9316 = pi3146 & ~pi3170;
  assign n9317 = ~pi3146 & pi3170;
  assign n9318 = ~n9316 & ~n9317;
  assign n9319 = ~pi3139 & pi3168;
  assign n9320 = pi3139 & ~pi3168;
  assign n9321 = ~n9319 & ~n9320;
  assign n9322 = ~n9318 & n9321;
  assign n9323 = n9318 & ~n9321;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = ~n9315 & n9324;
  assign n9326 = n9315 & ~n9324;
  assign n9327 = ~n9325 & ~n9326;
  assign n9328 = pi3142 & ~pi3166;
  assign n9329 = ~pi3142 & pi3166;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = ~pi3136 & pi3163;
  assign n9332 = pi3136 & ~pi3163;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = ~n9330 & n9333;
  assign n9335 = n9330 & ~n9333;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = pi3018 & ~pi3020;
  assign n9338 = ~pi3018 & pi3020;
  assign n9339 = ~n9337 & ~n9338;
  assign n9340 = ~pi2972 & pi3057;
  assign n9341 = ~n8031 & ~n9340;
  assign n9342 = ~n9339 & ~n9341;
  assign n9343 = n9339 & n9341;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = pi3133 & ~pi3158;
  assign n9346 = ~pi3133 & pi3158;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = ~pi3135 & pi3150;
  assign n9349 = pi3135 & ~pi3150;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n9347 & n9350;
  assign n9352 = n9347 & ~n9350;
  assign n9353 = ~n9351 & ~n9352;
  assign n9354 = ~n9344 & n9353;
  assign n9355 = n9344 & ~n9353;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = ~n9336 & n9356;
  assign n9358 = n9336 & ~n9356;
  assign n9359 = ~n9357 & ~n9358;
  assign n9360 = ~n9327 & n9359;
  assign n9361 = n9327 & ~n9359;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = ~n9306 & n9362;
  assign n9364 = n9306 & ~n9362;
  assign n9365 = ~n9363 & ~n9364;
  assign n9366 = ~n9261 & n9365;
  assign n9367 = n9261 & ~n9365;
  assign n9368 = ~n9366 & ~n9367;
  assign n9369 = n7257 & n9368;
  assign po0645 = ~pi0877 & pi0896;
  assign n9371 = pi1220 & ~pi3120;
  assign n9372 = ~pi3042 & pi3227;
  assign n9373 = ~n9371 & ~n9372;
  assign n9374 = pi0411 & ~n9373;
  assign n9375 = po0645 & n9374;
  assign po0405 = n9369 & n9375;
  assign po0335 = ~pi0202 & ~po0405;
  assign n9378 = ~pi1696 & ~pi1697;
  assign n9379 = pi1694 & n9378;
  assign n9380 = ~pi1695 & n9379;
  assign n9381 = ~pi1694 & n9378;
  assign n9382 = pi1695 & n9381;
  assign n9383 = pi3117 & pi3120;
  assign n9384 = ~pi3369 & n9383;
  assign n9385 = n9382 & n9384;
  assign n9386 = ~n9380 & ~n9385;
  assign n9387 = ~n8046 & n9386;
  assign n9388 = pi1220 & ~pi2969;
  assign n9389 = ~pi1694 & ~pi1695;
  assign n9390 = pi1696 & n9389;
  assign n9391 = ~pi1697 & n9390;
  assign n9392 = pi0307 & n9391;
  assign n9393 = ~n9388 & ~n9392;
  assign n9394 = ~pi1220 & pi3374;
  assign n9395 = ~pi0120 & pi1220;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = ~n9393 & n9396;
  assign n9398 = n8170 & n9397;
  assign n9399 = n9387 & ~n9398;
  assign n9400 = pi1696 & pi1697;
  assign n9401 = n9389 & ~n9400;
  assign n9402 = ~n9378 & n9401;
  assign n9403 = ~pi3042 & ~pi3118;
  assign n9404 = n9402 & n9403;
  assign n9405 = pi0426 & n9404;
  assign n9406 = ~pi0292 & ~n9404;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 = pi1676 & ~n9407;
  assign n9409 = ~pi1676 & pi1698;
  assign n9410 = ~pi0259 & n9409;
  assign n9411 = ~pi1676 & ~pi1698;
  assign n9412 = pi1667 & n9411;
  assign n9413 = ~n9410 & ~n9412;
  assign n9414 = ~n9408 & n9413;
  assign n9415 = pi0896 & ~n9414;
  assign n9416 = pi2920 & ~pi2982;
  assign n9417 = ~pi2995 & ~pi2997;
  assign n9418 = n9416 & n9417;
  assign n9419 = ~pi2966 & ~pi2996;
  assign n9420 = ~pi2981 & ~pi3001;
  assign n9421 = n9419 & n9420;
  assign n9422 = n9418 & n9421;
  assign n9423 = pi0133 & n9422;
  assign n9424 = pi2995 & ~pi2997;
  assign n9425 = pi2920 & n9424;
  assign n9426 = ~pi2982 & n9419;
  assign n9427 = n9420 & n9426;
  assign n9428 = n9425 & n9427;
  assign n9429 = n9100 & n9428;
  assign n9430 = ~n9423 & ~n9429;
  assign n9431 = pi2981 & ~pi3001;
  assign n9432 = pi2966 & ~pi2996;
  assign n9433 = n9431 & n9432;
  assign n9434 = ~pi2920 & ~pi2982;
  assign n9435 = n9417 & n9434;
  assign n9436 = n9433 & n9435;
  assign n9437 = pi2981 & pi3001;
  assign n9438 = n9432 & n9437;
  assign n9439 = ~pi2920 & pi2982;
  assign n9440 = n9417 & n9439;
  assign n9441 = n9438 & n9440;
  assign n9442 = pi2550 & n9441;
  assign n9443 = ~pi2966 & pi2996;
  assign n9444 = n9431 & n9443;
  assign n9445 = pi2920 & pi2982;
  assign n9446 = n9424 & n9445;
  assign n9447 = n9444 & n9446;
  assign n9448 = pi2555 & n9447;
  assign n9449 = ~n9442 & ~n9448;
  assign n9450 = n9419 & n9431;
  assign n9451 = n9418 & n9450;
  assign n9452 = pi1751 & n9451;
  assign n9453 = n9424 & n9434;
  assign n9454 = n9433 & n9453;
  assign n9455 = pi1793 & n9454;
  assign n9456 = ~n9452 & ~n9455;
  assign n9457 = n9444 & n9453;
  assign n9458 = pi1340 & n9457;
  assign n9459 = pi2966 & pi2996;
  assign n9460 = n9431 & n9459;
  assign n9461 = pi1334 & n9460;
  assign n9462 = n9418 & n9461;
  assign n9463 = ~n9458 & ~n9462;
  assign n9464 = pi1333 & pi1377;
  assign n9465 = n9453 & n9464;
  assign n9466 = ~pi2982 & n9425;
  assign n9467 = pi1333 & n9466;
  assign n9468 = ~n9465 & ~n9467;
  assign n9469 = n9460 & ~n9468;
  assign n9470 = n9463 & ~n9469;
  assign n9471 = n9456 & n9470;
  assign n9472 = n9449 & n9471;
  assign n9473 = n9446 & n9460;
  assign n9474 = pi2503 & n9473;
  assign n9475 = ~pi2982 & n9431;
  assign n9476 = n9432 & n9475;
  assign n9477 = n9425 & n9476;
  assign n9478 = pi1825 & n9477;
  assign n9479 = ~n9474 & ~n9478;
  assign n9480 = n9421 & n9453;
  assign n9481 = pi1751 & n9480;
  assign n9482 = n9479 & ~n9481;
  assign n9483 = n9424 & n9450;
  assign n9484 = n9416 & n9483;
  assign n9485 = n9100 & n9484;
  assign n9486 = n9482 & ~n9485;
  assign n9487 = n9437 & n9443;
  assign n9488 = pi1342 & n9487;
  assign n9489 = pi1334 & pi1378;
  assign n9490 = n9460 & n9489;
  assign n9491 = ~n9488 & ~n9490;
  assign n9492 = n9435 & ~n9491;
  assign n9493 = n9486 & ~n9492;
  assign n9494 = n9472 & n9493;
  assign n9495 = pi3001 & n9419;
  assign n9496 = pi2981 & n9495;
  assign n9497 = n9445 & n9496;
  assign n9498 = n9417 & n9497;
  assign n9499 = pi2537 & n9498;
  assign n9500 = n9419 & n9437;
  assign n9501 = n9440 & n9500;
  assign n9502 = pi2873 & n9501;
  assign n9503 = ~n9499 & ~n9502;
  assign n9504 = n9417 & n9445;
  assign n9505 = n9437 & n9504;
  assign n9506 = n9459 & n9505;
  assign n9507 = pi1677 & n9506;
  assign n9508 = n9424 & n9439;
  assign n9509 = n9460 & n9508;
  assign n9510 = pi2588 & n9509;
  assign n9511 = ~n9507 & ~n9510;
  assign n9512 = n9503 & n9511;
  assign n9513 = n9494 & n9512;
  assign n9514 = ~n9436 & n9513;
  assign n9515 = n9430 & n9514;
  assign n9516 = ~pi0896 & ~n7250;
  assign n9517 = ~n9515 & n9516;
  assign n9518 = ~n9415 & ~n9517;
  assign n9519 = pi0469 & n8059;
  assign n9520 = ~pi0397 & ~n8059;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = ~pi0896 & n7250;
  assign n9523 = ~n9521 & n9522;
  assign n9524 = n9518 & ~n9523;
  assign n9525 = ~n9399 & ~n9524;
  assign n9526 = pi0130 & n9399;
  assign po0333 = n9525 | n9526;
  assign n9528 = pi0131 & n9399;
  assign po0334 = n9525 | n9528;
  assign n9530 = ~pi3018 & pi3158;
  assign n9531 = n7247 & n9530;
  assign n9532 = n7254 & n9531;
  assign n9533 = pi0133 & ~n9532;
  assign n9534 = ~pi0223 & ~n9533;
  assign po0336 = ~pi0224 | ~n9534;
  assign n9536 = ~n8224 & n8229;
  assign po0337 = ~n8227 & n9536;
  assign n9538 = pi0434 & n9404;
  assign n9539 = ~pi0273 & ~n9404;
  assign n9540 = ~n9538 & ~n9539;
  assign n9541 = ~pi1337 & ~n9540;
  assign n9542 = pi0434 & ~pi2486;
  assign n9543 = ~pi1218 & ~pi1262;
  assign n9544 = pi2486 & n9543;
  assign n9545 = ~n9542 & ~n9544;
  assign n9546 = pi1337 & ~n9545;
  assign n9547 = ~n9541 & ~n9546;
  assign n9548 = pi1676 & ~n9547;
  assign n9549 = pi0307 & n9409;
  assign n9550 = ~n9548 & ~n9549;
  assign n9551 = pi0205 & n9411;
  assign n9552 = n9550 & ~n9551;
  assign n9553 = ~n9399 & ~n9552;
  assign n9554 = pi0135 & n9399;
  assign po0338 = n9553 | n9554;
  assign n9556 = pi0436 & n9404;
  assign n9557 = ~pi0332 & ~n9404;
  assign n9558 = ~n9556 & ~n9557;
  assign n9559 = ~pi1337 & ~n9558;
  assign n9560 = pi0436 & ~pi2486;
  assign n9561 = ~pi1218 & ~pi1268;
  assign n9562 = pi2486 & n9561;
  assign n9563 = ~n9560 & ~n9562;
  assign n9564 = pi1337 & ~n9563;
  assign n9565 = ~n9559 & ~n9564;
  assign n9566 = pi1676 & ~n9565;
  assign n9567 = pi0306 & n9409;
  assign n9568 = ~n9566 & ~n9567;
  assign n9569 = pi0207 & n9411;
  assign n9570 = n9568 & ~n9569;
  assign n9571 = ~n9399 & ~n9570;
  assign n9572 = pi0136 & n9399;
  assign po0339 = n9571 | n9572;
  assign n9574 = pi0137 & n9386;
  assign n9575 = ~n9386 & ~n9552;
  assign po0340 = n9574 | n9575;
  assign n9577 = pi0138 & n9386;
  assign n9578 = pi0435 & n9404;
  assign n9579 = ~pi0274 & ~n9404;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = ~pi1337 & ~n9580;
  assign n9582 = pi0435 & ~pi2486;
  assign n9583 = ~pi1218 & ~pi1264;
  assign n9584 = pi2486 & n9583;
  assign n9585 = ~n9582 & ~n9584;
  assign n9586 = pi1337 & ~n9585;
  assign n9587 = ~n9581 & ~n9586;
  assign n9588 = pi1676 & ~n9587;
  assign n9589 = pi0305 & n9409;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = pi0206 & n9411;
  assign n9592 = n9590 & ~n9591;
  assign n9593 = ~n9386 & ~n9592;
  assign po0341 = n9577 | n9593;
  assign n9595 = ~n9399 & ~n9592;
  assign n9596 = pi0139 & n9399;
  assign po0342 = n9595 | n9596;
  assign n9598 = pi0140 & n9386;
  assign n9599 = ~n9386 & ~n9570;
  assign po0343 = n9598 | n9599;
  assign n9601 = pi0141 & n9399;
  assign n9602 = pi1717 & n9451;
  assign n9603 = pi1757 & n9454;
  assign n9604 = ~n9602 & ~n9603;
  assign n9605 = pi2530 & n9498;
  assign n9606 = n9420 & n9432;
  assign n9607 = n9418 & n9606;
  assign n9608 = pi1705 & n9607;
  assign n9609 = ~n9605 & ~n9608;
  assign n9610 = n9132 & n9484;
  assign n9611 = pi2544 & n9441;
  assign n9612 = ~n9610 & ~n9611;
  assign n9613 = pi1717 & n9480;
  assign n9614 = pi2560 & n9473;
  assign n9615 = ~n9613 & ~n9614;
  assign n9616 = n9612 & n9615;
  assign n9617 = pi1847 & n9477;
  assign n9618 = n9616 & ~n9617;
  assign n9619 = n9609 & n9618;
  assign n9620 = n9604 & n9619;
  assign n9621 = ~n9436 & n9620;
  assign n9622 = pi2489 & n9509;
  assign n9623 = n9132 & n9428;
  assign n9624 = ~n9622 & ~n9623;
  assign n9625 = n9621 & n9624;
  assign n9626 = ~n7250 & ~n9625;
  assign n9627 = pi0450 & n8059;
  assign n9628 = ~pi0377 & ~n8059;
  assign n9629 = ~n9627 & ~n9628;
  assign n9630 = n7250 & ~n9629;
  assign n9631 = ~n9626 & ~n9630;
  assign n9632 = ~pi0896 & ~n9631;
  assign n9633 = pi0412 & n9404;
  assign n9634 = ~pi0281 & ~n9404;
  assign n9635 = ~n9633 & ~n9634;
  assign n9636 = pi1676 & ~n9635;
  assign n9637 = pi0299 & n9409;
  assign n9638 = pi1730 & n9411;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = ~n9636 & n9639;
  assign n9641 = pi0896 & ~n9640;
  assign n9642 = ~n9632 & ~n9641;
  assign n9643 = ~n9399 & ~n9642;
  assign po0344 = n9601 | n9643;
  assign n9645 = pi0142 & n9399;
  assign n9646 = pi0460 & n8059;
  assign n9647 = ~pi0406 & ~n8059;
  assign n9648 = ~n9646 & ~n9647;
  assign n9649 = n7250 & ~n9648;
  assign n9650 = ~n9451 & ~n9480;
  assign n9651 = pi1715 & ~n9650;
  assign n9652 = pi1822 & n9477;
  assign n9653 = pi1789 & n9454;
  assign n9654 = ~n9652 & ~n9653;
  assign n9655 = pi2779 & n9441;
  assign n9656 = pi2567 & n9473;
  assign n9657 = ~n9655 & ~n9656;
  assign n9658 = n9169 & n9484;
  assign n9659 = n9657 & ~n9658;
  assign n9660 = n9435 & n9606;
  assign n9661 = n9659 & ~n9660;
  assign n9662 = n9654 & n9661;
  assign n9663 = ~n9651 & n9662;
  assign n9664 = pi2865 & n9498;
  assign n9665 = pi2889 & n9509;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = n9169 & n9428;
  assign n9668 = ~n9436 & ~n9667;
  assign n9669 = n9666 & n9668;
  assign n9670 = ~n9422 & n9669;
  assign n9671 = n9663 & n9670;
  assign n9672 = ~n7250 & ~n9671;
  assign n9673 = ~n9649 & ~n9672;
  assign n9674 = ~pi0896 & ~n9673;
  assign n9675 = pi0420 & n9404;
  assign n9676 = ~pi0330 & ~n9404;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = pi1676 & ~n9677;
  assign n9679 = pi0254 & n9409;
  assign n9680 = pi1665 & n9411;
  assign n9681 = ~n9679 & ~n9680;
  assign n9682 = ~n9678 & n9681;
  assign n9683 = pi0896 & ~n9682;
  assign n9684 = ~n9674 & ~n9683;
  assign n9685 = ~n9399 & ~n9684;
  assign po0345 = n9645 | n9685;
  assign n9687 = pi0143 & n9399;
  assign n9688 = pi0461 & n8059;
  assign n9689 = ~pi0392 & ~n8059;
  assign n9690 = ~n9688 & ~n9689;
  assign n9691 = n7250 & ~n9690;
  assign n9692 = pi2795 & n9441;
  assign n9693 = pi2736 & n9447;
  assign n9694 = ~n9692 & ~n9693;
  assign n9695 = pi0002 & n9422;
  assign n9696 = n9219 & n9428;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = pi2866 & n9498;
  assign n9699 = pi2846 & n9501;
  assign n9700 = ~n9698 & ~n9699;
  assign n9701 = pi2584 & n9509;
  assign n9702 = n9700 & ~n9701;
  assign n9703 = n9697 & n9702;
  assign n9704 = ~n9436 & n9703;
  assign n9705 = n9694 & n9704;
  assign n9706 = pi1821 & n9477;
  assign n9707 = pi1758 & n9454;
  assign n9708 = ~n9706 & ~n9707;
  assign n9709 = pi2508 & n9473;
  assign n9710 = n9219 & n9484;
  assign n9711 = ~n9709 & ~n9710;
  assign n9712 = pi1753 & ~n9650;
  assign n9713 = n9711 & ~n9712;
  assign n9714 = n9708 & n9713;
  assign n9715 = n9705 & n9714;
  assign n9716 = ~n7250 & ~n9715;
  assign n9717 = ~n9691 & ~n9716;
  assign n9718 = ~pi0896 & ~n9717;
  assign n9719 = pi0421 & n9404;
  assign n9720 = ~pi0287 & ~n9404;
  assign n9721 = ~n9719 & ~n9720;
  assign n9722 = pi1676 & ~n9721;
  assign n9723 = pi0255 & n9409;
  assign n9724 = pi1736 & n9411;
  assign n9725 = ~n9723 & ~n9724;
  assign n9726 = ~n9722 & n9725;
  assign n9727 = pi0896 & ~n9726;
  assign n9728 = ~n9718 & ~n9727;
  assign n9729 = ~n9399 & ~n9728;
  assign po0346 = n9687 | n9729;
  assign n9731 = pi0144 & n9399;
  assign n9732 = pi0464 & n8059;
  assign n9733 = ~pi0405 & ~n8059;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = n7250 & ~n9734;
  assign n9736 = pi2819 & n9441;
  assign n9737 = pi2737 & n9447;
  assign n9738 = ~n9736 & ~n9737;
  assign n9739 = pi3001 & n9432;
  assign n9740 = ~pi2981 & n9739;
  assign n9741 = n9466 & n9740;
  assign n9742 = ~n9436 & ~n9741;
  assign n9743 = pi1368 & n9422;
  assign n9744 = n9095 & n9428;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = pi2861 & n9498;
  assign n9747 = pi2852 & n9501;
  assign n9748 = ~n9746 & ~n9747;
  assign n9749 = pi2904 & n9509;
  assign n9750 = n9748 & ~n9749;
  assign n9751 = n9745 & n9750;
  assign n9752 = n9742 & n9751;
  assign n9753 = n9738 & n9752;
  assign n9754 = pi1851 & n9477;
  assign n9755 = pi1810 & n9454;
  assign n9756 = ~n9754 & ~n9755;
  assign n9757 = pi2506 & n9473;
  assign n9758 = n9095 & n9484;
  assign n9759 = ~n9757 & ~n9758;
  assign n9760 = pi1720 & ~n9650;
  assign n9761 = n9759 & ~n9760;
  assign n9762 = n9756 & n9761;
  assign n9763 = n9753 & n9762;
  assign n9764 = ~n7250 & ~n9763;
  assign n9765 = ~n9735 & ~n9764;
  assign n9766 = ~pi0896 & ~n9765;
  assign n9767 = pi0422 & n9404;
  assign n9768 = ~pi0288 & ~n9404;
  assign n9769 = ~n9767 & ~n9768;
  assign n9770 = pi1676 & ~n9769;
  assign n9771 = pi0256 & n9409;
  assign n9772 = pi1669 & n9411;
  assign n9773 = ~n9771 & ~n9772;
  assign n9774 = ~n9770 & n9773;
  assign n9775 = pi0896 & ~n9774;
  assign n9776 = ~n9766 & ~n9775;
  assign n9777 = ~n9399 & ~n9776;
  assign po0347 = n9731 | n9777;
  assign n9779 = pi0145 & n9399;
  assign n9780 = pi0465 & n8059;
  assign n9781 = ~pi0394 & ~n8059;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = n7250 & ~n9782;
  assign n9784 = pi2535 & n9498;
  assign n9785 = pi2523 & n9501;
  assign n9786 = ~n9784 & ~n9785;
  assign n9787 = pi2586 & n9509;
  assign n9788 = n9786 & ~n9787;
  assign n9789 = pi2485 & n9441;
  assign n9790 = pi2488 & n9447;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = pi1370 & n9422;
  assign n9793 = n9116 & n9428;
  assign n9794 = ~n9792 & ~n9793;
  assign n9795 = n9791 & n9794;
  assign n9796 = n9742 & n9795;
  assign n9797 = n9788 & n9796;
  assign n9798 = pi1824 & n9477;
  assign n9799 = pi1795 & n9454;
  assign n9800 = ~n9798 & ~n9799;
  assign n9801 = pi2505 & n9473;
  assign n9802 = n9116 & n9484;
  assign n9803 = ~n9801 & ~n9802;
  assign n9804 = pi1721 & ~n9650;
  assign n9805 = n9803 & ~n9804;
  assign n9806 = n9800 & n9805;
  assign n9807 = n9797 & n9806;
  assign n9808 = ~n7250 & ~n9807;
  assign n9809 = ~n9783 & ~n9808;
  assign n9810 = ~pi0896 & ~n9809;
  assign n9811 = pi0423 & n9404;
  assign n9812 = ~pi0289 & ~n9404;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = pi1676 & ~n9813;
  assign n9815 = pi0257 & n9409;
  assign n9816 = pi1739 & n9411;
  assign n9817 = ~n9815 & ~n9816;
  assign n9818 = ~n9814 & n9817;
  assign n9819 = pi0896 & ~n9818;
  assign n9820 = ~n9810 & ~n9819;
  assign n9821 = ~n9399 & ~n9820;
  assign po0348 = n9779 | n9821;
  assign n9823 = pi0146 & n9399;
  assign n9824 = pi0466 & n8059;
  assign n9825 = ~pi0395 & ~n8059;
  assign n9826 = ~n9824 & ~n9825;
  assign n9827 = n7250 & ~n9826;
  assign n9828 = pi2549 & n9441;
  assign n9829 = pi2705 & n9447;
  assign n9830 = ~n9828 & ~n9829;
  assign n9831 = pi1372 & n9422;
  assign n9832 = n9111 & n9428;
  assign n9833 = ~n9831 & ~n9832;
  assign n9834 = pi2862 & n9498;
  assign n9835 = pi2524 & n9501;
  assign n9836 = ~n9834 & ~n9835;
  assign n9837 = pi2895 & n9509;
  assign n9838 = n9836 & ~n9837;
  assign n9839 = n9833 & n9838;
  assign n9840 = ~n9436 & n9839;
  assign n9841 = n9830 & n9840;
  assign n9842 = pi1814 & n9477;
  assign n9843 = pi1792 & n9454;
  assign n9844 = ~n9842 & ~n9843;
  assign n9845 = pi2570 & n9473;
  assign n9846 = n9111 & n9484;
  assign n9847 = ~n9845 & ~n9846;
  assign n9848 = pi1723 & ~n9650;
  assign n9849 = n9847 & ~n9848;
  assign n9850 = n9844 & n9849;
  assign n9851 = n9841 & n9850;
  assign n9852 = ~n7250 & ~n9851;
  assign n9853 = ~n9827 & ~n9852;
  assign n9854 = ~pi0896 & ~n9853;
  assign n9855 = pi0424 & n9404;
  assign n9856 = ~pi0290 & ~n9404;
  assign n9857 = ~n9855 & ~n9856;
  assign n9858 = pi1676 & ~n9857;
  assign n9859 = pi0258 & n9409;
  assign n9860 = pi1740 & n9411;
  assign n9861 = ~n9859 & ~n9860;
  assign n9862 = ~n9858 & n9861;
  assign n9863 = pi0896 & ~n9862;
  assign n9864 = ~n9854 & ~n9863;
  assign n9865 = ~n9399 & ~n9864;
  assign po0349 = n9823 | n9865;
  assign n9867 = pi0147 & n9399;
  assign n9868 = pi0467 & n8059;
  assign n9869 = ~pi0396 & ~n8059;
  assign n9870 = ~n9868 & ~n9869;
  assign n9871 = n7250 & ~n9870;
  assign n9872 = n9450 & n9453;
  assign n9873 = pi1339 & n9872;
  assign n9874 = pi2571 & n9473;
  assign n9875 = ~n9873 & ~n9874;
  assign n9876 = n9421 & n9435;
  assign n9877 = n9418 & n9740;
  assign n9878 = ~n9876 & ~n9877;
  assign n9879 = n9875 & n9878;
  assign n9880 = pi2752 & n9441;
  assign n9881 = n9879 & ~n9880;
  assign n9882 = n9444 & n9466;
  assign n9883 = pi1359 & n9882;
  assign n9884 = n9418 & n9444;
  assign n9885 = pi1349 & n9884;
  assign n9886 = ~n9883 & ~n9885;
  assign n9887 = pi2536 & n9498;
  assign n9888 = pi1352 & n9741;
  assign n9889 = ~n9887 & ~n9888;
  assign n9890 = pi1709 & n9607;
  assign n9891 = n9889 & ~n9890;
  assign n9892 = n9886 & n9891;
  assign n9893 = n9881 & n9892;
  assign n9894 = pi1397 & n9506;
  assign n9895 = pi2587 & n9509;
  assign n9896 = ~n9894 & ~n9895;
  assign n9897 = pi1362 & n9422;
  assign n9898 = n9487 & n9508;
  assign n9899 = pi3177 & n9898;
  assign n9900 = ~n9897 & ~n9899;
  assign n9901 = n9896 & n9900;
  assign n9902 = n9893 & n9901;
  assign n9903 = ~n7250 & ~n9902;
  assign n9904 = ~n9871 & ~n9903;
  assign n9905 = ~pi0896 & ~n9904;
  assign n9906 = pi0425 & n9404;
  assign n9907 = ~pi0291 & ~n9404;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = pi1676 & ~n9908;
  assign n9910 = pi0268 & n9409;
  assign n9911 = pi1741 & n9411;
  assign n9912 = ~n9910 & ~n9911;
  assign n9913 = ~n9909 & n9912;
  assign n9914 = pi0896 & ~n9913;
  assign n9915 = ~n9905 & ~n9914;
  assign n9916 = ~n9399 & ~n9915;
  assign po0350 = n9867 | n9916;
  assign n9918 = pi0148 & n9399;
  assign n9919 = pi2853 & n9498;
  assign n9920 = pi1399 & n9741;
  assign n9921 = ~n9919 & ~n9920;
  assign n9922 = pi1400 & n9607;
  assign n9923 = n9921 & ~n9922;
  assign n9924 = pi2551 & n9441;
  assign n9925 = n9923 & ~n9924;
  assign n9926 = pi2572 & n9473;
  assign n9927 = pi2888 & n9509;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = n9925 & n9928;
  assign n9930 = ~n7250 & ~n9929;
  assign n9931 = pi0470 & n8059;
  assign n9932 = ~pi0398 & ~n8059;
  assign n9933 = ~n9931 & ~n9932;
  assign n9934 = n7250 & ~n9933;
  assign n9935 = ~n9930 & ~n9934;
  assign n9936 = ~pi0896 & ~n9935;
  assign n9937 = pi0427 & n9404;
  assign n9938 = ~pi0293 & ~n9404;
  assign n9939 = ~n9937 & ~n9938;
  assign n9940 = pi1676 & ~n9939;
  assign n9941 = pi0301 & n9409;
  assign n9942 = pi1742 & n9411;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = ~n9940 & n9943;
  assign n9945 = pi0896 & ~n9944;
  assign n9946 = ~n9936 & ~n9945;
  assign n9947 = ~n9399 & ~n9946;
  assign po0351 = n9918 | n9947;
  assign n9949 = pi0149 & n9399;
  assign n9950 = pi0428 & n9404;
  assign n9951 = ~pi0294 & ~n9404;
  assign n9952 = ~n9950 & ~n9951;
  assign n9953 = pi1676 & ~n9952;
  assign n9954 = pi0260 & n9409;
  assign n9955 = pi1666 & n9411;
  assign n9956 = ~n9954 & ~n9955;
  assign n9957 = ~n9953 & n9956;
  assign n9958 = pi0896 & ~n9957;
  assign n9959 = pi1402 & n9741;
  assign n9960 = pi1404 & n9607;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = pi2767 & n9441;
  assign n9963 = pi2538 & n9498;
  assign n9964 = ~n9962 & ~n9963;
  assign n9965 = pi2502 & n9473;
  assign n9966 = pi2589 & n9509;
  assign n9967 = ~n9965 & ~n9966;
  assign n9968 = n9964 & n9967;
  assign n9969 = n9878 & n9968;
  assign n9970 = n9961 & n9969;
  assign n9971 = ~n7250 & ~n9970;
  assign n9972 = pi0471 & n8059;
  assign n9973 = ~pi0399 & ~n8059;
  assign n9974 = ~n9972 & ~n9973;
  assign n9975 = n7250 & ~n9974;
  assign n9976 = ~n9971 & ~n9975;
  assign n9977 = ~pi0896 & ~n9976;
  assign n9978 = ~n9958 & ~n9977;
  assign n9979 = ~n9399 & ~n9978;
  assign po0352 = n9949 | n9979;
  assign n9981 = pi0150 & n9399;
  assign n9982 = pi2858 & n9498;
  assign n9983 = pi1401 & n9741;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = pi1403 & n9607;
  assign n9986 = n9984 & ~n9985;
  assign n9987 = pi2765 & n9441;
  assign n9988 = n9986 & ~n9987;
  assign n9989 = pi2573 & n9473;
  assign n9990 = pi2885 & n9509;
  assign n9991 = ~n9989 & ~n9990;
  assign n9992 = n9988 & n9991;
  assign n9993 = ~n7250 & ~n9992;
  assign n9994 = pi0472 & n8059;
  assign n9995 = ~pi0403 & ~n8059;
  assign n9996 = ~n9994 & ~n9995;
  assign n9997 = n7250 & ~n9996;
  assign n9998 = ~n9993 & ~n9997;
  assign n9999 = ~pi0896 & ~n9998;
  assign n10000 = pi0429 & n9404;
  assign n10001 = ~pi0327 & ~n9404;
  assign n10002 = ~n10000 & ~n10001;
  assign n10003 = pi1676 & ~n10002;
  assign n10004 = pi0248 & n9409;
  assign n10005 = pi1662 & n9411;
  assign n10006 = ~n10004 & ~n10005;
  assign n10007 = ~n10003 & n10006;
  assign n10008 = pi0896 & ~n10007;
  assign n10009 = ~n9999 & ~n10008;
  assign n10010 = ~n9399 & ~n10009;
  assign po0353 = n9981 | n10010;
  assign n10012 = pi0151 & n9399;
  assign n10013 = pi2496 & n9473;
  assign n10014 = pi1379 & n9422;
  assign n10015 = ~n10013 & ~n10014;
  assign n10016 = pi2766 & n9441;
  assign n10017 = pi2590 & n9509;
  assign n10018 = ~n10016 & ~n10017;
  assign n10019 = n10015 & n10018;
  assign n10020 = pi1712 & n9607;
  assign n10021 = n10019 & ~n10020;
  assign n10022 = pi2539 & n9498;
  assign n10023 = pi1350 & n9741;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n10021 & n10024;
  assign n10026 = ~n7250 & ~n10025;
  assign n10027 = pi0473 & n8059;
  assign n10028 = ~pi0400 & ~n8059;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = n7250 & ~n10029;
  assign n10031 = ~n10026 & ~n10030;
  assign n10032 = ~pi0896 & ~n10031;
  assign n10033 = pi0430 & n9404;
  assign n10034 = ~pi0295 & ~n9404;
  assign n10035 = ~n10033 & ~n10034;
  assign n10036 = pi1676 & ~n10035;
  assign n10037 = pi0261 & n9409;
  assign n10038 = pi1743 & n9411;
  assign n10039 = ~n10037 & ~n10038;
  assign n10040 = ~n10036 & n10039;
  assign n10041 = pi0896 & ~n10040;
  assign n10042 = ~n10032 & ~n10041;
  assign n10043 = ~n9399 & ~n10042;
  assign po0354 = n10012 | n10043;
  assign n10045 = pi0152 & n9399;
  assign n10046 = pi0431 & n9404;
  assign n10047 = ~pi0296 & ~n9404;
  assign n10048 = ~n10046 & ~n10047;
  assign n10049 = pi1676 & ~n10048;
  assign n10050 = pi0262 & n9409;
  assign n10051 = pi1663 & n9411;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = ~n10049 & n10052;
  assign n10054 = pi0896 & ~n10053;
  assign n10055 = pi1595 & n9741;
  assign n10056 = pi1589 & n9607;
  assign n10057 = ~n10055 & ~n10056;
  assign n10058 = pi2552 & n9441;
  assign n10059 = pi2834 & n9498;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = pi2575 & n9473;
  assign n10062 = pi2591 & n9509;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = n10060 & n10063;
  assign n10065 = n9878 & n10064;
  assign n10066 = n10057 & n10065;
  assign n10067 = ~n7250 & ~n10066;
  assign n10068 = pi0451 & n8059;
  assign n10069 = ~pi0379 & ~n8059;
  assign n10070 = ~n10068 & ~n10069;
  assign n10071 = n7250 & ~n10070;
  assign n10072 = ~n10067 & ~n10071;
  assign n10073 = ~pi0896 & ~n10072;
  assign n10074 = ~n10054 & ~n10073;
  assign n10075 = ~n9399 & ~n10074;
  assign po0355 = n10045 | n10075;
  assign n10077 = pi0153 & n9399;
  assign n10078 = pi0474 & n8059;
  assign n10079 = ~pi0401 & ~n8059;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = n7250 & ~n10080;
  assign n10082 = pi2499 & n9473;
  assign n10083 = n9197 & n9484;
  assign n10084 = ~n10082 & ~n10083;
  assign n10085 = pi2540 & n9498;
  assign n10086 = pi1699 & n9607;
  assign n10087 = ~n10085 & ~n10086;
  assign n10088 = pi2760 & n9441;
  assign n10089 = pi1366 & n9447;
  assign n10090 = pi1808 & n9454;
  assign n10091 = ~n10089 & ~n10090;
  assign n10092 = ~n10088 & n10091;
  assign n10093 = pi1849 & n9477;
  assign n10094 = n10092 & ~n10093;
  assign n10095 = n10087 & n10094;
  assign n10096 = n10084 & n10095;
  assign n10097 = pi2592 & n9509;
  assign n10098 = n9197 & n9428;
  assign n10099 = ~n10097 & ~n10098;
  assign n10100 = pi3176 & n9501;
  assign n10101 = pi1365 & n9422;
  assign n10102 = ~n10100 & ~n10101;
  assign n10103 = n10099 & n10102;
  assign n10104 = ~n9741 & n10103;
  assign n10105 = n10096 & n10104;
  assign n10106 = ~n7250 & ~n10105;
  assign n10107 = ~n10081 & ~n10106;
  assign n10108 = ~pi0896 & ~n10107;
  assign n10109 = pi0432 & n9404;
  assign n10110 = ~pi0297 & ~n9404;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = pi1676 & ~n10111;
  assign n10113 = pi0302 & n9409;
  assign n10114 = pi1664 & n9411;
  assign n10115 = ~n10113 & ~n10114;
  assign n10116 = ~n10112 & n10115;
  assign n10117 = pi0896 & ~n10116;
  assign n10118 = ~n10108 & ~n10117;
  assign n10119 = ~n9399 & ~n10118;
  assign po0356 = n10077 | n10119;
  assign n10121 = pi0154 & n9399;
  assign n10122 = pi2542 & n9441;
  assign n10123 = pi1845 & n9477;
  assign n10124 = ~n10122 & ~n10123;
  assign n10125 = pi1782 & n9454;
  assign n10126 = pi2557 & n9473;
  assign n10127 = n9202 & n9484;
  assign n10128 = ~n10126 & ~n10127;
  assign n10129 = n9878 & n10128;
  assign n10130 = ~n10125 & n10129;
  assign n10131 = n10124 & n10130;
  assign n10132 = pi2479 & n9509;
  assign n10133 = n9202 & n9428;
  assign n10134 = ~n10132 & ~n10133;
  assign n10135 = n10131 & n10134;
  assign n10136 = pi2528 & n9498;
  assign n10137 = pi1701 & n9607;
  assign n10138 = ~n10136 & ~n10137;
  assign n10139 = n10135 & n10138;
  assign n10140 = ~n7250 & ~n10139;
  assign n10141 = pi0479 & n8059;
  assign n10142 = ~pi0383 & ~n8059;
  assign n10143 = ~n10141 & ~n10142;
  assign n10144 = n7250 & ~n10143;
  assign n10145 = ~n10140 & ~n10144;
  assign n10146 = ~pi0896 & ~n10145;
  assign n10147 = pi0439 & n9404;
  assign n10148 = ~pi0277 & ~n9404;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = pi1676 & ~n10149;
  assign n10151 = pi0325 & n9409;
  assign n10152 = pi1728 & n9411;
  assign n10153 = ~n10151 & ~n10152;
  assign n10154 = ~n10150 & n10153;
  assign n10155 = pi0896 & ~n10154;
  assign n10156 = ~n10146 & ~n10155;
  assign n10157 = ~n9399 & ~n10156;
  assign po0357 = n10121 | n10157;
  assign n10159 = pi0155 & n9399;
  assign n10160 = pi1668 & ~n9650;
  assign n10161 = pi1848 & n9477;
  assign n10162 = pi1781 & n9454;
  assign n10163 = ~n10161 & ~n10162;
  assign n10164 = pi2529 & n9498;
  assign n10165 = pi1702 & n9607;
  assign n10166 = ~n10164 & ~n10165;
  assign n10167 = pi2558 & n9473;
  assign n10168 = n9127 & n9484;
  assign n10169 = pi2850 & n9441;
  assign n10170 = ~n10168 & ~n10169;
  assign n10171 = ~n10167 & n10170;
  assign n10172 = n9878 & n10171;
  assign n10173 = n10166 & n10172;
  assign n10174 = n10163 & n10173;
  assign n10175 = ~n10160 & n10174;
  assign n10176 = ~n9436 & n10175;
  assign n10177 = pi2577 & n9509;
  assign n10178 = n9127 & n9428;
  assign n10179 = ~n10177 & ~n10178;
  assign n10180 = n10176 & n10179;
  assign n10181 = ~n7250 & ~n10180;
  assign n10182 = pi0480 & n8059;
  assign n10183 = ~pi0407 & ~n8059;
  assign n10184 = ~n10182 & ~n10183;
  assign n10185 = n7250 & ~n10184;
  assign n10186 = ~n10181 & ~n10185;
  assign n10187 = ~pi0896 & ~n10186;
  assign n10188 = pi0440 & n9404;
  assign n10189 = ~pi0278 & ~n9404;
  assign n10190 = ~n10188 & ~n10189;
  assign n10191 = pi1676 & ~n10190;
  assign n10192 = pi0304 & n9409;
  assign n10193 = pi1671 & n9411;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = ~n10191 & n10194;
  assign n10196 = pi0896 & ~n10195;
  assign n10197 = ~n10187 & ~n10196;
  assign n10198 = ~n9399 & ~n10197;
  assign po0358 = n10159 | n10198;
  assign n10200 = pi0156 & n9399;
  assign n10201 = pi1710 & n9451;
  assign n10202 = pi1783 & n9454;
  assign n10203 = ~n10201 & ~n10202;
  assign n10204 = pi2868 & n9498;
  assign n10205 = pi1703 & n9607;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = pi2543 & n9441;
  assign n10208 = pi1846 & n9477;
  assign n10209 = ~n10207 & ~n10208;
  assign n10210 = pi2733 & n9473;
  assign n10211 = n9122 & n9484;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = n10209 & n10212;
  assign n10214 = pi1710 & n9480;
  assign n10215 = n10213 & ~n10214;
  assign n10216 = n10206 & n10215;
  assign n10217 = n10203 & n10216;
  assign n10218 = ~n9436 & n10217;
  assign n10219 = pi2578 & n9509;
  assign n10220 = n9122 & n9428;
  assign n10221 = ~n10219 & ~n10220;
  assign n10222 = n10218 & n10221;
  assign n10223 = ~n7250 & ~n10222;
  assign n10224 = pi0481 & n8059;
  assign n10225 = ~pi0384 & ~n8059;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = n7250 & ~n10226;
  assign n10228 = ~n10223 & ~n10227;
  assign n10229 = ~pi0896 & ~n10228;
  assign n10230 = pi0441 & n9404;
  assign n10231 = ~pi0279 & ~n9404;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = pi1676 & ~n10232;
  assign n10234 = pi0298 & n9409;
  assign n10235 = pi1729 & n9411;
  assign n10236 = ~n10234 & ~n10235;
  assign n10237 = ~n10233 & n10236;
  assign n10238 = pi0896 & ~n10237;
  assign n10239 = ~n10229 & ~n10238;
  assign n10240 = ~n9399 & ~n10239;
  assign po0359 = n10200 | n10240;
  assign n10242 = pi0157 & n9399;
  assign n10243 = pi1707 & n9451;
  assign n10244 = pi1787 & n9454;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = pi2845 & n9441;
  assign n10247 = pi1707 & n9480;
  assign n10248 = pi2559 & n9473;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = n9137 & n9484;
  assign n10251 = n10249 & ~n10250;
  assign n10252 = ~n10246 & n10251;
  assign n10253 = pi1826 & n9477;
  assign n10254 = n10252 & ~n10253;
  assign n10255 = pi2871 & n9498;
  assign n10256 = pi1704 & n9607;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = n10254 & n10257;
  assign n10259 = n10245 & n10258;
  assign n10260 = ~n9436 & n10259;
  assign n10261 = pi2579 & n9509;
  assign n10262 = n9137 & n9428;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = n10260 & n10263;
  assign n10265 = ~n7250 & ~n10264;
  assign n10266 = pi0482 & n8059;
  assign n10267 = ~pi0385 & ~n8059;
  assign n10268 = ~n10266 & ~n10267;
  assign n10269 = n7250 & ~n10268;
  assign n10270 = ~n10265 & ~n10269;
  assign n10271 = ~pi0896 & ~n10270;
  assign n10272 = pi0442 & n9404;
  assign n10273 = ~pi0280 & ~n9404;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = pi1676 & ~n10274;
  assign n10276 = pi0249 & n9409;
  assign n10277 = pi1674 & n9411;
  assign n10278 = ~n10276 & ~n10277;
  assign n10279 = ~n10275 & n10278;
  assign n10280 = pi0896 & ~n10279;
  assign n10281 = ~n10271 & ~n10280;
  assign n10282 = ~n9399 & ~n10281;
  assign po0360 = n10242 | n10282;
  assign n10284 = pi0158 & n9399;
  assign po0361 = n9643 | n10284;
  assign n10286 = pi0159 & n9399;
  assign po0362 = n9729 | n10286;
  assign n10288 = pi0160 & n9399;
  assign po0363 = n9777 | n10288;
  assign n10290 = pi0161 & n9399;
  assign po0364 = n9865 | n10290;
  assign n10292 = pi0162 & n9399;
  assign po0365 = n9821 | n10292;
  assign n10294 = pi0163 & n9399;
  assign po0366 = n9916 | n10294;
  assign n10296 = pi0164 & n9399;
  assign po0367 = n9979 | n10296;
  assign n10298 = pi0165 & n9399;
  assign po0368 = n10010 | n10298;
  assign n10300 = pi0166 & n9399;
  assign po0369 = n10043 | n10300;
  assign n10302 = pi0167 & n9399;
  assign po0370 = n10075 | n10302;
  assign n10304 = pi0168 & n9399;
  assign po0371 = n9685 | n10304;
  assign n10306 = pi0169 & n9399;
  assign po0372 = n10119 | n10306;
  assign n10308 = pi0170 & n9399;
  assign po0373 = n9947 | n10308;
  assign n10310 = pi0171 & n9399;
  assign po0374 = n10240 | n10310;
  assign n10312 = pi0172 & n9399;
  assign po0375 = n10282 | n10312;
  assign n10314 = pi0173 & n9399;
  assign n10315 = pi1713 & ~n9650;
  assign n10316 = pi1815 & n9477;
  assign n10317 = pi1756 & n9454;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = pi2872 & n9498;
  assign n10320 = pi2580 & n9509;
  assign n10321 = ~n10319 & ~n10320;
  assign n10322 = pi2847 & n9441;
  assign n10323 = pi2561 & n9473;
  assign n10324 = ~n10322 & ~n10323;
  assign n10325 = n9150 & n9484;
  assign n10326 = n10324 & ~n10325;
  assign n10327 = n9878 & n10326;
  assign n10328 = n10321 & n10327;
  assign n10329 = n10318 & n10328;
  assign n10330 = ~n10315 & n10329;
  assign n10331 = n9150 & n9428;
  assign n10332 = n10330 & ~n10331;
  assign n10333 = ~n9436 & n10332;
  assign n10334 = ~n7250 & ~n10333;
  assign n10335 = pi0455 & n8059;
  assign n10336 = ~pi0409 & ~n8059;
  assign n10337 = ~n10335 & ~n10336;
  assign n10338 = n7250 & ~n10337;
  assign n10339 = ~n10334 & ~n10338;
  assign n10340 = ~pi0896 & ~n10339;
  assign n10341 = pi0413 & n9404;
  assign n10342 = ~pi0331 & ~n9404;
  assign n10343 = ~n10341 & ~n10342;
  assign n10344 = pi1676 & ~n10343;
  assign n10345 = pi0250 & n9409;
  assign n10346 = pi1675 & n9411;
  assign n10347 = ~n10345 & ~n10346;
  assign n10348 = ~n10344 & n10347;
  assign n10349 = pi0896 & ~n10348;
  assign n10350 = ~n10340 & ~n10349;
  assign n10351 = ~n9399 & ~n10350;
  assign po0376 = n10314 | n10351;
  assign n10353 = pi0174 & n9399;
  assign n10354 = pi2545 & n9441;
  assign n10355 = pi1817 & n9477;
  assign n10356 = ~n10354 & ~n10355;
  assign n10357 = pi2749 & n9473;
  assign n10358 = n9145 & n9484;
  assign n10359 = ~n10357 & ~n10358;
  assign n10360 = pi2870 & n9498;
  assign n10361 = pi1711 & n9480;
  assign n10362 = ~n10360 & ~n10361;
  assign n10363 = pi1711 & n9451;
  assign n10364 = pi1785 & n9454;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = n10362 & n10365;
  assign n10367 = n10359 & n10366;
  assign n10368 = n10356 & n10367;
  assign n10369 = ~n9436 & n10368;
  assign n10370 = pi2787 & n9509;
  assign n10371 = n9145 & n9428;
  assign n10372 = ~n10370 & ~n10371;
  assign n10373 = n10369 & n10372;
  assign n10374 = ~n7250 & ~n10373;
  assign n10375 = pi0453 & n8059;
  assign n10376 = ~pi0386 & ~n8059;
  assign n10377 = ~n10375 & ~n10376;
  assign n10378 = n7250 & ~n10377;
  assign n10379 = ~n10374 & ~n10378;
  assign n10380 = ~pi0896 & ~n10379;
  assign n10381 = pi0414 & n9404;
  assign n10382 = ~pi0282 & ~n9404;
  assign n10383 = ~n10381 & ~n10382;
  assign n10384 = pi1676 & ~n10383;
  assign n10385 = pi0300 & n9409;
  assign n10386 = pi1731 & n9411;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n10384 & n10387;
  assign n10389 = pi0896 & ~n10388;
  assign n10390 = ~n10380 & ~n10389;
  assign n10391 = ~n9399 & ~n10390;
  assign po0377 = n10353 | n10391;
  assign n10393 = pi0175 & n9399;
  assign n10394 = pi2840 & n9441;
  assign n10395 = pi1818 & n9477;
  assign n10396 = ~n10394 & ~n10395;
  assign n10397 = pi2562 & n9473;
  assign n10398 = n9160 & n9484;
  assign n10399 = ~n10397 & ~n10398;
  assign n10400 = pi2869 & n9498;
  assign n10401 = pi1716 & n9480;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = pi1716 & n9451;
  assign n10404 = pi1784 & n9454;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = n10402 & n10405;
  assign n10407 = n10399 & n10406;
  assign n10408 = n10396 & n10407;
  assign n10409 = ~n9436 & n10408;
  assign n10410 = pi2581 & n9509;
  assign n10411 = n9160 & n9428;
  assign n10412 = ~n10410 & ~n10411;
  assign n10413 = n10409 & n10412;
  assign n10414 = ~n7250 & ~n10413;
  assign n10415 = pi0454 & n8059;
  assign n10416 = ~pi0387 & ~n8059;
  assign n10417 = ~n10415 & ~n10416;
  assign n10418 = n7250 & ~n10417;
  assign n10419 = ~n10414 & ~n10418;
  assign n10420 = ~pi0896 & ~n10419;
  assign n10421 = pi0415 & n9404;
  assign n10422 = ~pi0283 & ~n9404;
  assign n10423 = ~n10421 & ~n10422;
  assign n10424 = pi1676 & ~n10423;
  assign n10425 = pi0272 & n9409;
  assign n10426 = pi1732 & n9411;
  assign n10427 = ~n10425 & ~n10426;
  assign n10428 = ~n10424 & n10427;
  assign n10429 = pi0896 & ~n10428;
  assign n10430 = ~n10420 & ~n10429;
  assign n10431 = ~n9399 & ~n10430;
  assign po0378 = n10393 | n10431;
  assign n10433 = pi0176 & n9399;
  assign n10434 = pi2546 & n9441;
  assign n10435 = pi1855 & n9477;
  assign n10436 = ~n10434 & ~n10435;
  assign n10437 = pi2563 & n9473;
  assign n10438 = n9155 & n9484;
  assign n10439 = ~n10437 & ~n10438;
  assign n10440 = n10436 & n10439;
  assign n10441 = pi1791 & n9454;
  assign n10442 = pi2483 & n9509;
  assign n10443 = pi2531 & n9498;
  assign n10444 = ~n10442 & ~n10443;
  assign n10445 = n9155 & n9428;
  assign n10446 = n10444 & ~n10445;
  assign n10447 = pi1718 & n9480;
  assign n10448 = n10446 & ~n10447;
  assign n10449 = pi1718 & n9451;
  assign n10450 = n10448 & ~n10449;
  assign n10451 = ~n10441 & n10450;
  assign n10452 = n10440 & n10451;
  assign n10453 = n9742 & n10452;
  assign n10454 = ~n7250 & ~n10453;
  assign n10455 = pi0456 & n8059;
  assign n10456 = ~pi0388 & ~n8059;
  assign n10457 = ~n10455 & ~n10456;
  assign n10458 = n7250 & ~n10457;
  assign n10459 = ~n10454 & ~n10458;
  assign n10460 = ~pi0896 & ~n10459;
  assign n10461 = pi0416 & n9404;
  assign n10462 = ~pi0284 & ~n9404;
  assign n10463 = ~n10461 & ~n10462;
  assign n10464 = pi1676 & ~n10463;
  assign n10465 = pi0251 & n9409;
  assign n10466 = pi1733 & n9411;
  assign n10467 = ~n10465 & ~n10466;
  assign n10468 = ~n10464 & n10467;
  assign n10469 = pi0896 & ~n10468;
  assign n10470 = ~n10460 & ~n10469;
  assign n10471 = ~n9399 & ~n10470;
  assign po0379 = n10433 | n10471;
  assign n10473 = pi0177 & n9399;
  assign n10474 = pi2842 & n9441;
  assign n10475 = pi1819 & n9477;
  assign n10476 = ~n10474 & ~n10475;
  assign n10477 = pi2518 & n9473;
  assign n10478 = n9174 & n9484;
  assign n10479 = ~n10477 & ~n10478;
  assign n10480 = pi2532 & n9498;
  assign n10481 = pi1714 & n9480;
  assign n10482 = ~n10480 & ~n10481;
  assign n10483 = pi1714 & n9451;
  assign n10484 = pi1786 & n9454;
  assign n10485 = ~n10483 & ~n10484;
  assign n10486 = n10482 & n10485;
  assign n10487 = n10479 & n10486;
  assign n10488 = n10476 & n10487;
  assign n10489 = ~n9436 & n10488;
  assign n10490 = pi2582 & n9509;
  assign n10491 = n9174 & n9428;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = n10489 & n10492;
  assign n10494 = ~n7250 & ~n10493;
  assign n10495 = pi0458 & n8059;
  assign n10496 = ~pi0391 & ~n8059;
  assign n10497 = ~n10495 & ~n10496;
  assign n10498 = n7250 & ~n10497;
  assign n10499 = ~n10494 & ~n10498;
  assign n10500 = ~pi0896 & ~n10499;
  assign n10501 = pi0418 & n9404;
  assign n10502 = ~pi0285 & ~n9404;
  assign n10503 = ~n10501 & ~n10502;
  assign n10504 = pi1676 & ~n10503;
  assign n10505 = pi0252 & n9409;
  assign n10506 = pi1734 & n9411;
  assign n10507 = ~n10505 & ~n10506;
  assign n10508 = ~n10504 & n10507;
  assign n10509 = pi0896 & ~n10508;
  assign n10510 = ~n10500 & ~n10509;
  assign n10511 = ~n9399 & ~n10510;
  assign po0380 = n10473 | n10511;
  assign n10513 = pi0178 & n9399;
  assign n10514 = pi2843 & n9441;
  assign n10515 = pi1854 & n9477;
  assign n10516 = ~n10514 & ~n10515;
  assign n10517 = pi2566 & n9473;
  assign n10518 = n9184 & n9484;
  assign n10519 = ~n10517 & ~n10518;
  assign n10520 = pi2533 & n9498;
  assign n10521 = pi1755 & n9480;
  assign n10522 = ~n10520 & ~n10521;
  assign n10523 = pi1755 & n9451;
  assign n10524 = pi1788 & n9454;
  assign n10525 = ~n10523 & ~n10524;
  assign n10526 = n10522 & n10525;
  assign n10527 = n10519 & n10526;
  assign n10528 = n10516 & n10527;
  assign n10529 = ~n9436 & n10528;
  assign n10530 = pi2583 & n9509;
  assign n10531 = n9184 & n9428;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = n10529 & n10532;
  assign n10534 = ~n7250 & ~n10533;
  assign n10535 = pi0462 & n8059;
  assign n10536 = ~pi0390 & ~n8059;
  assign n10537 = ~n10535 & ~n10536;
  assign n10538 = n7250 & ~n10537;
  assign n10539 = ~n10534 & ~n10538;
  assign n10540 = ~pi0896 & ~n10539;
  assign n10541 = pi0419 & n9404;
  assign n10542 = ~pi0286 & ~n9404;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = pi1676 & ~n10543;
  assign n10545 = pi0253 & n9409;
  assign n10546 = pi1735 & n9411;
  assign n10547 = ~n10545 & ~n10546;
  assign n10548 = ~n10544 & n10547;
  assign n10549 = pi0896 & ~n10548;
  assign n10550 = ~n10540 & ~n10549;
  assign n10551 = ~n9399 & ~n10550;
  assign po0381 = n10513 | n10551;
  assign n10553 = pi0179 & n9399;
  assign n10554 = n9192 & n9484;
  assign n10555 = pi2574 & n9473;
  assign n10556 = ~n10554 & ~n10555;
  assign n10557 = pi2520 & n9501;
  assign n10558 = pi1670 & n9607;
  assign n10559 = ~n10557 & ~n10558;
  assign n10560 = pi2762 & n9441;
  assign n10561 = pi1850 & n9477;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = pi1809 & n9454;
  assign n10564 = n10562 & ~n10563;
  assign n10565 = pi2285 & n9447;
  assign n10566 = n10564 & ~n10565;
  assign n10567 = n10559 & n10566;
  assign n10568 = n10556 & n10567;
  assign n10569 = pi2838 & n9498;
  assign n10570 = n10568 & ~n10569;
  assign n10571 = n9192 & n9428;
  assign n10572 = pi2884 & n9509;
  assign n10573 = ~n10571 & ~n10572;
  assign n10574 = n10570 & n10573;
  assign n10575 = ~n7250 & ~n10574;
  assign n10576 = pi0475 & n8059;
  assign n10577 = ~pi0402 & ~n8059;
  assign n10578 = ~n10576 & ~n10577;
  assign n10579 = n7250 & ~n10578;
  assign n10580 = ~n10575 & ~n10579;
  assign n10581 = ~pi0896 & ~n10580;
  assign n10582 = pi0433 & n9404;
  assign n10583 = ~pi0328 & ~n9404;
  assign n10584 = ~n10582 & ~n10583;
  assign n10585 = pi1676 & ~n10584;
  assign n10586 = pi0263 & n9409;
  assign n10587 = pi1744 & n9411;
  assign n10588 = ~n10586 & ~n10587;
  assign n10589 = ~n10585 & n10588;
  assign n10590 = pi0896 & ~n10589;
  assign n10591 = ~n10581 & ~n10590;
  assign n10592 = ~n9399 & ~n10591;
  assign po0382 = n10553 | n10592;
  assign n10594 = pi0180 & n9399;
  assign n10595 = pi1812 & n9477;
  assign n10596 = pi2849 & n9441;
  assign n10597 = pi1780 & n9454;
  assign n10598 = ~n10596 & ~n10597;
  assign n10599 = pi2521 & n9501;
  assign n10600 = pi1700 & n9607;
  assign n10601 = ~n10599 & ~n10600;
  assign n10602 = pi2556 & n9473;
  assign n10603 = n9207 & n9484;
  assign n10604 = ~n10602 & ~n10603;
  assign n10605 = n10601 & n10604;
  assign n10606 = n10598 & n10605;
  assign n10607 = ~n10595 & n10606;
  assign n10608 = pi2854 & n9498;
  assign n10609 = n10607 & ~n10608;
  assign n10610 = pi2576 & n9509;
  assign n10611 = n9207 & n9428;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = n10609 & n10612;
  assign n10614 = ~n7250 & ~n10613;
  assign n10615 = pi0478 & n8059;
  assign n10616 = ~pi0382 & ~n8059;
  assign n10617 = ~n10615 & ~n10616;
  assign n10618 = n7250 & ~n10617;
  assign n10619 = ~n10614 & ~n10618;
  assign n10620 = ~pi0896 & ~n10619;
  assign n10621 = pi0438 & n9404;
  assign n10622 = ~pi0276 & ~n9404;
  assign n10623 = ~n10621 & ~n10622;
  assign n10624 = pi1676 & ~n10623;
  assign n10625 = pi0303 & n9409;
  assign n10626 = pi1727 & n9411;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = ~n10624 & n10627;
  assign n10629 = pi0896 & ~n10628;
  assign n10630 = ~n10620 & ~n10629;
  assign n10631 = ~n9399 & ~n10630;
  assign po0383 = n10594 | n10631;
  assign n10633 = pi0181 & n9399;
  assign po0384 = n10351 | n10633;
  assign n10635 = pi0182 & n9399;
  assign po0385 = n10391 | n10635;
  assign n10637 = pi0183 & n9399;
  assign po0386 = n10431 | n10637;
  assign n10639 = pi0184 & n9399;
  assign po0387 = n10471 | n10639;
  assign n10641 = pi0185 & n9399;
  assign po0388 = n10551 | n10641;
  assign n10643 = pi0186 & n9399;
  assign po0389 = n10511 | n10643;
  assign n10645 = pi0187 & n9399;
  assign po0390 = n10631 | n10645;
  assign n10647 = pi0188 & n9399;
  assign po0391 = n10592 | n10647;
  assign n10649 = pi0189 & n9399;
  assign po0392 = n10157 | n10649;
  assign n10651 = pi0190 & n9399;
  assign po0393 = n10198 | n10651;
  assign n10653 = pi0191 & n9399;
  assign n10654 = pi2564 & n9473;
  assign n10655 = pi1338 & n9872;
  assign n10656 = ~n10654 & ~n10655;
  assign n10657 = pi1351 & n9882;
  assign n10658 = n10656 & ~n10657;
  assign n10659 = pi2841 & n9441;
  assign n10660 = pi1355 & n9884;
  assign n10661 = ~n10659 & ~n10660;
  assign n10662 = pi2864 & n9498;
  assign n10663 = pi1357 & n9741;
  assign n10664 = ~n10662 & ~n10663;
  assign n10665 = pi1708 & n9607;
  assign n10666 = n10664 & ~n10665;
  assign n10667 = n10661 & n10666;
  assign n10668 = n10658 & n10667;
  assign n10669 = pi1396 & n9506;
  assign n10670 = pi2755 & n9509;
  assign n10671 = ~n10669 & ~n10670;
  assign n10672 = pi1373 & n9898;
  assign n10673 = pi1361 & n9422;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = n10671 & n10674;
  assign n10676 = n10668 & n10675;
  assign n10677 = ~n7250 & n10676;
  assign n10678 = pi0457 & n8059;
  assign n10679 = ~pi0408 & ~n8059;
  assign n10680 = ~n10678 & ~n10679;
  assign n10681 = n7250 & n10680;
  assign n10682 = ~n10677 & ~n10681;
  assign n10683 = ~pi0896 & ~n10682;
  assign n10684 = pi1672 & n9411;
  assign n10685 = pi0305 & pi0306;
  assign n10686 = ~pi0307 & ~pi1683;
  assign n10687 = n10685 & n10686;
  assign n10688 = ~pi0307 & pi1683;
  assign n10689 = pi0307 & pi1683;
  assign n10690 = ~n10688 & ~n10689;
  assign n10691 = pi0305 & ~pi0306;
  assign n10692 = ~n10690 & n10691;
  assign n10693 = ~n10687 & ~n10692;
  assign n10694 = n10685 & ~n10690;
  assign n10695 = n10693 & ~n10694;
  assign n10696 = n9409 & n10695;
  assign n10697 = pi0205 & pi1902;
  assign n10698 = ~pi0305 & ~pi0306;
  assign n10699 = ~n10690 & n10698;
  assign n10700 = pi0206 & pi0207;
  assign n10701 = n10699 & ~n10700;
  assign n10702 = n10697 & n10701;
  assign n10703 = pi0326 & ~n10699;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = n10696 & ~n10704;
  assign n10706 = ~n10684 & ~n10705;
  assign n10707 = pi0417 & n9404;
  assign n10708 = ~pi0329 & ~n9404;
  assign n10709 = ~n10707 & ~n10708;
  assign n10710 = pi1676 & ~n10709;
  assign n10711 = n10706 & ~n10710;
  assign n10712 = pi0896 & n10711;
  assign n10713 = ~n10683 & ~n10712;
  assign n10714 = ~n9399 & n10713;
  assign po0394 = n10653 | n10714;
  assign n10716 = pi0192 & n9399;
  assign n10717 = pi0468 & n8059;
  assign n10718 = ~pi0404 & ~n8059;
  assign n10719 = ~n10717 & ~n10718;
  assign n10720 = n7250 & ~n10719;
  assign n10721 = pi2859 & n9498;
  assign n10722 = pi2522 & n9501;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = pi2894 & n9509;
  assign n10725 = n10723 & ~n10724;
  assign n10726 = pi2761 & n9441;
  assign n10727 = pi2482 & n9447;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = pi0197 & n9422;
  assign n10730 = n9106 & n9428;
  assign n10731 = ~n10729 & ~n10730;
  assign n10732 = n10728 & n10731;
  assign n10733 = ~n9436 & n10732;
  assign n10734 = n10725 & n10733;
  assign n10735 = pi1823 & n9477;
  assign n10736 = pi1794 & n9454;
  assign n10737 = ~n10735 & ~n10736;
  assign n10738 = pi2501 & n9473;
  assign n10739 = n9106 & n9484;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = pi1722 & ~n9650;
  assign n10742 = n10740 & ~n10741;
  assign n10743 = n10737 & n10742;
  assign n10744 = n10734 & n10743;
  assign n10745 = ~n7250 & ~n10744;
  assign n10746 = ~n10720 & ~n10745;
  assign n10747 = ~pi0896 & ~n10746;
  assign n10748 = pi0448 & n9404;
  assign n10749 = ~pi0352 & ~n9404;
  assign n10750 = ~n10748 & ~n10749;
  assign n10751 = pi1676 & ~n10750;
  assign n10752 = pi0271 & n9409;
  assign n10753 = pi1745 & n9411;
  assign n10754 = ~n10752 & ~n10753;
  assign n10755 = ~n10751 & n10754;
  assign n10756 = pi0896 & ~n10755;
  assign n10757 = ~n10747 & ~n10756;
  assign n10758 = ~n9399 & ~n10757;
  assign po0395 = n10716 | n10758;
  assign n10760 = pi0193 & n9399;
  assign po0396 = n10714 | n10760;
  assign n10762 = pi0194 & n9399;
  assign po0397 = n10758 | n10762;
  assign n10764 = pi0195 & n9399;
  assign n10765 = pi2547 & n9441;
  assign n10766 = pi1820 & n9477;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = pi2565 & n9473;
  assign n10769 = n9179 & n9484;
  assign n10770 = ~n10768 & ~n10769;
  assign n10771 = pi2867 & n9498;
  assign n10772 = pi1754 & n9480;
  assign n10773 = ~n10771 & ~n10772;
  assign n10774 = pi1754 & n9451;
  assign n10775 = pi1779 & n9454;
  assign n10776 = ~n10774 & ~n10775;
  assign n10777 = n10773 & n10776;
  assign n10778 = n10770 & n10777;
  assign n10779 = n10767 & n10778;
  assign n10780 = ~n9436 & n10779;
  assign n10781 = pi2856 & n9509;
  assign n10782 = n9179 & n9428;
  assign n10783 = ~n10781 & ~n10782;
  assign n10784 = n10780 & n10783;
  assign n10785 = ~n7250 & ~n10784;
  assign n10786 = pi0459 & n8059;
  assign n10787 = ~pi0389 & ~n8059;
  assign n10788 = ~n10786 & ~n10787;
  assign n10789 = n7250 & ~n10788;
  assign n10790 = ~n10785 & ~n10789;
  assign n10791 = ~pi0896 & ~n10790;
  assign n10792 = pi0446 & n9404;
  assign n10793 = ~pi0333 & ~n9404;
  assign n10794 = ~n10792 & ~n10793;
  assign n10795 = pi1676 & ~n10794;
  assign n10796 = pi0269 & n9409;
  assign n10797 = pi1673 & n9411;
  assign n10798 = ~n10796 & ~n10797;
  assign n10799 = ~n10795 & n10798;
  assign n10800 = pi0896 & ~n10799;
  assign n10801 = ~n10791 & ~n10800;
  assign n10802 = ~n9399 & ~n10801;
  assign po0398 = n10764 | n10802;
  assign n10804 = pi0196 & n9399;
  assign po0399 = n10802 | n10804;
  assign n10806 = ~pi3018 & pi3133;
  assign n10807 = n7247 & n10806;
  assign n10808 = n7254 & n10807;
  assign n10809 = pi0197 & ~n10808;
  assign po0400 = ~pi0230 | n10809;
  assign n10811 = pi0198 & n9399;
  assign n10812 = pi2534 & n9498;
  assign n10813 = pi2851 & n9501;
  assign n10814 = ~n10812 & ~n10813;
  assign n10815 = pi2585 & n9509;
  assign n10816 = pi2818 & n9441;
  assign n10817 = pi1807 & n9454;
  assign n10818 = ~n10816 & ~n10817;
  assign n10819 = ~n9660 & n10818;
  assign n10820 = pi2738 & n9447;
  assign n10821 = pi1752 & n9451;
  assign n10822 = ~n10820 & ~n10821;
  assign n10823 = pi1852 & n9477;
  assign n10824 = pi1752 & n9480;
  assign n10825 = ~n10823 & ~n10824;
  assign n10826 = pi2569 & n9473;
  assign n10827 = n9225 & n9484;
  assign n10828 = ~n10826 & ~n10827;
  assign n10829 = n10825 & n10828;
  assign n10830 = n10822 & n10829;
  assign n10831 = n10819 & n10830;
  assign n10832 = n9225 & n9428;
  assign n10833 = n10831 & ~n10832;
  assign n10834 = ~n9436 & n10833;
  assign n10835 = ~n10815 & n10834;
  assign n10836 = n10814 & n10835;
  assign n10837 = n9516 & ~n10836;
  assign n10838 = pi0463 & n8059;
  assign n10839 = ~pi0393 & ~n8059;
  assign n10840 = ~n10838 & ~n10839;
  assign n10841 = n9522 & ~n10840;
  assign n10842 = ~n10837 & ~n10841;
  assign n10843 = ~n9399 & ~n10842;
  assign n10844 = pi0896 & ~n9399;
  assign n10845 = pi0410 & n9404;
  assign n10846 = ~pi0264 & ~n9404;
  assign n10847 = ~n10845 & ~n10846;
  assign n10848 = pi1676 & ~n10847;
  assign n10849 = pi0247 & n9409;
  assign n10850 = pi1738 & n9411;
  assign n10851 = ~n10849 & ~n10850;
  assign n10852 = ~n10848 & n10851;
  assign n10853 = n10844 & ~n10852;
  assign n10854 = ~n10843 & ~n10853;
  assign po0401 = n10811 | ~n10854;
  assign n10856 = pi0199 & n9399;
  assign po0402 = ~n10854 | n10856;
  assign n10858 = pi0200 & n9399;
  assign n10859 = pi0477 & n8059;
  assign n10860 = ~pi0381 & ~n8059;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = n9522 & ~n10861;
  assign n10863 = pi1348 & n9501;
  assign n10864 = pi1356 & n9741;
  assign n10865 = ~n10863 & ~n10864;
  assign n10866 = pi3178 & n9898;
  assign n10867 = pi1360 & n9422;
  assign n10868 = ~n10866 & ~n10867;
  assign n10869 = pi2527 & n9498;
  assign n10870 = pi1970 & n9509;
  assign n10871 = ~n10869 & ~n10870;
  assign n10872 = pi1395 & n9506;
  assign n10873 = n10871 & ~n10872;
  assign n10874 = n10868 & n10873;
  assign n10875 = pi1341 & n9447;
  assign n10876 = pi1358 & n9882;
  assign n10877 = ~n10875 & ~n10876;
  assign n10878 = pi1354 & n9884;
  assign n10879 = pi1793 & n9484;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = n9453 & n9460;
  assign n10882 = pi1364 & n10881;
  assign n10883 = ~n9877 & ~n10882;
  assign n10884 = ~n9660 & n10883;
  assign n10885 = pi2541 & n9441;
  assign n10886 = n10884 & ~n10885;
  assign n10887 = n10880 & n10886;
  assign n10888 = n10877 & n10887;
  assign n10889 = pi2480 & n9473;
  assign n10890 = n10888 & ~n10889;
  assign n10891 = n9435 & n9460;
  assign n10892 = pi1363 & n10891;
  assign n10893 = n10890 & ~n10892;
  assign n10894 = ~n9876 & n10893;
  assign n10895 = n10874 & n10894;
  assign n10896 = pi1706 & n9607;
  assign n10897 = pi1793 & n9428;
  assign n10898 = ~n10896 & ~n10897;
  assign n10899 = n10895 & n10898;
  assign n10900 = n10865 & n10899;
  assign n10901 = n9516 & ~n10900;
  assign n10902 = ~n10862 & ~n10901;
  assign n10903 = ~n9399 & ~n10902;
  assign n10904 = pi0437 & n9404;
  assign n10905 = ~pi0275 & ~n9404;
  assign n10906 = ~n10904 & ~n10905;
  assign n10907 = pi1676 & ~n10906;
  assign n10908 = pi0205 & ~pi1902;
  assign n10909 = n10699 & n10908;
  assign n10910 = pi0206 & ~pi0207;
  assign n10911 = pi0205 & n10699;
  assign n10912 = n10910 & n10911;
  assign n10913 = ~n10909 & ~n10912;
  assign n10914 = n10695 & ~n10913;
  assign n10915 = pi0308 & n10695;
  assign n10916 = ~n10699 & n10915;
  assign n10917 = ~n10914 & ~n10916;
  assign n10918 = n9409 & ~n10917;
  assign n10919 = pi1726 & n9411;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = ~n10907 & n10920;
  assign n10922 = n10844 & ~n10921;
  assign n10923 = ~n10903 & ~n10922;
  assign po0403 = n10858 | ~n10923;
  assign n10925 = pi0201 & n9399;
  assign po0404 = ~n10923 | n10925;
  assign n10927 = pi0203 & n9399;
  assign n10928 = ~n9422 & ~n9741;
  assign n10929 = pi2863 & n9498;
  assign n10930 = pi2848 & n9501;
  assign n10931 = ~n10929 & ~n10930;
  assign n10932 = pi2901 & n9509;
  assign n10933 = n10931 & ~n10932;
  assign n10934 = n9090 & n9428;
  assign n10935 = n10933 & ~n10934;
  assign n10936 = ~n9436 & n10935;
  assign n10937 = pi2554 & n9447;
  assign n10938 = pi1719 & n9451;
  assign n10939 = ~n10937 & ~n10938;
  assign n10940 = pi1790 & n9454;
  assign n10941 = pi2548 & n9441;
  assign n10942 = pi1719 & n9480;
  assign n10943 = ~n10941 & ~n10942;
  assign n10944 = ~n9660 & n10943;
  assign n10945 = ~n10940 & n10944;
  assign n10946 = n10939 & n10945;
  assign n10947 = pi1853 & n9477;
  assign n10948 = n10946 & ~n10947;
  assign n10949 = pi2568 & n9473;
  assign n10950 = n9090 & n9484;
  assign n10951 = ~n10949 & ~n10950;
  assign n10952 = n10948 & n10951;
  assign n10953 = n10936 & n10952;
  assign n10954 = n10928 & n10953;
  assign n10955 = n9516 & ~n10954;
  assign n10956 = pi0449 & n8059;
  assign n10957 = ~pi0378 & ~n8059;
  assign n10958 = ~n10956 & ~n10957;
  assign n10959 = n9522 & ~n10958;
  assign n10960 = ~n10955 & ~n10959;
  assign n10961 = ~n9399 & ~n10960;
  assign n10962 = pi0447 & n9404;
  assign n10963 = ~pi0334 & ~n9404;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = pi1676 & ~n10964;
  assign n10966 = pi0270 & n9409;
  assign n10967 = pi1737 & n9411;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = ~n10965 & n10968;
  assign n10970 = n10844 & ~n10969;
  assign n10971 = ~n10961 & ~n10970;
  assign po0406 = n10927 | ~n10971;
  assign n10973 = pi0204 & n9399;
  assign po0407 = ~n10971 | n10973;
  assign n10975 = pi1858 & n9404;
  assign po3351 = pi1858 | pi2911;
  assign n10977 = ~pi1337 & ~po3351;
  assign n10978 = ~pi2989 & ~n10977;
  assign n10979 = ~n10975 & ~n10978;
  assign n10980 = pi0205 & n10979;
  assign n10981 = ~pi1858 & ~n9545;
  assign n10982 = ~pi0273 & pi1858;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = ~n10979 & ~n10983;
  assign po0408 = n10980 | n10984;
  assign n10986 = pi0206 & n10979;
  assign n10987 = ~pi1858 & ~n9585;
  assign n10988 = ~pi0274 & pi1858;
  assign n10989 = ~n10987 & ~n10988;
  assign n10990 = ~n10979 & ~n10989;
  assign po0409 = n10986 | n10990;
  assign n10992 = pi0207 & n10979;
  assign n10993 = ~pi1858 & ~n9563;
  assign n10994 = ~pi0332 & pi1858;
  assign n10995 = ~n10993 & ~n10994;
  assign n10996 = ~n10979 & ~n10995;
  assign po0410 = n10992 | n10996;
  assign n10998 = n8188 & n8296;
  assign n10999 = n8295 & n10998;
  assign n11000 = n8194 & n8300;
  assign n11001 = n8197 & n11000;
  assign n11002 = ~pi0359 & n8206;
  assign n11003 = ~n8298 & ~n11002;
  assign n11004 = n11001 & ~n11003;
  assign n11005 = pi0082 & n8196;
  assign n11006 = ~n8200 & n11005;
  assign n11007 = ~pi0359 & n8229;
  assign n11008 = n8187 & ~n8224;
  assign n11009 = n8200 & n11008;
  assign n11010 = n11007 & n11009;
  assign n11011 = pi0082 & pi1811;
  assign n11012 = ~pi0079 & n11011;
  assign n11013 = ~n8200 & n11012;
  assign n11014 = ~n11010 & ~n11013;
  assign n11015 = ~n11006 & n11014;
  assign n11016 = ~n11004 & n11015;
  assign n11017 = ~n10999 & n11016;
  assign n11018 = ~pi2960 & ~n11017;
  assign n11019 = pi0208 & ~n11018;
  assign n11020 = pi0341 & n11018;
  assign po0411 = n11019 | n11020;
  assign n11022 = pi0209 & ~n11018;
  assign n11023 = pi0342 & n11018;
  assign po0412 = n11022 | n11023;
  assign n11025 = pi0210 & ~n11018;
  assign n11026 = pi0343 & n11018;
  assign po0413 = n11025 | n11026;
  assign n11028 = pi0211 & ~n11018;
  assign n11029 = pi0344 & n11018;
  assign po0414 = n11028 | n11029;
  assign n11031 = pi0212 & ~n11018;
  assign n11032 = pi0345 & n11018;
  assign po0415 = n11031 | n11032;
  assign n11034 = pi0213 & ~n11018;
  assign n11035 = pi0346 & n11018;
  assign po0416 = n11034 | n11035;
  assign n11037 = pi0214 & ~n11018;
  assign n11038 = pi0347 & n11018;
  assign po0417 = n11037 | n11038;
  assign n11040 = pi0215 & ~n11018;
  assign n11041 = pi0348 & n11018;
  assign po0418 = n11040 | n11041;
  assign n11043 = pi0216 & ~n11018;
  assign n11044 = pi0349 & n11018;
  assign po0419 = n11043 | n11044;
  assign n11046 = pi0217 & ~n11018;
  assign n11047 = pi0350 & n11018;
  assign po0420 = n11046 | n11047;
  assign n11049 = pi0218 & ~n11018;
  assign n11050 = pi0351 & n11018;
  assign po0421 = n11049 | n11050;
  assign po0422 = ~n9368 | ~n9375;
  assign n11053 = pi3152 & n8008;
  assign n11054 = pi2950 & ~n11053;
  assign n11055 = n7257 & ~n11054;
  assign n11056 = pi3160 & n11055;
  assign n11057 = pi1365 & n11056;
  assign po0431 = n9368 & n11057;
  assign po0424 = ~n9368 | n11054;
  assign n11060 = pi0222 & ~pi3364;
  assign n11061 = ~pi3365 & n11060;
  assign po0425 = pi0339 | n11061;
  assign n11063 = pi0225 & ~n11018;
  assign n11064 = pi0353 & n11018;
  assign po0426 = n11063 | n11064;
  assign n11066 = pi0226 & ~n11018;
  assign n11067 = pi0354 & n11018;
  assign po0427 = n11066 | n11067;
  assign n11069 = pi0227 & ~n11018;
  assign n11070 = pi0355 & n11018;
  assign po0428 = n11069 | n11070;
  assign n11072 = pi0228 & ~n11018;
  assign n11073 = pi0356 & n11018;
  assign po0429 = n11072 | n11073;
  assign n11075 = pi0229 & ~n11018;
  assign n11076 = pi0357 & n11018;
  assign po0430 = n11075 | n11076;
  assign n11078 = pi0231 & ~n11018;
  assign n11079 = pi0361 & n11018;
  assign po0432 = n11078 | n11079;
  assign n11081 = pi0232 & ~n11018;
  assign n11082 = pi0362 & n11018;
  assign po0433 = n11081 | n11082;
  assign n11084 = pi0233 & ~n11018;
  assign n11085 = pi0363 & n11018;
  assign po0434 = n11084 | n11085;
  assign n11087 = pi0234 & ~n11018;
  assign n11088 = pi0364 & n11018;
  assign po0435 = n11087 | n11088;
  assign n11090 = pi0235 & ~n11018;
  assign n11091 = pi0365 & n11018;
  assign po0436 = n11090 | n11091;
  assign n11093 = pi0236 & ~n11018;
  assign n11094 = pi0366 & n11018;
  assign po0437 = n11093 | n11094;
  assign n11096 = pi0237 & ~n11018;
  assign n11097 = pi0367 & n11018;
  assign po0438 = n11096 | n11097;
  assign n11099 = pi0238 & ~n11018;
  assign n11100 = pi0368 & n11018;
  assign po0439 = n11099 | n11100;
  assign n11102 = pi0239 & ~n11018;
  assign n11103 = pi0369 & n11018;
  assign po0440 = n11102 | n11103;
  assign n11105 = pi0240 & ~n11018;
  assign n11106 = pi0370 & n11018;
  assign po0441 = n11105 | n11106;
  assign n11108 = pi0241 & ~n11018;
  assign n11109 = pi0371 & n11018;
  assign po0442 = n11108 | n11109;
  assign n11111 = pi0242 & ~n11018;
  assign n11112 = pi0372 & n11018;
  assign po0443 = n11111 | n11112;
  assign n11114 = pi0243 & ~n11018;
  assign n11115 = pi0373 & n11018;
  assign po0444 = n11114 | n11115;
  assign n11117 = pi0244 & ~n11018;
  assign n11118 = pi0374 & n11018;
  assign po0445 = n11117 | n11118;
  assign n11120 = pi0245 & ~n11018;
  assign n11121 = pi0375 & n11018;
  assign po0446 = n11120 | n11121;
  assign n11123 = pi0246 & ~n11018;
  assign n11124 = pi0376 & n11018;
  assign po0447 = n11123 | n11124;
  assign n11126 = ~pi1337 & ~pi1827;
  assign n11127 = ~po3351 & n11126;
  assign n11128 = ~pi1307 & ~pi3213;
  assign n11129 = pi1307 & pi3213;
  assign n11130 = ~n11128 & ~n11129;
  assign n11131 = ~pi1309 & pi3214;
  assign n11132 = pi1309 & ~pi3214;
  assign n11133 = ~n11131 & ~n11132;
  assign n11134 = ~pi1239 & pi3223;
  assign n11135 = pi1239 & ~pi3223;
  assign n11136 = ~n11134 & ~n11135;
  assign n11137 = n11133 & n11136;
  assign n11138 = n11130 & n11137;
  assign n11139 = n11127 & ~n11138;
  assign n11140 = ~pi1254 & ~pi3232;
  assign n11141 = pi1254 & pi3232;
  assign n11142 = ~n11140 & ~n11141;
  assign n11143 = ~pi1250 & ~pi3226;
  assign n11144 = pi1250 & pi3226;
  assign n11145 = ~n11143 & ~n11144;
  assign n11146 = ~n11142 & ~n11145;
  assign n11147 = ~pi1252 & ~pi3228;
  assign n11148 = pi1252 & pi3228;
  assign n11149 = ~n11147 & ~n11148;
  assign n11150 = ~pi1251 & ~pi3237;
  assign n11151 = pi1251 & pi3237;
  assign n11152 = ~n11150 & ~n11151;
  assign n11153 = ~n11149 & ~n11152;
  assign n11154 = n11146 & n11153;
  assign n11155 = n11139 & ~n11154;
  assign n11156 = pi0410 & n11155;
  assign n11157 = ~pi1144 & ~n11155;
  assign n11158 = ~n11156 & ~n11157;
  assign n11159 = n10977 & ~n11158;
  assign n11160 = pi0251 & pi0272;
  assign n11161 = pi0252 & pi0269;
  assign n11162 = n11160 & n11161;
  assign n11163 = pi0262 & pi0302;
  assign n11164 = pi0261 & n11163;
  assign n11165 = pi0263 & n11164;
  assign n11166 = pi0268 & pi0301;
  assign n11167 = pi0260 & n11166;
  assign n11168 = pi0248 & n11167;
  assign n11169 = n11165 & n11168;
  assign n11170 = pi0303 & pi0325;
  assign n11171 = pi0298 & pi0304;
  assign n11172 = n11170 & n11171;
  assign n11173 = pi0249 & pi0299;
  assign n11174 = pi0250 & pi0300;
  assign n11175 = n11173 & n11174;
  assign n11176 = n11172 & n11175;
  assign n11177 = pi0253 & pi0254;
  assign n11178 = pi0255 & pi0270;
  assign n11179 = n11177 & n11178;
  assign n11180 = n11176 & n11179;
  assign n11181 = n11169 & n11180;
  assign n11182 = n11162 & n11181;
  assign n11183 = pi0247 & n11182;
  assign n11184 = ~pi0247 & ~n11182;
  assign n11185 = ~n11183 & ~n11184;
  assign n11186 = n10975 & n11185;
  assign n11187 = pi0247 & ~n10975;
  assign n11188 = ~n11186 & ~n11187;
  assign n11189 = ~n10977 & ~n11188;
  assign po0448 = n11159 | n11189;
  assign n11191 = pi0429 & n11155;
  assign n11192 = ~pi1186 & ~n11155;
  assign n11193 = ~n11191 & ~n11192;
  assign n11194 = n10977 & ~n11193;
  assign n11195 = ~pi0248 & ~n11167;
  assign n11196 = ~n11168 & ~n11195;
  assign n11197 = n10975 & n11196;
  assign n11198 = pi0248 & ~n10975;
  assign n11199 = ~n11197 & ~n11198;
  assign n11200 = ~n10977 & ~n11199;
  assign po0449 = n11194 | n11200;
  assign n11202 = pi0442 & n11155;
  assign n11203 = ~pi1193 & ~n11155;
  assign n11204 = ~n11202 & ~n11203;
  assign n11205 = n10977 & ~n11204;
  assign n11206 = n11169 & n11172;
  assign n11207 = pi0249 & n11206;
  assign n11208 = ~pi0249 & ~n11206;
  assign n11209 = ~n11207 & ~n11208;
  assign n11210 = n10975 & n11209;
  assign n11211 = pi0249 & ~n10975;
  assign n11212 = ~n11210 & ~n11211;
  assign n11213 = ~n10977 & ~n11212;
  assign po0450 = n11205 | n11213;
  assign n11215 = pi0413 & n11155;
  assign n11216 = ~pi1137 & ~n11155;
  assign n11217 = ~n11215 & ~n11216;
  assign n11218 = n10977 & ~n11217;
  assign n11219 = pi0263 & pi0302;
  assign n11220 = n11170 & n11219;
  assign n11221 = pi0260 & pi0262;
  assign n11222 = pi0248 & pi0261;
  assign n11223 = n11221 & n11222;
  assign n11224 = n11166 & n11223;
  assign n11225 = n11220 & n11224;
  assign n11226 = n11171 & n11173;
  assign n11227 = n11225 & n11226;
  assign n11228 = pi0250 & n11227;
  assign n11229 = ~pi0250 & ~n11227;
  assign n11230 = ~n11228 & ~n11229;
  assign n11231 = n10975 & n11230;
  assign n11232 = pi0250 & ~n10975;
  assign n11233 = ~n11231 & ~n11232;
  assign n11234 = ~n10977 & ~n11233;
  assign po0451 = n11218 | n11234;
  assign n11236 = pi0416 & n11155;
  assign n11237 = ~pi1139 & ~n11155;
  assign n11238 = ~n11236 & ~n11237;
  assign n11239 = n10977 & ~n11238;
  assign n11240 = pi0260 & pi0301;
  assign n11241 = n11222 & n11240;
  assign n11242 = pi0263 & pi0303;
  assign n11243 = n11163 & n11242;
  assign n11244 = n11241 & n11243;
  assign n11245 = pi0249 & pi0325;
  assign n11246 = n11171 & n11245;
  assign n11247 = pi0250 & pi0299;
  assign n11248 = pi0272 & pi0300;
  assign n11249 = n11247 & n11248;
  assign n11250 = n11246 & n11249;
  assign n11251 = n11244 & n11250;
  assign n11252 = pi0268 & n11251;
  assign n11253 = pi0251 & n11252;
  assign n11254 = ~pi0251 & ~n11252;
  assign n11255 = ~n11253 & ~n11254;
  assign n11256 = n10975 & n11255;
  assign n11257 = pi0251 & ~n10975;
  assign n11258 = ~n11256 & ~n11257;
  assign n11259 = ~n10977 & ~n11258;
  assign po0452 = n11239 | n11259;
  assign n11261 = pi0418 & n11155;
  assign n11262 = ~pi1141 & ~n11155;
  assign n11263 = ~n11261 & ~n11262;
  assign n11264 = n10977 & ~n11263;
  assign n11265 = n11160 & n11174;
  assign n11266 = n11220 & n11226;
  assign n11267 = n11223 & n11266;
  assign n11268 = n11166 & n11267;
  assign n11269 = n11265 & n11268;
  assign n11270 = pi0252 & n11269;
  assign n11271 = ~pi0252 & ~n11269;
  assign n11272 = ~n11270 & ~n11271;
  assign n11273 = n10975 & n11272;
  assign n11274 = pi0252 & ~n10975;
  assign n11275 = ~n11273 & ~n11274;
  assign n11276 = ~n10977 & ~n11275;
  assign po0453 = n11264 | n11276;
  assign n11278 = pi0419 & n11155;
  assign n11279 = ~pi1184 & ~n11155;
  assign n11280 = ~n11278 & ~n11279;
  assign n11281 = n10977 & ~n11280;
  assign n11282 = n11165 & n11176;
  assign n11283 = n11162 & n11282;
  assign n11284 = n11168 & n11283;
  assign n11285 = pi0253 & n11284;
  assign n11286 = ~pi0253 & ~n11284;
  assign n11287 = ~n11285 & ~n11286;
  assign n11288 = n10975 & n11287;
  assign n11289 = pi0253 & ~n10975;
  assign n11290 = ~n11288 & ~n11289;
  assign n11291 = ~n10977 & ~n11290;
  assign po0454 = n11281 | n11291;
  assign n11293 = pi0420 & n11155;
  assign n11294 = ~pi1142 & ~n11155;
  assign n11295 = ~n11293 & ~n11294;
  assign n11296 = n10977 & ~n11295;
  assign n11297 = pi0251 & pi0252;
  assign n11298 = pi0253 & pi0269;
  assign n11299 = n11297 & n11298;
  assign n11300 = pi0268 & n11241;
  assign n11301 = n11243 & n11250;
  assign n11302 = n11300 & n11301;
  assign n11303 = n11299 & n11302;
  assign n11304 = pi0254 & n11303;
  assign n11305 = ~pi0254 & ~n11303;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = n10975 & n11306;
  assign n11308 = pi0254 & ~n10975;
  assign n11309 = ~n11307 & ~n11308;
  assign n11310 = ~n10977 & ~n11309;
  assign po0455 = n11296 | n11310;
  assign n11312 = pi0421 & n11155;
  assign n11313 = ~pi1143 & ~n11155;
  assign n11314 = ~n11312 & ~n11313;
  assign n11315 = n10977 & ~n11314;
  assign n11316 = n11161 & n11177;
  assign n11317 = n11266 & n11316;
  assign n11318 = n11224 & n11317;
  assign n11319 = n11265 & n11318;
  assign n11320 = pi0255 & n11319;
  assign n11321 = ~pi0255 & ~n11319;
  assign n11322 = ~n11320 & ~n11321;
  assign n11323 = n10975 & n11322;
  assign n11324 = pi0255 & ~n10975;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = ~n10977 & ~n11325;
  assign po0456 = n11315 | n11326;
  assign n11328 = pi0422 & n11155;
  assign n11329 = ~pi1145 & ~n11155;
  assign n11330 = ~n11328 & ~n11329;
  assign n11331 = n10977 & ~n11330;
  assign n11332 = n11243 & n11300;
  assign n11333 = pi0254 & pi0255;
  assign n11334 = pi0247 & pi0270;
  assign n11335 = n11333 & n11334;
  assign n11336 = n11250 & n11335;
  assign n11337 = n11332 & n11336;
  assign n11338 = n11299 & n11337;
  assign n11339 = pi0256 & n11338;
  assign n11340 = ~pi0256 & ~n11338;
  assign n11341 = ~n11339 & ~n11340;
  assign n11342 = n10975 & n11341;
  assign n11343 = pi0256 & ~n10975;
  assign n11344 = ~n11342 & ~n11343;
  assign n11345 = ~n10977 & ~n11344;
  assign po0457 = n11331 | n11345;
  assign n11347 = pi0423 & n11155;
  assign n11348 = ~pi1146 & ~n11155;
  assign n11349 = ~n11347 & ~n11348;
  assign n11350 = n10977 & ~n11349;
  assign n11351 = pi0247 & pi0256;
  assign n11352 = n11178 & n11351;
  assign n11353 = n11265 & n11352;
  assign n11354 = n11225 & n11353;
  assign n11355 = n11226 & n11354;
  assign n11356 = n11316 & n11355;
  assign n11357 = pi0257 & n11356;
  assign n11358 = ~pi0257 & ~n11356;
  assign n11359 = ~n11357 & ~n11358;
  assign n11360 = n10975 & n11359;
  assign n11361 = pi0257 & ~n10975;
  assign n11362 = ~n11360 & ~n11361;
  assign n11363 = ~n10977 & ~n11362;
  assign po0458 = n11350 | n11363;
  assign n11365 = pi0424 & n11155;
  assign n11366 = ~pi1156 & ~n11155;
  assign n11367 = ~n11365 & ~n11366;
  assign n11368 = n10977 & ~n11367;
  assign n11369 = pi0256 & pi0257;
  assign n11370 = pi0304 & n11170;
  assign n11371 = pi0263 & n11370;
  assign n11372 = n11167 & n11222;
  assign n11373 = n11163 & n11372;
  assign n11374 = n11371 & n11373;
  assign n11375 = n11298 & n11333;
  assign n11376 = n11374 & n11375;
  assign n11377 = pi0249 & pi0298;
  assign n11378 = n11247 & n11377;
  assign n11379 = n11376 & n11378;
  assign n11380 = n11248 & n11297;
  assign n11381 = n11379 & n11380;
  assign n11382 = n11369 & n11381;
  assign n11383 = n11334 & n11382;
  assign n11384 = pi0258 & n11383;
  assign n11385 = ~pi0258 & ~n11383;
  assign n11386 = ~n11384 & ~n11385;
  assign n11387 = n10975 & n11386;
  assign n11388 = pi0258 & ~n10975;
  assign n11389 = ~n11387 & ~n11388;
  assign n11390 = ~n10977 & ~n11389;
  assign po0459 = n11368 | n11390;
  assign n11392 = pi0426 & n11155;
  assign n11393 = ~pi1148 & ~n11155;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = n10977 & ~n11394;
  assign n11396 = n11335 & n11369;
  assign n11397 = pi0271 & n11396;
  assign n11398 = pi0258 & n11397;
  assign n11399 = n11246 & n11332;
  assign n11400 = n11398 & n11399;
  assign n11401 = n11249 & n11400;
  assign n11402 = n11299 & n11401;
  assign n11403 = ~pi0259 & n11402;
  assign n11404 = pi0259 & ~n11402;
  assign n11405 = ~n11403 & ~n11404;
  assign n11406 = n10975 & n11405;
  assign n11407 = ~pi0259 & ~n10975;
  assign n11408 = ~n11406 & ~n11407;
  assign n11409 = ~n10977 & ~n11408;
  assign po0460 = n11395 | n11409;
  assign n11411 = pi0428 & n11155;
  assign n11412 = ~pi1187 & ~n11155;
  assign n11413 = ~n11411 & ~n11412;
  assign n11414 = n10977 & ~n11413;
  assign n11415 = ~pi0260 & ~n11166;
  assign n11416 = ~n11167 & ~n11415;
  assign n11417 = n10975 & n11416;
  assign n11418 = pi0260 & ~n10975;
  assign n11419 = ~n11417 & ~n11418;
  assign n11420 = ~n10977 & ~n11419;
  assign po0461 = n11414 | n11420;
  assign n11422 = pi0430 & n11155;
  assign n11423 = ~pi1192 & ~n11155;
  assign n11424 = ~n11422 & ~n11423;
  assign n11425 = n10977 & ~n11424;
  assign n11426 = pi0261 & n11168;
  assign n11427 = ~pi0261 & ~n11168;
  assign n11428 = ~n11426 & ~n11427;
  assign n11429 = n10975 & n11428;
  assign n11430 = pi0261 & ~n10975;
  assign n11431 = ~n11429 & ~n11430;
  assign n11432 = ~n10977 & ~n11431;
  assign po0462 = n11425 | n11432;
  assign n11434 = pi0431 & n11155;
  assign n11435 = ~pi1149 & ~n11155;
  assign n11436 = ~n11434 & ~n11435;
  assign n11437 = n10977 & ~n11436;
  assign n11438 = pi0262 & n11300;
  assign n11439 = ~pi0262 & ~n11300;
  assign n11440 = ~n11438 & ~n11439;
  assign n11441 = n10975 & n11440;
  assign n11442 = pi0262 & ~n10975;
  assign n11443 = ~n11441 & ~n11442;
  assign n11444 = ~n10977 & ~n11443;
  assign po0463 = n11437 | n11444;
  assign n11446 = pi0433 & n11155;
  assign n11447 = ~pi1151 & ~n11155;
  assign n11448 = ~n11446 & ~n11447;
  assign n11449 = n10977 & ~n11448;
  assign n11450 = pi0263 & n11373;
  assign n11451 = ~pi0263 & ~n11373;
  assign n11452 = ~n11450 & ~n11451;
  assign n11453 = n10975 & n11452;
  assign n11454 = pi0263 & ~n10975;
  assign n11455 = ~n11453 & ~n11454;
  assign n11456 = ~n10977 & ~n11455;
  assign po0464 = n11449 | n11456;
  assign n11458 = pi2989 & ~n9404;
  assign n11459 = po3351 & ~n11458;
  assign n11460 = ~pi1692 & n11459;
  assign n11461 = ~pi3179 & po3351;
  assign n11462 = ~n11460 & ~n11461;
  assign n11463 = ~pi0264 & n11462;
  assign n11464 = pi0410 & ~pi2486;
  assign n11465 = pi2486 & pi3334;
  assign n11466 = ~n11464 & ~n11465;
  assign n11467 = ~n11462 & ~n11466;
  assign po0465 = n11463 | n11467;
  assign n11469 = pi0083 & n8309;
  assign n11470 = pi0265 & ~pi0309;
  assign n11471 = ~pi0265 & pi0309;
  assign n11472 = ~n11470 & ~n11471;
  assign n11473 = n11469 & ~n11472;
  assign n11474 = ~pi0265 & ~n11469;
  assign po0466 = n11473 | n11474;
  assign n11476 = ~pi0266 & ~n11469;
  assign po0467 = n11473 | n11476;
  assign n11478 = ~pi0267 & ~n8309;
  assign n11479 = pi0267 & n8309;
  assign po0468 = n11478 | n11479;
  assign n11481 = pi0268 & ~n10975;
  assign n11482 = ~pi0268 & n10975;
  assign n11483 = ~n11481 & ~n11482;
  assign n11484 = ~n10977 & ~n11483;
  assign n11485 = pi0425 & n11155;
  assign n11486 = ~pi1185 & ~n11155;
  assign n11487 = ~n11485 & ~n11486;
  assign n11488 = n10977 & ~n11487;
  assign po0469 = n11484 | n11488;
  assign n11490 = pi0446 & n11155;
  assign n11491 = ~pi1158 & ~n11155;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = n10977 & ~n11492;
  assign n11494 = n11371 & n11378;
  assign n11495 = n11373 & n11494;
  assign n11496 = n11380 & n11495;
  assign n11497 = pi0269 & n11496;
  assign n11498 = ~pi0269 & ~n11496;
  assign n11499 = ~n11497 & ~n11498;
  assign n11500 = n10975 & n11499;
  assign n11501 = pi0269 & ~n10975;
  assign n11502 = ~n11500 & ~n11501;
  assign n11503 = ~n10977 & ~n11502;
  assign po0470 = n11493 | n11503;
  assign n11505 = pi0447 & n11155;
  assign n11506 = ~pi1191 & ~n11155;
  assign n11507 = ~n11505 & ~n11506;
  assign n11508 = n10977 & ~n11507;
  assign n11509 = n11375 & n11494;
  assign n11510 = n11373 & n11509;
  assign n11511 = n11380 & n11510;
  assign n11512 = pi0270 & n11511;
  assign n11513 = ~pi0270 & ~n11511;
  assign n11514 = ~n11512 & ~n11513;
  assign n11515 = n10975 & n11514;
  assign n11516 = pi0270 & ~n10975;
  assign n11517 = ~n11515 & ~n11516;
  assign n11518 = ~n10977 & ~n11517;
  assign po0471 = n11508 | n11518;
  assign n11520 = pi0448 & n11155;
  assign n11521 = ~pi1147 & ~n11155;
  assign n11522 = ~n11520 & ~n11521;
  assign n11523 = n10977 & ~n11522;
  assign n11524 = n11179 & n11351;
  assign n11525 = pi0258 & n11524;
  assign n11526 = pi0257 & n11525;
  assign n11527 = n11206 & n11526;
  assign n11528 = n11175 & n11527;
  assign n11529 = n11162 & n11528;
  assign n11530 = pi0271 & n11529;
  assign n11531 = ~pi0271 & ~n11529;
  assign n11532 = ~n11530 & ~n11531;
  assign n11533 = n10975 & n11532;
  assign n11534 = pi0271 & ~n10975;
  assign n11535 = ~n11533 & ~n11534;
  assign n11536 = ~n10977 & ~n11535;
  assign po0472 = n11523 | n11536;
  assign n11538 = n11175 & n11206;
  assign n11539 = pi0272 & ~n11538;
  assign n11540 = ~pi0272 & n11538;
  assign n11541 = ~n11539 & ~n11540;
  assign n11542 = n10975 & ~n11541;
  assign n11543 = pi0272 & ~n10975;
  assign n11544 = ~n11542 & ~n11543;
  assign n11545 = ~n10977 & ~n11544;
  assign n11546 = pi0415 & n11155;
  assign n11547 = ~pi1157 & ~n11155;
  assign n11548 = ~n11546 & ~n11547;
  assign n11549 = n10977 & ~n11548;
  assign po0473 = n11545 | n11549;
  assign n11551 = ~pi0273 & n11462;
  assign n11552 = ~n9545 & ~n11462;
  assign po0474 = n11551 | n11552;
  assign n11554 = ~pi0274 & n11462;
  assign n11555 = ~n9585 & ~n11462;
  assign po0475 = n11554 | n11555;
  assign n11557 = ~pi0275 & n11462;
  assign n11558 = pi0437 & ~pi2486;
  assign n11559 = pi2486 & pi3292;
  assign n11560 = ~n11558 & ~n11559;
  assign n11561 = ~n11462 & ~n11560;
  assign po0476 = n11557 | n11561;
  assign n11563 = ~pi0276 & n11462;
  assign n11564 = pi0438 & ~pi2486;
  assign n11565 = pi2486 & pi3344;
  assign n11566 = ~n11564 & ~n11565;
  assign n11567 = ~n11462 & ~n11566;
  assign po0477 = n11563 | n11567;
  assign n11569 = ~pi0277 & n11462;
  assign n11570 = pi0439 & ~pi2486;
  assign n11571 = pi2486 & pi3279;
  assign n11572 = ~n11570 & ~n11571;
  assign n11573 = ~n11462 & ~n11572;
  assign po0478 = n11569 | n11573;
  assign n11575 = ~pi0278 & n11462;
  assign n11576 = pi0440 & ~pi2486;
  assign n11577 = pi2486 & pi3329;
  assign n11578 = ~n11576 & ~n11577;
  assign n11579 = ~n11462 & ~n11578;
  assign po0479 = n11575 | n11579;
  assign n11581 = ~pi0279 & n11462;
  assign n11582 = pi0441 & ~pi2486;
  assign n11583 = pi2486 & pi3312;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = ~n11462 & ~n11584;
  assign po0480 = n11581 | n11585;
  assign n11587 = ~pi0280 & n11462;
  assign n11588 = pi0442 & ~pi2486;
  assign n11589 = pi2486 & pi3283;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = ~n11462 & ~n11590;
  assign po0481 = n11587 | n11591;
  assign n11593 = ~pi0281 & n11462;
  assign n11594 = pi0412 & ~pi2486;
  assign n11595 = pi2486 & pi3282;
  assign n11596 = ~n11594 & ~n11595;
  assign n11597 = ~n11462 & ~n11596;
  assign po0482 = n11593 | n11597;
  assign n11599 = ~pi0282 & n11462;
  assign n11600 = pi0414 & ~pi2486;
  assign n11601 = pi2486 & pi3356;
  assign n11602 = ~n11600 & ~n11601;
  assign n11603 = ~n11462 & ~n11602;
  assign po0483 = n11599 | n11603;
  assign n11605 = ~pi0283 & n11462;
  assign n11606 = pi0415 & ~pi2486;
  assign n11607 = pi2486 & pi3272;
  assign n11608 = ~n11606 & ~n11607;
  assign n11609 = ~n11462 & ~n11608;
  assign po0484 = n11605 | n11609;
  assign n11611 = ~pi0284 & n11462;
  assign n11612 = pi0416 & ~pi2486;
  assign n11613 = pi2486 & pi3303;
  assign n11614 = ~n11612 & ~n11613;
  assign n11615 = ~n11462 & ~n11614;
  assign po0485 = n11611 | n11615;
  assign n11617 = ~pi0285 & n11462;
  assign n11618 = pi0418 & ~pi2486;
  assign n11619 = pi2486 & pi3327;
  assign n11620 = ~n11618 & ~n11619;
  assign n11621 = ~n11462 & ~n11620;
  assign po0486 = n11617 | n11621;
  assign n11623 = ~pi0286 & n11462;
  assign n11624 = pi0419 & ~pi2486;
  assign n11625 = pi2486 & pi3305;
  assign n11626 = ~n11624 & ~n11625;
  assign n11627 = ~n11462 & ~n11626;
  assign po0487 = n11623 | n11627;
  assign n11629 = ~pi0287 & n11462;
  assign n11630 = pi0421 & ~pi2486;
  assign n11631 = pi2486 & pi3307;
  assign n11632 = ~n11630 & ~n11631;
  assign n11633 = ~n11462 & ~n11632;
  assign po0488 = n11629 | n11633;
  assign n11635 = ~pi0288 & n11462;
  assign n11636 = pi0422 & ~pi2486;
  assign n11637 = pi2486 & pi3300;
  assign n11638 = ~n11636 & ~n11637;
  assign n11639 = ~n11462 & ~n11638;
  assign po0489 = n11635 | n11639;
  assign n11641 = ~pi0289 & n11462;
  assign n11642 = pi0423 & ~pi2486;
  assign n11643 = pi2486 & pi3306;
  assign n11644 = ~n11642 & ~n11643;
  assign n11645 = ~n11462 & ~n11644;
  assign po0490 = n11641 | n11645;
  assign n11647 = ~pi0290 & n11462;
  assign n11648 = pi0424 & ~pi2486;
  assign n11649 = pi2486 & pi3301;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = ~n11462 & ~n11650;
  assign po0491 = n11647 | n11651;
  assign n11653 = ~pi0291 & n11462;
  assign n11654 = pi0425 & ~pi2486;
  assign n11655 = pi2486 & pi3280;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = ~n11462 & ~n11656;
  assign po0492 = n11653 | n11657;
  assign n11659 = ~pi0292 & n11462;
  assign n11660 = pi0426 & ~pi2486;
  assign n11661 = pi2486 & pi3273;
  assign n11662 = ~n11660 & ~n11661;
  assign n11663 = ~n11462 & ~n11662;
  assign po0493 = n11659 | n11663;
  assign n11665 = ~pi0293 & n11462;
  assign n11666 = pi0427 & ~pi2486;
  assign n11667 = pi2486 & pi3274;
  assign n11668 = ~n11666 & ~n11667;
  assign n11669 = ~n11462 & ~n11668;
  assign po0494 = n11665 | n11669;
  assign n11671 = ~pi0294 & n11462;
  assign n11672 = pi0428 & ~pi2486;
  assign n11673 = pi2486 & pi3275;
  assign n11674 = ~n11672 & ~n11673;
  assign n11675 = ~n11462 & ~n11674;
  assign po0495 = n11671 | n11675;
  assign n11677 = ~pi0295 & n11462;
  assign n11678 = pi0430 & ~pi2486;
  assign n11679 = pi2486 & pi3277;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n11462 & ~n11680;
  assign po0496 = n11677 | n11681;
  assign n11683 = ~pi0296 & n11462;
  assign n11684 = pi0431 & ~pi2486;
  assign n11685 = pi2486 & pi3332;
  assign n11686 = ~n11684 & ~n11685;
  assign n11687 = ~n11462 & ~n11686;
  assign po0497 = n11683 | n11687;
  assign n11689 = ~pi0297 & n11462;
  assign n11690 = pi0432 & ~pi2486;
  assign n11691 = pi2486 & pi3291;
  assign n11692 = ~n11690 & ~n11691;
  assign n11693 = ~n11462 & ~n11692;
  assign po0498 = n11689 | n11693;
  assign n11695 = pi0298 & ~n11374;
  assign n11696 = ~pi0298 & n11374;
  assign n11697 = ~n11695 & ~n11696;
  assign n11698 = n10975 & ~n11697;
  assign n11699 = pi0298 & ~n10975;
  assign n11700 = ~n11698 & ~n11699;
  assign n11701 = ~n10977 & ~n11700;
  assign n11702 = pi0441 & n11155;
  assign n11703 = ~pi1135 & ~n11155;
  assign n11704 = ~n11702 & ~n11703;
  assign n11705 = n10977 & ~n11704;
  assign po0499 = n11701 | n11705;
  assign n11707 = pi0299 & ~n11399;
  assign n11708 = ~pi0299 & n11399;
  assign n11709 = ~n11707 & ~n11708;
  assign n11710 = n10975 & ~n11709;
  assign n11711 = pi0299 & ~n10975;
  assign n11712 = ~n11710 & ~n11711;
  assign n11713 = ~n10977 & ~n11712;
  assign n11714 = pi0412 & n11155;
  assign n11715 = ~pi1136 & ~n11155;
  assign n11716 = ~n11714 & ~n11715;
  assign n11717 = n10977 & ~n11716;
  assign po0500 = n11713 | n11717;
  assign n11719 = n11374 & n11378;
  assign n11720 = pi0300 & ~n11719;
  assign n11721 = ~pi0300 & n11719;
  assign n11722 = ~n11720 & ~n11721;
  assign n11723 = n10975 & ~n11722;
  assign n11724 = pi0300 & ~n10975;
  assign n11725 = ~n11723 & ~n11724;
  assign n11726 = ~n10977 & ~n11725;
  assign n11727 = pi0414 & n11155;
  assign n11728 = ~pi1138 & ~n11155;
  assign n11729 = ~n11727 & ~n11728;
  assign n11730 = n10977 & ~n11729;
  assign po0501 = n11726 | n11730;
  assign n11732 = pi0268 & ~pi0301;
  assign n11733 = ~pi0268 & pi0301;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = n10975 & ~n11734;
  assign n11736 = pi0301 & ~n10975;
  assign n11737 = ~n11735 & ~n11736;
  assign n11738 = ~n10977 & ~n11737;
  assign n11739 = pi0427 & n11155;
  assign n11740 = ~pi1155 & ~n11155;
  assign n11741 = ~n11739 & ~n11740;
  assign n11742 = n10977 & ~n11741;
  assign po0502 = n11738 | n11742;
  assign n11744 = pi0302 & ~n11224;
  assign n11745 = ~pi0302 & n11224;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = n10975 & ~n11746;
  assign n11748 = pi0302 & ~n10975;
  assign n11749 = ~n11747 & ~n11748;
  assign n11750 = ~n10977 & ~n11749;
  assign n11751 = pi0432 & n11155;
  assign n11752 = ~pi1150 & ~n11155;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = n10977 & ~n11753;
  assign po0503 = n11750 | n11754;
  assign n11756 = pi0303 & ~n11169;
  assign n11757 = ~pi0303 & n11169;
  assign n11758 = ~n11756 & ~n11757;
  assign n11759 = n10975 & ~n11758;
  assign n11760 = pi0303 & ~n10975;
  assign n11761 = ~n11759 & ~n11760;
  assign n11762 = ~n10977 & ~n11761;
  assign n11763 = pi0438 & n11155;
  assign n11764 = ~pi1133 & ~n11155;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = n10977 & ~n11765;
  assign po0504 = n11762 | n11766;
  assign n11768 = pi0304 & ~n11225;
  assign n11769 = ~pi0304 & n11225;
  assign n11770 = ~n11768 & ~n11769;
  assign n11771 = n10975 & ~n11770;
  assign n11772 = pi0304 & ~n10975;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = ~n10977 & ~n11773;
  assign n11775 = pi0440 & n11155;
  assign n11776 = ~pi1183 & ~n11155;
  assign n11777 = ~n11775 & ~n11776;
  assign n11778 = n10977 & ~n11777;
  assign po0505 = n11774 | n11778;
  assign n11780 = pi0305 & ~n10977;
  assign n11781 = pi0435 & n11155;
  assign n11782 = ~pi1235 & ~n11155;
  assign n11783 = ~n11781 & ~n11782;
  assign n11784 = n10977 & ~n11783;
  assign po0506 = n11780 | n11784;
  assign n11786 = pi0306 & ~n10977;
  assign n11787 = pi0436 & n11155;
  assign n11788 = ~pi1230 & ~n11155;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = n10977 & ~n11789;
  assign po0507 = n11786 | n11790;
  assign n11792 = pi0307 & ~n10977;
  assign n11793 = pi0434 & n11155;
  assign n11794 = ~pi1310 & ~n11155;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = n10977 & ~n11795;
  assign po0508 = n11792 | n11796;
  assign n11798 = pi0308 & ~n10977;
  assign n11799 = pi0437 & n11155;
  assign n11800 = ~pi1132 & ~n11155;
  assign n11801 = ~n11799 & ~n11800;
  assign n11802 = n10977 & ~n11801;
  assign po0509 = n11798 | n11802;
  assign n11804 = ~pi0309 & ~n11469;
  assign n11805 = pi0309 & n11469;
  assign po0510 = n11804 | n11805;
  assign n11807 = ~pi0310 & ~n11469;
  assign n11808 = ~pi0265 & n11469;
  assign po0511 = n11807 | n11808;
  assign n11810 = pi0267 & ~pi0311;
  assign n11811 = ~pi0267 & pi0311;
  assign n11812 = ~n11810 & ~n11811;
  assign n11813 = n8309 & ~n11812;
  assign n11814 = ~pi0311 & ~n8309;
  assign po0512 = n11813 | n11814;
  assign n11816 = ~pi0267 & ~pi0311;
  assign n11817 = ~pi0312 & ~n11816;
  assign n11818 = pi0312 & n11816;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = n8309 & ~n11819;
  assign n11821 = ~pi0312 & ~n8309;
  assign po0513 = n11820 | n11821;
  assign n11823 = ~pi0321 & n8309;
  assign n11824 = pi0313 & ~n8309;
  assign po0514 = n11823 | n11824;
  assign n11826 = ~pi0322 & n8309;
  assign n11827 = pi0314 & ~n8309;
  assign po0515 = n11826 | n11827;
  assign n11829 = ~pi0323 & n8309;
  assign n11830 = pi0315 & ~n8309;
  assign po0516 = n11829 | n11830;
  assign n11832 = pi0313 & n8309;
  assign n11833 = ~pi0316 & ~n8309;
  assign po0517 = n11832 | n11833;
  assign n11835 = pi0315 & n8309;
  assign n11836 = ~pi0317 & ~n8309;
  assign po0518 = n11835 | n11836;
  assign n11838 = ~pi0316 & n8309;
  assign n11839 = ~pi0318 & ~n8309;
  assign po0519 = n11838 | n11839;
  assign n11841 = ~pi0324 & n8309;
  assign n11842 = ~pi0319 & ~n8309;
  assign po0520 = n11841 | n11842;
  assign n11844 = ~pi0317 & n8309;
  assign n11845 = ~pi0320 & ~n8309;
  assign po0521 = n11844 | n11845;
  assign n11847 = ~pi0335 & pi0337;
  assign n11848 = pi0335 & ~pi0337;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = n8309 & ~n11849;
  assign n11851 = ~pi0321 & ~n8309;
  assign po0522 = n11850 | n11851;
  assign n11853 = pi0337 & ~pi0338;
  assign n11854 = ~pi0337 & pi0338;
  assign n11855 = ~n11853 & ~n11854;
  assign n11856 = n8309 & ~n11855;
  assign n11857 = ~pi0322 & ~n8309;
  assign po0523 = n11856 | n11857;
  assign n11859 = ~pi0338 & n8309;
  assign n11860 = ~pi0323 & ~n8309;
  assign po0524 = n11859 | n11860;
  assign n11862 = pi0314 & n8309;
  assign n11863 = ~pi0324 & ~n8309;
  assign po0525 = n11862 | n11863;
  assign n11865 = pi0325 & ~n11332;
  assign n11866 = ~pi0325 & n11332;
  assign n11867 = ~n11865 & ~n11866;
  assign n11868 = n10975 & ~n11867;
  assign n11869 = pi0325 & ~n10975;
  assign n11870 = ~n11868 & ~n11869;
  assign n11871 = ~n10977 & ~n11870;
  assign n11872 = pi0439 & n11155;
  assign n11873 = ~pi1134 & ~n11155;
  assign n11874 = ~n11872 & ~n11873;
  assign n11875 = n10977 & ~n11874;
  assign po0526 = n11871 | n11875;
  assign n11877 = pi0326 & ~n10977;
  assign n11878 = pi0417 & n11155;
  assign n11879 = ~pi1140 & ~n11155;
  assign n11880 = ~n11878 & ~n11879;
  assign n11881 = n10977 & ~n11880;
  assign po0527 = n11877 | n11881;
  assign n11883 = ~pi0327 & n11462;
  assign n11884 = pi0429 & ~pi2486;
  assign n11885 = pi2486 & pi3310;
  assign n11886 = ~n11884 & ~n11885;
  assign n11887 = ~n11462 & ~n11886;
  assign po0528 = n11883 | n11887;
  assign n11889 = ~pi0328 & n11462;
  assign n11890 = pi0433 & ~pi2486;
  assign n11891 = pi2486 & pi3357;
  assign n11892 = ~n11890 & ~n11891;
  assign n11893 = ~n11462 & ~n11892;
  assign po0529 = n11889 | n11893;
  assign n11895 = ~pi0329 & n11462;
  assign n11896 = pi0417 & ~pi2486;
  assign n11897 = pi2486 & pi3281;
  assign n11898 = ~n11896 & ~n11897;
  assign n11899 = ~n11462 & ~n11898;
  assign po0530 = n11895 | n11899;
  assign n11901 = ~pi0330 & n11462;
  assign n11902 = pi0420 & ~pi2486;
  assign n11903 = pi2486 & pi3304;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = ~n11462 & ~n11904;
  assign po0531 = n11901 | n11905;
  assign n11907 = ~pi0331 & n11462;
  assign n11908 = pi0413 & ~pi2486;
  assign n11909 = pi2486 & pi3278;
  assign n11910 = ~n11908 & ~n11909;
  assign n11911 = ~n11462 & ~n11910;
  assign po0532 = n11907 | n11911;
  assign n11913 = ~pi0332 & n11462;
  assign n11914 = ~n9563 & ~n11462;
  assign po0533 = n11913 | n11914;
  assign n11916 = ~pi0333 & n11462;
  assign n11917 = pi0446 & ~pi2486;
  assign n11918 = pi2486 & pi3294;
  assign n11919 = ~n11917 & ~n11918;
  assign n11920 = ~n11462 & ~n11919;
  assign po0534 = n11916 | n11920;
  assign n11922 = ~pi0334 & n11462;
  assign n11923 = pi0447 & ~pi2486;
  assign n11924 = pi2486 & pi3276;
  assign n11925 = ~n11923 & ~n11924;
  assign n11926 = ~n11462 & ~n11925;
  assign po0535 = n11922 | n11926;
  assign po0537 = ~po1399 & n7176;
  assign po0540 = ~po1399 & ~n7263;
  assign n11930 = ~n8193 & n8198;
  assign n11931 = ~n8188 & n11930;
  assign n11932 = ~n8189 & ~n8201;
  assign n11933 = n8206 & n11932;
  assign n11934 = n11931 & n11933;
  assign n11935 = n8200 & n8229;
  assign n11936 = ~n8224 & n11935;
  assign n11937 = n8187 & n11936;
  assign n11938 = ~n11934 & ~n11937;
  assign n11939 = ~n8224 & ~n11938;
  assign n11940 = ~pi1162 & n11939;
  assign n11941 = ~pi1131 & ~n11939;
  assign n11942 = ~n11940 & ~n11941;
  assign n11943 = pi1129 & n11939;
  assign n11944 = pi1128 & ~n11939;
  assign n11945 = ~n11943 & ~n11944;
  assign n11946 = ~n11942 & ~n11945;
  assign n11947 = ~n8193 & n8199;
  assign n11948 = n11932 & n11947;
  assign n11949 = ~n8204 & n11948;
  assign n11950 = ~n8205 & n11949;
  assign n11951 = ~n11937 & ~n11950;
  assign n11952 = ~n8224 & ~n11951;
  assign n11953 = ~pi1177 & n11952;
  assign n11954 = ~pi1130 & ~n11952;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = ~pi1181 & ~n11952;
  assign n11957 = ~pi1179 & n11939;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = n11955 & ~n11958;
  assign n11960 = n11946 & n11959;
  assign n11961 = ~pi1952 & n11960;
  assign n11962 = ~n11955 & ~n11958;
  assign n11963 = n11946 & n11962;
  assign n11964 = ~pi2224 & n11963;
  assign n11965 = ~n11961 & ~n11964;
  assign n11966 = ~pi1129 & n11939;
  assign n11967 = ~pi1128 & ~n11939;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = pi1162 & n11939;
  assign n11970 = pi1131 & ~n11939;
  assign n11971 = ~n11969 & ~n11970;
  assign n11972 = ~n11968 & ~n11971;
  assign n11973 = n11959 & n11972;
  assign n11974 = ~pi2333 & n11973;
  assign n11975 = ~n11945 & ~n11971;
  assign n11976 = n11962 & n11975;
  assign n11977 = ~pi1991 & n11976;
  assign n11978 = ~n11974 & ~n11977;
  assign n11979 = ~n11955 & n11958;
  assign n11980 = n11946 & n11979;
  assign n11981 = ~pi2125 & n11980;
  assign n11982 = ~n11942 & ~n11968;
  assign n11983 = n11979 & n11982;
  assign n11984 = ~pi2204 & n11983;
  assign n11985 = ~n11981 & ~n11984;
  assign n11986 = n11978 & n11985;
  assign n11987 = n11955 & n11958;
  assign n11988 = n11975 & n11987;
  assign n11989 = ~pi1988 & n11988;
  assign n11990 = n11946 & n11987;
  assign n11991 = ~pi2088 & n11990;
  assign n11992 = ~n11989 & ~n11991;
  assign n11993 = n11959 & n11982;
  assign n11994 = ~pi2175 & n11993;
  assign n11995 = n11962 & n11982;
  assign n11996 = ~pi1927 & n11995;
  assign n11997 = ~n11994 & ~n11996;
  assign n11998 = n11992 & n11997;
  assign n11999 = n11986 & n11998;
  assign n12000 = n11965 & n11999;
  assign n12001 = n11959 & n11975;
  assign n12002 = ~pi2133 & n12001;
  assign n12003 = n11962 & n11972;
  assign n12004 = ~pi2231 & n12003;
  assign n12005 = n11972 & n11979;
  assign n12006 = ~pi2270 & n12005;
  assign n12007 = n11982 & n11987;
  assign n12008 = ~pi2389 & n12007;
  assign n12009 = ~n12006 & ~n12008;
  assign n12010 = ~n12004 & n12009;
  assign n12011 = ~n12002 & n12010;
  assign n12012 = n11972 & n11987;
  assign n12013 = ~pi2426 & n12012;
  assign n12014 = n11975 & n11979;
  assign n12015 = ~pi2059 & n12014;
  assign n12016 = ~n12013 & ~n12015;
  assign n12017 = n12011 & n12016;
  assign po0541 = ~n12000 | ~n12017;
  assign n12019 = ~pi2040 & n12012;
  assign n12020 = ~pi2334 & n12014;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = ~pi2459 & n11973;
  assign n12023 = ~pi2007 & n11976;
  assign n12024 = ~n12022 & ~n12023;
  assign n12025 = ~pi1929 & n11995;
  assign n12026 = ~pi2455 & n11993;
  assign n12027 = ~n12025 & ~n12026;
  assign n12028 = n12024 & n12027;
  assign n12029 = ~pi2356 & n11988;
  assign n12030 = ~pi2354 & n11990;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = ~pi2300 & n11980;
  assign n12033 = ~pi2439 & n11983;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = n12031 & n12034;
  assign n12036 = n12028 & n12035;
  assign n12037 = n12021 & n12036;
  assign n12038 = ~pi2375 & n12001;
  assign n12039 = ~pi2229 & n12003;
  assign n12040 = ~pi2271 & n12005;
  assign n12041 = ~pi2108 & n12007;
  assign n12042 = ~n12040 & ~n12041;
  assign n12043 = ~n12039 & n12042;
  assign n12044 = ~n12038 & n12043;
  assign n12045 = ~pi2023 & n11960;
  assign n12046 = ~pi2233 & n11963;
  assign n12047 = ~n12045 & ~n12046;
  assign n12048 = n12044 & n12047;
  assign po0542 = ~n12037 | ~n12048;
  assign n12050 = ~pi2387 & n12007;
  assign n12051 = ~pi2320 & n11980;
  assign n12052 = ~pi2437 & n11983;
  assign n12053 = ~n12051 & ~n12052;
  assign n12054 = ~pi1940 & n12005;
  assign n12055 = ~pi1992 & n11988;
  assign n12056 = ~pi2092 & n11990;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = ~n12054 & n12057;
  assign n12059 = n12053 & n12058;
  assign n12060 = ~n12050 & n12059;
  assign n12061 = ~pi1916 & n11995;
  assign n12062 = ~pi2478 & n11993;
  assign n12063 = ~n12061 & ~n12062;
  assign n12064 = ~pi2269 & n11973;
  assign n12065 = ~pi1948 & n11976;
  assign n12066 = ~n12064 & ~n12065;
  assign n12067 = n12063 & n12066;
  assign n12068 = n12060 & n12067;
  assign n12069 = ~pi2424 & n12012;
  assign n12070 = ~pi2063 & n12014;
  assign n12071 = ~n12069 & ~n12070;
  assign n12072 = ~pi2136 & n12001;
  assign n12073 = ~pi2212 & n12003;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = n12071 & n12074;
  assign n12076 = ~pi1949 & n11960;
  assign n12077 = ~pi2234 & n11963;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = n12075 & n12078;
  assign po0543 = ~n12068 | ~n12079;
  assign n12081 = ~pi2194 & n11995;
  assign n12082 = ~pi2466 & n11993;
  assign n12083 = ~n12081 & ~n12082;
  assign n12084 = ~pi2307 & n11980;
  assign n12085 = ~pi2206 & n11983;
  assign n12086 = ~n12084 & ~n12085;
  assign n12087 = n12083 & n12086;
  assign n12088 = ~pi2280 & n11973;
  assign n12089 = ~pi1958 & n11976;
  assign n12090 = ~n12088 & ~n12089;
  assign n12091 = ~pi1993 & n11988;
  assign n12092 = ~pi2093 & n11990;
  assign n12093 = ~n12091 & ~n12092;
  assign n12094 = n12090 & n12093;
  assign n12095 = n12087 & n12094;
  assign n12096 = ~pi2028 & n11960;
  assign n12097 = ~pi2236 & n11963;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = n12095 & n12098;
  assign n12100 = ~pi2044 & n12012;
  assign n12101 = ~pi2359 & n12014;
  assign n12102 = ~n12100 & ~n12101;
  assign n12103 = ~pi2345 & n12005;
  assign n12104 = ~pi2113 & n12007;
  assign n12105 = ~n12103 & ~n12104;
  assign n12106 = n12102 & n12105;
  assign n12107 = ~pi2137 & n12001;
  assign n12108 = ~pi2213 & n12003;
  assign n12109 = ~n12107 & ~n12108;
  assign n12110 = n12106 & n12109;
  assign po0544 = ~n12099 | ~n12110;
  assign n12112 = ~pi1912 & n11995;
  assign n12113 = ~pi2472 & n11993;
  assign n12114 = ~n12112 & ~n12113;
  assign n12115 = ~pi2138 & n12001;
  assign n12116 = n12114 & ~n12115;
  assign n12117 = ~pi2168 & n12003;
  assign n12118 = ~pi2256 & n11973;
  assign n12119 = ~pi2011 & n11976;
  assign n12120 = ~n12118 & ~n12119;
  assign n12121 = ~pi2319 & n11988;
  assign n12122 = ~pi2094 & n11990;
  assign n12123 = ~n12121 & ~n12122;
  assign n12124 = ~pi2312 & n11980;
  assign n12125 = ~pi2428 & n11983;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = n12123 & n12126;
  assign n12128 = n12120 & n12127;
  assign n12129 = ~n12117 & n12128;
  assign n12130 = n12116 & n12129;
  assign n12131 = ~pi2045 & n12012;
  assign n12132 = ~pi2366 & n12014;
  assign n12133 = ~n12131 & ~n12132;
  assign n12134 = ~pi2074 & n12005;
  assign n12135 = ~pi2114 & n12007;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = n12133 & n12136;
  assign n12138 = ~pi2029 & n11960;
  assign n12139 = ~pi2186 & n11963;
  assign n12140 = ~n12138 & ~n12139;
  assign n12141 = n12137 & n12140;
  assign po0545 = ~n12130 | ~n12141;
  assign n12143 = ~pi2139 & n12001;
  assign n12144 = ~pi2218 & n12003;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = ~pi2262 & n11973;
  assign n12147 = ~pi1964 & n11976;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = ~pi2127 & n11980;
  assign n12150 = ~pi2207 & n11983;
  assign n12151 = ~n12149 & ~n12150;
  assign n12152 = n12148 & n12151;
  assign n12153 = ~pi2195 & n11995;
  assign n12154 = ~pi2177 & n11993;
  assign n12155 = ~n12153 & ~n12154;
  assign n12156 = ~pi1994 & n11988;
  assign n12157 = ~pi2095 & n11990;
  assign n12158 = ~n12156 & ~n12157;
  assign n12159 = n12155 & n12158;
  assign n12160 = n12152 & n12159;
  assign n12161 = n12145 & n12160;
  assign n12162 = ~pi1944 & n11960;
  assign n12163 = ~pi2219 & n11963;
  assign n12164 = ~pi2337 & n12005;
  assign n12165 = ~pi2362 & n12007;
  assign n12166 = ~n12164 & ~n12165;
  assign n12167 = ~n12163 & n12166;
  assign n12168 = ~n12162 & n12167;
  assign n12169 = ~pi2420 & n12012;
  assign n12170 = ~pi2064 & n12014;
  assign n12171 = ~n12169 & ~n12170;
  assign n12172 = n12168 & n12171;
  assign po0546 = ~n12161 | ~n12172;
  assign n12174 = ~pi2412 & n12012;
  assign n12175 = ~pi2348 & n12014;
  assign n12176 = ~n12174 & ~n12175;
  assign n12177 = ~pi2457 & n11995;
  assign n12178 = ~pi2458 & n11993;
  assign n12179 = ~n12177 & ~n12178;
  assign n12180 = ~pi2128 & n11980;
  assign n12181 = ~pi2421 & n11983;
  assign n12182 = ~n12180 & ~n12181;
  assign n12183 = n12179 & n12182;
  assign n12184 = ~pi2265 & n11973;
  assign n12185 = ~pi1961 & n11976;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = ~pi1995 & n11988;
  assign n12188 = ~pi2096 & n11990;
  assign n12189 = ~n12187 & ~n12188;
  assign n12190 = n12186 & n12189;
  assign n12191 = n12183 & n12190;
  assign n12192 = n12176 & n12191;
  assign n12193 = ~pi2031 & n11960;
  assign n12194 = ~pi2230 & n11963;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 = ~pi2140 & n12001;
  assign n12197 = ~pi2216 & n12003;
  assign n12198 = ~n12196 & ~n12197;
  assign n12199 = n12195 & n12198;
  assign n12200 = ~pi2400 & n12005;
  assign n12201 = ~pi2116 & n12007;
  assign n12202 = ~n12200 & ~n12201;
  assign n12203 = n12199 & n12202;
  assign po0547 = ~n12192 | ~n12203;
  assign n12205 = ~pi2047 & n12012;
  assign n12206 = ~pi2350 & n12014;
  assign n12207 = ~n12205 & ~n12206;
  assign n12208 = ~pi2266 & n11973;
  assign n12209 = ~pi2013 & n11976;
  assign n12210 = ~n12208 & ~n12209;
  assign n12211 = ~pi2464 & n11995;
  assign n12212 = ~pi2453 & n11993;
  assign n12213 = ~n12211 & ~n12212;
  assign n12214 = n12210 & n12213;
  assign n12215 = ~pi2316 & n11988;
  assign n12216 = ~pi2097 & n11990;
  assign n12217 = ~n12215 & ~n12216;
  assign n12218 = ~pi2247 & n11980;
  assign n12219 = ~pi2422 & n11983;
  assign n12220 = ~n12218 & ~n12219;
  assign n12221 = n12217 & n12220;
  assign n12222 = n12214 & n12221;
  assign n12223 = n12207 & n12222;
  assign n12224 = ~pi2032 & n11960;
  assign n12225 = ~pi2188 & n11963;
  assign n12226 = ~n12224 & ~n12225;
  assign n12227 = ~pi1957 & n12001;
  assign n12228 = ~pi2215 & n12003;
  assign n12229 = ~n12227 & ~n12228;
  assign n12230 = n12226 & n12229;
  assign n12231 = ~pi2076 & n12005;
  assign n12232 = ~pi2117 & n12007;
  assign n12233 = ~n12231 & ~n12232;
  assign n12234 = n12230 & n12233;
  assign po0548 = ~n12223 | ~n12234;
  assign n12236 = ~pi2408 & n12012;
  assign n12237 = ~pi2067 & n12014;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = ~pi2200 & n11995;
  assign n12240 = ~pi2410 & n11993;
  assign n12241 = ~n12239 & ~n12240;
  assign n12242 = ~pi2002 & n11988;
  assign n12243 = ~pi2103 & n11990;
  assign n12244 = ~n12242 & ~n12243;
  assign n12245 = ~pi2131 & n11980;
  assign n12246 = ~pi2364 & n11983;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = n12244 & n12247;
  assign n12249 = ~pi2259 & n11973;
  assign n12250 = ~pi2017 & n11976;
  assign n12251 = ~n12249 & ~n12250;
  assign n12252 = n12248 & n12251;
  assign n12253 = n12241 & n12252;
  assign n12254 = n12238 & n12253;
  assign n12255 = ~pi2409 & n11960;
  assign n12256 = ~pi2214 & n11963;
  assign n12257 = ~n12255 & ~n12256;
  assign n12258 = ~pi2081 & n12005;
  assign n12259 = ~pi2360 & n12007;
  assign n12260 = ~n12258 & ~n12259;
  assign n12261 = n12257 & n12260;
  assign n12262 = ~pi2302 & n12001;
  assign n12263 = ~pi1920 & n12003;
  assign n12264 = ~n12262 & ~n12263;
  assign n12265 = n12261 & n12264;
  assign po0549 = ~n12254 | ~n12265;
  assign n12267 = ~pi2036 & n11960;
  assign n12268 = ~pi2192 & n11963;
  assign n12269 = ~n12267 & ~n12268;
  assign n12270 = ~pi2250 & n11988;
  assign n12271 = ~pi2249 & n11990;
  assign n12272 = ~n12270 & ~n12271;
  assign n12273 = ~pi2385 & n11980;
  assign n12274 = ~pi2286 & n11983;
  assign n12275 = ~n12273 & ~n12274;
  assign n12276 = n12272 & n12275;
  assign n12277 = ~pi2153 & n11973;
  assign n12278 = ~pi2020 & n11976;
  assign n12279 = ~n12277 & ~n12278;
  assign n12280 = ~pi2278 & n11993;
  assign n12281 = ~pi2448 & n11995;
  assign n12282 = ~n12280 & ~n12281;
  assign n12283 = n12279 & n12282;
  assign n12284 = n12276 & n12283;
  assign n12285 = n12269 & n12284;
  assign n12286 = ~pi2248 & n12001;
  assign n12287 = ~pi2173 & n12003;
  assign n12288 = ~pi2084 & n12005;
  assign n12289 = ~pi2351 & n12007;
  assign n12290 = ~n12288 & ~n12289;
  assign n12291 = ~n12287 & n12290;
  assign n12292 = ~n12286 & n12291;
  assign n12293 = ~pi2055 & n12012;
  assign n12294 = ~pi2304 & n12014;
  assign n12295 = ~n12293 & ~n12294;
  assign n12296 = n12292 & n12295;
  assign po0550 = ~n12285 | ~n12296;
  assign n12298 = ~pi2361 & n12005;
  assign n12299 = ~pi2346 & n12007;
  assign n12300 = ~n12298 & ~n12299;
  assign n12301 = ~pi2154 & n11973;
  assign n12302 = ~pi1939 & n11976;
  assign n12303 = ~n12301 & ~n12302;
  assign n12304 = ~pi2332 & n11980;
  assign n12305 = ~pi2211 & n11983;
  assign n12306 = ~n12304 & ~n12305;
  assign n12307 = n12303 & n12306;
  assign n12308 = ~pi2004 & n11988;
  assign n12309 = ~pi2105 & n11990;
  assign n12310 = ~n12308 & ~n12309;
  assign n12311 = ~pi2443 & n11995;
  assign n12312 = ~pi2183 & n11993;
  assign n12313 = ~n12311 & ~n12312;
  assign n12314 = n12310 & n12313;
  assign n12315 = n12307 & n12314;
  assign n12316 = n12300 & n12315;
  assign n12317 = ~pi2433 & n11960;
  assign n12318 = ~pi1905 & n11963;
  assign n12319 = ~n12317 & ~n12318;
  assign n12320 = ~pi2253 & n12001;
  assign n12321 = ~pi1913 & n12003;
  assign n12322 = ~n12320 & ~n12321;
  assign n12323 = n12319 & n12322;
  assign n12324 = ~pi2069 & n12014;
  assign n12325 = ~pi2056 & n12012;
  assign n12326 = ~n12324 & ~n12325;
  assign n12327 = n12323 & n12326;
  assign po0551 = ~n12316 | ~n12327;
  assign n12329 = ~pi0352 & n11462;
  assign n12330 = pi0448 & ~pi2486;
  assign n12331 = pi2486 & pi3358;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = ~n11462 & ~n12332;
  assign po0552 = n12329 | n12333;
  assign n12335 = ~pi2073 & n12005;
  assign n12336 = ~pi2111 & n12007;
  assign n12337 = ~n12335 & ~n12336;
  assign n12338 = ~pi2042 & n12012;
  assign n12339 = ~pi2379 & n12014;
  assign n12340 = ~n12338 & ~n12339;
  assign n12341 = n12337 & n12340;
  assign n12342 = ~pi2026 & n11960;
  assign n12343 = ~pi2239 & n11963;
  assign n12344 = ~n12342 & ~n12343;
  assign n12345 = ~pi2368 & n12001;
  assign n12346 = ~pi2167 & n12003;
  assign n12347 = ~n12345 & ~n12346;
  assign n12348 = n12344 & n12347;
  assign n12349 = ~pi2275 & n11988;
  assign n12350 = ~pi2091 & n11990;
  assign n12351 = ~n12349 & ~n12350;
  assign n12352 = ~pi2281 & n11973;
  assign n12353 = ~pi2009 & n11976;
  assign n12354 = ~n12352 & ~n12353;
  assign n12355 = n12351 & n12354;
  assign n12356 = ~pi2477 & n11993;
  assign n12357 = ~pi1914 & n11995;
  assign n12358 = ~n12356 & ~n12357;
  assign n12359 = n12355 & n12358;
  assign n12360 = ~pi2314 & n11980;
  assign n12361 = ~pi2435 & n11983;
  assign n12362 = ~n12360 & ~n12361;
  assign n12363 = n12359 & n12362;
  assign n12364 = n12348 & n12363;
  assign po0553 = ~n12341 | ~n12364;
  assign n12366 = ~pi2048 & n12012;
  assign n12367 = ~pi2274 & n12014;
  assign n12368 = ~n12366 & ~n12367;
  assign n12369 = ~pi2305 & n12001;
  assign n12370 = ~pi2170 & n12003;
  assign n12371 = ~n12369 & ~n12370;
  assign n12372 = n12368 & n12371;
  assign n12373 = ~pi2078 & n12005;
  assign n12374 = ~pi2118 & n12007;
  assign n12375 = ~n12373 & ~n12374;
  assign n12376 = ~pi2033 & n11960;
  assign n12377 = ~pi2226 & n11963;
  assign n12378 = ~n12376 & ~n12377;
  assign n12379 = n12375 & n12378;
  assign n12380 = ~pi1997 & n11988;
  assign n12381 = ~pi2321 & n11990;
  assign n12382 = ~n12380 & ~n12381;
  assign n12383 = ~pi2147 & n11973;
  assign n12384 = ~pi2014 & n11976;
  assign n12385 = ~n12383 & ~n12384;
  assign n12386 = n12382 & n12385;
  assign n12387 = ~pi2085 & n11980;
  assign n12388 = ~pi2418 & n11983;
  assign n12389 = ~n12387 & ~n12388;
  assign n12390 = n12386 & n12389;
  assign n12391 = ~pi2456 & n11993;
  assign n12392 = ~pi2473 & n11995;
  assign n12393 = ~n12391 & ~n12392;
  assign n12394 = n12390 & n12393;
  assign n12395 = n12379 & n12394;
  assign po0554 = ~n12372 | ~n12395;
  assign n12397 = ~pi2264 & n11973;
  assign n12398 = ~pi2049 & n12012;
  assign n12399 = ~pi2299 & n12014;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = ~n12397 & n12400;
  assign n12402 = ~pi1921 & n12003;
  assign n12403 = ~pi2142 & n12001;
  assign n12404 = ~n12402 & ~n12403;
  assign n12405 = ~pi1945 & n11960;
  assign n12406 = ~pi2399 & n11993;
  assign n12407 = ~pi2196 & n11995;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = ~pi1954 & n11976;
  assign n12410 = ~pi2227 & n11963;
  assign n12411 = ~n12409 & ~n12410;
  assign n12412 = n12408 & n12411;
  assign n12413 = ~n12405 & n12412;
  assign n12414 = n12404 & n12413;
  assign n12415 = ~pi2390 & n12005;
  assign n12416 = ~pi2378 & n12007;
  assign n12417 = ~n12415 & ~n12416;
  assign n12418 = ~pi1998 & n11988;
  assign n12419 = ~pi2099 & n11990;
  assign n12420 = ~n12418 & ~n12419;
  assign n12421 = ~pi1936 & n11980;
  assign n12422 = ~pi2415 & n11983;
  assign n12423 = ~n12421 & ~n12422;
  assign n12424 = n12420 & n12423;
  assign n12425 = n12417 & n12424;
  assign n12426 = n12414 & n12425;
  assign po0555 = ~n12401 | ~n12426;
  assign n12428 = ~pi1941 & n11960;
  assign n12429 = ~pi2222 & n11963;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = ~pi2402 & n12012;
  assign n12432 = ~pi2065 & n12014;
  assign n12433 = ~n12431 & ~n12432;
  assign n12434 = ~pi2322 & n12001;
  assign n12435 = ~pi1962 & n12003;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = n12433 & n12436;
  assign n12438 = ~pi2339 & n12005;
  assign n12439 = ~pi2373 & n12007;
  assign n12440 = ~n12438 & ~n12439;
  assign n12441 = n12437 & n12440;
  assign n12442 = ~pi1999 & n11988;
  assign n12443 = ~pi2100 & n11990;
  assign n12444 = ~pi2130 & n11980;
  assign n12445 = ~pi2394 & n11983;
  assign n12446 = ~n12444 & ~n12445;
  assign n12447 = ~n12443 & n12446;
  assign n12448 = ~n12442 & n12447;
  assign n12449 = ~pi2197 & n11995;
  assign n12450 = ~pi2180 & n11993;
  assign n12451 = ~pi2255 & n11973;
  assign n12452 = ~pi1959 & n11976;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = ~n12450 & n12453;
  assign n12455 = ~n12449 & n12454;
  assign n12456 = n12448 & n12455;
  assign n12457 = n12441 & n12456;
  assign po0556 = ~n12430 | ~n12457;
  assign n12459 = ~pi2315 & n12001;
  assign n12460 = ~pi1931 & n12003;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = ~pi2034 & n11960;
  assign n12463 = ~pi2189 & n11963;
  assign n12464 = ~n12462 & ~n12463;
  assign n12465 = n12461 & n12464;
  assign n12466 = ~pi2082 & n12005;
  assign n12467 = ~pi2122 & n12007;
  assign n12468 = ~n12466 & ~n12467;
  assign n12469 = ~pi2052 & n12012;
  assign n12470 = ~pi2327 & n12014;
  assign n12471 = ~n12469 & ~n12470;
  assign n12472 = n12468 & n12471;
  assign n12473 = ~pi2277 & n11988;
  assign n12474 = ~pi2102 & n11990;
  assign n12475 = ~n12473 & ~n12474;
  assign n12476 = ~pi2151 & n11973;
  assign n12477 = ~pi2018 & n11976;
  assign n12478 = ~n12476 & ~n12477;
  assign n12479 = n12475 & n12478;
  assign n12480 = ~pi2450 & n11993;
  assign n12481 = ~pi2413 & n11995;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = n12479 & n12482;
  assign n12484 = ~pi2382 & n11980;
  assign n12485 = ~pi2406 & n11983;
  assign n12486 = ~n12484 & ~n12485;
  assign n12487 = n12483 & n12486;
  assign n12488 = n12472 & n12487;
  assign po0557 = ~n12465 | ~n12488;
  assign n12490 = ~pi2159 & n12005;
  assign n12491 = ~pi2160 & n12007;
  assign n12492 = ~n12490 & ~n12491;
  assign n12493 = ~pi2468 & n11960;
  assign n12494 = ~pi2217 & n11963;
  assign n12495 = ~pi2297 & n12001;
  assign n12496 = ~pi1928 & n12003;
  assign n12497 = ~n12495 & ~n12496;
  assign n12498 = ~n12494 & n12497;
  assign n12499 = ~n12493 & n12498;
  assign n12500 = ~pi2202 & n12012;
  assign n12501 = ~pi2441 & n12014;
  assign n12502 = ~n12500 & ~n12501;
  assign n12503 = n12499 & n12502;
  assign n12504 = ~pi2165 & n11988;
  assign n12505 = ~pi2203 & n11990;
  assign n12506 = ~pi2201 & n11995;
  assign n12507 = ~pi2393 & n11993;
  assign n12508 = ~n12506 & ~n12507;
  assign n12509 = ~n12505 & n12508;
  assign n12510 = ~n12504 & n12509;
  assign n12511 = ~pi2475 & n11980;
  assign n12512 = ~pi2210 & n11983;
  assign n12513 = ~pi2161 & n11973;
  assign n12514 = ~pi2474 & n11976;
  assign n12515 = ~n12513 & ~n12514;
  assign n12516 = ~n12512 & n12515;
  assign n12517 = ~n12511 & n12516;
  assign n12518 = n12510 & n12517;
  assign n12519 = n12503 & n12518;
  assign po0558 = ~n12492 | ~n12519;
  assign n12521 = ~pi1836 & n12005;
  assign n12522 = ~pi1842 & n12007;
  assign n12523 = ~n12521 & ~n12522;
  assign n12524 = ~pi1831 & n11960;
  assign n12525 = ~pi1833 & n11963;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = n12523 & n12526;
  assign n12528 = ~pi1834 & n12012;
  assign n12529 = ~pi1835 & n12014;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = ~pi1839 & n12001;
  assign n12532 = ~pi1830 & n12003;
  assign n12533 = ~n12531 & ~n12532;
  assign n12534 = n12530 & n12533;
  assign n12535 = ~pi1841 & n11988;
  assign n12536 = ~pi1837 & n11990;
  assign n12537 = ~pi1840 & n11973;
  assign n12538 = ~pi1829 & n11976;
  assign n12539 = ~n12537 & ~n12538;
  assign n12540 = ~n12536 & n12539;
  assign n12541 = ~n12535 & n12540;
  assign n12542 = ~pi1844 & n11995;
  assign n12543 = ~pi1832 & n11993;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = n12541 & n12544;
  assign n12546 = ~pi1843 & n11980;
  assign n12547 = ~pi1838 & n11983;
  assign n12548 = ~n12546 & ~n12547;
  assign n12549 = n12545 & n12548;
  assign n12550 = n12534 & n12549;
  assign po0559 = ~n12527 | ~n12550;
  assign n12552 = pi2553 & ~pi2984;
  assign n12553 = ~pi3042 & n9371;
  assign n12554 = n12552 & n12553;
  assign n12555 = ~pi2969 & n12554;
  assign n12556 = pi2963 & n12555;
  assign po3339 = pi2943 & ~pi3123;
  assign n12558 = pi3167 & po3339;
  assign n12559 = pi2963 & ~n8036;
  assign n12560 = ~pi2969 & n8046;
  assign n12561 = n12559 & n12560;
  assign n12562 = n12552 & n12561;
  assign n12563 = ~n12558 & ~n12562;
  assign n12564 = ~n12556 & n12563;
  assign n12565 = pi0360 & n12564;
  assign n12566 = n8058 & ~n12564;
  assign po0560 = n12565 | n12566;
  assign n12568 = ~pi2381 & n12001;
  assign n12569 = ~pi2228 & n12003;
  assign n12570 = ~n12568 & ~n12569;
  assign n12571 = ~pi2039 & n12012;
  assign n12572 = ~pi2392 & n12014;
  assign n12573 = ~n12571 & ~n12572;
  assign n12574 = n12570 & n12573;
  assign n12575 = ~pi2072 & n12005;
  assign n12576 = ~pi2107 & n12007;
  assign n12577 = ~n12575 & ~n12576;
  assign n12578 = ~pi2022 & n11960;
  assign n12579 = ~pi2185 & n11963;
  assign n12580 = ~n12578 & ~n12579;
  assign n12581 = n12577 & n12580;
  assign n12582 = ~pi2145 & n11973;
  assign n12583 = ~pi2006 & n11976;
  assign n12584 = ~pi2288 & n11980;
  assign n12585 = ~pi2440 & n11983;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = ~n12583 & n12586;
  assign n12588 = ~n12582 & n12587;
  assign n12589 = ~pi1987 & n11988;
  assign n12590 = ~pi2342 & n11990;
  assign n12591 = ~n12589 & ~n12590;
  assign n12592 = n12588 & n12591;
  assign n12593 = ~pi1911 & n11993;
  assign n12594 = ~pi1922 & n11995;
  assign n12595 = ~n12593 & ~n12594;
  assign n12596 = n12592 & n12595;
  assign n12597 = n12581 & n12596;
  assign po0561 = ~n12574 | ~n12597;
  assign n12599 = ~pi2272 & n12005;
  assign n12600 = ~pi2403 & n12007;
  assign n12601 = ~n12599 & ~n12600;
  assign n12602 = ~pi1951 & n11960;
  assign n12603 = ~pi2238 & n11963;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = n12601 & n12604;
  assign n12606 = ~pi2134 & n12001;
  assign n12607 = ~pi2225 & n12003;
  assign n12608 = ~n12606 & ~n12607;
  assign n12609 = ~pi2419 & n12012;
  assign n12610 = ~pi2060 & n12014;
  assign n12611 = ~n12609 & ~n12610;
  assign n12612 = n12608 & n12611;
  assign n12613 = ~pi1926 & n11995;
  assign n12614 = ~pi2462 & n11993;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = ~pi2126 & n11980;
  assign n12617 = ~pi2417 & n11983;
  assign n12618 = ~n12616 & ~n12617;
  assign n12619 = n12615 & n12618;
  assign n12620 = ~pi1989 & n11988;
  assign n12621 = ~pi2089 & n11990;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = n12619 & n12622;
  assign n12624 = ~pi2460 & n11973;
  assign n12625 = ~pi1924 & n11976;
  assign n12626 = ~n12624 & ~n12625;
  assign n12627 = n12623 & n12626;
  assign n12628 = n12612 & n12627;
  assign po0562 = ~n12605 | ~n12628;
  assign n12630 = ~pi2041 & n12012;
  assign n12631 = ~pi2061 & n12014;
  assign n12632 = ~n12630 & ~n12631;
  assign n12633 = ~pi1942 & n12005;
  assign n12634 = ~pi2109 & n12007;
  assign n12635 = ~n12633 & ~n12634;
  assign n12636 = n12632 & n12635;
  assign n12637 = ~pi2365 & n12001;
  assign n12638 = ~pi2166 & n12003;
  assign n12639 = ~n12637 & ~n12638;
  assign n12640 = ~pi2024 & n11960;
  assign n12641 = ~pi2240 & n11963;
  assign n12642 = ~n12640 & ~n12641;
  assign n12643 = n12639 & n12642;
  assign n12644 = ~pi2349 & n11988;
  assign n12645 = ~pi2352 & n11990;
  assign n12646 = ~pi2146 & n11973;
  assign n12647 = ~pi2008 & n11976;
  assign n12648 = ~n12646 & ~n12647;
  assign n12649 = ~n12645 & n12648;
  assign n12650 = ~n12644 & n12649;
  assign n12651 = ~pi1907 & n11995;
  assign n12652 = ~pi2471 & n11993;
  assign n12653 = ~n12651 & ~n12652;
  assign n12654 = n12650 & n12653;
  assign n12655 = ~pi2325 & n11980;
  assign n12656 = ~pi2427 & n11983;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = n12654 & n12657;
  assign n12659 = n12643 & n12658;
  assign po0563 = ~n12636 | ~n12659;
  assign n12661 = ~pi2244 & n12005;
  assign n12662 = ~pi2110 & n12007;
  assign n12663 = ~n12661 & ~n12662;
  assign n12664 = ~pi2025 & n11960;
  assign n12665 = ~pi2237 & n11963;
  assign n12666 = ~n12664 & ~n12665;
  assign n12667 = n12663 & n12666;
  assign n12668 = ~pi2423 & n12012;
  assign n12669 = ~pi2062 & n12014;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = ~pi2135 & n12001;
  assign n12672 = ~pi2221 & n12003;
  assign n12673 = ~n12671 & ~n12672;
  assign n12674 = n12670 & n12673;
  assign n12675 = ~pi1990 & n11988;
  assign n12676 = ~pi2090 & n11990;
  assign n12677 = ~n12675 & ~n12676;
  assign n12678 = ~pi2193 & n11995;
  assign n12679 = ~pi2176 & n11993;
  assign n12680 = ~n12678 & ~n12679;
  assign n12681 = n12677 & n12680;
  assign n12682 = ~pi2326 & n11980;
  assign n12683 = ~pi2205 & n11983;
  assign n12684 = ~n12682 & ~n12683;
  assign n12685 = n12681 & n12684;
  assign n12686 = ~pi2162 & n11973;
  assign n12687 = ~pi1938 & n11976;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = n12685 & n12688;
  assign n12690 = n12674 & n12689;
  assign po0564 = ~n12667 | ~n12690;
  assign n12692 = ~pi2355 & n12005;
  assign n12693 = ~pi2112 & n12007;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = ~pi2338 & n12001;
  assign n12696 = ~pi2129 & n12003;
  assign n12697 = ~n12695 & ~n12696;
  assign n12698 = n12694 & n12697;
  assign n12699 = ~pi2043 & n12012;
  assign n12700 = ~pi2371 & n12014;
  assign n12701 = ~n12699 & ~n12700;
  assign n12702 = ~pi2027 & n11960;
  assign n12703 = ~pi2235 & n11963;
  assign n12704 = ~n12702 & ~n12703;
  assign n12705 = n12701 & n12704;
  assign n12706 = ~pi2282 & n11973;
  assign n12707 = ~pi2010 & n11976;
  assign n12708 = ~pi2301 & n11980;
  assign n12709 = ~pi2430 & n11983;
  assign n12710 = ~n12708 & ~n12709;
  assign n12711 = ~n12707 & n12710;
  assign n12712 = ~n12706 & n12711;
  assign n12713 = ~pi1918 & n11995;
  assign n12714 = ~pi2476 & n11993;
  assign n12715 = ~n12713 & ~n12714;
  assign n12716 = n12712 & n12715;
  assign n12717 = ~pi2290 & n11988;
  assign n12718 = ~pi2273 & n11990;
  assign n12719 = ~n12717 & ~n12718;
  assign n12720 = n12716 & n12719;
  assign n12721 = n12705 & n12720;
  assign po0565 = ~n12698 | ~n12721;
  assign n12723 = ~pi2046 & n12012;
  assign n12724 = ~pi2335 & n12014;
  assign n12725 = ~n12723 & ~n12724;
  assign n12726 = ~pi2030 & n11960;
  assign n12727 = ~pi2187 & n11963;
  assign n12728 = ~n12726 & ~n12727;
  assign n12729 = n12725 & n12728;
  assign n12730 = ~pi2075 & n12005;
  assign n12731 = ~pi2115 & n12007;
  assign n12732 = ~n12730 & ~n12731;
  assign n12733 = ~pi2347 & n12001;
  assign n12734 = ~pi2169 & n12003;
  assign n12735 = ~n12733 & ~n12734;
  assign n12736 = n12732 & n12735;
  assign n12737 = ~pi2261 & n11973;
  assign n12738 = ~pi2012 & n11976;
  assign n12739 = ~pi2245 & n11980;
  assign n12740 = ~pi2414 & n11983;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = ~n12738 & n12741;
  assign n12743 = ~n12737 & n12742;
  assign n12744 = ~pi2397 & n11995;
  assign n12745 = ~pi2469 & n11993;
  assign n12746 = ~n12744 & ~n12745;
  assign n12747 = n12743 & n12746;
  assign n12748 = ~pi2329 & n11988;
  assign n12749 = ~pi2313 & n11990;
  assign n12750 = ~n12748 & ~n12749;
  assign n12751 = n12747 & n12750;
  assign n12752 = n12736 & n12751;
  assign po0566 = ~n12729 | ~n12752;
  assign n12754 = ~pi2077 & n12005;
  assign n12755 = ~pi2380 & n12007;
  assign n12756 = ~n12754 & ~n12755;
  assign n12757 = ~pi2416 & n12012;
  assign n12758 = ~pi2287 & n12014;
  assign n12759 = ~n12757 & ~n12758;
  assign n12760 = n12756 & n12759;
  assign n12761 = ~pi2141 & n12001;
  assign n12762 = ~pi2123 & n12003;
  assign n12763 = ~n12761 & ~n12762;
  assign n12764 = ~pi1947 & n11960;
  assign n12765 = ~pi2232 & n11963;
  assign n12766 = ~n12764 & ~n12765;
  assign n12767 = n12763 & n12766;
  assign n12768 = ~pi1937 & n11980;
  assign n12769 = ~pi2208 & n11983;
  assign n12770 = ~n12768 & ~n12769;
  assign n12771 = ~pi2470 & n11995;
  assign n12772 = ~pi2178 & n11993;
  assign n12773 = ~n12771 & ~n12772;
  assign n12774 = n12770 & n12773;
  assign n12775 = ~pi2263 & n11973;
  assign n12776 = ~pi1963 & n11976;
  assign n12777 = ~n12775 & ~n12776;
  assign n12778 = n12774 & n12777;
  assign n12779 = ~pi1996 & n11988;
  assign n12780 = ~pi2098 & n11990;
  assign n12781 = ~n12779 & ~n12780;
  assign n12782 = n12778 & n12781;
  assign n12783 = n12767 & n12782;
  assign po0567 = ~n12760 | ~n12783;
  assign n12785 = ~pi2079 & n12005;
  assign n12786 = ~pi2119 & n12007;
  assign n12787 = ~n12785 & ~n12786;
  assign n12788 = ~pi2298 & n12001;
  assign n12789 = ~pi2425 & n12003;
  assign n12790 = ~n12788 & ~n12789;
  assign n12791 = n12787 & n12790;
  assign n12792 = ~pi1946 & n11960;
  assign n12793 = ~pi2220 & n11963;
  assign n12794 = ~n12792 & ~n12793;
  assign n12795 = ~pi2050 & n12012;
  assign n12796 = ~pi2291 & n12014;
  assign n12797 = ~n12795 & ~n12796;
  assign n12798 = n12794 & n12797;
  assign n12799 = ~pi2454 & n11995;
  assign n12800 = ~pi2446 & n11993;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = ~pi2310 & n11988;
  assign n12803 = ~pi2309 & n11990;
  assign n12804 = ~n12802 & ~n12803;
  assign n12805 = n12801 & n12804;
  assign n12806 = ~pi2148 & n11973;
  assign n12807 = ~pi2015 & n11976;
  assign n12808 = ~n12806 & ~n12807;
  assign n12809 = n12805 & n12808;
  assign n12810 = ~pi2341 & n11980;
  assign n12811 = ~pi2340 & n11983;
  assign n12812 = ~n12810 & ~n12811;
  assign n12813 = n12809 & n12812;
  assign n12814 = n12798 & n12813;
  assign po0568 = ~n12791 | ~n12814;
  assign n12816 = ~pi1943 & n11960;
  assign n12817 = ~pi2223 & n11963;
  assign n12818 = ~n12816 & ~n12817;
  assign n12819 = ~pi2328 & n12001;
  assign n12820 = ~pi2171 & n12003;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = n12818 & n12821;
  assign n12823 = ~pi2051 & n12012;
  assign n12824 = ~pi2317 & n12014;
  assign n12825 = ~n12823 & ~n12824;
  assign n12826 = ~pi2080 & n12005;
  assign n12827 = ~pi2120 & n12007;
  assign n12828 = ~n12826 & ~n12827;
  assign n12829 = n12825 & n12828;
  assign n12830 = ~pi2452 & n11995;
  assign n12831 = ~pi2445 & n11993;
  assign n12832 = ~n12830 & ~n12831;
  assign n12833 = ~pi2344 & n11980;
  assign n12834 = ~pi2398 & n11983;
  assign n12835 = ~n12833 & ~n12834;
  assign n12836 = n12832 & n12835;
  assign n12837 = ~pi2000 & n11988;
  assign n12838 = ~pi2306 & n11990;
  assign n12839 = ~n12837 & ~n12838;
  assign n12840 = n12836 & n12839;
  assign n12841 = ~pi2149 & n11973;
  assign n12842 = ~pi2016 & n11976;
  assign n12843 = ~n12841 & ~n12842;
  assign n12844 = n12840 & n12843;
  assign n12845 = n12829 & n12844;
  assign po0569 = ~n12822 | ~n12845;
  assign n12847 = ~pi2143 & n12001;
  assign n12848 = ~pi1932 & n12003;
  assign n12849 = ~n12847 & ~n12848;
  assign n12850 = ~pi2407 & n12012;
  assign n12851 = ~pi2324 & n12014;
  assign n12852 = ~n12850 & ~n12851;
  assign n12853 = n12849 & n12852;
  assign n12854 = ~pi2372 & n12005;
  assign n12855 = ~pi2121 & n12007;
  assign n12856 = ~n12854 & ~n12855;
  assign n12857 = ~pi2330 & n11960;
  assign n12858 = ~pi2198 & n11963;
  assign n12859 = ~n12857 & ~n12858;
  assign n12860 = n12856 & n12859;
  assign n12861 = ~pi2001 & n11988;
  assign n12862 = ~pi2101 & n11990;
  assign n12863 = ~n12861 & ~n12862;
  assign n12864 = ~pi2391 & n11980;
  assign n12865 = ~pi2209 & n11983;
  assign n12866 = ~n12864 & ~n12865;
  assign n12867 = n12863 & n12866;
  assign n12868 = ~pi2150 & n11973;
  assign n12869 = ~pi1960 & n11976;
  assign n12870 = ~n12868 & ~n12869;
  assign n12871 = n12867 & n12870;
  assign n12872 = ~pi2181 & n11993;
  assign n12873 = ~pi2199 & n11995;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = n12871 & n12874;
  assign n12876 = n12860 & n12875;
  assign po0570 = ~n12853 | ~n12876;
  assign n12878 = ~pi2308 & n12001;
  assign n12879 = ~pi2172 & n12003;
  assign n12880 = ~n12878 & ~n12879;
  assign n12881 = ~pi2377 & n12005;
  assign n12882 = ~pi2336 & n12007;
  assign n12883 = ~n12881 & ~n12882;
  assign n12884 = n12880 & n12883;
  assign n12885 = ~pi2053 & n12012;
  assign n12886 = ~pi2066 & n12014;
  assign n12887 = ~n12885 & ~n12886;
  assign n12888 = ~pi2411 & n11960;
  assign n12889 = ~pi2190 & n11963;
  assign n12890 = ~n12888 & ~n12889;
  assign n12891 = n12887 & n12890;
  assign n12892 = ~pi2442 & n11995;
  assign n12893 = ~pi2383 & n11993;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = ~pi2260 & n11973;
  assign n12896 = ~pi1955 & n11976;
  assign n12897 = ~n12895 & ~n12896;
  assign n12898 = n12894 & n12897;
  assign n12899 = ~pi2395 & n11980;
  assign n12900 = ~pi2374 & n11983;
  assign n12901 = ~n12899 & ~n12900;
  assign n12902 = n12898 & n12901;
  assign n12903 = ~pi2267 & n11988;
  assign n12904 = ~pi2276 & n11990;
  assign n12905 = ~n12903 & ~n12904;
  assign n12906 = n12902 & n12905;
  assign n12907 = n12891 & n12906;
  assign po0571 = ~n12884 | ~n12907;
  assign n12909 = ~pi2083 & n12005;
  assign n12910 = ~pi2353 & n12007;
  assign n12911 = ~n12909 & ~n12910;
  assign n12912 = ~pi2054 & n12012;
  assign n12913 = ~pi2323 & n12014;
  assign n12914 = ~n12912 & ~n12913;
  assign n12915 = n12911 & n12914;
  assign n12916 = ~pi2035 & n11960;
  assign n12917 = ~pi2191 & n11963;
  assign n12918 = ~n12916 & ~n12917;
  assign n12919 = ~pi2279 & n12001;
  assign n12920 = ~pi1925 & n12003;
  assign n12921 = ~n12919 & ~n12920;
  assign n12922 = n12918 & n12921;
  assign n12923 = ~pi2268 & n11988;
  assign n12924 = ~pi2241 & n11990;
  assign n12925 = ~pi2152 & n11973;
  assign n12926 = ~pi2019 & n11976;
  assign n12927 = ~n12925 & ~n12926;
  assign n12928 = ~n12924 & n12927;
  assign n12929 = ~n12923 & n12928;
  assign n12930 = ~pi2449 & n11995;
  assign n12931 = ~pi2401 & n11993;
  assign n12932 = ~n12930 & ~n12931;
  assign n12933 = n12929 & n12932;
  assign n12934 = ~pi2386 & n11980;
  assign n12935 = ~pi1908 & n11983;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = n12933 & n12936;
  assign n12938 = n12922 & n12937;
  assign po0572 = ~n12915 | ~n12938;
  assign n12940 = ~pi2431 & n11960;
  assign n12941 = ~pi2179 & n11963;
  assign n12942 = ~n12940 & ~n12941;
  assign n12943 = ~pi2144 & n12001;
  assign n12944 = ~pi1906 & n12003;
  assign n12945 = ~n12943 & ~n12944;
  assign n12946 = n12942 & n12945;
  assign n12947 = ~pi2396 & n12012;
  assign n12948 = ~pi2068 & n12014;
  assign n12949 = ~n12947 & ~n12948;
  assign n12950 = ~pi2369 & n12005;
  assign n12951 = ~pi2357 & n12007;
  assign n12952 = ~n12950 & ~n12951;
  assign n12953 = n12949 & n12952;
  assign n12954 = ~pi2258 & n11973;
  assign n12955 = ~pi1956 & n11976;
  assign n12956 = ~n12954 & ~n12955;
  assign n12957 = ~pi2451 & n11995;
  assign n12958 = ~pi2182 & n11993;
  assign n12959 = ~n12957 & ~n12958;
  assign n12960 = n12956 & n12959;
  assign n12961 = ~pi2003 & n11988;
  assign n12962 = ~pi2104 & n11990;
  assign n12963 = ~n12961 & ~n12962;
  assign n12964 = n12960 & n12963;
  assign n12965 = ~pi2132 & n11980;
  assign n12966 = ~pi2283 & n11983;
  assign n12967 = ~n12965 & ~n12966;
  assign n12968 = n12964 & n12967;
  assign n12969 = n12953 & n12968;
  assign po0573 = ~n12946 | ~n12969;
  assign n12971 = ~pi2254 & n12001;
  assign n12972 = ~pi1915 & n12003;
  assign n12973 = ~n12971 & ~n12972;
  assign n12974 = ~pi2086 & n12005;
  assign n12975 = ~pi2331 & n12007;
  assign n12976 = ~n12974 & ~n12975;
  assign n12977 = n12973 & n12976;
  assign n12978 = ~pi2057 & n12012;
  assign n12979 = ~pi2311 & n12014;
  assign n12980 = ~n12978 & ~n12979;
  assign n12981 = ~pi2037 & n11960;
  assign n12982 = ~pi1919 & n11963;
  assign n12983 = ~n12981 & ~n12982;
  assign n12984 = n12980 & n12983;
  assign n12985 = ~pi2363 & n11980;
  assign n12986 = ~pi2303 & n11983;
  assign n12987 = ~n12985 & ~n12986;
  assign n12988 = ~pi2444 & n11995;
  assign n12989 = ~pi1909 & n11993;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = n12987 & n12990;
  assign n12992 = ~pi2155 & n11973;
  assign n12993 = ~pi2021 & n11976;
  assign n12994 = ~n12992 & ~n12993;
  assign n12995 = n12991 & n12994;
  assign n12996 = ~pi2251 & n11988;
  assign n12997 = ~pi1934 & n11990;
  assign n12998 = ~n12996 & ~n12997;
  assign n12999 = n12995 & n12998;
  assign n13000 = n12984 & n12999;
  assign po0574 = ~n12977 | ~n13000;
  assign n13002 = ~pi2367 & n12005;
  assign n13003 = ~pi1935 & n12007;
  assign n13004 = ~n13002 & ~n13003;
  assign n13005 = ~pi2429 & n11960;
  assign n13006 = ~pi1933 & n11963;
  assign n13007 = ~n13005 & ~n13006;
  assign n13008 = n13004 & n13007;
  assign n13009 = ~pi2242 & n12001;
  assign n13010 = ~pi1917 & n12003;
  assign n13011 = ~n13009 & ~n13010;
  assign n13012 = ~pi2388 & n12012;
  assign n13013 = ~pi2070 & n12014;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = n13011 & n13014;
  assign n13016 = ~pi2370 & n11980;
  assign n13017 = ~pi2318 & n11983;
  assign n13018 = ~n13016 & ~n13017;
  assign n13019 = ~pi2447 & n11995;
  assign n13020 = ~pi2184 & n11993;
  assign n13021 = ~n13019 & ~n13020;
  assign n13022 = n13018 & n13021;
  assign n13023 = ~pi2005 & n11988;
  assign n13024 = ~pi2106 & n11990;
  assign n13025 = ~n13023 & ~n13024;
  assign n13026 = n13022 & n13025;
  assign n13027 = ~pi2257 & n11973;
  assign n13028 = ~pi1950 & n11976;
  assign n13029 = ~n13027 & ~n13028;
  assign n13030 = n13026 & n13029;
  assign n13031 = n13015 & n13030;
  assign po0575 = ~n13008 | ~n13031;
  assign n13033 = ~pi2058 & n12012;
  assign n13034 = ~pi2071 & n12014;
  assign n13035 = ~n13033 & ~n13034;
  assign n13036 = ~pi2038 & n11960;
  assign n13037 = ~pi1930 & n11963;
  assign n13038 = ~n13036 & ~n13037;
  assign n13039 = n13035 & n13038;
  assign n13040 = ~pi2087 & n12005;
  assign n13041 = ~pi2124 & n12007;
  assign n13042 = ~n13040 & ~n13041;
  assign n13043 = ~pi2243 & n12001;
  assign n13044 = ~pi2174 & n12003;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = n13042 & n13045;
  assign n13047 = ~pi2246 & n11988;
  assign n13048 = ~pi2343 & n11990;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = ~pi2438 & n11995;
  assign n13051 = ~pi1910 & n11993;
  assign n13052 = ~n13050 & ~n13051;
  assign n13053 = n13049 & n13052;
  assign n13054 = ~pi2156 & n11973;
  assign n13055 = ~pi1953 & n11976;
  assign n13056 = ~n13054 & ~n13055;
  assign n13057 = n13053 & n13056;
  assign n13058 = ~pi2376 & n11980;
  assign n13059 = ~pi2296 & n11983;
  assign n13060 = ~n13058 & ~n13059;
  assign n13061 = n13057 & n13060;
  assign n13062 = n13046 & n13061;
  assign po0576 = ~n13039 | ~n13062;
  assign n13064 = ~pi0377 & n12564;
  assign n13065 = pi0450 & ~n12564;
  assign po0577 = n13064 | n13065;
  assign n13067 = ~pi0378 & n12564;
  assign n13068 = pi0449 & ~n12564;
  assign po0578 = n13067 | n13068;
  assign n13070 = ~pi0379 & n12564;
  assign n13071 = pi0451 & ~n12564;
  assign po0579 = n13070 | n13071;
  assign n13073 = ~pi0381 & n12564;
  assign n13074 = pi0477 & ~n12564;
  assign po0581 = n13073 | n13074;
  assign n13076 = ~pi0382 & n12564;
  assign n13077 = pi0478 & ~n12564;
  assign po0582 = n13076 | n13077;
  assign n13079 = ~pi0383 & n12564;
  assign n13080 = pi0479 & ~n12564;
  assign po0583 = n13079 | n13080;
  assign n13082 = ~pi0384 & n12564;
  assign n13083 = pi0481 & ~n12564;
  assign po0584 = n13082 | n13083;
  assign n13085 = ~pi0385 & n12564;
  assign n13086 = pi0482 & ~n12564;
  assign po0585 = n13085 | n13086;
  assign n13088 = ~pi0386 & n12564;
  assign n13089 = pi0453 & ~n12564;
  assign po0586 = n13088 | n13089;
  assign n13091 = ~pi0387 & n12564;
  assign n13092 = pi0454 & ~n12564;
  assign po0587 = n13091 | n13092;
  assign n13094 = ~pi0388 & n12564;
  assign n13095 = pi0456 & ~n12564;
  assign po0588 = n13094 | n13095;
  assign n13097 = ~pi0389 & n12564;
  assign n13098 = pi0459 & ~n12564;
  assign po0589 = n13097 | n13098;
  assign n13100 = ~pi0390 & n12564;
  assign n13101 = pi0462 & ~n12564;
  assign po0590 = n13100 | n13101;
  assign n13103 = ~pi0391 & n12564;
  assign n13104 = pi0458 & ~n12564;
  assign po0591 = n13103 | n13104;
  assign n13106 = ~pi0392 & n12564;
  assign n13107 = pi0461 & ~n12564;
  assign po0592 = n13106 | n13107;
  assign n13109 = ~pi0393 & n12564;
  assign n13110 = pi0463 & ~n12564;
  assign po0593 = n13109 | n13110;
  assign n13112 = ~pi0394 & n12564;
  assign n13113 = pi0465 & ~n12564;
  assign po0594 = n13112 | n13113;
  assign n13115 = ~pi0395 & n12564;
  assign n13116 = pi0466 & ~n12564;
  assign po0595 = n13115 | n13116;
  assign n13118 = ~pi0396 & n12564;
  assign n13119 = pi0467 & ~n12564;
  assign po0596 = n13118 | n13119;
  assign n13121 = ~pi0397 & n12564;
  assign n13122 = pi0469 & ~n12564;
  assign po0597 = n13121 | n13122;
  assign n13124 = ~pi0398 & n12564;
  assign n13125 = pi0470 & ~n12564;
  assign po0598 = n13124 | n13125;
  assign n13127 = ~pi0399 & n12564;
  assign n13128 = pi0471 & ~n12564;
  assign po0599 = n13127 | n13128;
  assign n13130 = ~pi0400 & n12564;
  assign n13131 = pi0473 & ~n12564;
  assign po0600 = n13130 | n13131;
  assign n13133 = ~pi0401 & n12564;
  assign n13134 = pi0474 & ~n12564;
  assign po0601 = n13133 | n13134;
  assign n13136 = ~pi0402 & n12564;
  assign n13137 = pi0475 & ~n12564;
  assign po0602 = n13136 | n13137;
  assign n13139 = ~pi0403 & n12564;
  assign n13140 = pi0472 & ~n12564;
  assign po0603 = n13139 | n13140;
  assign n13142 = ~pi0404 & n12564;
  assign n13143 = pi0468 & ~n12564;
  assign po0604 = n13142 | n13143;
  assign n13145 = ~pi0405 & n12564;
  assign n13146 = pi0464 & ~n12564;
  assign po0605 = n13145 | n13146;
  assign n13148 = ~pi0406 & n12564;
  assign n13149 = pi0460 & ~n12564;
  assign po0606 = n13148 | n13149;
  assign n13151 = ~pi0407 & n12564;
  assign n13152 = pi0480 & ~n12564;
  assign po0607 = n13151 | n13152;
  assign n13154 = ~pi0408 & n12564;
  assign n13155 = pi0457 & ~n12564;
  assign po0608 = n13154 | n13155;
  assign n13157 = ~pi0409 & n12564;
  assign n13158 = pi0455 & ~n12564;
  assign po0609 = n13157 | n13158;
  assign n13160 = pi1827 & n10977;
  assign n13161 = ~pi1692 & ~pi2989;
  assign n13162 = pi3179 & ~n13161;
  assign n13163 = ~pi1692 & ~pi3118;
  assign n13164 = n9401 & n13163;
  assign n13165 = ~n9378 & n13164;
  assign n13166 = ~pi3042 & n13165;
  assign n13167 = n13162 & ~n13166;
  assign n13168 = pi1858 & ~n13167;
  assign n13169 = ~n13160 & ~n13168;
  assign n13170 = ~n11139 & n13169;
  assign n13171 = ~n11154 & ~n13170;
  assign n13172 = ~pi1241 & n13171;
  assign n13173 = ~pi1256 & ~n13171;
  assign po1434 = ~n13172 & ~n13173;
  assign n13175 = ~pi1242 & n13171;
  assign n13176 = ~pi1267 & ~n13171;
  assign po1445 = ~n13175 & ~n13176;
  assign n13178 = ~po1434 & po1445;
  assign n13179 = pi1240 & n13171;
  assign n13180 = pi1243 & ~n13171;
  assign po1421 = n13179 | n13180;
  assign n13182 = pi1229 & n13171;
  assign n13183 = pi1231 & ~n13171;
  assign po1409 = n13182 | n13183;
  assign n13185 = po1421 & po1409;
  assign n13186 = n13178 & n13185;
  assign n13187 = ~pi0886 & n13186;
  assign n13188 = po1421 & ~po1409;
  assign n13189 = n13178 & n13188;
  assign n13190 = ~pi0647 & n13189;
  assign n13191 = ~n13187 & ~n13190;
  assign n13192 = ~po1434 & ~po1445;
  assign n13193 = n13188 & n13192;
  assign n13194 = ~pi0751 & n13193;
  assign n13195 = ~po1421 & ~po1409;
  assign n13196 = n13192 & n13195;
  assign n13197 = ~pi0690 & n13196;
  assign n13198 = ~n13194 & ~n13197;
  assign n13199 = n13185 & n13192;
  assign n13200 = ~pi0626 & n13199;
  assign n13201 = ~po1421 & po1409;
  assign n13202 = n13178 & n13201;
  assign n13203 = ~pi0605 & n13202;
  assign n13204 = ~n13200 & ~n13203;
  assign n13205 = po1434 & po1445;
  assign n13206 = n13201 & n13205;
  assign n13207 = ~pi0792 & n13206;
  assign n13208 = po1434 & ~po1445;
  assign n13209 = n13195 & n13208;
  assign n13210 = ~pi0771 & n13209;
  assign n13211 = ~n13207 & ~n13210;
  assign n13212 = n13178 & n13195;
  assign n13213 = ~pi0729 & n13212;
  assign n13214 = n13192 & n13201;
  assign n13215 = ~pi0710 & n13214;
  assign n13216 = ~n13213 & ~n13215;
  assign n13217 = n13188 & n13205;
  assign n13218 = ~pi0839 & n13217;
  assign n13219 = n13188 & n13208;
  assign n13220 = ~pi0584 & n13219;
  assign n13221 = ~n13218 & ~n13220;
  assign n13222 = n13216 & n13221;
  assign n13223 = n13211 & n13222;
  assign n13224 = n13204 & n13223;
  assign n13225 = n13195 & n13205;
  assign n13226 = ~pi0565 & n13225;
  assign n13227 = n13201 & n13208;
  assign n13228 = ~pi0669 & n13227;
  assign n13229 = ~n13226 & ~n13228;
  assign n13230 = n13224 & n13229;
  assign n13231 = n13185 & n13208;
  assign n13232 = ~pi0815 & n13231;
  assign n13233 = n13185 & n13205;
  assign n13234 = ~pi0862 & n13233;
  assign n13235 = ~n13232 & ~n13234;
  assign n13236 = n13230 & n13235;
  assign n13237 = n13198 & n13236;
  assign po0610 = ~n13191 | ~n13237;
  assign n13239 = ~pi0556 & n13225;
  assign n13240 = ~pi0660 & n13227;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = ~pi0806 & n13231;
  assign n13243 = ~pi0853 & n13233;
  assign n13244 = ~n13242 & ~n13243;
  assign n13245 = ~pi0830 & n13217;
  assign n13246 = ~pi0577 & n13219;
  assign n13247 = ~n13245 & ~n13246;
  assign n13248 = ~pi0721 & n13212;
  assign n13249 = ~pi0701 & n13214;
  assign n13250 = ~n13248 & ~n13249;
  assign n13251 = ~pi0617 & n13199;
  assign n13252 = ~pi0596 & n13202;
  assign n13253 = ~n13251 & ~n13252;
  assign n13254 = ~pi0783 & n13206;
  assign n13255 = ~pi0762 & n13209;
  assign n13256 = ~n13254 & ~n13255;
  assign n13257 = n13253 & n13256;
  assign n13258 = n13250 & n13257;
  assign n13259 = n13247 & n13258;
  assign n13260 = ~pi0878 & n13186;
  assign n13261 = ~pi0639 & n13189;
  assign n13262 = ~n13260 & ~n13261;
  assign n13263 = n13259 & n13262;
  assign n13264 = ~pi0743 & n13193;
  assign n13265 = ~pi0681 & n13196;
  assign n13266 = ~n13264 & ~n13265;
  assign n13267 = n13263 & n13266;
  assign n13268 = n13244 & n13267;
  assign po0612 = ~n13241 | ~n13268;
  assign n13270 = ~pi0831 & n13217;
  assign n13271 = ~pi0578 & n13219;
  assign n13272 = ~n13270 & ~n13271;
  assign n13273 = ~pi0618 & n13199;
  assign n13274 = ~pi0597 & n13202;
  assign n13275 = ~n13273 & ~n13274;
  assign n13276 = ~pi0879 & n13186;
  assign n13277 = ~pi0945 & n13189;
  assign n13278 = ~n13276 & ~n13277;
  assign n13279 = ~pi0557 & n13225;
  assign n13280 = ~pi0661 & n13227;
  assign n13281 = ~n13279 & ~n13280;
  assign n13282 = ~pi0807 & n13231;
  assign n13283 = ~pi0854 & n13233;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = ~pi0744 & n13193;
  assign n13286 = ~pi0682 & n13196;
  assign n13287 = ~n13285 & ~n13286;
  assign n13288 = n13284 & n13287;
  assign n13289 = n13281 & n13288;
  assign n13290 = n13278 & n13289;
  assign n13291 = ~pi0722 & n13212;
  assign n13292 = ~pi0702 & n13214;
  assign n13293 = ~n13291 & ~n13292;
  assign n13294 = n13290 & n13293;
  assign n13295 = ~pi0784 & n13206;
  assign n13296 = ~pi0763 & n13209;
  assign n13297 = ~n13295 & ~n13296;
  assign n13298 = n13294 & n13297;
  assign n13299 = n13275 & n13298;
  assign po0613 = ~n13272 | ~n13299;
  assign n13301 = ~pi0785 & n13206;
  assign n13302 = ~pi0764 & n13209;
  assign n13303 = ~n13301 & ~n13302;
  assign n13304 = ~pi0619 & n13199;
  assign n13305 = ~pi0598 & n13202;
  assign n13306 = ~n13304 & ~n13305;
  assign n13307 = ~pi0880 & n13186;
  assign n13308 = ~pi0640 & n13189;
  assign n13309 = ~n13307 & ~n13308;
  assign n13310 = ~pi0558 & n13225;
  assign n13311 = ~pi0662 & n13227;
  assign n13312 = ~n13310 & ~n13311;
  assign n13313 = ~pi0745 & n13193;
  assign n13314 = ~pi0683 & n13196;
  assign n13315 = ~n13313 & ~n13314;
  assign n13316 = ~pi0808 & n13231;
  assign n13317 = ~pi0855 & n13233;
  assign n13318 = ~n13316 & ~n13317;
  assign n13319 = n13315 & n13318;
  assign n13320 = n13312 & n13319;
  assign n13321 = n13309 & n13320;
  assign n13322 = ~pi0832 & n13217;
  assign n13323 = ~pi0907 & n13219;
  assign n13324 = ~n13322 & ~n13323;
  assign n13325 = n13321 & n13324;
  assign n13326 = ~pi0738 & n13212;
  assign n13327 = ~pi0703 & n13214;
  assign n13328 = ~n13326 & ~n13327;
  assign n13329 = n13325 & n13328;
  assign n13330 = n13306 & n13329;
  assign po0614 = ~n13303 | ~n13330;
  assign n13332 = ~pi0809 & n13231;
  assign n13333 = ~pi0856 & n13233;
  assign n13334 = ~n13332 & ~n13333;
  assign n13335 = ~pi0786 & n13206;
  assign n13336 = ~pi0915 & n13209;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = ~pi0833 & n13217;
  assign n13339 = ~pi0579 & n13219;
  assign n13340 = ~n13338 & ~n13339;
  assign n13341 = n13337 & n13340;
  assign n13342 = ~pi0940 & n13196;
  assign n13343 = n13341 & ~n13342;
  assign n13344 = ~pi0663 & n13227;
  assign n13345 = ~pi0723 & n13212;
  assign n13346 = ~pi0932 & n13214;
  assign n13347 = ~n13345 & ~n13346;
  assign n13348 = ~n13344 & n13347;
  assign n13349 = ~pi0641 & n13189;
  assign n13350 = ~pi0949 & n13186;
  assign n13351 = ~n13349 & ~n13350;
  assign n13352 = n13348 & n13351;
  assign n13353 = ~pi0620 & n13199;
  assign n13354 = ~pi0599 & n13202;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = ~pi0921 & n13193;
  assign n13357 = n13355 & ~n13356;
  assign n13358 = ~pi0559 & n13225;
  assign n13359 = n13357 & ~n13358;
  assign n13360 = n13352 & n13359;
  assign n13361 = n13343 & n13360;
  assign po0615 = ~n13334 | ~n13361;
  assign n13363 = ~pi0881 & n13186;
  assign n13364 = ~pi0642 & n13189;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = ~pi0560 & n13225;
  assign n13367 = ~pi0664 & n13227;
  assign n13368 = ~n13366 & ~n13367;
  assign n13369 = ~pi0517 & n13199;
  assign n13370 = ~pi0600 & n13202;
  assign n13371 = ~n13369 & ~n13370;
  assign n13372 = ~pi0898 & n13217;
  assign n13373 = ~pi0580 & n13219;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = ~pi0908 & n13206;
  assign n13376 = ~pi0765 & n13209;
  assign n13377 = ~n13375 & ~n13376;
  assign n13378 = ~pi0925 & n13212;
  assign n13379 = ~pi0704 & n13214;
  assign n13380 = ~n13378 & ~n13379;
  assign n13381 = n13377 & n13380;
  assign n13382 = n13374 & n13381;
  assign n13383 = n13371 & n13382;
  assign n13384 = ~pi0902 & n13231;
  assign n13385 = ~pi0518 & n13233;
  assign n13386 = ~n13384 & ~n13385;
  assign n13387 = n13383 & n13386;
  assign n13388 = ~pi0746 & n13193;
  assign n13389 = ~pi0684 & n13196;
  assign n13390 = ~n13388 & ~n13389;
  assign n13391 = n13387 & n13390;
  assign n13392 = n13368 & n13391;
  assign po0616 = ~n13365 | ~n13392;
  assign n13394 = ~pi0724 & n13212;
  assign n13395 = ~pi0705 & n13214;
  assign n13396 = ~n13394 & ~n13395;
  assign n13397 = ~pi0834 & n13217;
  assign n13398 = ~pi0586 & n13219;
  assign n13399 = ~n13397 & ~n13398;
  assign n13400 = ~pi0747 & n13193;
  assign n13401 = ~pi0685 & n13196;
  assign n13402 = ~n13400 & ~n13401;
  assign n13403 = ~pi0810 & n13231;
  assign n13404 = ~pi0857 & n13233;
  assign n13405 = ~n13403 & ~n13404;
  assign n13406 = ~pi0916 & n13225;
  assign n13407 = ~pi0665 & n13227;
  assign n13408 = ~n13406 & ~n13407;
  assign n13409 = ~pi0882 & n13186;
  assign n13410 = ~pi0944 & n13189;
  assign n13411 = ~n13409 & ~n13410;
  assign n13412 = n13408 & n13411;
  assign n13413 = n13405 & n13412;
  assign n13414 = n13402 & n13413;
  assign n13415 = ~pi0621 & n13199;
  assign n13416 = ~pi0601 & n13202;
  assign n13417 = ~n13415 & ~n13416;
  assign n13418 = n13414 & n13417;
  assign n13419 = ~pi0787 & n13206;
  assign n13420 = ~pi0766 & n13209;
  assign n13421 = ~n13419 & ~n13420;
  assign n13422 = n13418 & n13421;
  assign n13423 = n13399 & n13422;
  assign po0617 = ~n13396 | ~n13423;
  assign n13425 = ~pi0561 & n13225;
  assign n13426 = ~pi0942 & n13227;
  assign n13427 = ~n13425 & ~n13426;
  assign n13428 = ~pi0811 & n13231;
  assign n13429 = ~pi0858 & n13233;
  assign n13430 = ~n13428 & ~n13429;
  assign n13431 = ~pi0725 & n13212;
  assign n13432 = ~pi0706 & n13214;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = ~pi0788 & n13206;
  assign n13435 = ~pi0767 & n13209;
  assign n13436 = ~n13434 & ~n13435;
  assign n13437 = ~pi0835 & n13217;
  assign n13438 = ~pi0581 & n13219;
  assign n13439 = ~n13437 & ~n13438;
  assign n13440 = ~pi0622 & n13199;
  assign n13441 = ~pi0602 & n13202;
  assign n13442 = ~n13440 & ~n13441;
  assign n13443 = n13439 & n13442;
  assign n13444 = n13436 & n13443;
  assign n13445 = n13433 & n13444;
  assign n13446 = ~pi0883 & n13186;
  assign n13447 = ~pi0643 & n13189;
  assign n13448 = ~n13446 & ~n13447;
  assign n13449 = n13445 & n13448;
  assign n13450 = ~pi0748 & n13193;
  assign n13451 = ~pi0686 & n13196;
  assign n13452 = ~n13450 & ~n13451;
  assign n13453 = n13449 & n13452;
  assign n13454 = n13430 & n13453;
  assign po0618 = ~n13427 | ~n13454;
  assign n13456 = ~pi1031 & n13193;
  assign n13457 = ~pi1018 & n13196;
  assign n13458 = ~n13456 & ~n13457;
  assign n13459 = ~pi1054 & n13186;
  assign n13460 = ~pi1119 & n13189;
  assign n13461 = ~n13459 & ~n13460;
  assign n13462 = ~pi1112 & n13199;
  assign n13463 = ~pi1000 & n13202;
  assign n13464 = ~n13462 & ~n13463;
  assign n13465 = ~pi1103 & n13212;
  assign n13466 = ~pi1024 & n13214;
  assign n13467 = ~n13465 & ~n13466;
  assign n13468 = ~pi1066 & n13217;
  assign n13469 = ~pi0995 & n13219;
  assign n13470 = ~n13468 & ~n13469;
  assign n13471 = ~pi1087 & n13206;
  assign n13472 = ~pi1036 & n13209;
  assign n13473 = ~n13471 & ~n13472;
  assign n13474 = n13470 & n13473;
  assign n13475 = n13467 & n13474;
  assign n13476 = n13464 & n13475;
  assign n13477 = ~pi1071 & n13231;
  assign n13478 = ~pi1049 & n13233;
  assign n13479 = ~n13477 & ~n13478;
  assign n13480 = n13476 & n13479;
  assign n13481 = ~pi0990 & n13225;
  assign n13482 = ~pi1012 & n13227;
  assign n13483 = ~n13481 & ~n13482;
  assign n13484 = n13480 & n13483;
  assign n13485 = n13461 & n13484;
  assign po0619 = ~n13458 | ~n13485;
  assign n13487 = ~pi0749 & n13193;
  assign n13488 = ~pi0688 & n13196;
  assign n13489 = ~n13487 & ~n13488;
  assign n13490 = ~pi0884 & n13186;
  assign n13491 = ~pi0645 & n13189;
  assign n13492 = ~n13490 & ~n13491;
  assign n13493 = ~pi0563 & n13225;
  assign n13494 = ~pi0667 & n13227;
  assign n13495 = ~n13493 & ~n13494;
  assign n13496 = ~pi0790 & n13206;
  assign n13497 = ~pi0769 & n13209;
  assign n13498 = ~n13496 & ~n13497;
  assign n13499 = ~pi0624 & n13199;
  assign n13500 = ~pi0603 & n13202;
  assign n13501 = ~n13499 & ~n13500;
  assign n13502 = ~pi0837 & n13217;
  assign n13503 = ~pi0582 & n13219;
  assign n13504 = ~n13502 & ~n13503;
  assign n13505 = ~pi0727 & n13212;
  assign n13506 = ~pi0708 & n13214;
  assign n13507 = ~n13505 & ~n13506;
  assign n13508 = n13504 & n13507;
  assign n13509 = n13501 & n13508;
  assign n13510 = n13498 & n13509;
  assign n13511 = n13495 & n13510;
  assign n13512 = ~pi0813 & n13231;
  assign n13513 = ~pi0860 & n13233;
  assign n13514 = ~n13512 & ~n13513;
  assign n13515 = n13511 & n13514;
  assign n13516 = n13492 & n13515;
  assign po0620 = ~n13489 | ~n13516;
  assign n13518 = ~pi0838 & n13217;
  assign n13519 = ~pi0583 & n13219;
  assign n13520 = ~n13518 & ~n13519;
  assign n13521 = ~pi0791 & n13206;
  assign n13522 = ~pi0770 & n13209;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = ~pi0625 & n13199;
  assign n13525 = ~pi0604 & n13202;
  assign n13526 = ~n13524 & ~n13525;
  assign n13527 = ~pi0728 & n13212;
  assign n13528 = ~pi0709 & n13214;
  assign n13529 = ~n13527 & ~n13528;
  assign n13530 = n13526 & n13529;
  assign n13531 = n13523 & n13530;
  assign n13532 = n13520 & n13531;
  assign n13533 = ~pi0750 & n13193;
  assign n13534 = ~pi0689 & n13196;
  assign n13535 = ~n13533 & ~n13534;
  assign n13536 = n13532 & n13535;
  assign n13537 = ~pi0814 & n13231;
  assign n13538 = ~pi0861 & n13233;
  assign n13539 = ~pi0668 & n13227;
  assign n13540 = ~pi0564 & n13225;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = ~pi0646 & n13189;
  assign n13543 = ~pi0885 & n13186;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = n13541 & n13544;
  assign n13546 = ~n13538 & n13545;
  assign n13547 = ~n13537 & n13546;
  assign po0621 = ~n13536 | ~n13547;
  assign n13549 = ~pi0752 & n13193;
  assign n13550 = ~pi0691 & n13196;
  assign n13551 = ~n13549 & ~n13550;
  assign n13552 = ~pi0913 & n13225;
  assign n13553 = ~pi0670 & n13227;
  assign n13554 = ~n13552 & ~n13553;
  assign n13555 = ~pi0627 & n13199;
  assign n13556 = ~pi0606 & n13202;
  assign n13557 = ~n13555 & ~n13556;
  assign n13558 = ~pi0840 & n13217;
  assign n13559 = ~pi0585 & n13219;
  assign n13560 = ~n13558 & ~n13559;
  assign n13561 = ~pi0793 & n13206;
  assign n13562 = ~pi0772 & n13209;
  assign n13563 = ~n13561 & ~n13562;
  assign n13564 = ~pi0730 & n13212;
  assign n13565 = ~pi0711 & n13214;
  assign n13566 = ~n13564 & ~n13565;
  assign n13567 = n13563 & n13566;
  assign n13568 = n13560 & n13567;
  assign n13569 = n13557 & n13568;
  assign n13570 = ~pi0816 & n13231;
  assign n13571 = ~pi0863 & n13233;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = n13569 & n13572;
  assign n13574 = ~pi0887 & n13186;
  assign n13575 = ~pi0648 & n13189;
  assign n13576 = ~n13574 & ~n13575;
  assign n13577 = n13573 & n13576;
  assign n13578 = n13554 & n13577;
  assign po0622 = ~n13551 | ~n13578;
  assign n13580 = ~pi0566 & n13225;
  assign n13581 = ~pi0912 & n13227;
  assign n13582 = ~n13580 & ~n13581;
  assign n13583 = ~pi0888 & n13186;
  assign n13584 = ~pi0649 & n13189;
  assign n13585 = ~n13583 & ~n13584;
  assign n13586 = ~pi0628 & n13199;
  assign n13587 = ~pi0607 & n13202;
  assign n13588 = ~n13586 & ~n13587;
  assign n13589 = ~pi0794 & n13206;
  assign n13590 = ~pi0773 & n13209;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = ~pi0731 & n13212;
  assign n13593 = ~pi0712 & n13214;
  assign n13594 = ~n13592 & ~n13593;
  assign n13595 = ~pi0841 & n13217;
  assign n13596 = ~pi0904 & n13219;
  assign n13597 = ~n13595 & ~n13596;
  assign n13598 = n13594 & n13597;
  assign n13599 = n13591 & n13598;
  assign n13600 = n13588 & n13599;
  assign n13601 = ~pi0753 & n13193;
  assign n13602 = ~pi0692 & n13196;
  assign n13603 = ~n13601 & ~n13602;
  assign n13604 = n13600 & n13603;
  assign n13605 = ~pi0817 & n13231;
  assign n13606 = ~pi0864 & n13233;
  assign n13607 = ~n13605 & ~n13606;
  assign n13608 = n13604 & n13607;
  assign n13609 = n13585 & n13608;
  assign po0623 = ~n13582 | ~n13609;
  assign n13611 = ~pi0818 & n13231;
  assign n13612 = ~pi0865 & n13233;
  assign n13613 = ~n13611 & ~n13612;
  assign n13614 = ~pi0567 & n13225;
  assign n13615 = ~pi0671 & n13227;
  assign n13616 = ~n13614 & ~n13615;
  assign n13617 = ~pi0842 & n13217;
  assign n13618 = ~pi0905 & n13219;
  assign n13619 = ~n13617 & ~n13618;
  assign n13620 = ~pi0629 & n13199;
  assign n13621 = ~pi0900 & n13202;
  assign n13622 = ~n13620 & ~n13621;
  assign n13623 = ~pi0795 & n13206;
  assign n13624 = ~pi0910 & n13209;
  assign n13625 = ~n13623 & ~n13624;
  assign n13626 = ~pi0732 & n13212;
  assign n13627 = ~pi0929 & n13214;
  assign n13628 = ~n13626 & ~n13627;
  assign n13629 = n13625 & n13628;
  assign n13630 = n13622 & n13629;
  assign n13631 = n13619 & n13630;
  assign n13632 = ~pi0919 & n13193;
  assign n13633 = ~pi0926 & n13196;
  assign n13634 = ~n13632 & ~n13633;
  assign n13635 = n13631 & n13634;
  assign n13636 = ~pi0947 & n13186;
  assign n13637 = ~pi0650 & n13189;
  assign n13638 = ~n13636 & ~n13637;
  assign n13639 = n13635 & n13638;
  assign n13640 = n13616 & n13639;
  assign po0624 = ~n13613 | ~n13640;
  assign n13642 = ~pi1127 & n13199;
  assign n13643 = ~pi1001 & n13202;
  assign n13644 = ~n13642 & ~n13643;
  assign n13645 = ~pi1101 & n13212;
  assign n13646 = ~pi1025 & n13214;
  assign n13647 = ~n13645 & ~n13646;
  assign n13648 = ~pi1032 & n13193;
  assign n13649 = ~pi1019 & n13196;
  assign n13650 = ~n13648 & ~n13649;
  assign n13651 = ~pi1120 & n13186;
  assign n13652 = ~pi1118 & n13189;
  assign n13653 = ~n13651 & ~n13652;
  assign n13654 = ~pi1072 & n13231;
  assign n13655 = ~pi0986 & n13233;
  assign n13656 = ~n13654 & ~n13655;
  assign n13657 = ~pi1078 & n13225;
  assign n13658 = ~pi1111 & n13227;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = n13656 & n13659;
  assign n13661 = n13653 & n13660;
  assign n13662 = n13650 & n13661;
  assign n13663 = ~pi1063 & n13217;
  assign n13664 = ~pi0996 & n13219;
  assign n13665 = ~n13663 & ~n13664;
  assign n13666 = n13662 & n13665;
  assign n13667 = ~pi1085 & n13206;
  assign n13668 = ~pi1037 & n13209;
  assign n13669 = ~n13667 & ~n13668;
  assign n13670 = n13666 & n13669;
  assign n13671 = n13647 & n13670;
  assign po0625 = ~n13644 | ~n13671;
  assign n13673 = ~pi0569 & n13225;
  assign n13674 = ~pi0673 & n13227;
  assign n13675 = ~n13673 & ~n13674;
  assign n13676 = ~pi0890 & n13186;
  assign n13677 = ~pi0652 & n13189;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = ~pi0844 & n13217;
  assign n13680 = ~pi0588 & n13219;
  assign n13681 = ~n13679 & ~n13680;
  assign n13682 = ~pi0734 & n13212;
  assign n13683 = ~pi0714 & n13214;
  assign n13684 = ~n13682 & ~n13683;
  assign n13685 = ~pi0631 & n13199;
  assign n13686 = ~pi0609 & n13202;
  assign n13687 = ~n13685 & ~n13686;
  assign n13688 = ~pi0797 & n13206;
  assign n13689 = ~pi0775 & n13209;
  assign n13690 = ~n13688 & ~n13689;
  assign n13691 = n13687 & n13690;
  assign n13692 = n13684 & n13691;
  assign n13693 = n13681 & n13692;
  assign n13694 = ~pi0755 & n13193;
  assign n13695 = ~pi0694 & n13196;
  assign n13696 = ~n13694 & ~n13695;
  assign n13697 = n13693 & n13696;
  assign n13698 = ~pi0820 & n13231;
  assign n13699 = ~pi0867 & n13233;
  assign n13700 = ~n13698 & ~n13699;
  assign n13701 = n13697 & n13700;
  assign n13702 = n13678 & n13701;
  assign po0626 = ~n13675 | ~n13702;
  assign n13704 = ~pi0799 & n13206;
  assign n13705 = ~pi0911 & n13209;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = ~pi0735 & n13212;
  assign n13708 = ~pi0927 & n13214;
  assign n13709 = ~n13707 & ~n13708;
  assign n13710 = ~pi0917 & n13193;
  assign n13711 = ~pi0937 & n13196;
  assign n13712 = ~n13710 & ~n13711;
  assign n13713 = ~pi0570 & n13225;
  assign n13714 = ~pi0674 & n13227;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = ~pi0892 & n13186;
  assign n13717 = ~pi0653 & n13189;
  assign n13718 = ~n13716 & ~n13717;
  assign n13719 = ~pi0822 & n13231;
  assign n13720 = ~pi0869 & n13233;
  assign n13721 = ~n13719 & ~n13720;
  assign n13722 = n13718 & n13721;
  assign n13723 = n13715 & n13722;
  assign n13724 = n13712 & n13723;
  assign n13725 = ~pi0846 & n13217;
  assign n13726 = ~pi0589 & n13219;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = n13724 & n13727;
  assign n13729 = ~pi0632 & n13199;
  assign n13730 = ~pi0610 & n13202;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = n13728 & n13731;
  assign n13733 = n13709 & n13732;
  assign po0627 = ~n13706 | ~n13733;
  assign n13735 = ~pi1083 & n13206;
  assign n13736 = ~pi1038 & n13209;
  assign n13737 = ~n13735 & ~n13736;
  assign n13738 = ~pi1060 & n13217;
  assign n13739 = ~pi0998 & n13219;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = ~pi1056 & n13186;
  assign n13742 = ~pi1010 & n13189;
  assign n13743 = ~n13741 & ~n13742;
  assign n13744 = ~pi1033 & n13193;
  assign n13745 = ~pi1020 & n13196;
  assign n13746 = ~n13744 & ~n13745;
  assign n13747 = ~pi1067 & n13231;
  assign n13748 = ~pi0985 & n13233;
  assign n13749 = ~n13747 & ~n13748;
  assign n13750 = ~pi0992 & n13225;
  assign n13751 = ~pi1014 & n13227;
  assign n13752 = ~n13750 & ~n13751;
  assign n13753 = n13749 & n13752;
  assign n13754 = n13746 & n13753;
  assign n13755 = n13743 & n13754;
  assign n13756 = ~pi1006 & n13199;
  assign n13757 = ~pi1065 & n13202;
  assign n13758 = ~n13756 & ~n13757;
  assign n13759 = n13755 & n13758;
  assign n13760 = ~pi1099 & n13212;
  assign n13761 = ~pi1026 & n13214;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = n13759 & n13762;
  assign n13764 = n13740 & n13763;
  assign po0628 = ~n13737 | ~n13764;
  assign n13766 = ~pi0993 & n13225;
  assign n13767 = ~pi1015 & n13227;
  assign n13768 = ~n13766 & ~n13767;
  assign n13769 = ~pi1070 & n13231;
  assign n13770 = ~pi0984 & n13233;
  assign n13771 = ~n13769 & ~n13770;
  assign n13772 = ~pi1122 & n13199;
  assign n13773 = ~pi1003 & n13202;
  assign n13774 = ~n13772 & ~n13773;
  assign n13775 = ~pi1041 & n13206;
  assign n13776 = ~pi1039 & n13209;
  assign n13777 = ~n13775 & ~n13776;
  assign n13778 = ~pi1029 & n13212;
  assign n13779 = ~pi1027 & n13214;
  assign n13780 = ~n13778 & ~n13779;
  assign n13781 = ~pi1046 & n13217;
  assign n13782 = ~pi0997 & n13219;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = n13780 & n13783;
  assign n13785 = n13777 & n13784;
  assign n13786 = n13774 & n13785;
  assign n13787 = ~pi1057 & n13186;
  assign n13788 = ~pi1011 & n13189;
  assign n13789 = ~n13787 & ~n13788;
  assign n13790 = n13786 & n13789;
  assign n13791 = ~pi1034 & n13193;
  assign n13792 = ~pi1022 & n13196;
  assign n13793 = ~n13791 & ~n13792;
  assign n13794 = n13790 & n13793;
  assign n13795 = n13771 & n13794;
  assign po0629 = ~n13768 | ~n13795;
  assign n13797 = ~pi1047 & n13217;
  assign n13798 = ~pi1076 & n13219;
  assign n13799 = ~n13797 & ~n13798;
  assign n13800 = ~pi1077 & n13206;
  assign n13801 = ~pi1091 & n13209;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~pi1090 & n13225;
  assign n13804 = ~pi1109 & n13227;
  assign n13805 = ~n13803 & ~n13804;
  assign n13806 = ~pi1121 & n13186;
  assign n13807 = ~pi1117 & n13189;
  assign n13808 = ~n13806 & ~n13807;
  assign n13809 = ~pi1044 & n13231;
  assign n13810 = ~pi1051 & n13233;
  assign n13811 = ~n13809 & ~n13810;
  assign n13812 = ~pi1094 & n13193;
  assign n13813 = ~pi1021 & n13196;
  assign n13814 = ~n13812 & ~n13813;
  assign n13815 = n13811 & n13814;
  assign n13816 = n13808 & n13815;
  assign n13817 = n13805 & n13816;
  assign n13818 = ~pi1007 & n13199;
  assign n13819 = ~pi1062 & n13202;
  assign n13820 = ~n13818 & ~n13819;
  assign n13821 = n13817 & n13820;
  assign n13822 = ~pi1100 & n13212;
  assign n13823 = ~pi1105 & n13214;
  assign n13824 = ~n13822 & ~n13823;
  assign n13825 = n13821 & n13824;
  assign n13826 = n13802 & n13825;
  assign po0630 = ~n13799 | ~n13826;
  assign n13828 = ~pi0736 & n13212;
  assign n13829 = ~pi0715 & n13214;
  assign n13830 = ~n13828 & ~n13829;
  assign n13831 = ~pi0633 & n13199;
  assign n13832 = ~pi0611 & n13202;
  assign n13833 = ~n13831 & ~n13832;
  assign n13834 = ~pi0893 & n13186;
  assign n13835 = ~pi0654 & n13189;
  assign n13836 = ~n13834 & ~n13835;
  assign n13837 = ~pi0571 & n13225;
  assign n13838 = ~pi0675 & n13227;
  assign n13839 = ~n13837 & ~n13838;
  assign n13840 = ~pi0823 & n13231;
  assign n13841 = ~pi0870 & n13233;
  assign n13842 = ~n13840 & ~n13841;
  assign n13843 = ~pi0756 & n13193;
  assign n13844 = ~pi0695 & n13196;
  assign n13845 = ~n13843 & ~n13844;
  assign n13846 = n13842 & n13845;
  assign n13847 = n13839 & n13846;
  assign n13848 = n13836 & n13847;
  assign n13849 = ~pi0847 & n13217;
  assign n13850 = ~pi0590 & n13219;
  assign n13851 = ~n13849 & ~n13850;
  assign n13852 = n13848 & n13851;
  assign n13853 = ~pi0800 & n13206;
  assign n13854 = ~pi0776 & n13209;
  assign n13855 = ~n13853 & ~n13854;
  assign n13856 = n13852 & n13855;
  assign n13857 = n13833 & n13856;
  assign po0631 = ~n13830 | ~n13857;
  assign n13859 = ~pi0737 & n13212;
  assign n13860 = ~pi0716 & n13214;
  assign n13861 = ~n13859 & ~n13860;
  assign n13862 = ~pi0848 & n13217;
  assign n13863 = ~pi0591 & n13219;
  assign n13864 = ~n13862 & ~n13863;
  assign n13865 = ~pi0894 & n13186;
  assign n13866 = ~pi0655 & n13189;
  assign n13867 = ~n13865 & ~n13866;
  assign n13868 = ~pi0572 & n13225;
  assign n13869 = ~pi0676 & n13227;
  assign n13870 = ~n13868 & ~n13869;
  assign n13871 = ~pi0824 & n13231;
  assign n13872 = ~pi0871 & n13233;
  assign n13873 = ~n13871 & ~n13872;
  assign n13874 = ~pi0757 & n13193;
  assign n13875 = ~pi0696 & n13196;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = n13873 & n13876;
  assign n13878 = n13870 & n13877;
  assign n13879 = n13867 & n13878;
  assign n13880 = ~pi0634 & n13199;
  assign n13881 = ~pi0612 & n13202;
  assign n13882 = ~n13880 & ~n13881;
  assign n13883 = n13879 & n13882;
  assign n13884 = ~pi0802 & n13206;
  assign n13885 = ~pi0777 & n13209;
  assign n13886 = ~n13884 & ~n13885;
  assign n13887 = n13883 & n13886;
  assign n13888 = n13864 & n13887;
  assign po0632 = ~n13861 | ~n13888;
  assign n13890 = ~pi0825 & n13231;
  assign n13891 = ~pi0872 & n13233;
  assign n13892 = ~n13890 & ~n13891;
  assign n13893 = ~pi0573 & n13225;
  assign n13894 = ~pi0677 & n13227;
  assign n13895 = ~n13893 & ~n13894;
  assign n13896 = ~pi0849 & n13217;
  assign n13897 = ~pi0592 & n13219;
  assign n13898 = ~n13896 & ~n13897;
  assign n13899 = ~pi0801 & n13206;
  assign n13900 = ~pi0778 & n13209;
  assign n13901 = ~n13899 & ~n13900;
  assign n13902 = ~pi0946 & n13199;
  assign n13903 = ~pi0613 & n13202;
  assign n13904 = ~n13902 & ~n13903;
  assign n13905 = ~pi0739 & n13212;
  assign n13906 = ~pi0717 & n13214;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = n13904 & n13907;
  assign n13909 = n13901 & n13908;
  assign n13910 = n13898 & n13909;
  assign n13911 = ~pi0895 & n13186;
  assign n13912 = ~pi0656 & n13189;
  assign n13913 = ~n13911 & ~n13912;
  assign n13914 = n13910 & n13913;
  assign n13915 = ~pi0758 & n13193;
  assign n13916 = ~pi0697 & n13196;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = n13914 & n13917;
  assign n13919 = n13895 & n13918;
  assign po0633 = ~n13892 | ~n13919;
  assign n13921 = ~pi0969 & n13212;
  assign n13922 = ~pi0967 & n13214;
  assign n13923 = ~n13921 & ~n13922;
  assign n13924 = ~pi0963 & n13206;
  assign n13925 = ~pi0974 & n13209;
  assign n13926 = ~n13924 & ~n13925;
  assign n13927 = ~pi0973 & n13186;
  assign n13928 = ~pi0958 & n13189;
  assign n13929 = ~n13927 & ~n13928;
  assign n13930 = ~pi0964 & n13231;
  assign n13931 = ~pi0966 & n13233;
  assign n13932 = ~n13930 & ~n13931;
  assign n13933 = ~pi0971 & n13193;
  assign n13934 = ~pi0962 & n13196;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = ~pi0951 & n13225;
  assign n13937 = ~pi0961 & n13227;
  assign n13938 = ~n13936 & ~n13937;
  assign n13939 = n13935 & n13938;
  assign n13940 = n13932 & n13939;
  assign n13941 = n13929 & n13940;
  assign n13942 = ~pi0965 & n13217;
  assign n13943 = ~pi0954 & n13219;
  assign n13944 = ~n13942 & ~n13943;
  assign n13945 = n13941 & n13944;
  assign n13946 = ~pi0957 & n13199;
  assign n13947 = ~pi0955 & n13202;
  assign n13948 = ~n13946 & ~n13947;
  assign n13949 = n13945 & n13948;
  assign n13950 = n13926 & n13949;
  assign po0634 = ~n13923 | ~n13950;
  assign n13952 = ~pi1059 & n13217;
  assign n13953 = ~pi1080 & n13219;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = ~pi1005 & n13199;
  assign n13956 = ~pi1002 & n13202;
  assign n13957 = ~n13955 & ~n13956;
  assign n13958 = ~pi1092 & n13225;
  assign n13959 = ~pi1110 & n13227;
  assign n13960 = ~n13958 & ~n13959;
  assign n13961 = ~pi1052 & n13193;
  assign n13962 = ~pi1086 & n13196;
  assign n13963 = ~n13961 & ~n13962;
  assign n13964 = ~pi1043 & n13231;
  assign n13965 = ~pi1050 & n13233;
  assign n13966 = ~n13964 & ~n13965;
  assign n13967 = ~pi1055 & n13186;
  assign n13968 = ~pi1116 & n13189;
  assign n13969 = ~n13967 & ~n13968;
  assign n13970 = n13966 & n13969;
  assign n13971 = n13963 & n13970;
  assign n13972 = n13960 & n13971;
  assign n13973 = ~pi1123 & n13212;
  assign n13974 = ~pi0983 & n13214;
  assign n13975 = ~n13973 & ~n13974;
  assign n13976 = n13972 & n13975;
  assign n13977 = ~pi1082 & n13206;
  assign n13978 = ~pi1058 & n13209;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = n13976 & n13979;
  assign n13981 = n13957 & n13980;
  assign po0635 = ~n13954 | ~n13981;
  assign n13983 = ~pi0549 & n13199;
  assign n13984 = ~pi0548 & n13202;
  assign n13985 = ~n13983 & ~n13984;
  assign n13986 = ~pi0798 & n13206;
  assign n13987 = ~pi0551 & n13209;
  assign n13988 = ~n13986 & ~n13987;
  assign n13989 = ~pi0891 & n13186;
  assign n13990 = ~pi0550 & n13189;
  assign n13991 = ~n13989 & ~n13990;
  assign n13992 = ~pi0923 & n13193;
  assign n13993 = ~pi0543 & n13196;
  assign n13994 = ~n13992 & ~n13993;
  assign n13995 = ~pi0821 & n13231;
  assign n13996 = ~pi0868 & n13233;
  assign n13997 = ~n13995 & ~n13996;
  assign n13998 = ~pi0544 & n13225;
  assign n13999 = ~pi0920 & n13227;
  assign n14000 = ~n13998 & ~n13999;
  assign n14001 = n13997 & n14000;
  assign n14002 = n13994 & n14001;
  assign n14003 = n13991 & n14002;
  assign n14004 = ~pi0547 & n13212;
  assign n14005 = ~pi0546 & n13214;
  assign n14006 = ~n14004 & ~n14005;
  assign n14007 = n14003 & n14006;
  assign n14008 = ~pi0845 & n13217;
  assign n14009 = ~pi0545 & n13219;
  assign n14010 = ~n14008 & ~n14009;
  assign n14011 = n14007 & n14010;
  assign n14012 = n13988 & n14011;
  assign po0636 = ~n13985 | ~n14012;
  assign n14014 = ~pi0826 & n13217;
  assign n14015 = ~pi0909 & n13219;
  assign n14016 = ~n14014 & ~n14015;
  assign n14017 = ~pi0614 & n13199;
  assign n14018 = ~pi0593 & n13202;
  assign n14019 = ~n14017 & ~n14018;
  assign n14020 = ~pi0873 & n13186;
  assign n14021 = ~pi0635 & n13189;
  assign n14022 = ~n14020 & ~n14021;
  assign n14023 = ~pi0552 & n13225;
  assign n14024 = ~pi0943 & n13227;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = ~pi0803 & n13231;
  assign n14027 = ~pi0850 & n13233;
  assign n14028 = ~n14026 & ~n14027;
  assign n14029 = ~pi0740 & n13193;
  assign n14030 = ~pi0678 & n13196;
  assign n14031 = ~n14029 & ~n14030;
  assign n14032 = n14028 & n14031;
  assign n14033 = n14025 & n14032;
  assign n14034 = n14022 & n14033;
  assign n14035 = ~pi0718 & n13212;
  assign n14036 = ~pi0698 & n13214;
  assign n14037 = ~n14035 & ~n14036;
  assign n14038 = n14034 & n14037;
  assign n14039 = ~pi0779 & n13206;
  assign n14040 = ~pi0759 & n13209;
  assign n14041 = ~n14039 & ~n14040;
  assign n14042 = n14038 & n14041;
  assign n14043 = n14019 & n14042;
  assign po0637 = ~n14016 | ~n14043;
  assign n14045 = ~pi0924 & n13193;
  assign n14046 = ~pi0941 & n13196;
  assign n14047 = ~n14045 & ~n14046;
  assign n14048 = ~pi0874 & n13186;
  assign n14049 = ~pi0636 & n13189;
  assign n14050 = ~n14048 & ~n14049;
  assign n14051 = ~pi0922 & n13212;
  assign n14052 = ~pi0936 & n13214;
  assign n14053 = ~n14051 & ~n14052;
  assign n14054 = ~pi0780 & n13206;
  assign n14055 = ~pi0914 & n13209;
  assign n14056 = ~n14054 & ~n14055;
  assign n14057 = ~pi0827 & n13217;
  assign n14058 = ~pi0574 & n13219;
  assign n14059 = ~n14057 & ~n14058;
  assign n14060 = ~pi0615 & n13199;
  assign n14061 = ~pi0897 & n13202;
  assign n14062 = ~n14060 & ~n14061;
  assign n14063 = n14059 & n14062;
  assign n14064 = n14056 & n14063;
  assign n14065 = n14053 & n14064;
  assign n14066 = ~pi0804 & n13231;
  assign n14067 = ~pi0851 & n13233;
  assign n14068 = ~n14066 & ~n14067;
  assign n14069 = n14065 & n14068;
  assign n14070 = ~pi0553 & n13225;
  assign n14071 = ~pi0657 & n13227;
  assign n14072 = ~n14070 & ~n14071;
  assign n14073 = n14069 & n14072;
  assign n14074 = n14050 & n14073;
  assign po0638 = ~n14047 | ~n14074;
  assign n14076 = ~pi0741 & n13193;
  assign n14077 = ~pi0679 & n13196;
  assign n14078 = ~n14076 & ~n14077;
  assign n14079 = ~pi0875 & n13186;
  assign n14080 = ~pi0637 & n13189;
  assign n14081 = ~n14079 & ~n14080;
  assign n14082 = ~pi0828 & n13217;
  assign n14083 = ~pi0575 & n13219;
  assign n14084 = ~n14082 & ~n14083;
  assign n14085 = ~pi0899 & n13199;
  assign n14086 = ~pi0594 & n13202;
  assign n14087 = ~n14085 & ~n14086;
  assign n14088 = ~pi0781 & n13206;
  assign n14089 = ~pi0760 & n13209;
  assign n14090 = ~n14088 & ~n14089;
  assign n14091 = ~pi0719 & n13212;
  assign n14092 = ~pi0699 & n13214;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = n14090 & n14093;
  assign n14095 = n14087 & n14094;
  assign n14096 = n14084 & n14095;
  assign n14097 = ~pi0903 & n13231;
  assign n14098 = ~pi0516 & n13233;
  assign n14099 = ~n14097 & ~n14098;
  assign n14100 = n14096 & n14099;
  assign n14101 = ~pi0554 & n13225;
  assign n14102 = ~pi0658 & n13227;
  assign n14103 = ~n14101 & ~n14102;
  assign n14104 = n14100 & n14103;
  assign n14105 = n14081 & n14104;
  assign po0639 = ~n14078 | ~n14105;
  assign n14107 = ~pi1028 & n13212;
  assign n14108 = ~pi1023 & n13214;
  assign n14109 = ~n14107 & ~n14108;
  assign n14110 = ~pi1004 & n13199;
  assign n14111 = ~pi0999 & n13202;
  assign n14112 = ~n14110 & ~n14111;
  assign n14113 = ~pi1096 & n13225;
  assign n14114 = ~pi1115 & n13227;
  assign n14115 = ~n14113 & ~n14114;
  assign n14116 = ~pi1030 & n13193;
  assign n14117 = ~pi1016 & n13196;
  assign n14118 = ~n14116 & ~n14117;
  assign n14119 = ~pi1042 & n13231;
  assign n14120 = ~pi1048 & n13233;
  assign n14121 = ~n14119 & ~n14120;
  assign n14122 = ~pi1053 & n13186;
  assign n14123 = ~pi1008 & n13189;
  assign n14124 = ~n14122 & ~n14123;
  assign n14125 = n14121 & n14124;
  assign n14126 = n14118 & n14125;
  assign n14127 = n14115 & n14126;
  assign n14128 = ~pi1045 & n13217;
  assign n14129 = ~pi1088 & n13219;
  assign n14130 = ~n14128 & ~n14129;
  assign n14131 = n14127 & n14130;
  assign n14132 = ~pi1040 & n13206;
  assign n14133 = ~pi1035 & n13209;
  assign n14134 = ~n14132 & ~n14133;
  assign n14135 = n14131 & n14134;
  assign n14136 = n14112 & n14135;
  assign po0640 = ~n14109 | ~n14136;
  assign n14138 = ~pi0742 & n13193;
  assign n14139 = ~pi0680 & n13196;
  assign n14140 = ~n14138 & ~n14139;
  assign n14141 = ~pi0805 & n13231;
  assign n14142 = ~pi0852 & n13233;
  assign n14143 = ~n14141 & ~n14142;
  assign n14144 = ~pi0720 & n13212;
  assign n14145 = ~pi0700 & n13214;
  assign n14146 = ~n14144 & ~n14145;
  assign n14147 = ~pi0782 & n13206;
  assign n14148 = ~pi0761 & n13209;
  assign n14149 = ~n14147 & ~n14148;
  assign n14150 = ~pi0829 & n13217;
  assign n14151 = ~pi0576 & n13219;
  assign n14152 = ~n14150 & ~n14151;
  assign n14153 = ~pi0616 & n13199;
  assign n14154 = ~pi0595 & n13202;
  assign n14155 = ~n14153 & ~n14154;
  assign n14156 = n14152 & n14155;
  assign n14157 = n14149 & n14156;
  assign n14158 = n14146 & n14157;
  assign n14159 = ~pi0876 & n13186;
  assign n14160 = ~pi0638 & n13189;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = n14158 & n14161;
  assign n14163 = ~pi0555 & n13225;
  assign n14164 = ~pi0659 & n13227;
  assign n14165 = ~n14163 & ~n14164;
  assign n14166 = n14162 & n14165;
  assign n14167 = n14143 & n14166;
  assign po0641 = ~n14140 | ~n14167;
  assign n14169 = ~pi1125 & n13186;
  assign n14170 = ~pi1009 & n13189;
  assign n14171 = ~n14169 & ~n14170;
  assign n14172 = ~pi1098 & n13193;
  assign n14173 = ~pi1017 & n13196;
  assign n14174 = ~n14172 & ~n14173;
  assign n14175 = ~pi1068 & n13217;
  assign n14176 = ~pi0994 & n13219;
  assign n14177 = ~n14175 & ~n14176;
  assign n14178 = ~pi1061 & n13199;
  assign n14179 = ~pi1073 & n13202;
  assign n14180 = ~n14178 & ~n14179;
  assign n14181 = ~pi1104 & n13212;
  assign n14182 = ~pi1107 & n13214;
  assign n14183 = ~n14181 & ~n14182;
  assign n14184 = ~pi1089 & n13206;
  assign n14185 = ~pi1093 & n13209;
  assign n14186 = ~n14184 & ~n14185;
  assign n14187 = n14183 & n14186;
  assign n14188 = n14180 & n14187;
  assign n14189 = n14177 & n14188;
  assign n14190 = ~pi1079 & n13231;
  assign n14191 = ~pi0989 & n13233;
  assign n14192 = ~n14190 & ~n14191;
  assign n14193 = n14189 & n14192;
  assign n14194 = ~pi1095 & n13225;
  assign n14195 = ~pi1114 & n13227;
  assign n14196 = ~n14194 & ~n14195;
  assign n14197 = n14193 & n14196;
  assign n14198 = n14174 & n14197;
  assign po0642 = ~n14171 | ~n14198;
  assign n14200 = ~pi0977 & n13231;
  assign n14201 = ~pi0950 & n13233;
  assign n14202 = ~n14200 & ~n14201;
  assign n14203 = ~pi0952 & n13225;
  assign n14204 = ~pi0960 & n13227;
  assign n14205 = ~n14203 & ~n14204;
  assign n14206 = ~pi0976 & n13217;
  assign n14207 = ~pi0953 & n13219;
  assign n14208 = ~n14206 & ~n14207;
  assign n14209 = ~pi0982 & n13199;
  assign n14210 = ~pi0956 & n13202;
  assign n14211 = ~n14209 & ~n14210;
  assign n14212 = ~pi0978 & n13206;
  assign n14213 = ~pi0980 & n13209;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = ~pi0970 & n13212;
  assign n14216 = ~pi0968 & n13214;
  assign n14217 = ~n14215 & ~n14216;
  assign n14218 = n14214 & n14217;
  assign n14219 = n14211 & n14218;
  assign n14220 = n14208 & n14219;
  assign n14221 = ~pi0981 & n13186;
  assign n14222 = ~pi0959 & n13189;
  assign n14223 = ~n14221 & ~n14222;
  assign n14224 = n14220 & n14223;
  assign n14225 = ~pi0972 & n13193;
  assign n14226 = ~pi0979 & n13196;
  assign n14227 = ~n14225 & ~n14226;
  assign n14228 = n14224 & n14227;
  assign n14229 = n14205 & n14228;
  assign po0643 = ~n14202 | ~n14229;
  assign n14231 = ~pi1203 & n13217;
  assign n14232 = ~pi1204 & n13219;
  assign n14233 = ~n14231 & ~n14232;
  assign n14234 = ~pi1199 & n13212;
  assign n14235 = ~pi1198 & n13214;
  assign n14236 = ~n14234 & ~n14235;
  assign n14237 = ~pi1207 & n13193;
  assign n14238 = ~pi1188 & n13196;
  assign n14239 = ~n14237 & ~n14238;
  assign n14240 = ~pi1197 & n13225;
  assign n14241 = ~pi1173 & n13227;
  assign n14242 = ~n14240 & ~n14241;
  assign n14243 = ~pi1202 & n13231;
  assign n14244 = ~pi1205 & n13233;
  assign n14245 = ~n14243 & ~n14244;
  assign n14246 = ~pi1174 & n13186;
  assign n14247 = ~pi1201 & n13189;
  assign n14248 = ~n14246 & ~n14247;
  assign n14249 = n14245 & n14248;
  assign n14250 = n14242 & n14249;
  assign n14251 = n14239 & n14250;
  assign n14252 = ~pi1190 & n13206;
  assign n14253 = ~pi1189 & n13209;
  assign n14254 = ~n14252 & ~n14253;
  assign n14255 = n14251 & n14254;
  assign n14256 = ~pi1206 & n13199;
  assign n14257 = ~pi1200 & n13202;
  assign n14258 = ~n14256 & ~n14257;
  assign n14259 = n14255 & n14258;
  assign n14260 = n14236 & n14259;
  assign po0644 = ~n14233 | ~n14260;
  assign n14262 = ~pi0623 & n13199;
  assign n14263 = ~pi0901 & n13202;
  assign n14264 = ~n14262 & ~n14263;
  assign n14265 = ~pi0836 & n13217;
  assign n14266 = ~pi0906 & n13219;
  assign n14267 = ~n14265 & ~n14266;
  assign n14268 = ~pi0948 & n13186;
  assign n14269 = ~pi0644 & n13189;
  assign n14270 = ~n14268 & ~n14269;
  assign n14271 = ~pi0918 & n13193;
  assign n14272 = ~pi0687 & n13196;
  assign n14273 = ~n14271 & ~n14272;
  assign n14274 = ~pi0562 & n13225;
  assign n14275 = ~pi0666 & n13227;
  assign n14276 = ~n14274 & ~n14275;
  assign n14277 = ~pi0812 & n13231;
  assign n14278 = ~pi0859 & n13233;
  assign n14279 = ~n14277 & ~n14278;
  assign n14280 = n14276 & n14279;
  assign n14281 = n14273 & n14280;
  assign n14282 = n14270 & n14281;
  assign n14283 = ~pi0789 & n13206;
  assign n14284 = ~pi0768 & n13209;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = n14282 & n14285;
  assign n14287 = ~pi0726 & n13212;
  assign n14288 = ~pi0707 & n13214;
  assign n14289 = ~n14287 & ~n14288;
  assign n14290 = n14286 & n14289;
  assign n14291 = n14267 & n14290;
  assign po0646 = ~n14264 | ~n14291;
  assign n14293 = ~pi1126 & n13199;
  assign n14294 = ~pi1069 & n13202;
  assign n14295 = ~n14293 & ~n14294;
  assign n14296 = ~pi1081 & n13206;
  assign n14297 = ~pi1075 & n13209;
  assign n14298 = ~n14296 & ~n14297;
  assign n14299 = ~pi1097 & n13193;
  assign n14300 = ~pi1108 & n13196;
  assign n14301 = ~n14299 & ~n14300;
  assign n14302 = ~pi1124 & n13186;
  assign n14303 = ~pi1113 & n13189;
  assign n14304 = ~n14302 & ~n14303;
  assign n14305 = ~pi0991 & n13225;
  assign n14306 = ~pi1013 & n13227;
  assign n14307 = ~n14305 & ~n14306;
  assign n14308 = ~pi1074 & n13231;
  assign n14309 = ~pi0987 & n13233;
  assign n14310 = ~n14308 & ~n14309;
  assign n14311 = n14307 & n14310;
  assign n14312 = n14304 & n14311;
  assign n14313 = n14301 & n14312;
  assign n14314 = ~pi1064 & n13217;
  assign n14315 = ~pi1084 & n13219;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = n14313 & n14316;
  assign n14318 = ~pi1102 & n13212;
  assign n14319 = ~pi1106 & n13214;
  assign n14320 = ~n14318 & ~n14319;
  assign n14321 = n14317 & n14320;
  assign n14322 = n14298 & n14321;
  assign po0647 = ~n14295 | ~n14322;
  assign n14324 = ~pi0843 & n13217;
  assign n14325 = ~pi0587 & n13219;
  assign n14326 = ~n14324 & ~n14325;
  assign n14327 = ~pi0733 & n13212;
  assign n14328 = ~pi0713 & n13214;
  assign n14329 = ~n14327 & ~n14328;
  assign n14330 = ~pi0889 & n13186;
  assign n14331 = ~pi0651 & n13189;
  assign n14332 = ~n14330 & ~n14331;
  assign n14333 = ~pi0754 & n13193;
  assign n14334 = ~pi0693 & n13196;
  assign n14335 = ~n14333 & ~n14334;
  assign n14336 = ~pi0568 & n13225;
  assign n14337 = ~pi0672 & n13227;
  assign n14338 = ~n14336 & ~n14337;
  assign n14339 = ~pi0819 & n13231;
  assign n14340 = ~pi0866 & n13233;
  assign n14341 = ~n14339 & ~n14340;
  assign n14342 = n14338 & n14341;
  assign n14343 = n14335 & n14342;
  assign n14344 = n14332 & n14343;
  assign n14345 = ~pi0630 & n13199;
  assign n14346 = ~pi0608 & n13202;
  assign n14347 = ~n14345 & ~n14346;
  assign n14348 = n14344 & n14347;
  assign n14349 = ~pi0796 & n13206;
  assign n14350 = ~pi0774 & n13209;
  assign n14351 = ~n14349 & ~n14350;
  assign n14352 = n14348 & n14351;
  assign n14353 = n14329 & n14352;
  assign po0648 = ~n14326 | ~n14353;
  assign n14355 = n8038 & n12553;
  assign n14356 = pi2553 & n14355;
  assign n14357 = pi2963 & n14356;
  assign n14358 = ~n12558 & ~n14357;
  assign n14359 = pi2963 & n8038;
  assign n14360 = pi2553 & n14359;
  assign n14361 = n8046 & n14360;
  assign n14362 = ~n8036 & n14361;
  assign n14363 = n14358 & ~n14362;
  assign n14364 = ~n8057 & ~n14363;
  assign n14365 = ~pi1180 & n14364;
  assign n14366 = ~pi1221 & ~n14364;
  assign n14367 = ~n14365 & ~n14366;
  assign n14368 = ~pi1213 & ~n14364;
  assign n14369 = ~pi1211 & n14364;
  assign n14370 = ~n14368 & ~n14369;
  assign n14371 = ~pi1212 & ~n14364;
  assign n14372 = pi1224 & n14364;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = ~n14370 & n14373;
  assign n14375 = ~n14367 & n14374;
  assign n14376 = ~pi1635 & n14375;
  assign n14377 = n14367 & n14374;
  assign n14378 = ~pi1421 & n14377;
  assign n14379 = ~n14376 & ~n14378;
  assign n14380 = n14370 & ~n14373;
  assign n14381 = ~n14367 & n14380;
  assign n14382 = ~pi1543 & n14381;
  assign n14383 = n14367 & n14380;
  assign n14384 = ~pi1578 & n14383;
  assign n14385 = ~n14382 & ~n14384;
  assign n14386 = ~n14370 & ~n14373;
  assign n14387 = ~n14367 & n14386;
  assign n14388 = ~pi1484 & n14387;
  assign n14389 = n14367 & n14386;
  assign n14390 = ~pi1462 & n14389;
  assign n14391 = ~n14388 & ~n14390;
  assign n14392 = n14370 & n14373;
  assign n14393 = ~n14367 & n14392;
  assign n14394 = ~pi1503 & n14393;
  assign n14395 = n14367 & n14392;
  assign n14396 = ~pi1633 & n14395;
  assign n14397 = ~n14394 & ~n14396;
  assign n14398 = n14391 & n14397;
  assign n14399 = n14385 & n14398;
  assign po0649 = ~n14379 | ~n14399;
  assign n14401 = ~pi1496 & n14393;
  assign n14402 = ~pi1557 & n14395;
  assign n14403 = ~n14401 & ~n14402;
  assign n14404 = ~pi1434 & n14375;
  assign n14405 = ~pi1660 & n14377;
  assign n14406 = ~n14404 & ~n14405;
  assign n14407 = ~pi1477 & n14387;
  assign n14408 = ~pi1623 & n14389;
  assign n14409 = ~n14407 & ~n14408;
  assign n14410 = ~pi1394 & n14381;
  assign n14411 = ~pi1517 & n14383;
  assign n14412 = ~n14410 & ~n14411;
  assign n14413 = n14409 & n14412;
  assign n14414 = n14406 & n14413;
  assign po0650 = ~n14403 | ~n14414;
  assign n14416 = ~pi1648 & n14381;
  assign n14417 = ~pi1531 & n14383;
  assign n14418 = ~n14416 & ~n14417;
  assign n14419 = ~pi1449 & n14375;
  assign n14420 = ~pi1649 & n14377;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = ~pi1493 & n14387;
  assign n14423 = ~pi1471 & n14389;
  assign n14424 = ~n14422 & ~n14423;
  assign n14425 = ~pi1511 & n14393;
  assign n14426 = ~pi1572 & n14395;
  assign n14427 = ~n14425 & ~n14426;
  assign n14428 = n14424 & n14427;
  assign n14429 = n14421 & n14428;
  assign po0651 = ~n14418 | ~n14429;
  assign n14431 = ~pi1538 & n14381;
  assign n14432 = ~pi1518 & n14383;
  assign n14433 = ~n14431 & ~n14432;
  assign n14434 = ~pi1598 & n14393;
  assign n14435 = ~pi1558 & n14395;
  assign n14436 = ~n14434 & ~n14435;
  assign n14437 = ~pi1478 & n14387;
  assign n14438 = ~pi1621 & n14389;
  assign n14439 = ~n14437 & ~n14438;
  assign n14440 = ~pi1436 & n14375;
  assign n14441 = ~pi1659 & n14377;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = n14439 & n14442;
  assign n14444 = n14436 & n14443;
  assign po0653 = ~n14433 | ~n14444;
  assign n14446 = ~pi1539 & n14381;
  assign n14447 = ~pi1519 & n14383;
  assign n14448 = ~n14446 & ~n14447;
  assign n14449 = ~pi1498 & n14393;
  assign n14450 = ~pi1637 & n14395;
  assign n14451 = ~n14449 & ~n14450;
  assign n14452 = ~pi1640 & n14375;
  assign n14453 = ~pi1416 & n14377;
  assign n14454 = ~n14452 & ~n14453;
  assign n14455 = ~pi1479 & n14387;
  assign n14456 = ~pi1457 & n14389;
  assign n14457 = ~n14455 & ~n14456;
  assign n14458 = n14454 & n14457;
  assign n14459 = n14451 & n14458;
  assign po0654 = ~n14448 | ~n14459;
  assign n14461 = ~pi1609 & n14387;
  assign n14462 = ~pi1456 & n14389;
  assign n14463 = ~n14461 & ~n14462;
  assign n14464 = ~pi1537 & n14381;
  assign n14465 = ~pi1583 & n14383;
  assign n14466 = ~n14464 & ~n14465;
  assign n14467 = ~pi1497 & n14393;
  assign n14468 = ~pi1639 & n14395;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = ~pi1435 & n14375;
  assign n14471 = ~pi1415 & n14377;
  assign n14472 = ~n14470 & ~n14471;
  assign n14473 = n14469 & n14472;
  assign n14474 = n14466 & n14473;
  assign po0655 = ~n14463 | ~n14474;
  assign n14476 = ~pi1437 & n14375;
  assign n14477 = ~pi1658 & n14377;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = ~pi1389 & n14381;
  assign n14480 = ~pi1520 & n14383;
  assign n14481 = ~n14479 & ~n14480;
  assign n14482 = ~pi1596 & n14393;
  assign n14483 = ~pi1559 & n14395;
  assign n14484 = ~n14482 & ~n14483;
  assign n14485 = ~pi1480 & n14387;
  assign n14486 = ~pi1458 & n14389;
  assign n14487 = ~n14485 & ~n14486;
  assign n14488 = n14484 & n14487;
  assign n14489 = n14481 & n14488;
  assign po0656 = ~n14478 | ~n14489;
  assign n14491 = ~pi1540 & n14381;
  assign n14492 = ~pi1582 & n14383;
  assign n14493 = ~n14491 & ~n14492;
  assign n14494 = ~pi1380 & n14387;
  assign n14495 = ~pi1459 & n14389;
  assign n14496 = ~n14494 & ~n14495;
  assign n14497 = ~pi1499 & n14393;
  assign n14498 = ~pi1560 & n14395;
  assign n14499 = ~n14497 & ~n14498;
  assign n14500 = ~pi1438 & n14375;
  assign n14501 = ~pi1417 & n14377;
  assign n14502 = ~n14500 & ~n14501;
  assign n14503 = n14499 & n14502;
  assign n14504 = n14496 & n14503;
  assign po0657 = ~n14493 | ~n14504;
  assign n14506 = ~pi1481 & n14387;
  assign n14507 = ~pi1618 & n14389;
  assign n14508 = ~n14506 & ~n14507;
  assign n14509 = ~pi1597 & n14393;
  assign n14510 = ~pi1561 & n14395;
  assign n14511 = ~n14509 & ~n14510;
  assign n14512 = ~pi1390 & n14381;
  assign n14513 = ~pi1521 & n14383;
  assign n14514 = ~n14512 & ~n14513;
  assign n14515 = ~pi1439 & n14375;
  assign n14516 = ~pi1418 & n14377;
  assign n14517 = ~n14515 & ~n14516;
  assign n14518 = n14514 & n14517;
  assign n14519 = n14511 & n14518;
  assign po0658 = ~n14508 | ~n14519;
  assign n14521 = ~pi1588 & n14387;
  assign n14522 = ~pi1460 & n14389;
  assign n14523 = ~n14521 & ~n14522;
  assign n14524 = ~pi1644 & n14375;
  assign n14525 = ~pi1419 & n14377;
  assign n14526 = ~n14524 & ~n14525;
  assign n14527 = ~pi1500 & n14393;
  assign n14528 = ~pi1628 & n14395;
  assign n14529 = ~n14527 & ~n14528;
  assign n14530 = ~pi1541 & n14381;
  assign n14531 = ~pi1581 & n14383;
  assign n14532 = ~n14530 & ~n14531;
  assign n14533 = n14529 & n14532;
  assign n14534 = n14526 & n14533;
  assign po0659 = ~n14523 | ~n14534;
  assign n14536 = ~pi1542 & n14381;
  assign n14537 = ~pi1580 & n14383;
  assign n14538 = ~n14536 & ~n14537;
  assign n14539 = ~pi1502 & n14393;
  assign n14540 = ~pi1634 & n14395;
  assign n14541 = ~n14539 & ~n14540;
  assign n14542 = ~pi1641 & n14375;
  assign n14543 = ~pi1420 & n14377;
  assign n14544 = ~n14542 & ~n14543;
  assign n14545 = ~pi1604 & n14387;
  assign n14546 = ~pi1461 & n14389;
  assign n14547 = ~n14545 & ~n14546;
  assign n14548 = n14544 & n14547;
  assign n14549 = n14541 & n14548;
  assign po0660 = ~n14538 | ~n14549;
  assign n14551 = ~pi1388 & n14381;
  assign n14552 = ~pi1523 & n14383;
  assign n14553 = ~n14551 & ~n14552;
  assign n14554 = ~pi1594 & n14393;
  assign n14555 = ~pi1563 & n14395;
  assign n14556 = ~n14554 & ~n14555;
  assign n14557 = ~pi1483 & n14387;
  assign n14558 = ~pi1614 & n14389;
  assign n14559 = ~n14557 & ~n14558;
  assign n14560 = ~pi1441 & n14375;
  assign n14561 = ~pi1656 & n14377;
  assign n14562 = ~n14560 & ~n14561;
  assign n14563 = n14559 & n14562;
  assign n14564 = n14556 & n14563;
  assign po0661 = ~n14553 | ~n14564;
  assign n14566 = ~pi1440 & n14375;
  assign n14567 = ~pi1655 & n14377;
  assign n14568 = ~n14566 & ~n14567;
  assign n14569 = ~pi1482 & n14387;
  assign n14570 = ~pi1615 & n14389;
  assign n14571 = ~n14569 & ~n14570;
  assign n14572 = ~pi1387 & n14381;
  assign n14573 = ~pi1522 & n14383;
  assign n14574 = ~n14572 & ~n14573;
  assign n14575 = ~pi1501 & n14393;
  assign n14576 = ~pi1562 & n14395;
  assign n14577 = ~n14575 & ~n14576;
  assign n14578 = n14574 & n14577;
  assign n14579 = n14571 & n14578;
  assign po0662 = ~n14568 | ~n14579;
  assign n14581 = ~pi1485 & n14387;
  assign n14582 = ~pi1463 & n14389;
  assign n14583 = ~n14581 & ~n14582;
  assign n14584 = ~pi1587 & n14393;
  assign n14585 = ~pi1564 & n14395;
  assign n14586 = ~n14584 & ~n14585;
  assign n14587 = ~pi1384 & n14381;
  assign n14588 = ~pi1524 & n14383;
  assign n14589 = ~n14587 & ~n14588;
  assign n14590 = ~pi1442 & n14375;
  assign n14591 = ~pi1654 & n14377;
  assign n14592 = ~n14590 & ~n14591;
  assign n14593 = n14589 & n14592;
  assign n14594 = n14586 & n14593;
  assign po0663 = ~n14583 | ~n14594;
  assign n14596 = ~pi1603 & n14387;
  assign n14597 = ~pi1464 & n14389;
  assign n14598 = ~n14596 & ~n14597;
  assign n14599 = ~pi1544 & n14381;
  assign n14600 = ~pi1579 & n14383;
  assign n14601 = ~n14599 & ~n14600;
  assign n14602 = ~pi1504 & n14393;
  assign n14603 = ~pi1565 & n14395;
  assign n14604 = ~n14602 & ~n14603;
  assign n14605 = ~pi1638 & n14375;
  assign n14606 = ~pi1422 & n14377;
  assign n14607 = ~n14605 & ~n14606;
  assign n14608 = n14604 & n14607;
  assign n14609 = n14601 & n14608;
  assign po0664 = ~n14598 | ~n14609;
  assign n14611 = ~pi1545 & n14381;
  assign n14612 = ~pi1525 & n14383;
  assign n14613 = ~n14611 & ~n14612;
  assign n14614 = ~pi1486 & n14387;
  assign n14615 = ~pi1607 & n14389;
  assign n14616 = ~n14614 & ~n14615;
  assign n14617 = ~pi1443 & n14375;
  assign n14618 = ~pi1650 & n14377;
  assign n14619 = ~n14617 & ~n14618;
  assign n14620 = ~pi1593 & n14393;
  assign n14621 = ~pi1566 & n14395;
  assign n14622 = ~n14620 & ~n14621;
  assign n14623 = n14619 & n14622;
  assign n14624 = n14616 & n14623;
  assign po0665 = ~n14613 | ~n14624;
  assign n14626 = ~pi1505 & n14393;
  assign n14627 = ~pi1630 & n14395;
  assign n14628 = ~n14626 & ~n14627;
  assign n14629 = ~pi1487 & n14387;
  assign n14630 = ~pi1465 & n14389;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~pi1624 & n14375;
  assign n14633 = ~pi1423 & n14377;
  assign n14634 = ~n14632 & ~n14633;
  assign n14635 = ~pi1546 & n14381;
  assign n14636 = ~pi1526 & n14383;
  assign n14637 = ~n14635 & ~n14636;
  assign n14638 = n14634 & n14637;
  assign n14639 = n14631 & n14638;
  assign po0666 = ~n14628 | ~n14639;
  assign n14641 = ~pi1444 & n14375;
  assign n14642 = ~pi1651 & n14377;
  assign n14643 = ~n14641 & ~n14642;
  assign n14644 = ~pi1488 & n14387;
  assign n14645 = ~pi1612 & n14389;
  assign n14646 = ~n14644 & ~n14645;
  assign n14647 = ~pi1386 & n14381;
  assign n14648 = ~pi1527 & n14383;
  assign n14649 = ~n14647 & ~n14648;
  assign n14650 = ~pi1506 & n14393;
  assign n14651 = ~pi1567 & n14395;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = n14649 & n14652;
  assign n14654 = n14646 & n14653;
  assign po0667 = ~n14643 | ~n14654;
  assign n14656 = ~pi1547 & n14381;
  assign n14657 = ~pi1576 & n14383;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~pi1507 & n14393;
  assign n14660 = ~pi1629 & n14395;
  assign n14661 = ~n14659 & ~n14660;
  assign n14662 = ~pi1602 & n14387;
  assign n14663 = ~pi1466 & n14389;
  assign n14664 = ~n14662 & ~n14663;
  assign n14665 = ~pi1631 & n14375;
  assign n14666 = ~pi1424 & n14377;
  assign n14667 = ~n14665 & ~n14666;
  assign n14668 = n14664 & n14667;
  assign n14669 = n14661 & n14668;
  assign po0668 = ~n14658 | ~n14669;
  assign n14671 = ~pi1592 & n14393;
  assign n14672 = ~pi1568 & n14395;
  assign n14673 = ~n14671 & ~n14672;
  assign n14674 = ~pi1489 & n14387;
  assign n14675 = ~pi1613 & n14389;
  assign n14676 = ~n14674 & ~n14675;
  assign n14677 = ~pi1445 & n14375;
  assign n14678 = ~pi1653 & n14377;
  assign n14679 = ~n14677 & ~n14678;
  assign n14680 = ~pi1385 & n14381;
  assign n14681 = ~pi1528 & n14383;
  assign n14682 = ~n14680 & ~n14681;
  assign n14683 = n14679 & n14682;
  assign n14684 = n14676 & n14683;
  assign po0669 = ~n14673 | ~n14684;
  assign n14686 = ~pi1446 & n14375;
  assign n14687 = ~pi1652 & n14377;
  assign n14688 = ~n14686 & ~n14687;
  assign n14689 = ~pi1590 & n14393;
  assign n14690 = ~pi1569 & n14395;
  assign n14691 = ~n14689 & ~n14690;
  assign n14692 = ~pi1382 & n14381;
  assign n14693 = ~pi1529 & n14383;
  assign n14694 = ~n14692 & ~n14693;
  assign n14695 = ~pi1491 & n14387;
  assign n14696 = ~pi1468 & n14389;
  assign n14697 = ~n14695 & ~n14696;
  assign n14698 = n14694 & n14697;
  assign n14699 = n14691 & n14698;
  assign po0670 = ~n14688 | ~n14699;
  assign n14701 = ~pi1447 & n14375;
  assign n14702 = ~pi1426 & n14377;
  assign n14703 = ~n14701 & ~n14702;
  assign n14704 = ~pi1599 & n14387;
  assign n14705 = ~pi1469 & n14389;
  assign n14706 = ~n14704 & ~n14705;
  assign n14707 = ~pi1509 & n14393;
  assign n14708 = ~pi1570 & n14395;
  assign n14709 = ~n14707 & ~n14708;
  assign n14710 = ~pi1549 & n14381;
  assign n14711 = ~pi1398 & n14383;
  assign n14712 = ~n14710 & ~n14711;
  assign n14713 = n14709 & n14712;
  assign n14714 = n14706 & n14713;
  assign po0671 = ~n14703 | ~n14714;
  assign n14716 = ~pi1591 & n14393;
  assign n14717 = ~pi1571 & n14395;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = ~pi1448 & n14375;
  assign n14720 = ~pi1427 & n14377;
  assign n14721 = ~n14719 & ~n14720;
  assign n14722 = ~pi1550 & n14381;
  assign n14723 = ~pi1530 & n14383;
  assign n14724 = ~n14722 & ~n14723;
  assign n14725 = ~pi1492 & n14387;
  assign n14726 = ~pi1611 & n14389;
  assign n14727 = ~n14725 & ~n14726;
  assign n14728 = n14724 & n14727;
  assign n14729 = n14721 & n14728;
  assign po0672 = ~n14718 | ~n14729;
  assign n14731 = ~pi1601 & n14387;
  assign n14732 = ~pi1470 & n14389;
  assign n14733 = ~n14731 & ~n14732;
  assign n14734 = ~pi1510 & n14393;
  assign n14735 = ~pi1625 & n14395;
  assign n14736 = ~n14734 & ~n14735;
  assign n14737 = ~pi1551 & n14381;
  assign n14738 = ~pi1381 & n14383;
  assign n14739 = ~n14737 & ~n14738;
  assign n14740 = ~pi1626 & n14375;
  assign n14741 = ~pi1428 & n14377;
  assign n14742 = ~n14740 & ~n14741;
  assign n14743 = n14739 & n14742;
  assign n14744 = n14736 & n14743;
  assign po0673 = ~n14733 | ~n14744;
  assign n14746 = ~pi1450 & n14375;
  assign n14747 = ~pi1429 & n14377;
  assign n14748 = ~n14746 & ~n14747;
  assign n14749 = ~pi1512 & n14393;
  assign n14750 = ~pi1605 & n14395;
  assign n14751 = ~n14749 & ~n14750;
  assign n14752 = ~pi1552 & n14381;
  assign n14753 = ~pi1393 & n14383;
  assign n14754 = ~n14752 & ~n14753;
  assign n14755 = ~pi1600 & n14387;
  assign n14756 = ~pi1472 & n14389;
  assign n14757 = ~n14755 & ~n14756;
  assign n14758 = n14754 & n14757;
  assign n14759 = n14751 & n14758;
  assign po0674 = ~n14748 | ~n14759;
  assign n14761 = ~pi1494 & n14387;
  assign n14762 = ~pi1606 & n14389;
  assign n14763 = ~n14761 & ~n14762;
  assign n14764 = ~pi1451 & n14375;
  assign n14765 = ~pi1647 & n14377;
  assign n14766 = ~n14764 & ~n14765;
  assign n14767 = ~pi1584 & n14393;
  assign n14768 = ~pi1573 & n14395;
  assign n14769 = ~n14767 & ~n14768;
  assign n14770 = ~pi1553 & n14381;
  assign n14771 = ~pi1532 & n14383;
  assign n14772 = ~n14770 & ~n14771;
  assign n14773 = n14769 & n14772;
  assign n14774 = n14766 & n14773;
  assign po0675 = ~n14763 | ~n14774;
  assign n14776 = ~pi1490 & n14387;
  assign n14777 = ~pi1467 & n14389;
  assign n14778 = ~n14776 & ~n14777;
  assign n14779 = ~pi1548 & n14381;
  assign n14780 = ~pi1577 & n14383;
  assign n14781 = ~n14779 & ~n14780;
  assign n14782 = ~pi1632 & n14375;
  assign n14783 = ~pi1425 & n14377;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = ~pi1508 & n14393;
  assign n14786 = ~pi1627 & n14395;
  assign n14787 = ~n14785 & ~n14786;
  assign n14788 = n14784 & n14787;
  assign n14789 = n14781 & n14788;
  assign po0676 = ~n14778 | ~n14789;
  assign n14791 = ~pi1430 & n14375;
  assign n14792 = ~pi1411 & n14377;
  assign n14793 = ~n14791 & ~n14792;
  assign n14794 = ~pi1617 & n14393;
  assign n14795 = ~pi1554 & n14395;
  assign n14796 = ~n14794 & ~n14795;
  assign n14797 = ~pi1392 & n14381;
  assign n14798 = ~pi1513 & n14383;
  assign n14799 = ~n14797 & ~n14798;
  assign n14800 = ~pi1473 & n14387;
  assign n14801 = ~pi1616 & n14389;
  assign n14802 = ~n14800 & ~n14801;
  assign n14803 = n14799 & n14802;
  assign n14804 = n14796 & n14803;
  assign po0677 = ~n14793 | ~n14804;
  assign n14806 = ~pi1574 & n14393;
  assign n14807 = ~pi1636 & n14395;
  assign n14808 = ~n14806 & ~n14807;
  assign n14809 = ~pi1533 & n14381;
  assign n14810 = ~pi1585 & n14383;
  assign n14811 = ~n14809 & ~n14810;
  assign n14812 = ~pi1646 & n14375;
  assign n14813 = ~pi1412 & n14377;
  assign n14814 = ~n14812 & ~n14813;
  assign n14815 = ~pi1474 & n14387;
  assign n14816 = ~pi1452 & n14389;
  assign n14817 = ~n14815 & ~n14816;
  assign n14818 = n14814 & n14817;
  assign n14819 = n14811 & n14818;
  assign po0678 = ~n14808 | ~n14819;
  assign n14821 = ~pi1475 & n14387;
  assign n14822 = ~pi1453 & n14389;
  assign n14823 = ~n14821 & ~n14822;
  assign n14824 = ~pi1391 & n14381;
  assign n14825 = ~pi1514 & n14383;
  assign n14826 = ~n14824 & ~n14825;
  assign n14827 = ~pi1431 & n14375;
  assign n14828 = ~pi1661 & n14377;
  assign n14829 = ~n14827 & ~n14828;
  assign n14830 = ~pi1619 & n14393;
  assign n14831 = ~pi1555 & n14395;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = n14829 & n14832;
  assign n14834 = n14826 & n14833;
  assign po0679 = ~n14823 | ~n14834;
  assign n14836 = ~pi1610 & n14387;
  assign n14837 = ~pi1454 & n14389;
  assign n14838 = ~n14836 & ~n14837;
  assign n14839 = ~pi1534 & n14381;
  assign n14840 = ~pi1586 & n14383;
  assign n14841 = ~n14839 & ~n14840;
  assign n14842 = ~pi1575 & n14393;
  assign n14843 = ~pi1642 & n14395;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = ~pi1432 & n14375;
  assign n14846 = ~pi1413 & n14377;
  assign n14847 = ~n14845 & ~n14846;
  assign n14848 = n14844 & n14847;
  assign n14849 = n14841 & n14848;
  assign po0680 = ~n14838 | ~n14849;
  assign n14851 = ~pi1476 & n14387;
  assign n14852 = ~pi1620 & n14389;
  assign n14853 = ~n14851 & ~n14852;
  assign n14854 = ~pi1535 & n14381;
  assign n14855 = ~pi1515 & n14383;
  assign n14856 = ~n14854 & ~n14855;
  assign n14857 = ~pi1622 & n14393;
  assign n14858 = ~pi1556 & n14395;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = ~pi1433 & n14375;
  assign n14861 = ~pi1657 & n14377;
  assign n14862 = ~n14860 & ~n14861;
  assign n14863 = n14859 & n14862;
  assign n14864 = n14856 & n14863;
  assign po0681 = ~n14853 | ~n14864;
  assign n14866 = ~pi1645 & n14375;
  assign n14867 = ~pi1414 & n14377;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = ~pi1536 & n14381;
  assign n14870 = ~pi1516 & n14383;
  assign n14871 = ~n14869 & ~n14870;
  assign n14872 = ~pi1495 & n14393;
  assign n14873 = ~pi1643 & n14395;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = ~pi1608 & n14387;
  assign n14876 = ~pi1455 & n14389;
  assign n14877 = ~n14875 & ~n14876;
  assign n14878 = n14874 & n14877;
  assign n14879 = n14871 & n14878;
  assign po0682 = ~n14868 | ~n14879;
  assign n14881 = pi3361 & pi3362;
  assign n14882 = n8177 & n14881;
  assign n14883 = pi2465 & n14882;
  assign n14884 = pi0988 & n14883;
  assign n14885 = n8200 & n8296;
  assign n14886 = ~n8277 & ~n8294;
  assign n14887 = n14885 & ~n14886;
  assign n14888 = n8194 & ~n8206;
  assign n14889 = n8198 & n14888;
  assign n14890 = ~n8201 & n14889;
  assign n14891 = ~n14887 & ~n14890;
  assign n14892 = ~pi2465 & n14881;
  assign n14893 = ~n11017 & n14892;
  assign n14894 = n14891 & ~n14893;
  assign n14895 = ~n11005 & ~n11012;
  assign n14896 = n8200 & ~n14895;
  assign n14897 = ~pi1969 & n8201;
  assign n14898 = n8194 & n14897;
  assign n14899 = n8194 & n8206;
  assign n14900 = pi0359 & n14899;
  assign n14901 = n8243 & n14900;
  assign n14902 = ~n14898 & ~n14901;
  assign n14903 = n8197 & ~n14902;
  assign n14904 = ~n14896 & ~n14903;
  assign n14905 = pi0359 & n8229;
  assign n14906 = n11009 & n14905;
  assign n14907 = n14904 & ~n14906;
  assign n14908 = n14894 & n14907;
  assign n14909 = pi0483 & n14908;
  assign n14910 = ~n14884 & n14909;
  assign n14911 = ~pi0483 & ~pi0988;
  assign n14912 = pi3149 & pi3361;
  assign n14913 = ~pi1210 & ~pi1312;
  assign n14914 = n14912 & n14913;
  assign n14915 = pi3362 & n14914;
  assign n14916 = n14911 & n14915;
  assign po0683 = n14910 | n14916;
  assign n14918 = pi0484 & ~po1484;
  assign n14919 = ~pi0484 & po1484;
  assign n14920 = ~n8150 & ~n8157;
  assign n14921 = n14919 & ~n14920;
  assign po0684 = n14918 | n14921;
  assign n14923 = pi3389 & n14916;
  assign n14924 = pi0485 & n11017;
  assign n14925 = pi0486 & pi0507;
  assign n14926 = pi0506 & pi0512;
  assign n14927 = n14925 & n14926;
  assign n14928 = pi0503 & pi0514;
  assign n14929 = pi0504 & pi0505;
  assign n14930 = n14928 & n14929;
  assign n14931 = pi0515 & n14930;
  assign n14932 = n14927 & n14931;
  assign n14933 = pi0485 & ~n14932;
  assign n14934 = ~pi0485 & n14932;
  assign n14935 = ~n14933 & ~n14934;
  assign n14936 = ~n11017 & ~n14935;
  assign n14937 = ~n14924 & ~n14936;
  assign n14938 = ~n14916 & ~n14937;
  assign po0685 = n14923 | n14938;
  assign n14940 = pi3388 & n14916;
  assign n14941 = pi0486 & n11017;
  assign n14942 = pi0507 & pi0512;
  assign n14943 = pi0505 & pi0506;
  assign n14944 = n14942 & n14943;
  assign n14945 = pi0503 & pi0515;
  assign n14946 = pi0514 & n14945;
  assign n14947 = pi0504 & n14946;
  assign n14948 = n14944 & n14947;
  assign n14949 = pi0486 & ~n14948;
  assign n14950 = ~pi0486 & n14948;
  assign n14951 = ~n14949 & ~n14950;
  assign n14952 = ~n11017 & ~n14951;
  assign n14953 = ~n14941 & ~n14952;
  assign n14954 = ~n14916 & ~n14953;
  assign po0686 = n14940 | n14954;
  assign n14956 = pi3391 & n14916;
  assign n14957 = pi0487 & n11017;
  assign n14958 = pi0485 & pi0499;
  assign n14959 = n14925 & n14958;
  assign n14960 = n14926 & n14929;
  assign n14961 = n14946 & n14960;
  assign n14962 = n14959 & n14961;
  assign n14963 = pi0487 & ~n14962;
  assign n14964 = ~pi0487 & n14962;
  assign n14965 = ~n14963 & ~n14964;
  assign n14966 = ~n11017 & ~n14965;
  assign n14967 = ~n14957 & ~n14966;
  assign n14968 = ~n14916 & ~n14967;
  assign po0687 = n14956 | n14968;
  assign n14970 = pi3392 & n14916;
  assign n14971 = pi0488 & n11017;
  assign n14972 = pi0485 & pi0486;
  assign n14973 = pi0487 & pi0499;
  assign n14974 = n14972 & n14973;
  assign n14975 = n14948 & n14974;
  assign n14976 = pi0488 & ~n14975;
  assign n14977 = ~pi0488 & n14975;
  assign n14978 = ~n14976 & ~n14977;
  assign n14979 = ~n11017 & ~n14978;
  assign n14980 = ~n14971 & ~n14979;
  assign n14981 = ~n14916 & ~n14980;
  assign po0688 = n14970 | n14981;
  assign n14983 = pi3393 & n14916;
  assign n14984 = pi0489 & n11017;
  assign n14985 = pi0487 & pi0488;
  assign n14986 = n14958 & n14985;
  assign n14987 = n14932 & n14986;
  assign n14988 = pi0489 & ~n14987;
  assign n14989 = ~pi0489 & n14987;
  assign n14990 = ~n14988 & ~n14989;
  assign n14991 = ~n11017 & ~n14990;
  assign n14992 = ~n14984 & ~n14991;
  assign n14993 = ~n14916 & ~n14992;
  assign po0689 = n14983 | n14993;
  assign n14995 = pi3394 & n14916;
  assign n14996 = pi0490 & n11017;
  assign n14997 = n14942 & n14972;
  assign n14998 = pi0504 & pi0514;
  assign n14999 = n14943 & n14998;
  assign n15000 = n14945 & n14999;
  assign n15001 = n14997 & n15000;
  assign n15002 = pi0488 & pi0489;
  assign n15003 = n14973 & n15002;
  assign n15004 = n15001 & n15003;
  assign n15005 = pi0490 & ~n15004;
  assign n15006 = ~pi0490 & n15004;
  assign n15007 = ~n15005 & ~n15006;
  assign n15008 = ~n11017 & ~n15007;
  assign n15009 = ~n14996 & ~n15008;
  assign n15010 = ~n14916 & ~n15009;
  assign po0690 = n14995 | n15010;
  assign n15012 = pi3395 & n14916;
  assign n15013 = pi0491 & n11017;
  assign n15014 = pi0487 & pi0490;
  assign n15015 = n15002 & n15014;
  assign n15016 = n14962 & n15015;
  assign n15017 = pi0491 & ~n15016;
  assign n15018 = ~pi0491 & n15016;
  assign n15019 = ~n15017 & ~n15018;
  assign n15020 = ~n11017 & ~n15019;
  assign n15021 = ~n15013 & ~n15020;
  assign n15022 = ~n14916 & ~n15021;
  assign po0691 = n15012 | n15022;
  assign n15024 = pi3397 & n14916;
  assign n15025 = pi0492 & n11017;
  assign n15026 = pi0489 & pi0511;
  assign n15027 = pi0490 & pi0491;
  assign n15028 = n15026 & n15027;
  assign n15029 = n14930 & n15028;
  assign n15030 = n14927 & n14986;
  assign n15031 = n15029 & n15030;
  assign n15032 = pi0515 & n15031;
  assign n15033 = pi0492 & ~n15032;
  assign n15034 = ~pi0492 & n15032;
  assign n15035 = ~n15033 & ~n15034;
  assign n15036 = ~n11017 & ~n15035;
  assign n15037 = ~n15025 & ~n15036;
  assign n15038 = ~n14916 & ~n15037;
  assign po0692 = n15024 | n15038;
  assign n15040 = pi3398 & n14916;
  assign n15041 = pi0493 & n11017;
  assign n15042 = pi0492 & pi0511;
  assign n15043 = n15027 & n15042;
  assign n15044 = n14997 & n15003;
  assign n15045 = n14999 & n15044;
  assign n15046 = n14945 & n15045;
  assign n15047 = n15043 & n15046;
  assign n15048 = pi0493 & ~n15047;
  assign n15049 = ~pi0493 & n15047;
  assign n15050 = ~n15048 & ~n15049;
  assign n15051 = ~n11017 & ~n15050;
  assign n15052 = ~n15041 & ~n15051;
  assign n15053 = ~n14916 & ~n15052;
  assign po0693 = n15040 | n15053;
  assign n15055 = pi3399 & n14916;
  assign n15056 = pi0494 & n11017;
  assign n15057 = pi0491 & pi0511;
  assign n15058 = pi0492 & pi0493;
  assign n15059 = n15057 & n15058;
  assign n15060 = n14959 & n15015;
  assign n15061 = n15059 & n15060;
  assign n15062 = n14961 & n15061;
  assign n15063 = pi0494 & ~n15062;
  assign n15064 = ~pi0494 & n15062;
  assign n15065 = ~n15063 & ~n15064;
  assign n15066 = ~n11017 & ~n15065;
  assign n15067 = ~n15056 & ~n15066;
  assign n15068 = ~n14916 & ~n15067;
  assign po0694 = n15055 | n15068;
  assign n15070 = pi3401 & n14916;
  assign n15071 = pi0495 & n11017;
  assign n15072 = pi0494 & pi0510;
  assign n15073 = n15058 & n15072;
  assign n15074 = n15028 & n15073;
  assign n15075 = n15030 & n15074;
  assign n15076 = n14931 & n15075;
  assign n15077 = pi0495 & ~n15076;
  assign n15078 = ~pi0495 & n15076;
  assign n15079 = ~n15077 & ~n15078;
  assign n15080 = ~n11017 & ~n15079;
  assign n15081 = ~n15071 & ~n15080;
  assign n15082 = ~n14916 & ~n15081;
  assign po0695 = n15070 | n15082;
  assign n15084 = pi3402 & n14916;
  assign n15085 = pi0496 & n11017;
  assign n15086 = pi0493 & pi0494;
  assign n15087 = pi0495 & pi0510;
  assign n15088 = n15086 & n15087;
  assign n15089 = n15044 & n15088;
  assign n15090 = n15000 & n15089;
  assign n15091 = n15043 & n15090;
  assign n15092 = pi0496 & ~n15091;
  assign n15093 = ~pi0496 & n15091;
  assign n15094 = ~n15092 & ~n15093;
  assign n15095 = ~n11017 & ~n15094;
  assign n15096 = ~n15085 & ~n15095;
  assign n15097 = ~n14916 & ~n15096;
  assign po0696 = n15084 | n15097;
  assign n15099 = pi3403 & n14916;
  assign n15100 = pi0497 & n11017;
  assign n15101 = pi0495 & pi0496;
  assign n15102 = n15072 & n15101;
  assign n15103 = n15061 & n15102;
  assign n15104 = n14961 & n15103;
  assign n15105 = pi0497 & ~n15104;
  assign n15106 = ~pi0497 & n15104;
  assign n15107 = ~n15105 & ~n15106;
  assign n15108 = ~n11017 & ~n15107;
  assign n15109 = ~n15100 & ~n15108;
  assign n15110 = ~n14916 & ~n15109;
  assign po0697 = n15099 | n15110;
  assign n15112 = pi3405 & n14916;
  assign n15113 = pi0498 & n11017;
  assign n15114 = pi0497 & pi0513;
  assign n15115 = n15101 & n15114;
  assign n15116 = n14986 & n15028;
  assign n15117 = n14932 & n15116;
  assign n15118 = n15115 & n15117;
  assign n15119 = n15073 & n15118;
  assign n15120 = pi0498 & ~n15119;
  assign n15121 = ~pi0498 & n15119;
  assign n15122 = ~n15120 & ~n15121;
  assign n15123 = ~n11017 & ~n15122;
  assign n15124 = ~n15113 & ~n15123;
  assign n15125 = ~n14916 & ~n15124;
  assign po0698 = n15112 | n15125;
  assign n15127 = pi3390 & n14916;
  assign n15128 = pi0499 & n11017;
  assign n15129 = pi0499 & ~n15001;
  assign n15130 = ~pi0499 & n15001;
  assign n15131 = ~n15129 & ~n15130;
  assign n15132 = ~n11017 & ~n15131;
  assign n15133 = ~n15128 & ~n15132;
  assign n15134 = ~n14916 & ~n15133;
  assign po0699 = n15127 | n15134;
  assign n15136 = pi3407 & n14916;
  assign n15137 = ~pi0500 & n11017;
  assign n15138 = pi0498 & pi0508;
  assign n15139 = n15114 & n15138;
  assign n15140 = n14962 & n15059;
  assign n15141 = n15015 & n15140;
  assign n15142 = n15102 & n15141;
  assign n15143 = n15139 & n15142;
  assign n15144 = ~pi0500 & n15143;
  assign n15145 = pi0500 & ~n15143;
  assign n15146 = ~n15144 & ~n15145;
  assign n15147 = ~n11017 & n15146;
  assign n15148 = ~n15137 & ~n15147;
  assign n15149 = ~n14916 & ~n15148;
  assign po0700 = n15136 | n15149;
  assign n15151 = pi3408 & n14916;
  assign n15152 = pi0501 & n11017;
  assign n15153 = pi0496 & pi0497;
  assign n15154 = n15087 & n15153;
  assign n15155 = n15002 & n15027;
  assign n15156 = n15042 & n15086;
  assign n15157 = n15155 & n15156;
  assign n15158 = n14975 & n15157;
  assign n15159 = n15154 & n15158;
  assign n15160 = pi0498 & pi0513;
  assign n15161 = ~pi0500 & n15160;
  assign n15162 = pi0508 & n15161;
  assign n15163 = n15159 & n15162;
  assign n15164 = pi0501 & ~n15163;
  assign n15165 = ~pi0501 & n15163;
  assign n15166 = ~n15164 & ~n15165;
  assign n15167 = ~n11017 & ~n15166;
  assign n15168 = ~n15152 & ~n15167;
  assign n15169 = ~n14916 & ~n15168;
  assign po0701 = n15151 | n15169;
  assign n15171 = pi3409 & n14916;
  assign n15172 = ~pi0502 & n11017;
  assign n15173 = ~pi0500 & pi0501;
  assign n15174 = n15138 & n15173;
  assign n15175 = n14987 & n15174;
  assign n15176 = n15115 & n15175;
  assign n15177 = n15074 & n15176;
  assign n15178 = ~pi0502 & n15177;
  assign n15179 = pi0502 & ~n15177;
  assign n15180 = ~n15178 & ~n15179;
  assign n15181 = ~n11017 & n15180;
  assign n15182 = ~n15172 & ~n15181;
  assign n15183 = ~n14916 & ~n15182;
  assign po0702 = n15171 | n15183;
  assign n15185 = pi3381 & n14916;
  assign n15186 = pi0503 & n11017;
  assign n15187 = pi0503 & ~pi0515;
  assign n15188 = ~pi0503 & pi0515;
  assign n15189 = ~n15187 & ~n15188;
  assign n15190 = ~n11017 & ~n15189;
  assign n15191 = ~n15186 & ~n15190;
  assign n15192 = ~n14916 & ~n15191;
  assign po0703 = n15185 | n15192;
  assign n15194 = pi3383 & n14916;
  assign n15195 = pi0504 & n11017;
  assign n15196 = pi0504 & ~n14946;
  assign n15197 = ~pi0504 & n14946;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = ~n11017 & ~n15198;
  assign n15200 = ~n15195 & ~n15199;
  assign n15201 = ~n14916 & ~n15200;
  assign po0704 = n15194 | n15201;
  assign n15203 = pi3384 & n14916;
  assign n15204 = pi0505 & n11017;
  assign n15205 = pi0505 & ~n14947;
  assign n15206 = ~pi0505 & n14947;
  assign n15207 = ~n15205 & ~n15206;
  assign n15208 = ~n11017 & ~n15207;
  assign n15209 = ~n15204 & ~n15208;
  assign n15210 = ~n14916 & ~n15209;
  assign po0705 = n15203 | n15210;
  assign n15212 = pi3385 & n14916;
  assign n15213 = pi0506 & n11017;
  assign n15214 = pi0506 & ~n14931;
  assign n15215 = ~pi0506 & n14931;
  assign n15216 = ~n15214 & ~n15215;
  assign n15217 = ~n11017 & ~n15216;
  assign n15218 = ~n15213 & ~n15217;
  assign n15219 = ~n14916 & ~n15218;
  assign po0706 = n15212 | n15219;
  assign n15221 = pi3387 & n14916;
  assign n15222 = pi0507 & n11017;
  assign n15223 = pi0507 & ~n14961;
  assign n15224 = ~pi0507 & n14961;
  assign n15225 = ~n15223 & ~n15224;
  assign n15226 = ~n11017 & ~n15225;
  assign n15227 = ~n15222 & ~n15226;
  assign n15228 = ~n14916 & ~n15227;
  assign po0707 = n15221 | n15228;
  assign n15230 = pi3406 & n14916;
  assign n15231 = pi0508 & n11017;
  assign n15232 = n15001 & n15088;
  assign n15233 = n15003 & n15232;
  assign n15234 = n15043 & n15153;
  assign n15235 = n15160 & n15234;
  assign n15236 = n15233 & n15235;
  assign n15237 = pi0508 & ~n15236;
  assign n15238 = ~pi0508 & n15236;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = ~n11017 & ~n15239;
  assign n15241 = ~n15231 & ~n15240;
  assign n15242 = ~n14916 & ~n15241;
  assign po0708 = n15230 | n15242;
  assign n15244 = n11017 & n14891;
  assign n15245 = pi0509 & n15244;
  assign n15246 = n14907 & n15245;
  assign n15247 = ~pi0988 & pi3149;
  assign n15248 = pi3363 & n14881;
  assign n15249 = n14913 & n15248;
  assign n15250 = n15247 & n15249;
  assign n15251 = ~pi0509 & n15250;
  assign po0709 = n15246 | n15251;
  assign n15253 = pi3400 & n14916;
  assign n15254 = pi0510 & n11017;
  assign n15255 = n14944 & n14974;
  assign n15256 = n14947 & n15255;
  assign n15257 = n15157 & n15256;
  assign n15258 = pi0510 & ~n15257;
  assign n15259 = ~pi0510 & n15257;
  assign n15260 = ~n15258 & ~n15259;
  assign n15261 = ~n11017 & ~n15260;
  assign n15262 = ~n15254 & ~n15261;
  assign n15263 = ~n14916 & ~n15262;
  assign po0710 = n15253 | n15263;
  assign n15265 = pi3396 & n14916;
  assign n15266 = pi0511 & n11017;
  assign n15267 = n14975 & n15155;
  assign n15268 = pi0511 & ~n15267;
  assign n15269 = ~pi0511 & n15267;
  assign n15270 = ~n15268 & ~n15269;
  assign n15271 = ~n11017 & ~n15270;
  assign n15272 = ~n15266 & ~n15271;
  assign n15273 = ~n14916 & ~n15272;
  assign po0711 = n15265 | n15273;
  assign n15275 = pi3386 & n14916;
  assign n15276 = pi0512 & n11017;
  assign n15277 = pi0512 & ~n15000;
  assign n15278 = ~pi0512 & n15000;
  assign n15279 = ~n15277 & ~n15278;
  assign n15280 = ~n11017 & ~n15279;
  assign n15281 = ~n15276 & ~n15280;
  assign n15282 = ~n14916 & ~n15281;
  assign po0712 = n15275 | n15282;
  assign n15284 = pi3404 & n14916;
  assign n15285 = pi0513 & n11017;
  assign n15286 = n15154 & n15267;
  assign n15287 = n15156 & n15286;
  assign n15288 = pi0513 & ~n15287;
  assign n15289 = ~pi0513 & n15287;
  assign n15290 = ~n15288 & ~n15289;
  assign n15291 = ~n11017 & ~n15290;
  assign n15292 = ~n15285 & ~n15291;
  assign n15293 = ~n14916 & ~n15292;
  assign po0713 = n15284 | n15293;
  assign n15295 = pi3382 & n14916;
  assign n15296 = pi0514 & n11017;
  assign n15297 = pi0514 & ~n14945;
  assign n15298 = ~pi0514 & n14945;
  assign n15299 = ~n15297 & ~n15298;
  assign n15300 = ~n11017 & ~n15299;
  assign n15301 = ~n15296 & ~n15300;
  assign n15302 = ~n14916 & ~n15301;
  assign po0714 = n15295 | n15302;
  assign n15304 = pi3380 & n14916;
  assign n15305 = pi0515 & n11017;
  assign n15306 = ~pi0515 & ~n11017;
  assign n15307 = ~n15305 & ~n15306;
  assign n15308 = ~n14916 & ~n15307;
  assign po0715 = n15304 | n15308;
  assign n15310 = pi1152 & pi1176;
  assign n15311 = pi1154 & pi1167;
  assign n15312 = n15310 & n15311;
  assign n15313 = ~pi0516 & ~n15312;
  assign n15314 = pi0485 & ~pi1345;
  assign n15315 = ~pi1274 & pi1345;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = n15312 & ~n15316;
  assign n15318 = ~n15313 & ~n15317;
  assign n15319 = n8194 & ~n8201;
  assign n15320 = n8206 & n15319;
  assign n15321 = n8188 & n15320;
  assign n15322 = n8198 & n15321;
  assign n15323 = ~n8295 & n8296;
  assign n15324 = ~n15322 & ~n15323;
  assign n15325 = ~n10998 & n15324;
  assign n15326 = ~n8276 & ~n15325;
  assign n15327 = ~n15318 & n15326;
  assign n15328 = ~pi0516 & ~n15326;
  assign po0716 = n15327 | n15328;
  assign n15330 = pi0492 & ~pi1345;
  assign n15331 = ~pi1329 & pi1345;
  assign n15332 = ~n15330 & ~n15331;
  assign n15333 = ~pi1152 & pi1176;
  assign n15334 = pi1154 & ~pi1167;
  assign n15335 = n15333 & n15334;
  assign n15336 = ~n15332 & n15335;
  assign n15337 = ~pi0517 & ~n15335;
  assign n15338 = ~n15336 & ~n15337;
  assign n15339 = n15326 & ~n15338;
  assign n15340 = ~pi0517 & ~n15326;
  assign po0717 = n15339 | n15340;
  assign n15342 = ~pi0518 & ~n15312;
  assign n15343 = n15312 & ~n15332;
  assign n15344 = ~n15342 & ~n15343;
  assign n15345 = n15326 & ~n15344;
  assign n15346 = ~pi0518 & ~n15326;
  assign po0718 = n15345 | n15346;
  assign n15348 = ~n8990 & ~n12560;
  assign n15349 = ~pi2972 & ~n9242;
  assign n15350 = ~pi3117 & po3257;
  assign n15351 = ~pi2969 & n15350;
  assign n15352 = ~n15349 & ~n15351;
  assign n15353 = pi1232 & pi3027;
  assign n15354 = ~pi3201 & ~n15353;
  assign n15355 = n9391 & n15354;
  assign n15356 = ~n9380 & ~n15355;
  assign n15357 = pi0307 & ~n15356;
  assign n15358 = ~n9385 & ~n15357;
  assign n15359 = pi1697 & n9389;
  assign n15360 = ~pi1696 & n15359;
  assign n15361 = ~pi3369 & n15360;
  assign n15362 = n15358 & ~n15361;
  assign n15363 = n15352 & n15362;
  assign n15364 = n15348 & n15363;
  assign n15365 = ~pi1220 & pi3375;
  assign n15366 = ~pi0126 & pi1220;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~n9396 & ~n15367;
  assign n15369 = ~n8078 & ~n15368;
  assign po0719 = n15364 | n15369;
  assign n15371 = ~pi0543 & ~n15326;
  assign n15372 = ~pi1154 & ~pi1167;
  assign n15373 = ~pi1152 & ~pi1176;
  assign n15374 = n15372 & n15373;
  assign n15375 = pi1321 & pi1345;
  assign n15376 = ~pi1345 & pi1762;
  assign n15377 = n15375 & ~n15376;
  assign n15378 = n15374 & n15377;
  assign n15379 = ~pi0543 & ~n15374;
  assign n15380 = ~n15378 & ~n15379;
  assign n15381 = n15326 & ~n15380;
  assign po0731 = n15371 | n15381;
  assign n15383 = ~pi0544 & ~n15326;
  assign n15384 = pi1152 & ~pi1176;
  assign n15385 = ~pi1154 & pi1167;
  assign n15386 = n15384 & n15385;
  assign n15387 = n15377 & n15386;
  assign n15388 = ~pi0544 & ~n15386;
  assign n15389 = ~n15387 & ~n15388;
  assign n15390 = n15326 & ~n15389;
  assign po0732 = n15383 | n15390;
  assign n15392 = ~pi0545 & ~n15326;
  assign n15393 = n15333 & n15385;
  assign n15394 = n15377 & n15393;
  assign n15395 = ~pi0545 & ~n15393;
  assign n15396 = ~n15394 & ~n15395;
  assign n15397 = n15326 & ~n15396;
  assign po0733 = n15392 | n15397;
  assign n15399 = ~pi0546 & ~n15326;
  assign n15400 = n15334 & n15373;
  assign n15401 = n15377 & n15400;
  assign n15402 = ~pi0546 & ~n15400;
  assign n15403 = ~n15401 & ~n15402;
  assign n15404 = n15326 & ~n15403;
  assign po0734 = n15399 | n15404;
  assign n15406 = ~pi0547 & ~n15326;
  assign n15407 = n15372 & n15384;
  assign n15408 = n15377 & n15407;
  assign n15409 = ~pi0547 & ~n15407;
  assign n15410 = ~n15408 & ~n15409;
  assign n15411 = n15326 & ~n15410;
  assign po0735 = n15406 | n15411;
  assign n15413 = ~pi0548 & ~n15326;
  assign n15414 = n15334 & n15384;
  assign n15415 = n15377 & n15414;
  assign n15416 = ~pi0548 & ~n15414;
  assign n15417 = ~n15415 & ~n15416;
  assign n15418 = n15326 & ~n15417;
  assign po0736 = n15413 | n15418;
  assign n15420 = ~pi0549 & ~n15326;
  assign n15421 = n15335 & n15377;
  assign n15422 = ~pi0549 & ~n15335;
  assign n15423 = ~n15421 & ~n15422;
  assign n15424 = n15326 & ~n15423;
  assign po0737 = n15420 | n15424;
  assign n15426 = ~pi0550 & ~n15326;
  assign n15427 = n15310 & n15372;
  assign n15428 = n15377 & n15427;
  assign n15429 = ~pi0550 & ~n15427;
  assign n15430 = ~n15428 & ~n15429;
  assign n15431 = n15326 & ~n15430;
  assign po0738 = n15426 | n15431;
  assign n15433 = ~pi0551 & ~n15326;
  assign n15434 = n15373 & n15385;
  assign n15435 = n15377 & n15434;
  assign n15436 = ~pi0551 & ~n15434;
  assign n15437 = ~n15435 & ~n15436;
  assign n15438 = n15326 & ~n15437;
  assign po0739 = n15433 | n15438;
  assign n15440 = ~pi1345 & pi2938;
  assign n15441 = ~pi1272 & pi1345;
  assign n15442 = ~n15440 & ~n15441;
  assign n15443 = n15386 & ~n15442;
  assign n15444 = ~pi0552 & ~n15386;
  assign n15445 = ~n15443 & ~n15444;
  assign n15446 = n15326 & ~n15445;
  assign n15447 = ~pi0552 & ~n15326;
  assign po0740 = n15446 | n15447;
  assign n15449 = pi0486 & ~pi1345;
  assign n15450 = ~pi1273 & pi1345;
  assign n15451 = ~n15449 & ~n15450;
  assign n15452 = n15386 & ~n15451;
  assign n15453 = ~pi0553 & ~n15386;
  assign n15454 = ~n15452 & ~n15453;
  assign n15455 = n15326 & ~n15454;
  assign n15456 = ~pi0553 & ~n15326;
  assign po0741 = n15455 | n15456;
  assign n15458 = ~n15316 & n15386;
  assign n15459 = ~pi0554 & ~n15386;
  assign n15460 = ~n15458 & ~n15459;
  assign n15461 = n15326 & ~n15460;
  assign n15462 = ~pi0554 & ~n15326;
  assign po0742 = n15461 | n15462;
  assign n15464 = pi0487 & ~pi1345;
  assign n15465 = ~pi1275 & pi1345;
  assign n15466 = ~n15464 & ~n15465;
  assign n15467 = n15386 & ~n15466;
  assign n15468 = ~pi0555 & ~n15386;
  assign n15469 = ~n15467 & ~n15468;
  assign n15470 = n15326 & ~n15469;
  assign n15471 = ~pi0555 & ~n15326;
  assign po0743 = n15470 | n15471;
  assign n15473 = pi0489 & ~pi1345;
  assign n15474 = ~pi1277 & pi1345;
  assign n15475 = ~n15473 & ~n15474;
  assign n15476 = n15386 & ~n15475;
  assign n15477 = ~pi0556 & ~n15386;
  assign n15478 = ~n15476 & ~n15477;
  assign n15479 = n15326 & ~n15478;
  assign n15480 = ~pi0556 & ~n15326;
  assign po0744 = n15479 | n15480;
  assign n15482 = pi0490 & ~pi1345;
  assign n15483 = ~pi1326 & pi1345;
  assign n15484 = ~n15482 & ~n15483;
  assign n15485 = n15386 & ~n15484;
  assign n15486 = ~pi0557 & ~n15386;
  assign n15487 = ~n15485 & ~n15486;
  assign n15488 = n15326 & ~n15487;
  assign n15489 = ~pi0557 & ~n15326;
  assign po0745 = n15488 | n15489;
  assign n15491 = pi0491 & ~pi1345;
  assign n15492 = ~pi1278 & pi1345;
  assign n15493 = ~n15491 & ~n15492;
  assign n15494 = n15386 & ~n15493;
  assign n15495 = ~pi0558 & ~n15386;
  assign n15496 = ~n15494 & ~n15495;
  assign n15497 = n15326 & ~n15496;
  assign n15498 = ~pi0558 & ~n15326;
  assign po0746 = n15497 | n15498;
  assign n15500 = pi0511 & ~pi1345;
  assign n15501 = ~pi1279 & pi1345;
  assign n15502 = ~n15500 & ~n15501;
  assign n15503 = n15386 & ~n15502;
  assign n15504 = ~pi0559 & ~n15386;
  assign n15505 = ~n15503 & ~n15504;
  assign n15506 = n15326 & ~n15505;
  assign n15507 = ~pi0559 & ~n15326;
  assign po0747 = n15506 | n15507;
  assign n15509 = ~n15332 & n15386;
  assign n15510 = ~pi0560 & ~n15386;
  assign n15511 = ~n15509 & ~n15510;
  assign n15512 = n15326 & ~n15511;
  assign n15513 = ~pi0560 & ~n15326;
  assign po0748 = n15512 | n15513;
  assign n15515 = pi0493 & ~pi1345;
  assign n15516 = ~pi1327 & pi1345;
  assign n15517 = ~n15515 & ~n15516;
  assign n15518 = n15386 & ~n15517;
  assign n15519 = ~pi0561 & ~n15386;
  assign n15520 = ~n15518 & ~n15519;
  assign n15521 = n15326 & ~n15520;
  assign n15522 = ~pi0561 & ~n15326;
  assign po0749 = n15521 | n15522;
  assign n15524 = pi0494 & ~pi1345;
  assign n15525 = ~pi1281 & pi1345;
  assign n15526 = ~n15524 & ~n15525;
  assign n15527 = n15386 & ~n15526;
  assign n15528 = ~pi0562 & ~n15386;
  assign n15529 = ~n15527 & ~n15528;
  assign n15530 = n15326 & ~n15529;
  assign n15531 = ~pi0562 & ~n15326;
  assign po0750 = n15530 | n15531;
  assign n15533 = pi0495 & ~pi1345;
  assign n15534 = ~pi1282 & pi1345;
  assign n15535 = ~n15533 & ~n15534;
  assign n15536 = n15386 & ~n15535;
  assign n15537 = ~pi0563 & ~n15386;
  assign n15538 = ~n15536 & ~n15537;
  assign n15539 = n15326 & ~n15538;
  assign n15540 = ~pi0563 & ~n15326;
  assign po0751 = n15539 | n15540;
  assign n15542 = pi0496 & ~pi1345;
  assign n15543 = ~pi1325 & pi1345;
  assign n15544 = ~n15542 & ~n15543;
  assign n15545 = n15386 & ~n15544;
  assign n15546 = ~pi0564 & ~n15386;
  assign n15547 = ~n15545 & ~n15546;
  assign n15548 = n15326 & ~n15547;
  assign n15549 = ~pi0564 & ~n15326;
  assign po0752 = n15548 | n15549;
  assign n15551 = pi0513 & ~pi1345;
  assign n15552 = ~pi1284 & pi1345;
  assign n15553 = ~n15551 & ~n15552;
  assign n15554 = n15386 & ~n15553;
  assign n15555 = ~pi0565 & ~n15386;
  assign n15556 = ~n15554 & ~n15555;
  assign n15557 = n15326 & ~n15556;
  assign n15558 = ~pi0565 & ~n15326;
  assign po0753 = n15557 | n15558;
  assign n15560 = pi0508 & ~pi1345;
  assign n15561 = ~pi1324 & pi1345;
  assign n15562 = ~n15560 & ~n15561;
  assign n15563 = n15386 & ~n15562;
  assign n15564 = ~pi0566 & ~n15386;
  assign n15565 = ~n15563 & ~n15564;
  assign n15566 = n15326 & ~n15565;
  assign n15567 = ~pi0566 & ~n15326;
  assign po0754 = n15566 | n15567;
  assign n15569 = ~pi0500 & ~pi1345;
  assign n15570 = ~pi1286 & pi1345;
  assign n15571 = ~n15569 & ~n15570;
  assign n15572 = n15386 & ~n15571;
  assign n15573 = ~pi0567 & ~n15386;
  assign n15574 = ~n15572 & ~n15573;
  assign n15575 = n15326 & ~n15574;
  assign n15576 = ~pi0567 & ~n15326;
  assign po0755 = n15575 | n15576;
  assign n15578 = pi0501 & ~pi1345;
  assign n15579 = ~pi1288 & pi1345;
  assign n15580 = ~n15578 & ~n15579;
  assign n15581 = n15386 & ~n15580;
  assign n15582 = ~pi0568 & ~n15386;
  assign n15583 = ~n15581 & ~n15582;
  assign n15584 = n15326 & ~n15583;
  assign n15585 = ~pi0568 & ~n15326;
  assign po0756 = n15584 | n15585;
  assign n15587 = ~pi0502 & ~pi1345;
  assign n15588 = ~pi1322 & pi1345;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = n15386 & ~n15589;
  assign n15591 = ~pi0569 & ~n15386;
  assign n15592 = ~n15590 & ~n15591;
  assign n15593 = n15326 & ~n15592;
  assign n15594 = ~pi0569 & ~n15326;
  assign po0757 = n15593 | n15594;
  assign n15596 = pi0503 & ~pi1345;
  assign n15597 = ~pi1292 & pi1345;
  assign n15598 = ~n15596 & ~n15597;
  assign n15599 = n15386 & ~n15598;
  assign n15600 = ~pi0570 & ~n15386;
  assign n15601 = ~n15599 & ~n15600;
  assign n15602 = n15326 & ~n15601;
  assign n15603 = ~pi0570 & ~n15326;
  assign po0758 = n15602 | n15603;
  assign n15605 = pi0506 & ~pi1345;
  assign n15606 = ~pi1295 & pi1345;
  assign n15607 = ~n15605 & ~n15606;
  assign n15608 = n15386 & ~n15607;
  assign n15609 = ~pi0571 & ~n15386;
  assign n15610 = ~n15608 & ~n15609;
  assign n15611 = n15326 & ~n15610;
  assign n15612 = ~pi0571 & ~n15326;
  assign po0759 = n15611 | n15612;
  assign n15614 = pi0512 & ~pi1345;
  assign n15615 = ~pi1294 & pi1345;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = n15386 & ~n15616;
  assign n15618 = ~pi0572 & ~n15386;
  assign n15619 = ~n15617 & ~n15618;
  assign n15620 = n15326 & ~n15619;
  assign n15621 = ~pi0572 & ~n15326;
  assign po0760 = n15620 | n15621;
  assign n15623 = pi0507 & ~pi1345;
  assign n15624 = ~pi1319 & pi1345;
  assign n15625 = ~n15623 & ~n15624;
  assign n15626 = n15386 & ~n15625;
  assign n15627 = ~pi0573 & ~n15386;
  assign n15628 = ~n15626 & ~n15627;
  assign n15629 = n15326 & ~n15628;
  assign n15630 = ~pi0573 & ~n15326;
  assign po0761 = n15629 | n15630;
  assign n15632 = n15393 & ~n15451;
  assign n15633 = ~pi0574 & ~n15393;
  assign n15634 = ~n15632 & ~n15633;
  assign n15635 = n15326 & ~n15634;
  assign n15636 = ~pi0574 & ~n15326;
  assign po0762 = n15635 | n15636;
  assign n15638 = ~n15316 & n15393;
  assign n15639 = ~pi0575 & ~n15393;
  assign n15640 = ~n15638 & ~n15639;
  assign n15641 = n15326 & ~n15640;
  assign n15642 = ~pi0575 & ~n15326;
  assign po0763 = n15641 | n15642;
  assign n15644 = n15393 & ~n15466;
  assign n15645 = ~pi0576 & ~n15393;
  assign n15646 = ~n15644 & ~n15645;
  assign n15647 = n15326 & ~n15646;
  assign n15648 = ~pi0576 & ~n15326;
  assign po0764 = n15647 | n15648;
  assign n15650 = n15393 & ~n15475;
  assign n15651 = ~pi0577 & ~n15393;
  assign n15652 = ~n15650 & ~n15651;
  assign n15653 = n15326 & ~n15652;
  assign n15654 = ~pi0577 & ~n15326;
  assign po0765 = n15653 | n15654;
  assign n15656 = n15393 & ~n15484;
  assign n15657 = ~pi0578 & ~n15393;
  assign n15658 = ~n15656 & ~n15657;
  assign n15659 = n15326 & ~n15658;
  assign n15660 = ~pi0578 & ~n15326;
  assign po0766 = n15659 | n15660;
  assign n15662 = n15393 & ~n15502;
  assign n15663 = ~pi0579 & ~n15393;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = n15326 & ~n15664;
  assign n15666 = ~pi0579 & ~n15326;
  assign po0767 = n15665 | n15666;
  assign n15668 = ~n15332 & n15393;
  assign n15669 = ~pi0580 & ~n15393;
  assign n15670 = ~n15668 & ~n15669;
  assign n15671 = n15326 & ~n15670;
  assign n15672 = ~pi0580 & ~n15326;
  assign po0768 = n15671 | n15672;
  assign n15674 = n15393 & ~n15517;
  assign n15675 = ~pi0581 & ~n15393;
  assign n15676 = ~n15674 & ~n15675;
  assign n15677 = n15326 & ~n15676;
  assign n15678 = ~pi0581 & ~n15326;
  assign po0769 = n15677 | n15678;
  assign n15680 = n15393 & ~n15535;
  assign n15681 = ~pi0582 & ~n15393;
  assign n15682 = ~n15680 & ~n15681;
  assign n15683 = n15326 & ~n15682;
  assign n15684 = ~pi0582 & ~n15326;
  assign po0770 = n15683 | n15684;
  assign n15686 = n15393 & ~n15544;
  assign n15687 = ~pi0583 & ~n15393;
  assign n15688 = ~n15686 & ~n15687;
  assign n15689 = n15326 & ~n15688;
  assign n15690 = ~pi0583 & ~n15326;
  assign po0771 = n15689 | n15690;
  assign n15692 = n15393 & ~n15553;
  assign n15693 = ~pi0584 & ~n15393;
  assign n15694 = ~n15692 & ~n15693;
  assign n15695 = n15326 & ~n15694;
  assign n15696 = ~pi0584 & ~n15326;
  assign po0772 = n15695 | n15696;
  assign n15698 = pi0498 & ~pi1345;
  assign n15699 = ~pi1285 & pi1345;
  assign n15700 = ~n15698 & ~n15699;
  assign n15701 = n15393 & ~n15700;
  assign n15702 = ~pi0585 & ~n15393;
  assign n15703 = ~n15701 & ~n15702;
  assign n15704 = n15326 & ~n15703;
  assign n15705 = ~pi0585 & ~n15326;
  assign po0773 = n15704 | n15705;
  assign n15707 = ~pi1345 & pi2941;
  assign n15708 = ~pi1280 & pi1345;
  assign n15709 = ~n15707 & ~n15708;
  assign n15710 = n15393 & ~n15709;
  assign n15711 = ~pi0586 & ~n15393;
  assign n15712 = ~n15710 & ~n15711;
  assign n15713 = n15326 & ~n15712;
  assign n15714 = ~pi0586 & ~n15326;
  assign po0774 = n15713 | n15714;
  assign n15716 = n15393 & ~n15580;
  assign n15717 = ~pi0587 & ~n15393;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = n15326 & ~n15718;
  assign n15720 = ~pi0587 & ~n15326;
  assign po0775 = n15719 | n15720;
  assign n15722 = n15393 & ~n15589;
  assign n15723 = ~pi0588 & ~n15393;
  assign n15724 = ~n15722 & ~n15723;
  assign n15725 = n15326 & ~n15724;
  assign n15726 = ~pi0588 & ~n15326;
  assign po0776 = n15725 | n15726;
  assign n15728 = n15393 & ~n15598;
  assign n15729 = ~pi0589 & ~n15393;
  assign n15730 = ~n15728 & ~n15729;
  assign n15731 = n15326 & ~n15730;
  assign n15732 = ~pi0589 & ~n15326;
  assign po0777 = n15731 | n15732;
  assign n15734 = n15393 & ~n15607;
  assign n15735 = ~pi0590 & ~n15393;
  assign n15736 = ~n15734 & ~n15735;
  assign n15737 = n15326 & ~n15736;
  assign n15738 = ~pi0590 & ~n15326;
  assign po0778 = n15737 | n15738;
  assign n15740 = n15393 & ~n15616;
  assign n15741 = ~pi0591 & ~n15393;
  assign n15742 = ~n15740 & ~n15741;
  assign n15743 = n15326 & ~n15742;
  assign n15744 = ~pi0591 & ~n15326;
  assign po0779 = n15743 | n15744;
  assign n15746 = n15393 & ~n15625;
  assign n15747 = ~pi0592 & ~n15393;
  assign n15748 = ~n15746 & ~n15747;
  assign n15749 = n15326 & ~n15748;
  assign n15750 = ~pi0592 & ~n15326;
  assign po0780 = n15749 | n15750;
  assign n15752 = n15414 & ~n15442;
  assign n15753 = ~pi0593 & ~n15414;
  assign n15754 = ~n15752 & ~n15753;
  assign n15755 = n15326 & ~n15754;
  assign n15756 = ~pi0593 & ~n15326;
  assign po0781 = n15755 | n15756;
  assign n15758 = ~n15316 & n15414;
  assign n15759 = ~pi0594 & ~n15414;
  assign n15760 = ~n15758 & ~n15759;
  assign n15761 = n15326 & ~n15760;
  assign n15762 = ~pi0594 & ~n15326;
  assign po0782 = n15761 | n15762;
  assign n15764 = n15414 & ~n15466;
  assign n15765 = ~pi0595 & ~n15414;
  assign n15766 = ~n15764 & ~n15765;
  assign n15767 = n15326 & ~n15766;
  assign n15768 = ~pi0595 & ~n15326;
  assign po0783 = n15767 | n15768;
  assign n15770 = n15414 & ~n15475;
  assign n15771 = ~pi0596 & ~n15414;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = n15326 & ~n15772;
  assign n15774 = ~pi0596 & ~n15326;
  assign po0784 = n15773 | n15774;
  assign n15776 = n15414 & ~n15484;
  assign n15777 = ~pi0597 & ~n15414;
  assign n15778 = ~n15776 & ~n15777;
  assign n15779 = n15326 & ~n15778;
  assign n15780 = ~pi0597 & ~n15326;
  assign po0785 = n15779 | n15780;
  assign n15782 = n15414 & ~n15493;
  assign n15783 = ~pi0598 & ~n15414;
  assign n15784 = ~n15782 & ~n15783;
  assign n15785 = n15326 & ~n15784;
  assign n15786 = ~pi0598 & ~n15326;
  assign po0786 = n15785 | n15786;
  assign n15788 = n15414 & ~n15502;
  assign n15789 = ~pi0599 & ~n15414;
  assign n15790 = ~n15788 & ~n15789;
  assign n15791 = n15326 & ~n15790;
  assign n15792 = ~pi0599 & ~n15326;
  assign po0787 = n15791 | n15792;
  assign n15794 = ~n15332 & n15414;
  assign n15795 = ~pi0600 & ~n15414;
  assign n15796 = ~n15794 & ~n15795;
  assign n15797 = n15326 & ~n15796;
  assign n15798 = ~pi0600 & ~n15326;
  assign po0788 = n15797 | n15798;
  assign n15800 = n15414 & ~n15709;
  assign n15801 = ~pi0601 & ~n15414;
  assign n15802 = ~n15800 & ~n15801;
  assign n15803 = n15326 & ~n15802;
  assign n15804 = ~pi0601 & ~n15326;
  assign po0789 = n15803 | n15804;
  assign n15806 = n15414 & ~n15517;
  assign n15807 = ~pi0602 & ~n15414;
  assign n15808 = ~n15806 & ~n15807;
  assign n15809 = n15326 & ~n15808;
  assign n15810 = ~pi0602 & ~n15326;
  assign po0790 = n15809 | n15810;
  assign n15812 = n15414 & ~n15535;
  assign n15813 = ~pi0603 & ~n15414;
  assign n15814 = ~n15812 & ~n15813;
  assign n15815 = n15326 & ~n15814;
  assign n15816 = ~pi0603 & ~n15326;
  assign po0791 = n15815 | n15816;
  assign n15818 = n15414 & ~n15544;
  assign n15819 = ~pi0604 & ~n15414;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = n15326 & ~n15820;
  assign n15822 = ~pi0604 & ~n15326;
  assign po0792 = n15821 | n15822;
  assign n15824 = n15414 & ~n15553;
  assign n15825 = ~pi0605 & ~n15414;
  assign n15826 = ~n15824 & ~n15825;
  assign n15827 = n15326 & ~n15826;
  assign n15828 = ~pi0605 & ~n15326;
  assign po0793 = n15827 | n15828;
  assign n15830 = n15414 & ~n15700;
  assign n15831 = ~pi0606 & ~n15414;
  assign n15832 = ~n15830 & ~n15831;
  assign n15833 = n15326 & ~n15832;
  assign n15834 = ~pi0606 & ~n15326;
  assign po0794 = n15833 | n15834;
  assign n15836 = n15414 & ~n15562;
  assign n15837 = ~pi0607 & ~n15414;
  assign n15838 = ~n15836 & ~n15837;
  assign n15839 = n15326 & ~n15838;
  assign n15840 = ~pi0607 & ~n15326;
  assign po0795 = n15839 | n15840;
  assign n15842 = n15414 & ~n15580;
  assign n15843 = ~pi0608 & ~n15414;
  assign n15844 = ~n15842 & ~n15843;
  assign n15845 = n15326 & ~n15844;
  assign n15846 = ~pi0608 & ~n15326;
  assign po0796 = n15845 | n15846;
  assign n15848 = n15414 & ~n15589;
  assign n15849 = ~pi0609 & ~n15414;
  assign n15850 = ~n15848 & ~n15849;
  assign n15851 = n15326 & ~n15850;
  assign n15852 = ~pi0609 & ~n15326;
  assign po0797 = n15851 | n15852;
  assign n15854 = n15414 & ~n15598;
  assign n15855 = ~pi0610 & ~n15414;
  assign n15856 = ~n15854 & ~n15855;
  assign n15857 = n15326 & ~n15856;
  assign n15858 = ~pi0610 & ~n15326;
  assign po0798 = n15857 | n15858;
  assign n15860 = n15414 & ~n15607;
  assign n15861 = ~pi0611 & ~n15414;
  assign n15862 = ~n15860 & ~n15861;
  assign n15863 = n15326 & ~n15862;
  assign n15864 = ~pi0611 & ~n15326;
  assign po0799 = n15863 | n15864;
  assign n15866 = n15414 & ~n15616;
  assign n15867 = ~pi0612 & ~n15414;
  assign n15868 = ~n15866 & ~n15867;
  assign n15869 = n15326 & ~n15868;
  assign n15870 = ~pi0612 & ~n15326;
  assign po0800 = n15869 | n15870;
  assign n15872 = n15414 & ~n15625;
  assign n15873 = ~pi0613 & ~n15414;
  assign n15874 = ~n15872 & ~n15873;
  assign n15875 = n15326 & ~n15874;
  assign n15876 = ~pi0613 & ~n15326;
  assign po0801 = n15875 | n15876;
  assign n15878 = n15335 & ~n15442;
  assign n15879 = ~pi0614 & ~n15335;
  assign n15880 = ~n15878 & ~n15879;
  assign n15881 = n15326 & ~n15880;
  assign n15882 = ~pi0614 & ~n15326;
  assign po0802 = n15881 | n15882;
  assign n15884 = n15335 & ~n15451;
  assign n15885 = ~pi0615 & ~n15335;
  assign n15886 = ~n15884 & ~n15885;
  assign n15887 = n15326 & ~n15886;
  assign n15888 = ~pi0615 & ~n15326;
  assign po0803 = n15887 | n15888;
  assign n15890 = n15335 & ~n15466;
  assign n15891 = ~pi0616 & ~n15335;
  assign n15892 = ~n15890 & ~n15891;
  assign n15893 = n15326 & ~n15892;
  assign n15894 = ~pi0616 & ~n15326;
  assign po0804 = n15893 | n15894;
  assign n15896 = n15335 & ~n15475;
  assign n15897 = ~pi0617 & ~n15335;
  assign n15898 = ~n15896 & ~n15897;
  assign n15899 = n15326 & ~n15898;
  assign n15900 = ~pi0617 & ~n15326;
  assign po0805 = n15899 | n15900;
  assign n15902 = n15335 & ~n15484;
  assign n15903 = ~pi0618 & ~n15335;
  assign n15904 = ~n15902 & ~n15903;
  assign n15905 = n15326 & ~n15904;
  assign n15906 = ~pi0618 & ~n15326;
  assign po0806 = n15905 | n15906;
  assign n15908 = n15335 & ~n15493;
  assign n15909 = ~pi0619 & ~n15335;
  assign n15910 = ~n15908 & ~n15909;
  assign n15911 = n15326 & ~n15910;
  assign n15912 = ~pi0619 & ~n15326;
  assign po0807 = n15911 | n15912;
  assign n15914 = n15335 & ~n15502;
  assign n15915 = ~pi0620 & ~n15335;
  assign n15916 = ~n15914 & ~n15915;
  assign n15917 = n15326 & ~n15916;
  assign n15918 = ~pi0620 & ~n15326;
  assign po0808 = n15917 | n15918;
  assign n15920 = n15335 & ~n15709;
  assign n15921 = ~pi0621 & ~n15335;
  assign n15922 = ~n15920 & ~n15921;
  assign n15923 = n15326 & ~n15922;
  assign n15924 = ~pi0621 & ~n15326;
  assign po0809 = n15923 | n15924;
  assign n15926 = n15335 & ~n15517;
  assign n15927 = ~pi0622 & ~n15335;
  assign n15928 = ~n15926 & ~n15927;
  assign n15929 = n15326 & ~n15928;
  assign n15930 = ~pi0622 & ~n15326;
  assign po0810 = n15929 | n15930;
  assign n15932 = n15335 & ~n15526;
  assign n15933 = ~pi0623 & ~n15335;
  assign n15934 = ~n15932 & ~n15933;
  assign n15935 = n15326 & ~n15934;
  assign n15936 = ~pi0623 & ~n15326;
  assign po0811 = n15935 | n15936;
  assign n15938 = n15335 & ~n15535;
  assign n15939 = ~pi0624 & ~n15335;
  assign n15940 = ~n15938 & ~n15939;
  assign n15941 = n15326 & ~n15940;
  assign n15942 = ~pi0624 & ~n15326;
  assign po0812 = n15941 | n15942;
  assign n15944 = n15335 & ~n15544;
  assign n15945 = ~pi0625 & ~n15335;
  assign n15946 = ~n15944 & ~n15945;
  assign n15947 = n15326 & ~n15946;
  assign n15948 = ~pi0625 & ~n15326;
  assign po0813 = n15947 | n15948;
  assign n15950 = n15335 & ~n15553;
  assign n15951 = ~pi0626 & ~n15335;
  assign n15952 = ~n15950 & ~n15951;
  assign n15953 = n15326 & ~n15952;
  assign n15954 = ~pi0626 & ~n15326;
  assign po0814 = n15953 | n15954;
  assign n15956 = n15335 & ~n15700;
  assign n15957 = ~pi0627 & ~n15335;
  assign n15958 = ~n15956 & ~n15957;
  assign n15959 = n15326 & ~n15958;
  assign n15960 = ~pi0627 & ~n15326;
  assign po0815 = n15959 | n15960;
  assign n15962 = n15335 & ~n15562;
  assign n15963 = ~pi0628 & ~n15335;
  assign n15964 = ~n15962 & ~n15963;
  assign n15965 = n15326 & ~n15964;
  assign n15966 = ~pi0628 & ~n15326;
  assign po0816 = n15965 | n15966;
  assign n15968 = n15335 & ~n15571;
  assign n15969 = ~pi0629 & ~n15335;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = n15326 & ~n15970;
  assign n15972 = ~pi0629 & ~n15326;
  assign po0817 = n15971 | n15972;
  assign n15974 = n15335 & ~n15580;
  assign n15975 = ~pi0630 & ~n15335;
  assign n15976 = ~n15974 & ~n15975;
  assign n15977 = n15326 & ~n15976;
  assign n15978 = ~pi0630 & ~n15326;
  assign po0818 = n15977 | n15978;
  assign n15980 = n15335 & ~n15589;
  assign n15981 = ~pi0631 & ~n15335;
  assign n15982 = ~n15980 & ~n15981;
  assign n15983 = n15326 & ~n15982;
  assign n15984 = ~pi0631 & ~n15326;
  assign po0819 = n15983 | n15984;
  assign n15986 = n15335 & ~n15598;
  assign n15987 = ~pi0632 & ~n15335;
  assign n15988 = ~n15986 & ~n15987;
  assign n15989 = n15326 & ~n15988;
  assign n15990 = ~pi0632 & ~n15326;
  assign po0820 = n15989 | n15990;
  assign n15992 = n15335 & ~n15607;
  assign n15993 = ~pi0633 & ~n15335;
  assign n15994 = ~n15992 & ~n15993;
  assign n15995 = n15326 & ~n15994;
  assign n15996 = ~pi0633 & ~n15326;
  assign po0821 = n15995 | n15996;
  assign n15998 = n15335 & ~n15616;
  assign n15999 = ~pi0634 & ~n15335;
  assign n16000 = ~n15998 & ~n15999;
  assign n16001 = n15326 & ~n16000;
  assign n16002 = ~pi0634 & ~n15326;
  assign po0822 = n16001 | n16002;
  assign n16004 = n15427 & ~n15442;
  assign n16005 = ~pi0635 & ~n15427;
  assign n16006 = ~n16004 & ~n16005;
  assign n16007 = n15326 & ~n16006;
  assign n16008 = ~pi0635 & ~n15326;
  assign po0823 = n16007 | n16008;
  assign n16010 = n15427 & ~n15451;
  assign n16011 = ~pi0636 & ~n15427;
  assign n16012 = ~n16010 & ~n16011;
  assign n16013 = n15326 & ~n16012;
  assign n16014 = ~pi0636 & ~n15326;
  assign po0824 = n16013 | n16014;
  assign n16016 = ~n15316 & n15427;
  assign n16017 = ~pi0637 & ~n15427;
  assign n16018 = ~n16016 & ~n16017;
  assign n16019 = n15326 & ~n16018;
  assign n16020 = ~pi0637 & ~n15326;
  assign po0825 = n16019 | n16020;
  assign n16022 = n15427 & ~n15466;
  assign n16023 = ~pi0638 & ~n15427;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = n15326 & ~n16024;
  assign n16026 = ~pi0638 & ~n15326;
  assign po0826 = n16025 | n16026;
  assign n16028 = n15427 & ~n15475;
  assign n16029 = ~pi0639 & ~n15427;
  assign n16030 = ~n16028 & ~n16029;
  assign n16031 = n15326 & ~n16030;
  assign n16032 = ~pi0639 & ~n15326;
  assign po0827 = n16031 | n16032;
  assign n16034 = n15427 & ~n15493;
  assign n16035 = ~pi0640 & ~n15427;
  assign n16036 = ~n16034 & ~n16035;
  assign n16037 = n15326 & ~n16036;
  assign n16038 = ~pi0640 & ~n15326;
  assign po0828 = n16037 | n16038;
  assign n16040 = n15427 & ~n15502;
  assign n16041 = ~pi0641 & ~n15427;
  assign n16042 = ~n16040 & ~n16041;
  assign n16043 = n15326 & ~n16042;
  assign n16044 = ~pi0641 & ~n15326;
  assign po0829 = n16043 | n16044;
  assign n16046 = ~n15332 & n15427;
  assign n16047 = ~pi0642 & ~n15427;
  assign n16048 = ~n16046 & ~n16047;
  assign n16049 = n15326 & ~n16048;
  assign n16050 = ~pi0642 & ~n15326;
  assign po0830 = n16049 | n16050;
  assign n16052 = n15427 & ~n15517;
  assign n16053 = ~pi0643 & ~n15427;
  assign n16054 = ~n16052 & ~n16053;
  assign n16055 = n15326 & ~n16054;
  assign n16056 = ~pi0643 & ~n15326;
  assign po0831 = n16055 | n16056;
  assign n16058 = n15427 & ~n15526;
  assign n16059 = ~pi0644 & ~n15427;
  assign n16060 = ~n16058 & ~n16059;
  assign n16061 = n15326 & ~n16060;
  assign n16062 = ~pi0644 & ~n15326;
  assign po0832 = n16061 | n16062;
  assign n16064 = n15427 & ~n15535;
  assign n16065 = ~pi0645 & ~n15427;
  assign n16066 = ~n16064 & ~n16065;
  assign n16067 = n15326 & ~n16066;
  assign n16068 = ~pi0645 & ~n15326;
  assign po0833 = n16067 | n16068;
  assign n16070 = n15427 & ~n15544;
  assign n16071 = ~pi0646 & ~n15427;
  assign n16072 = ~n16070 & ~n16071;
  assign n16073 = n15326 & ~n16072;
  assign n16074 = ~pi0646 & ~n15326;
  assign po0834 = n16073 | n16074;
  assign n16076 = n15427 & ~n15553;
  assign n16077 = ~pi0647 & ~n15427;
  assign n16078 = ~n16076 & ~n16077;
  assign n16079 = n15326 & ~n16078;
  assign n16080 = ~pi0647 & ~n15326;
  assign po0835 = n16079 | n16080;
  assign n16082 = n15427 & ~n15700;
  assign n16083 = ~pi0648 & ~n15427;
  assign n16084 = ~n16082 & ~n16083;
  assign n16085 = n15326 & ~n16084;
  assign n16086 = ~pi0648 & ~n15326;
  assign po0836 = n16085 | n16086;
  assign n16088 = n15427 & ~n15562;
  assign n16089 = ~pi0649 & ~n15427;
  assign n16090 = ~n16088 & ~n16089;
  assign n16091 = n15326 & ~n16090;
  assign n16092 = ~pi0649 & ~n15326;
  assign po0837 = n16091 | n16092;
  assign n16094 = n15427 & ~n15571;
  assign n16095 = ~pi0650 & ~n15427;
  assign n16096 = ~n16094 & ~n16095;
  assign n16097 = n15326 & ~n16096;
  assign n16098 = ~pi0650 & ~n15326;
  assign po0838 = n16097 | n16098;
  assign n16100 = n15427 & ~n15580;
  assign n16101 = ~pi0651 & ~n15427;
  assign n16102 = ~n16100 & ~n16101;
  assign n16103 = n15326 & ~n16102;
  assign n16104 = ~pi0651 & ~n15326;
  assign po0839 = n16103 | n16104;
  assign n16106 = n15427 & ~n15589;
  assign n16107 = ~pi0652 & ~n15427;
  assign n16108 = ~n16106 & ~n16107;
  assign n16109 = n15326 & ~n16108;
  assign n16110 = ~pi0652 & ~n15326;
  assign po0840 = n16109 | n16110;
  assign n16112 = n15427 & ~n15598;
  assign n16113 = ~pi0653 & ~n15427;
  assign n16114 = ~n16112 & ~n16113;
  assign n16115 = n15326 & ~n16114;
  assign n16116 = ~pi0653 & ~n15326;
  assign po0841 = n16115 | n16116;
  assign n16118 = n15427 & ~n15607;
  assign n16119 = ~pi0654 & ~n15427;
  assign n16120 = ~n16118 & ~n16119;
  assign n16121 = n15326 & ~n16120;
  assign n16122 = ~pi0654 & ~n15326;
  assign po0842 = n16121 | n16122;
  assign n16124 = n15427 & ~n15616;
  assign n16125 = ~pi0655 & ~n15427;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = n15326 & ~n16126;
  assign n16128 = ~pi0655 & ~n15326;
  assign po0843 = n16127 | n16128;
  assign n16130 = n15427 & ~n15625;
  assign n16131 = ~pi0656 & ~n15427;
  assign n16132 = ~n16130 & ~n16131;
  assign n16133 = n15326 & ~n16132;
  assign n16134 = ~pi0656 & ~n15326;
  assign po0844 = n16133 | n16134;
  assign n16136 = n15311 & n15373;
  assign n16137 = ~n15451 & n16136;
  assign n16138 = ~pi0657 & ~n16136;
  assign n16139 = ~n16137 & ~n16138;
  assign n16140 = n15326 & ~n16139;
  assign n16141 = ~pi0657 & ~n15326;
  assign po0845 = n16140 | n16141;
  assign n16143 = ~n15316 & n16136;
  assign n16144 = ~pi0658 & ~n16136;
  assign n16145 = ~n16143 & ~n16144;
  assign n16146 = n15326 & ~n16145;
  assign n16147 = ~pi0658 & ~n15326;
  assign po0846 = n16146 | n16147;
  assign n16149 = ~n15466 & n16136;
  assign n16150 = ~pi0659 & ~n16136;
  assign n16151 = ~n16149 & ~n16150;
  assign n16152 = n15326 & ~n16151;
  assign n16153 = ~pi0659 & ~n15326;
  assign po0847 = n16152 | n16153;
  assign n16155 = ~n15475 & n16136;
  assign n16156 = ~pi0660 & ~n16136;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = n15326 & ~n16157;
  assign n16159 = ~pi0660 & ~n15326;
  assign po0848 = n16158 | n16159;
  assign n16161 = ~n15484 & n16136;
  assign n16162 = ~pi0661 & ~n16136;
  assign n16163 = ~n16161 & ~n16162;
  assign n16164 = n15326 & ~n16163;
  assign n16165 = ~pi0661 & ~n15326;
  assign po0849 = n16164 | n16165;
  assign n16167 = ~n15493 & n16136;
  assign n16168 = ~pi0662 & ~n16136;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = n15326 & ~n16169;
  assign n16171 = ~pi0662 & ~n15326;
  assign po0850 = n16170 | n16171;
  assign n16173 = ~n15502 & n16136;
  assign n16174 = ~pi0663 & ~n16136;
  assign n16175 = ~n16173 & ~n16174;
  assign n16176 = n15326 & ~n16175;
  assign n16177 = ~pi0663 & ~n15326;
  assign po0851 = n16176 | n16177;
  assign n16179 = ~n15332 & n16136;
  assign n16180 = ~pi0664 & ~n16136;
  assign n16181 = ~n16179 & ~n16180;
  assign n16182 = n15326 & ~n16181;
  assign n16183 = ~pi0664 & ~n15326;
  assign po0852 = n16182 | n16183;
  assign n16185 = ~n15709 & n16136;
  assign n16186 = ~pi0665 & ~n16136;
  assign n16187 = ~n16185 & ~n16186;
  assign n16188 = n15326 & ~n16187;
  assign n16189 = ~pi0665 & ~n15326;
  assign po0853 = n16188 | n16189;
  assign n16191 = ~n15526 & n16136;
  assign n16192 = ~pi0666 & ~n16136;
  assign n16193 = ~n16191 & ~n16192;
  assign n16194 = n15326 & ~n16193;
  assign n16195 = ~pi0666 & ~n15326;
  assign po0854 = n16194 | n16195;
  assign n16197 = ~n15535 & n16136;
  assign n16198 = ~pi0667 & ~n16136;
  assign n16199 = ~n16197 & ~n16198;
  assign n16200 = n15326 & ~n16199;
  assign n16201 = ~pi0667 & ~n15326;
  assign po0855 = n16200 | n16201;
  assign n16203 = ~n15544 & n16136;
  assign n16204 = ~pi0668 & ~n16136;
  assign n16205 = ~n16203 & ~n16204;
  assign n16206 = n15326 & ~n16205;
  assign n16207 = ~pi0668 & ~n15326;
  assign po0856 = n16206 | n16207;
  assign n16209 = ~n15553 & n16136;
  assign n16210 = ~pi0669 & ~n16136;
  assign n16211 = ~n16209 & ~n16210;
  assign n16212 = n15326 & ~n16211;
  assign n16213 = ~pi0669 & ~n15326;
  assign po0857 = n16212 | n16213;
  assign n16215 = ~n15700 & n16136;
  assign n16216 = ~pi0670 & ~n16136;
  assign n16217 = ~n16215 & ~n16216;
  assign n16218 = n15326 & ~n16217;
  assign n16219 = ~pi0670 & ~n15326;
  assign po0858 = n16218 | n16219;
  assign n16221 = ~n15571 & n16136;
  assign n16222 = ~pi0671 & ~n16136;
  assign n16223 = ~n16221 & ~n16222;
  assign n16224 = n15326 & ~n16223;
  assign n16225 = ~pi0671 & ~n15326;
  assign po0859 = n16224 | n16225;
  assign n16227 = ~n15580 & n16136;
  assign n16228 = ~pi0672 & ~n16136;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = n15326 & ~n16229;
  assign n16231 = ~pi0672 & ~n15326;
  assign po0860 = n16230 | n16231;
  assign n16233 = ~n15589 & n16136;
  assign n16234 = ~pi0673 & ~n16136;
  assign n16235 = ~n16233 & ~n16234;
  assign n16236 = n15326 & ~n16235;
  assign n16237 = ~pi0673 & ~n15326;
  assign po0861 = n16236 | n16237;
  assign n16239 = ~n15598 & n16136;
  assign n16240 = ~pi0674 & ~n16136;
  assign n16241 = ~n16239 & ~n16240;
  assign n16242 = n15326 & ~n16241;
  assign n16243 = ~pi0674 & ~n15326;
  assign po0862 = n16242 | n16243;
  assign n16245 = ~n15607 & n16136;
  assign n16246 = ~pi0675 & ~n16136;
  assign n16247 = ~n16245 & ~n16246;
  assign n16248 = n15326 & ~n16247;
  assign n16249 = ~pi0675 & ~n15326;
  assign po0863 = n16248 | n16249;
  assign n16251 = ~n15616 & n16136;
  assign n16252 = ~pi0676 & ~n16136;
  assign n16253 = ~n16251 & ~n16252;
  assign n16254 = n15326 & ~n16253;
  assign n16255 = ~pi0676 & ~n15326;
  assign po0864 = n16254 | n16255;
  assign n16257 = ~n15625 & n16136;
  assign n16258 = ~pi0677 & ~n16136;
  assign n16259 = ~n16257 & ~n16258;
  assign n16260 = n15326 & ~n16259;
  assign n16261 = ~pi0677 & ~n15326;
  assign po0865 = n16260 | n16261;
  assign n16263 = n15374 & ~n15442;
  assign n16264 = ~pi0678 & ~n15374;
  assign n16265 = ~n16263 & ~n16264;
  assign n16266 = n15326 & ~n16265;
  assign n16267 = ~pi0678 & ~n15326;
  assign po0866 = n16266 | n16267;
  assign n16269 = ~n15316 & n15374;
  assign n16270 = ~pi0679 & ~n15374;
  assign n16271 = ~n16269 & ~n16270;
  assign n16272 = n15326 & ~n16271;
  assign n16273 = ~pi0679 & ~n15326;
  assign po0867 = n16272 | n16273;
  assign n16275 = n15374 & ~n15466;
  assign n16276 = ~pi0680 & ~n15374;
  assign n16277 = ~n16275 & ~n16276;
  assign n16278 = n15326 & ~n16277;
  assign n16279 = ~pi0680 & ~n15326;
  assign po0868 = n16278 | n16279;
  assign n16281 = n15374 & ~n15475;
  assign n16282 = ~pi0681 & ~n15374;
  assign n16283 = ~n16281 & ~n16282;
  assign n16284 = n15326 & ~n16283;
  assign n16285 = ~pi0681 & ~n15326;
  assign po0869 = n16284 | n16285;
  assign n16287 = n15374 & ~n15484;
  assign n16288 = ~pi0682 & ~n15374;
  assign n16289 = ~n16287 & ~n16288;
  assign n16290 = n15326 & ~n16289;
  assign n16291 = ~pi0682 & ~n15326;
  assign po0870 = n16290 | n16291;
  assign n16293 = n15374 & ~n15493;
  assign n16294 = ~pi0683 & ~n15374;
  assign n16295 = ~n16293 & ~n16294;
  assign n16296 = n15326 & ~n16295;
  assign n16297 = ~pi0683 & ~n15326;
  assign po0871 = n16296 | n16297;
  assign n16299 = ~n15332 & n15374;
  assign n16300 = ~pi0684 & ~n15374;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = n15326 & ~n16301;
  assign n16303 = ~pi0684 & ~n15326;
  assign po0872 = n16302 | n16303;
  assign n16305 = n15374 & ~n15709;
  assign n16306 = ~pi0685 & ~n15374;
  assign n16307 = ~n16305 & ~n16306;
  assign n16308 = n15326 & ~n16307;
  assign n16309 = ~pi0685 & ~n15326;
  assign po0873 = n16308 | n16309;
  assign n16311 = n15374 & ~n15517;
  assign n16312 = ~pi0686 & ~n15374;
  assign n16313 = ~n16311 & ~n16312;
  assign n16314 = n15326 & ~n16313;
  assign n16315 = ~pi0686 & ~n15326;
  assign po0874 = n16314 | n16315;
  assign n16317 = n15374 & ~n15526;
  assign n16318 = ~pi0687 & ~n15374;
  assign n16319 = ~n16317 & ~n16318;
  assign n16320 = n15326 & ~n16319;
  assign n16321 = ~pi0687 & ~n15326;
  assign po0875 = n16320 | n16321;
  assign n16323 = n15374 & ~n15535;
  assign n16324 = ~pi0688 & ~n15374;
  assign n16325 = ~n16323 & ~n16324;
  assign n16326 = n15326 & ~n16325;
  assign n16327 = ~pi0688 & ~n15326;
  assign po0876 = n16326 | n16327;
  assign n16329 = n15374 & ~n15544;
  assign n16330 = ~pi0689 & ~n15374;
  assign n16331 = ~n16329 & ~n16330;
  assign n16332 = n15326 & ~n16331;
  assign n16333 = ~pi0689 & ~n15326;
  assign po0877 = n16332 | n16333;
  assign n16335 = n15374 & ~n15553;
  assign n16336 = ~pi0690 & ~n15374;
  assign n16337 = ~n16335 & ~n16336;
  assign n16338 = n15326 & ~n16337;
  assign n16339 = ~pi0690 & ~n15326;
  assign po0878 = n16338 | n16339;
  assign n16341 = n15374 & ~n15700;
  assign n16342 = ~pi0691 & ~n15374;
  assign n16343 = ~n16341 & ~n16342;
  assign n16344 = n15326 & ~n16343;
  assign n16345 = ~pi0691 & ~n15326;
  assign po0879 = n16344 | n16345;
  assign n16347 = n15374 & ~n15562;
  assign n16348 = ~pi0692 & ~n15374;
  assign n16349 = ~n16347 & ~n16348;
  assign n16350 = n15326 & ~n16349;
  assign n16351 = ~pi0692 & ~n15326;
  assign po0880 = n16350 | n16351;
  assign n16353 = n15374 & ~n15580;
  assign n16354 = ~pi0693 & ~n15374;
  assign n16355 = ~n16353 & ~n16354;
  assign n16356 = n15326 & ~n16355;
  assign n16357 = ~pi0693 & ~n15326;
  assign po0881 = n16356 | n16357;
  assign n16359 = n15374 & ~n15589;
  assign n16360 = ~pi0694 & ~n15374;
  assign n16361 = ~n16359 & ~n16360;
  assign n16362 = n15326 & ~n16361;
  assign n16363 = ~pi0694 & ~n15326;
  assign po0882 = n16362 | n16363;
  assign n16365 = n15374 & ~n15607;
  assign n16366 = ~pi0695 & ~n15374;
  assign n16367 = ~n16365 & ~n16366;
  assign n16368 = n15326 & ~n16367;
  assign n16369 = ~pi0695 & ~n15326;
  assign po0883 = n16368 | n16369;
  assign n16371 = n15374 & ~n15616;
  assign n16372 = ~pi0696 & ~n15374;
  assign n16373 = ~n16371 & ~n16372;
  assign n16374 = n15326 & ~n16373;
  assign n16375 = ~pi0696 & ~n15326;
  assign po0884 = n16374 | n16375;
  assign n16377 = n15374 & ~n15625;
  assign n16378 = ~pi0697 & ~n15374;
  assign n16379 = ~n16377 & ~n16378;
  assign n16380 = n15326 & ~n16379;
  assign n16381 = ~pi0697 & ~n15326;
  assign po0885 = n16380 | n16381;
  assign n16383 = n15400 & ~n15442;
  assign n16384 = ~pi0698 & ~n15400;
  assign n16385 = ~n16383 & ~n16384;
  assign n16386 = n15326 & ~n16385;
  assign n16387 = ~pi0698 & ~n15326;
  assign po0886 = n16386 | n16387;
  assign n16389 = ~n15316 & n15400;
  assign n16390 = ~pi0699 & ~n15400;
  assign n16391 = ~n16389 & ~n16390;
  assign n16392 = n15326 & ~n16391;
  assign n16393 = ~pi0699 & ~n15326;
  assign po0887 = n16392 | n16393;
  assign n16395 = n15400 & ~n15466;
  assign n16396 = ~pi0700 & ~n15400;
  assign n16397 = ~n16395 & ~n16396;
  assign n16398 = n15326 & ~n16397;
  assign n16399 = ~pi0700 & ~n15326;
  assign po0888 = n16398 | n16399;
  assign n16401 = n15400 & ~n15475;
  assign n16402 = ~pi0701 & ~n15400;
  assign n16403 = ~n16401 & ~n16402;
  assign n16404 = n15326 & ~n16403;
  assign n16405 = ~pi0701 & ~n15326;
  assign po0889 = n16404 | n16405;
  assign n16407 = n15400 & ~n15484;
  assign n16408 = ~pi0702 & ~n15400;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = n15326 & ~n16409;
  assign n16411 = ~pi0702 & ~n15326;
  assign po0890 = n16410 | n16411;
  assign n16413 = n15400 & ~n15493;
  assign n16414 = ~pi0703 & ~n15400;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = n15326 & ~n16415;
  assign n16417 = ~pi0703 & ~n15326;
  assign po0891 = n16416 | n16417;
  assign n16419 = ~n15332 & n15400;
  assign n16420 = ~pi0704 & ~n15400;
  assign n16421 = ~n16419 & ~n16420;
  assign n16422 = n15326 & ~n16421;
  assign n16423 = ~pi0704 & ~n15326;
  assign po0892 = n16422 | n16423;
  assign n16425 = n15400 & ~n15709;
  assign n16426 = ~pi0705 & ~n15400;
  assign n16427 = ~n16425 & ~n16426;
  assign n16428 = n15326 & ~n16427;
  assign n16429 = ~pi0705 & ~n15326;
  assign po0893 = n16428 | n16429;
  assign n16431 = n15400 & ~n15517;
  assign n16432 = ~pi0706 & ~n15400;
  assign n16433 = ~n16431 & ~n16432;
  assign n16434 = n15326 & ~n16433;
  assign n16435 = ~pi0706 & ~n15326;
  assign po0894 = n16434 | n16435;
  assign n16437 = n15400 & ~n15526;
  assign n16438 = ~pi0707 & ~n15400;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = n15326 & ~n16439;
  assign n16441 = ~pi0707 & ~n15326;
  assign po0895 = n16440 | n16441;
  assign n16443 = n15400 & ~n15535;
  assign n16444 = ~pi0708 & ~n15400;
  assign n16445 = ~n16443 & ~n16444;
  assign n16446 = n15326 & ~n16445;
  assign n16447 = ~pi0708 & ~n15326;
  assign po0896 = n16446 | n16447;
  assign n16449 = n15400 & ~n15544;
  assign n16450 = ~pi0709 & ~n15400;
  assign n16451 = ~n16449 & ~n16450;
  assign n16452 = n15326 & ~n16451;
  assign n16453 = ~pi0709 & ~n15326;
  assign po0897 = n16452 | n16453;
  assign n16455 = n15400 & ~n15553;
  assign n16456 = ~pi0710 & ~n15400;
  assign n16457 = ~n16455 & ~n16456;
  assign n16458 = n15326 & ~n16457;
  assign n16459 = ~pi0710 & ~n15326;
  assign po0898 = n16458 | n16459;
  assign n16461 = n15400 & ~n15700;
  assign n16462 = ~pi0711 & ~n15400;
  assign n16463 = ~n16461 & ~n16462;
  assign n16464 = n15326 & ~n16463;
  assign n16465 = ~pi0711 & ~n15326;
  assign po0899 = n16464 | n16465;
  assign n16467 = n15400 & ~n15562;
  assign n16468 = ~pi0712 & ~n15400;
  assign n16469 = ~n16467 & ~n16468;
  assign n16470 = n15326 & ~n16469;
  assign n16471 = ~pi0712 & ~n15326;
  assign po0900 = n16470 | n16471;
  assign n16473 = n15400 & ~n15580;
  assign n16474 = ~pi0713 & ~n15400;
  assign n16475 = ~n16473 & ~n16474;
  assign n16476 = n15326 & ~n16475;
  assign n16477 = ~pi0713 & ~n15326;
  assign po0901 = n16476 | n16477;
  assign n16479 = n15400 & ~n15589;
  assign n16480 = ~pi0714 & ~n15400;
  assign n16481 = ~n16479 & ~n16480;
  assign n16482 = n15326 & ~n16481;
  assign n16483 = ~pi0714 & ~n15326;
  assign po0902 = n16482 | n16483;
  assign n16485 = n15400 & ~n15607;
  assign n16486 = ~pi0715 & ~n15400;
  assign n16487 = ~n16485 & ~n16486;
  assign n16488 = n15326 & ~n16487;
  assign n16489 = ~pi0715 & ~n15326;
  assign po0903 = n16488 | n16489;
  assign n16491 = n15400 & ~n15616;
  assign n16492 = ~pi0716 & ~n15400;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = n15326 & ~n16493;
  assign n16495 = ~pi0716 & ~n15326;
  assign po0904 = n16494 | n16495;
  assign n16497 = n15400 & ~n15625;
  assign n16498 = ~pi0717 & ~n15400;
  assign n16499 = ~n16497 & ~n16498;
  assign n16500 = n15326 & ~n16499;
  assign n16501 = ~pi0717 & ~n15326;
  assign po0905 = n16500 | n16501;
  assign n16503 = n15407 & ~n15442;
  assign n16504 = ~pi0718 & ~n15407;
  assign n16505 = ~n16503 & ~n16504;
  assign n16506 = n15326 & ~n16505;
  assign n16507 = ~pi0718 & ~n15326;
  assign po0906 = n16506 | n16507;
  assign n16509 = ~n15316 & n15407;
  assign n16510 = ~pi0719 & ~n15407;
  assign n16511 = ~n16509 & ~n16510;
  assign n16512 = n15326 & ~n16511;
  assign n16513 = ~pi0719 & ~n15326;
  assign po0907 = n16512 | n16513;
  assign n16515 = n15407 & ~n15466;
  assign n16516 = ~pi0720 & ~n15407;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = n15326 & ~n16517;
  assign n16519 = ~pi0720 & ~n15326;
  assign po0908 = n16518 | n16519;
  assign n16521 = n15407 & ~n15475;
  assign n16522 = ~pi0721 & ~n15407;
  assign n16523 = ~n16521 & ~n16522;
  assign n16524 = n15326 & ~n16523;
  assign n16525 = ~pi0721 & ~n15326;
  assign po0909 = n16524 | n16525;
  assign n16527 = n15407 & ~n15484;
  assign n16528 = ~pi0722 & ~n15407;
  assign n16529 = ~n16527 & ~n16528;
  assign n16530 = n15326 & ~n16529;
  assign n16531 = ~pi0722 & ~n15326;
  assign po0910 = n16530 | n16531;
  assign n16533 = n15407 & ~n15502;
  assign n16534 = ~pi0723 & ~n15407;
  assign n16535 = ~n16533 & ~n16534;
  assign n16536 = n15326 & ~n16535;
  assign n16537 = ~pi0723 & ~n15326;
  assign po0911 = n16536 | n16537;
  assign n16539 = n15407 & ~n15709;
  assign n16540 = ~pi0724 & ~n15407;
  assign n16541 = ~n16539 & ~n16540;
  assign n16542 = n15326 & ~n16541;
  assign n16543 = ~pi0724 & ~n15326;
  assign po0912 = n16542 | n16543;
  assign n16545 = n15407 & ~n15517;
  assign n16546 = ~pi0725 & ~n15407;
  assign n16547 = ~n16545 & ~n16546;
  assign n16548 = n15326 & ~n16547;
  assign n16549 = ~pi0725 & ~n15326;
  assign po0913 = n16548 | n16549;
  assign n16551 = n15407 & ~n15526;
  assign n16552 = ~pi0726 & ~n15407;
  assign n16553 = ~n16551 & ~n16552;
  assign n16554 = n15326 & ~n16553;
  assign n16555 = ~pi0726 & ~n15326;
  assign po0914 = n16554 | n16555;
  assign n16557 = n15407 & ~n15535;
  assign n16558 = ~pi0727 & ~n15407;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = n15326 & ~n16559;
  assign n16561 = ~pi0727 & ~n15326;
  assign po0915 = n16560 | n16561;
  assign n16563 = n15407 & ~n15544;
  assign n16564 = ~pi0728 & ~n15407;
  assign n16565 = ~n16563 & ~n16564;
  assign n16566 = n15326 & ~n16565;
  assign n16567 = ~pi0728 & ~n15326;
  assign po0916 = n16566 | n16567;
  assign n16569 = n15407 & ~n15553;
  assign n16570 = ~pi0729 & ~n15407;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = n15326 & ~n16571;
  assign n16573 = ~pi0729 & ~n15326;
  assign po0917 = n16572 | n16573;
  assign n16575 = n15407 & ~n15700;
  assign n16576 = ~pi0730 & ~n15407;
  assign n16577 = ~n16575 & ~n16576;
  assign n16578 = n15326 & ~n16577;
  assign n16579 = ~pi0730 & ~n15326;
  assign po0918 = n16578 | n16579;
  assign n16581 = n15407 & ~n15562;
  assign n16582 = ~pi0731 & ~n15407;
  assign n16583 = ~n16581 & ~n16582;
  assign n16584 = n15326 & ~n16583;
  assign n16585 = ~pi0731 & ~n15326;
  assign po0919 = n16584 | n16585;
  assign n16587 = n15407 & ~n15571;
  assign n16588 = ~pi0732 & ~n15407;
  assign n16589 = ~n16587 & ~n16588;
  assign n16590 = n15326 & ~n16589;
  assign n16591 = ~pi0732 & ~n15326;
  assign po0920 = n16590 | n16591;
  assign n16593 = n15407 & ~n15580;
  assign n16594 = ~pi0733 & ~n15407;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = n15326 & ~n16595;
  assign n16597 = ~pi0733 & ~n15326;
  assign po0921 = n16596 | n16597;
  assign n16599 = n15407 & ~n15589;
  assign n16600 = ~pi0734 & ~n15407;
  assign n16601 = ~n16599 & ~n16600;
  assign n16602 = n15326 & ~n16601;
  assign n16603 = ~pi0734 & ~n15326;
  assign po0922 = n16602 | n16603;
  assign n16605 = n15407 & ~n15598;
  assign n16606 = ~pi0735 & ~n15407;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = n15326 & ~n16607;
  assign n16609 = ~pi0735 & ~n15326;
  assign po0923 = n16608 | n16609;
  assign n16611 = n15407 & ~n15607;
  assign n16612 = ~pi0736 & ~n15407;
  assign n16613 = ~n16611 & ~n16612;
  assign n16614 = n15326 & ~n16613;
  assign n16615 = ~pi0736 & ~n15326;
  assign po0924 = n16614 | n16615;
  assign n16617 = n15407 & ~n15616;
  assign n16618 = ~pi0737 & ~n15407;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = n15326 & ~n16619;
  assign n16621 = ~pi0737 & ~n15326;
  assign po0925 = n16620 | n16621;
  assign n16623 = n15407 & ~n15493;
  assign n16624 = ~pi0738 & ~n15407;
  assign n16625 = ~n16623 & ~n16624;
  assign n16626 = n15326 & ~n16625;
  assign n16627 = ~pi0738 & ~n15326;
  assign po0926 = n16626 | n16627;
  assign n16629 = n15407 & ~n15625;
  assign n16630 = ~pi0739 & ~n15407;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = n15326 & ~n16631;
  assign n16633 = ~pi0739 & ~n15326;
  assign po0927 = n16632 | n16633;
  assign n16635 = n15333 & n15372;
  assign n16636 = ~n15442 & n16635;
  assign n16637 = ~pi0740 & ~n16635;
  assign n16638 = ~n16636 & ~n16637;
  assign n16639 = n15326 & ~n16638;
  assign n16640 = ~pi0740 & ~n15326;
  assign po0928 = n16639 | n16640;
  assign n16642 = ~n15316 & n16635;
  assign n16643 = ~pi0741 & ~n16635;
  assign n16644 = ~n16642 & ~n16643;
  assign n16645 = n15326 & ~n16644;
  assign n16646 = ~pi0741 & ~n15326;
  assign po0929 = n16645 | n16646;
  assign n16648 = ~n15466 & n16635;
  assign n16649 = ~pi0742 & ~n16635;
  assign n16650 = ~n16648 & ~n16649;
  assign n16651 = n15326 & ~n16650;
  assign n16652 = ~pi0742 & ~n15326;
  assign po0930 = n16651 | n16652;
  assign n16654 = ~n15475 & n16635;
  assign n16655 = ~pi0743 & ~n16635;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = n15326 & ~n16656;
  assign n16658 = ~pi0743 & ~n15326;
  assign po0931 = n16657 | n16658;
  assign n16660 = ~n15484 & n16635;
  assign n16661 = ~pi0744 & ~n16635;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = n15326 & ~n16662;
  assign n16664 = ~pi0744 & ~n15326;
  assign po0932 = n16663 | n16664;
  assign n16666 = ~n15493 & n16635;
  assign n16667 = ~pi0745 & ~n16635;
  assign n16668 = ~n16666 & ~n16667;
  assign n16669 = n15326 & ~n16668;
  assign n16670 = ~pi0745 & ~n15326;
  assign po0933 = n16669 | n16670;
  assign n16672 = ~n15332 & n16635;
  assign n16673 = ~pi0746 & ~n16635;
  assign n16674 = ~n16672 & ~n16673;
  assign n16675 = n15326 & ~n16674;
  assign n16676 = ~pi0746 & ~n15326;
  assign po0934 = n16675 | n16676;
  assign n16678 = ~n15709 & n16635;
  assign n16679 = ~pi0747 & ~n16635;
  assign n16680 = ~n16678 & ~n16679;
  assign n16681 = n15326 & ~n16680;
  assign n16682 = ~pi0747 & ~n15326;
  assign po0935 = n16681 | n16682;
  assign n16684 = ~n15517 & n16635;
  assign n16685 = ~pi0748 & ~n16635;
  assign n16686 = ~n16684 & ~n16685;
  assign n16687 = n15326 & ~n16686;
  assign n16688 = ~pi0748 & ~n15326;
  assign po0936 = n16687 | n16688;
  assign n16690 = ~n15535 & n16635;
  assign n16691 = ~pi0749 & ~n16635;
  assign n16692 = ~n16690 & ~n16691;
  assign n16693 = n15326 & ~n16692;
  assign n16694 = ~pi0749 & ~n15326;
  assign po0937 = n16693 | n16694;
  assign n16696 = ~n15544 & n16635;
  assign n16697 = ~pi0750 & ~n16635;
  assign n16698 = ~n16696 & ~n16697;
  assign n16699 = n15326 & ~n16698;
  assign n16700 = ~pi0750 & ~n15326;
  assign po0938 = n16699 | n16700;
  assign n16702 = ~n15553 & n16635;
  assign n16703 = ~pi0751 & ~n16635;
  assign n16704 = ~n16702 & ~n16703;
  assign n16705 = n15326 & ~n16704;
  assign n16706 = ~pi0751 & ~n15326;
  assign po0939 = n16705 | n16706;
  assign n16708 = ~n15700 & n16635;
  assign n16709 = ~pi0752 & ~n16635;
  assign n16710 = ~n16708 & ~n16709;
  assign n16711 = n15326 & ~n16710;
  assign n16712 = ~pi0752 & ~n15326;
  assign po0940 = n16711 | n16712;
  assign n16714 = ~n15562 & n16635;
  assign n16715 = ~pi0753 & ~n16635;
  assign n16716 = ~n16714 & ~n16715;
  assign n16717 = n15326 & ~n16716;
  assign n16718 = ~pi0753 & ~n15326;
  assign po0941 = n16717 | n16718;
  assign n16720 = ~n15580 & n16635;
  assign n16721 = ~pi0754 & ~n16635;
  assign n16722 = ~n16720 & ~n16721;
  assign n16723 = n15326 & ~n16722;
  assign n16724 = ~pi0754 & ~n15326;
  assign po0942 = n16723 | n16724;
  assign n16726 = ~n15589 & n16635;
  assign n16727 = ~pi0755 & ~n16635;
  assign n16728 = ~n16726 & ~n16727;
  assign n16729 = n15326 & ~n16728;
  assign n16730 = ~pi0755 & ~n15326;
  assign po0943 = n16729 | n16730;
  assign n16732 = ~n15607 & n16635;
  assign n16733 = ~pi0756 & ~n16635;
  assign n16734 = ~n16732 & ~n16733;
  assign n16735 = n15326 & ~n16734;
  assign n16736 = ~pi0756 & ~n15326;
  assign po0944 = n16735 | n16736;
  assign n16738 = ~n15616 & n16635;
  assign n16739 = ~pi0757 & ~n16635;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = n15326 & ~n16740;
  assign n16742 = ~pi0757 & ~n15326;
  assign po0945 = n16741 | n16742;
  assign n16744 = ~n15625 & n16635;
  assign n16745 = ~pi0758 & ~n16635;
  assign n16746 = ~n16744 & ~n16745;
  assign n16747 = n15326 & ~n16746;
  assign n16748 = ~pi0758 & ~n15326;
  assign po0946 = n16747 | n16748;
  assign n16750 = n15434 & ~n15442;
  assign n16751 = ~pi0759 & ~n15434;
  assign n16752 = ~n16750 & ~n16751;
  assign n16753 = n15326 & ~n16752;
  assign n16754 = ~pi0759 & ~n15326;
  assign po0947 = n16753 | n16754;
  assign n16756 = ~n15316 & n15434;
  assign n16757 = ~pi0760 & ~n15434;
  assign n16758 = ~n16756 & ~n16757;
  assign n16759 = n15326 & ~n16758;
  assign n16760 = ~pi0760 & ~n15326;
  assign po0948 = n16759 | n16760;
  assign n16762 = n15434 & ~n15466;
  assign n16763 = ~pi0761 & ~n15434;
  assign n16764 = ~n16762 & ~n16763;
  assign n16765 = n15326 & ~n16764;
  assign n16766 = ~pi0761 & ~n15326;
  assign po0949 = n16765 | n16766;
  assign n16768 = n15434 & ~n15475;
  assign n16769 = ~pi0762 & ~n15434;
  assign n16770 = ~n16768 & ~n16769;
  assign n16771 = n15326 & ~n16770;
  assign n16772 = ~pi0762 & ~n15326;
  assign po0950 = n16771 | n16772;
  assign n16774 = n15434 & ~n15484;
  assign n16775 = ~pi0763 & ~n15434;
  assign n16776 = ~n16774 & ~n16775;
  assign n16777 = n15326 & ~n16776;
  assign n16778 = ~pi0763 & ~n15326;
  assign po0951 = n16777 | n16778;
  assign n16780 = n15434 & ~n15493;
  assign n16781 = ~pi0764 & ~n15434;
  assign n16782 = ~n16780 & ~n16781;
  assign n16783 = n15326 & ~n16782;
  assign n16784 = ~pi0764 & ~n15326;
  assign po0952 = n16783 | n16784;
  assign n16786 = ~n15332 & n15434;
  assign n16787 = ~pi0765 & ~n15434;
  assign n16788 = ~n16786 & ~n16787;
  assign n16789 = n15326 & ~n16788;
  assign n16790 = ~pi0765 & ~n15326;
  assign po0953 = n16789 | n16790;
  assign n16792 = n15434 & ~n15709;
  assign n16793 = ~pi0766 & ~n15434;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = n15326 & ~n16794;
  assign n16796 = ~pi0766 & ~n15326;
  assign po0954 = n16795 | n16796;
  assign n16798 = n15434 & ~n15517;
  assign n16799 = ~pi0767 & ~n15434;
  assign n16800 = ~n16798 & ~n16799;
  assign n16801 = n15326 & ~n16800;
  assign n16802 = ~pi0767 & ~n15326;
  assign po0955 = n16801 | n16802;
  assign n16804 = n15434 & ~n15526;
  assign n16805 = ~pi0768 & ~n15434;
  assign n16806 = ~n16804 & ~n16805;
  assign n16807 = n15326 & ~n16806;
  assign n16808 = ~pi0768 & ~n15326;
  assign po0956 = n16807 | n16808;
  assign n16810 = n15434 & ~n15535;
  assign n16811 = ~pi0769 & ~n15434;
  assign n16812 = ~n16810 & ~n16811;
  assign n16813 = n15326 & ~n16812;
  assign n16814 = ~pi0769 & ~n15326;
  assign po0957 = n16813 | n16814;
  assign n16816 = n15434 & ~n15544;
  assign n16817 = ~pi0770 & ~n15434;
  assign n16818 = ~n16816 & ~n16817;
  assign n16819 = n15326 & ~n16818;
  assign n16820 = ~pi0770 & ~n15326;
  assign po0958 = n16819 | n16820;
  assign n16822 = n15434 & ~n15553;
  assign n16823 = ~pi0771 & ~n15434;
  assign n16824 = ~n16822 & ~n16823;
  assign n16825 = n15326 & ~n16824;
  assign n16826 = ~pi0771 & ~n15326;
  assign po0959 = n16825 | n16826;
  assign n16828 = n15434 & ~n15700;
  assign n16829 = ~pi0772 & ~n15434;
  assign n16830 = ~n16828 & ~n16829;
  assign n16831 = n15326 & ~n16830;
  assign n16832 = ~pi0772 & ~n15326;
  assign po0960 = n16831 | n16832;
  assign n16834 = n15434 & ~n15562;
  assign n16835 = ~pi0773 & ~n15434;
  assign n16836 = ~n16834 & ~n16835;
  assign n16837 = n15326 & ~n16836;
  assign n16838 = ~pi0773 & ~n15326;
  assign po0961 = n16837 | n16838;
  assign n16840 = n15434 & ~n15580;
  assign n16841 = ~pi0774 & ~n15434;
  assign n16842 = ~n16840 & ~n16841;
  assign n16843 = n15326 & ~n16842;
  assign n16844 = ~pi0774 & ~n15326;
  assign po0962 = n16843 | n16844;
  assign n16846 = n15434 & ~n15589;
  assign n16847 = ~pi0775 & ~n15434;
  assign n16848 = ~n16846 & ~n16847;
  assign n16849 = n15326 & ~n16848;
  assign n16850 = ~pi0775 & ~n15326;
  assign po0963 = n16849 | n16850;
  assign n16852 = n15434 & ~n15607;
  assign n16853 = ~pi0776 & ~n15434;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = n15326 & ~n16854;
  assign n16856 = ~pi0776 & ~n15326;
  assign po0964 = n16855 | n16856;
  assign n16858 = n15434 & ~n15616;
  assign n16859 = ~pi0777 & ~n15434;
  assign n16860 = ~n16858 & ~n16859;
  assign n16861 = n15326 & ~n16860;
  assign n16862 = ~pi0777 & ~n15326;
  assign po0965 = n16861 | n16862;
  assign n16864 = n15434 & ~n15625;
  assign n16865 = ~pi0778 & ~n15434;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = n15326 & ~n16866;
  assign n16868 = ~pi0778 & ~n15326;
  assign po0966 = n16867 | n16868;
  assign n16870 = n15311 & n15384;
  assign n16871 = ~pi0779 & ~n16870;
  assign n16872 = ~n15442 & n16870;
  assign n16873 = ~n16871 & ~n16872;
  assign n16874 = n15326 & ~n16873;
  assign n16875 = ~pi0779 & ~n15326;
  assign po0967 = n16874 | n16875;
  assign n16877 = ~pi0780 & ~n16870;
  assign n16878 = ~n15451 & n16870;
  assign n16879 = ~n16877 & ~n16878;
  assign n16880 = n15326 & ~n16879;
  assign n16881 = ~pi0780 & ~n15326;
  assign po0968 = n16880 | n16881;
  assign n16883 = ~pi0781 & ~n16870;
  assign n16884 = ~n15316 & n16870;
  assign n16885 = ~n16883 & ~n16884;
  assign n16886 = n15326 & ~n16885;
  assign n16887 = ~pi0781 & ~n15326;
  assign po0969 = n16886 | n16887;
  assign n16889 = ~pi0782 & ~n16870;
  assign n16890 = ~n15466 & n16870;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = n15326 & ~n16891;
  assign n16893 = ~pi0782 & ~n15326;
  assign po0970 = n16892 | n16893;
  assign n16895 = ~pi0783 & ~n16870;
  assign n16896 = ~n15475 & n16870;
  assign n16897 = ~n16895 & ~n16896;
  assign n16898 = n15326 & ~n16897;
  assign n16899 = ~pi0783 & ~n15326;
  assign po0971 = n16898 | n16899;
  assign n16901 = ~pi0784 & ~n16870;
  assign n16902 = ~n15484 & n16870;
  assign n16903 = ~n16901 & ~n16902;
  assign n16904 = n15326 & ~n16903;
  assign n16905 = ~pi0784 & ~n15326;
  assign po0972 = n16904 | n16905;
  assign n16907 = ~pi0785 & ~n16870;
  assign n16908 = ~n15493 & n16870;
  assign n16909 = ~n16907 & ~n16908;
  assign n16910 = n15326 & ~n16909;
  assign n16911 = ~pi0785 & ~n15326;
  assign po0973 = n16910 | n16911;
  assign n16913 = ~pi0786 & ~n16870;
  assign n16914 = ~n15502 & n16870;
  assign n16915 = ~n16913 & ~n16914;
  assign n16916 = n15326 & ~n16915;
  assign n16917 = ~pi0786 & ~n15326;
  assign po0974 = n16916 | n16917;
  assign n16919 = ~pi0787 & ~n16870;
  assign n16920 = ~n15709 & n16870;
  assign n16921 = ~n16919 & ~n16920;
  assign n16922 = n15326 & ~n16921;
  assign n16923 = ~pi0787 & ~n15326;
  assign po0975 = n16922 | n16923;
  assign n16925 = ~pi0788 & ~n16870;
  assign n16926 = ~n15517 & n16870;
  assign n16927 = ~n16925 & ~n16926;
  assign n16928 = n15326 & ~n16927;
  assign n16929 = ~pi0788 & ~n15326;
  assign po0976 = n16928 | n16929;
  assign n16931 = ~pi0789 & ~n16870;
  assign n16932 = ~n15526 & n16870;
  assign n16933 = ~n16931 & ~n16932;
  assign n16934 = n15326 & ~n16933;
  assign n16935 = ~pi0789 & ~n15326;
  assign po0977 = n16934 | n16935;
  assign n16937 = ~pi0790 & ~n16870;
  assign n16938 = ~n15535 & n16870;
  assign n16939 = ~n16937 & ~n16938;
  assign n16940 = n15326 & ~n16939;
  assign n16941 = ~pi0790 & ~n15326;
  assign po0978 = n16940 | n16941;
  assign n16943 = ~pi0791 & ~n16870;
  assign n16944 = ~n15544 & n16870;
  assign n16945 = ~n16943 & ~n16944;
  assign n16946 = n15326 & ~n16945;
  assign n16947 = ~pi0791 & ~n15326;
  assign po0979 = n16946 | n16947;
  assign n16949 = ~pi0792 & ~n16870;
  assign n16950 = ~n15553 & n16870;
  assign n16951 = ~n16949 & ~n16950;
  assign n16952 = n15326 & ~n16951;
  assign n16953 = ~pi0792 & ~n15326;
  assign po0980 = n16952 | n16953;
  assign n16955 = ~pi0793 & ~n16870;
  assign n16956 = ~n15700 & n16870;
  assign n16957 = ~n16955 & ~n16956;
  assign n16958 = n15326 & ~n16957;
  assign n16959 = ~pi0793 & ~n15326;
  assign po0981 = n16958 | n16959;
  assign n16961 = ~pi0794 & ~n16870;
  assign n16962 = ~n15562 & n16870;
  assign n16963 = ~n16961 & ~n16962;
  assign n16964 = n15326 & ~n16963;
  assign n16965 = ~pi0794 & ~n15326;
  assign po0982 = n16964 | n16965;
  assign n16967 = ~pi0795 & ~n16870;
  assign n16968 = ~n15571 & n16870;
  assign n16969 = ~n16967 & ~n16968;
  assign n16970 = n15326 & ~n16969;
  assign n16971 = ~pi0795 & ~n15326;
  assign po0983 = n16970 | n16971;
  assign n16973 = ~pi0796 & ~n16870;
  assign n16974 = ~n15580 & n16870;
  assign n16975 = ~n16973 & ~n16974;
  assign n16976 = n15326 & ~n16975;
  assign n16977 = ~pi0796 & ~n15326;
  assign po0984 = n16976 | n16977;
  assign n16979 = ~pi0797 & ~n16870;
  assign n16980 = ~n15589 & n16870;
  assign n16981 = ~n16979 & ~n16980;
  assign n16982 = n15326 & ~n16981;
  assign n16983 = ~pi0797 & ~n15326;
  assign po0985 = n16982 | n16983;
  assign n16985 = ~pi0798 & ~n16870;
  assign n16986 = n15377 & n16870;
  assign n16987 = ~n16985 & ~n16986;
  assign n16988 = n15326 & ~n16987;
  assign n16989 = ~pi0798 & ~n15326;
  assign po0986 = n16988 | n16989;
  assign n16991 = ~pi0799 & ~n16870;
  assign n16992 = ~n15598 & n16870;
  assign n16993 = ~n16991 & ~n16992;
  assign n16994 = n15326 & ~n16993;
  assign n16995 = ~pi0799 & ~n15326;
  assign po0987 = n16994 | n16995;
  assign n16997 = ~pi0800 & ~n16870;
  assign n16998 = ~n15607 & n16870;
  assign n16999 = ~n16997 & ~n16998;
  assign n17000 = n15326 & ~n16999;
  assign n17001 = ~pi0800 & ~n15326;
  assign po0988 = n17000 | n17001;
  assign n17003 = ~pi0801 & ~n16870;
  assign n17004 = ~n15625 & n16870;
  assign n17005 = ~n17003 & ~n17004;
  assign n17006 = n15326 & ~n17005;
  assign n17007 = ~pi0801 & ~n15326;
  assign po0989 = n17006 | n17007;
  assign n17009 = ~pi0802 & ~n16870;
  assign n17010 = ~n15616 & n16870;
  assign n17011 = ~n17009 & ~n17010;
  assign n17012 = n15326 & ~n17011;
  assign n17013 = ~pi0802 & ~n15326;
  assign po0990 = n17012 | n17013;
  assign n17015 = n15311 & n15333;
  assign n17016 = ~pi0803 & ~n17015;
  assign n17017 = ~n15442 & n17015;
  assign n17018 = ~n17016 & ~n17017;
  assign n17019 = n15326 & ~n17018;
  assign n17020 = ~pi0803 & ~n15326;
  assign po0991 = n17019 | n17020;
  assign n17022 = ~pi0804 & ~n17015;
  assign n17023 = ~n15451 & n17015;
  assign n17024 = ~n17022 & ~n17023;
  assign n17025 = n15326 & ~n17024;
  assign n17026 = ~pi0804 & ~n15326;
  assign po0992 = n17025 | n17026;
  assign n17028 = ~pi0805 & ~n17015;
  assign n17029 = ~n15466 & n17015;
  assign n17030 = ~n17028 & ~n17029;
  assign n17031 = n15326 & ~n17030;
  assign n17032 = ~pi0805 & ~n15326;
  assign po0993 = n17031 | n17032;
  assign n17034 = ~pi0806 & ~n17015;
  assign n17035 = ~n15475 & n17015;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = n15326 & ~n17036;
  assign n17038 = ~pi0806 & ~n15326;
  assign po0994 = n17037 | n17038;
  assign n17040 = ~pi0807 & ~n17015;
  assign n17041 = ~n15484 & n17015;
  assign n17042 = ~n17040 & ~n17041;
  assign n17043 = n15326 & ~n17042;
  assign n17044 = ~pi0807 & ~n15326;
  assign po0995 = n17043 | n17044;
  assign n17046 = ~pi0808 & ~n17015;
  assign n17047 = ~n15493 & n17015;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = n15326 & ~n17048;
  assign n17050 = ~pi0808 & ~n15326;
  assign po0996 = n17049 | n17050;
  assign n17052 = ~pi0809 & ~n17015;
  assign n17053 = ~n15502 & n17015;
  assign n17054 = ~n17052 & ~n17053;
  assign n17055 = n15326 & ~n17054;
  assign n17056 = ~pi0809 & ~n15326;
  assign po0997 = n17055 | n17056;
  assign n17058 = ~pi0810 & ~n17015;
  assign n17059 = ~n15709 & n17015;
  assign n17060 = ~n17058 & ~n17059;
  assign n17061 = n15326 & ~n17060;
  assign n17062 = ~pi0810 & ~n15326;
  assign po0998 = n17061 | n17062;
  assign n17064 = ~pi0811 & ~n17015;
  assign n17065 = ~n15517 & n17015;
  assign n17066 = ~n17064 & ~n17065;
  assign n17067 = n15326 & ~n17066;
  assign n17068 = ~pi0811 & ~n15326;
  assign po0999 = n17067 | n17068;
  assign n17070 = ~pi0812 & ~n17015;
  assign n17071 = ~n15526 & n17015;
  assign n17072 = ~n17070 & ~n17071;
  assign n17073 = n15326 & ~n17072;
  assign n17074 = ~pi0812 & ~n15326;
  assign po1000 = n17073 | n17074;
  assign n17076 = ~pi0813 & ~n17015;
  assign n17077 = ~n15535 & n17015;
  assign n17078 = ~n17076 & ~n17077;
  assign n17079 = n15326 & ~n17078;
  assign n17080 = ~pi0813 & ~n15326;
  assign po1001 = n17079 | n17080;
  assign n17082 = ~pi0814 & ~n17015;
  assign n17083 = ~n15544 & n17015;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = n15326 & ~n17084;
  assign n17086 = ~pi0814 & ~n15326;
  assign po1002 = n17085 | n17086;
  assign n17088 = ~pi0815 & ~n17015;
  assign n17089 = ~n15553 & n17015;
  assign n17090 = ~n17088 & ~n17089;
  assign n17091 = n15326 & ~n17090;
  assign n17092 = ~pi0815 & ~n15326;
  assign po1003 = n17091 | n17092;
  assign n17094 = ~pi0816 & ~n17015;
  assign n17095 = ~n15700 & n17015;
  assign n17096 = ~n17094 & ~n17095;
  assign n17097 = n15326 & ~n17096;
  assign n17098 = ~pi0816 & ~n15326;
  assign po1004 = n17097 | n17098;
  assign n17100 = ~pi0817 & ~n17015;
  assign n17101 = ~n15562 & n17015;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = n15326 & ~n17102;
  assign n17104 = ~pi0817 & ~n15326;
  assign po1005 = n17103 | n17104;
  assign n17106 = ~pi0818 & ~n17015;
  assign n17107 = ~n15571 & n17015;
  assign n17108 = ~n17106 & ~n17107;
  assign n17109 = n15326 & ~n17108;
  assign n17110 = ~pi0818 & ~n15326;
  assign po1006 = n17109 | n17110;
  assign n17112 = ~pi0819 & ~n17015;
  assign n17113 = ~n15580 & n17015;
  assign n17114 = ~n17112 & ~n17113;
  assign n17115 = n15326 & ~n17114;
  assign n17116 = ~pi0819 & ~n15326;
  assign po1007 = n17115 | n17116;
  assign n17118 = ~pi0820 & ~n17015;
  assign n17119 = ~n15589 & n17015;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = n15326 & ~n17120;
  assign n17122 = ~pi0820 & ~n15326;
  assign po1008 = n17121 | n17122;
  assign n17124 = ~pi0821 & ~n17015;
  assign n17125 = n15377 & n17015;
  assign n17126 = ~n17124 & ~n17125;
  assign n17127 = n15326 & ~n17126;
  assign n17128 = ~pi0821 & ~n15326;
  assign po1009 = n17127 | n17128;
  assign n17130 = ~pi0822 & ~n17015;
  assign n17131 = ~n15598 & n17015;
  assign n17132 = ~n17130 & ~n17131;
  assign n17133 = n15326 & ~n17132;
  assign n17134 = ~pi0822 & ~n15326;
  assign po1010 = n17133 | n17134;
  assign n17136 = ~pi0823 & ~n17015;
  assign n17137 = ~n15607 & n17015;
  assign n17138 = ~n17136 & ~n17137;
  assign n17139 = n15326 & ~n17138;
  assign n17140 = ~pi0823 & ~n15326;
  assign po1011 = n17139 | n17140;
  assign n17142 = ~pi0824 & ~n17015;
  assign n17143 = ~n15616 & n17015;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 = n15326 & ~n17144;
  assign n17146 = ~pi0824 & ~n15326;
  assign po1012 = n17145 | n17146;
  assign n17148 = ~pi0825 & ~n17015;
  assign n17149 = ~n15625 & n17015;
  assign n17150 = ~n17148 & ~n17149;
  assign n17151 = n15326 & ~n17150;
  assign n17152 = ~pi0825 & ~n15326;
  assign po1013 = n17151 | n17152;
  assign n17154 = n15310 & n15385;
  assign n17155 = ~pi0826 & ~n17154;
  assign n17156 = ~n15442 & n17154;
  assign n17157 = ~n17155 & ~n17156;
  assign n17158 = n15326 & ~n17157;
  assign n17159 = ~pi0826 & ~n15326;
  assign po1014 = n17158 | n17159;
  assign n17161 = ~pi0827 & ~n17154;
  assign n17162 = ~n15451 & n17154;
  assign n17163 = ~n17161 & ~n17162;
  assign n17164 = n15326 & ~n17163;
  assign n17165 = ~pi0827 & ~n15326;
  assign po1015 = n17164 | n17165;
  assign n17167 = ~pi0828 & ~n17154;
  assign n17168 = ~n15316 & n17154;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = n15326 & ~n17169;
  assign n17171 = ~pi0828 & ~n15326;
  assign po1016 = n17170 | n17171;
  assign n17173 = ~pi0829 & ~n17154;
  assign n17174 = ~n15466 & n17154;
  assign n17175 = ~n17173 & ~n17174;
  assign n17176 = n15326 & ~n17175;
  assign n17177 = ~pi0829 & ~n15326;
  assign po1017 = n17176 | n17177;
  assign n17179 = ~pi0830 & ~n17154;
  assign n17180 = ~n15475 & n17154;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = n15326 & ~n17181;
  assign n17183 = ~pi0830 & ~n15326;
  assign po1018 = n17182 | n17183;
  assign n17185 = ~pi0831 & ~n17154;
  assign n17186 = ~n15484 & n17154;
  assign n17187 = ~n17185 & ~n17186;
  assign n17188 = n15326 & ~n17187;
  assign n17189 = ~pi0831 & ~n15326;
  assign po1019 = n17188 | n17189;
  assign n17191 = ~pi0832 & ~n17154;
  assign n17192 = ~n15493 & n17154;
  assign n17193 = ~n17191 & ~n17192;
  assign n17194 = n15326 & ~n17193;
  assign n17195 = ~pi0832 & ~n15326;
  assign po1020 = n17194 | n17195;
  assign n17197 = ~pi0833 & ~n17154;
  assign n17198 = ~n15502 & n17154;
  assign n17199 = ~n17197 & ~n17198;
  assign n17200 = n15326 & ~n17199;
  assign n17201 = ~pi0833 & ~n15326;
  assign po1021 = n17200 | n17201;
  assign n17203 = ~pi0834 & ~n17154;
  assign n17204 = ~n15709 & n17154;
  assign n17205 = ~n17203 & ~n17204;
  assign n17206 = n15326 & ~n17205;
  assign n17207 = ~pi0834 & ~n15326;
  assign po1022 = n17206 | n17207;
  assign n17209 = ~pi0835 & ~n17154;
  assign n17210 = ~n15517 & n17154;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = n15326 & ~n17211;
  assign n17213 = ~pi0835 & ~n15326;
  assign po1023 = n17212 | n17213;
  assign n17215 = ~pi0836 & ~n17154;
  assign n17216 = ~n15526 & n17154;
  assign n17217 = ~n17215 & ~n17216;
  assign n17218 = n15326 & ~n17217;
  assign n17219 = ~pi0836 & ~n15326;
  assign po1024 = n17218 | n17219;
  assign n17221 = ~pi0837 & ~n17154;
  assign n17222 = ~n15535 & n17154;
  assign n17223 = ~n17221 & ~n17222;
  assign n17224 = n15326 & ~n17223;
  assign n17225 = ~pi0837 & ~n15326;
  assign po1025 = n17224 | n17225;
  assign n17227 = ~pi0838 & ~n17154;
  assign n17228 = ~n15544 & n17154;
  assign n17229 = ~n17227 & ~n17228;
  assign n17230 = n15326 & ~n17229;
  assign n17231 = ~pi0838 & ~n15326;
  assign po1026 = n17230 | n17231;
  assign n17233 = ~pi0839 & ~n17154;
  assign n17234 = ~n15553 & n17154;
  assign n17235 = ~n17233 & ~n17234;
  assign n17236 = n15326 & ~n17235;
  assign n17237 = ~pi0839 & ~n15326;
  assign po1027 = n17236 | n17237;
  assign n17239 = ~pi0840 & ~n17154;
  assign n17240 = ~n15700 & n17154;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = n15326 & ~n17241;
  assign n17243 = ~pi0840 & ~n15326;
  assign po1028 = n17242 | n17243;
  assign n17245 = ~pi0841 & ~n17154;
  assign n17246 = ~n15562 & n17154;
  assign n17247 = ~n17245 & ~n17246;
  assign n17248 = n15326 & ~n17247;
  assign n17249 = ~pi0841 & ~n15326;
  assign po1029 = n17248 | n17249;
  assign n17251 = ~pi0842 & ~n17154;
  assign n17252 = ~n15571 & n17154;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = n15326 & ~n17253;
  assign n17255 = ~pi0842 & ~n15326;
  assign po1030 = n17254 | n17255;
  assign n17257 = ~pi0843 & ~n17154;
  assign n17258 = ~n15580 & n17154;
  assign n17259 = ~n17257 & ~n17258;
  assign n17260 = n15326 & ~n17259;
  assign n17261 = ~pi0843 & ~n15326;
  assign po1031 = n17260 | n17261;
  assign n17263 = ~pi0844 & ~n17154;
  assign n17264 = ~n15589 & n17154;
  assign n17265 = ~n17263 & ~n17264;
  assign n17266 = n15326 & ~n17265;
  assign n17267 = ~pi0844 & ~n15326;
  assign po1032 = n17266 | n17267;
  assign n17269 = ~pi0845 & ~n17154;
  assign n17270 = n15377 & n17154;
  assign n17271 = ~n17269 & ~n17270;
  assign n17272 = n15326 & ~n17271;
  assign n17273 = ~pi0845 & ~n15326;
  assign po1033 = n17272 | n17273;
  assign n17275 = ~pi0846 & ~n17154;
  assign n17276 = ~n15598 & n17154;
  assign n17277 = ~n17275 & ~n17276;
  assign n17278 = n15326 & ~n17277;
  assign n17279 = ~pi0846 & ~n15326;
  assign po1034 = n17278 | n17279;
  assign n17281 = ~pi0847 & ~n17154;
  assign n17282 = ~n15607 & n17154;
  assign n17283 = ~n17281 & ~n17282;
  assign n17284 = n15326 & ~n17283;
  assign n17285 = ~pi0847 & ~n15326;
  assign po1035 = n17284 | n17285;
  assign n17287 = ~pi0848 & ~n17154;
  assign n17288 = ~n15616 & n17154;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = n15326 & ~n17289;
  assign n17291 = ~pi0848 & ~n15326;
  assign po1036 = n17290 | n17291;
  assign n17293 = ~pi0849 & ~n17154;
  assign n17294 = ~n15625 & n17154;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = n15326 & ~n17295;
  assign n17297 = ~pi0849 & ~n15326;
  assign po1037 = n17296 | n17297;
  assign n17299 = ~pi0850 & ~n15312;
  assign n17300 = n15312 & ~n15442;
  assign n17301 = ~n17299 & ~n17300;
  assign n17302 = n15326 & ~n17301;
  assign n17303 = ~pi0850 & ~n15326;
  assign po1038 = n17302 | n17303;
  assign n17305 = ~pi0851 & ~n15312;
  assign n17306 = n15312 & ~n15451;
  assign n17307 = ~n17305 & ~n17306;
  assign n17308 = n15326 & ~n17307;
  assign n17309 = ~pi0851 & ~n15326;
  assign po1039 = n17308 | n17309;
  assign n17311 = ~pi0852 & ~n15312;
  assign n17312 = n15312 & ~n15466;
  assign n17313 = ~n17311 & ~n17312;
  assign n17314 = n15326 & ~n17313;
  assign n17315 = ~pi0852 & ~n15326;
  assign po1040 = n17314 | n17315;
  assign n17317 = ~pi0853 & ~n15312;
  assign n17318 = n15312 & ~n15475;
  assign n17319 = ~n17317 & ~n17318;
  assign n17320 = n15326 & ~n17319;
  assign n17321 = ~pi0853 & ~n15326;
  assign po1041 = n17320 | n17321;
  assign n17323 = ~pi0854 & ~n15312;
  assign n17324 = n15312 & ~n15484;
  assign n17325 = ~n17323 & ~n17324;
  assign n17326 = n15326 & ~n17325;
  assign n17327 = ~pi0854 & ~n15326;
  assign po1042 = n17326 | n17327;
  assign n17329 = ~pi0855 & ~n15312;
  assign n17330 = n15312 & ~n15493;
  assign n17331 = ~n17329 & ~n17330;
  assign n17332 = n15326 & ~n17331;
  assign n17333 = ~pi0855 & ~n15326;
  assign po1043 = n17332 | n17333;
  assign n17335 = ~pi0856 & ~n15312;
  assign n17336 = n15312 & ~n15502;
  assign n17337 = ~n17335 & ~n17336;
  assign n17338 = n15326 & ~n17337;
  assign n17339 = ~pi0856 & ~n15326;
  assign po1044 = n17338 | n17339;
  assign n17341 = ~pi0857 & ~n15312;
  assign n17342 = n15312 & ~n15709;
  assign n17343 = ~n17341 & ~n17342;
  assign n17344 = n15326 & ~n17343;
  assign n17345 = ~pi0857 & ~n15326;
  assign po1045 = n17344 | n17345;
  assign n17347 = ~pi0858 & ~n15312;
  assign n17348 = n15312 & ~n15517;
  assign n17349 = ~n17347 & ~n17348;
  assign n17350 = n15326 & ~n17349;
  assign n17351 = ~pi0858 & ~n15326;
  assign po1046 = n17350 | n17351;
  assign n17353 = ~pi0859 & ~n15312;
  assign n17354 = n15312 & ~n15526;
  assign n17355 = ~n17353 & ~n17354;
  assign n17356 = n15326 & ~n17355;
  assign n17357 = ~pi0859 & ~n15326;
  assign po1047 = n17356 | n17357;
  assign n17359 = ~pi0860 & ~n15312;
  assign n17360 = n15312 & ~n15535;
  assign n17361 = ~n17359 & ~n17360;
  assign n17362 = n15326 & ~n17361;
  assign n17363 = ~pi0860 & ~n15326;
  assign po1048 = n17362 | n17363;
  assign n17365 = ~pi0861 & ~n15312;
  assign n17366 = n15312 & ~n15544;
  assign n17367 = ~n17365 & ~n17366;
  assign n17368 = n15326 & ~n17367;
  assign n17369 = ~pi0861 & ~n15326;
  assign po1049 = n17368 | n17369;
  assign n17371 = ~pi0862 & ~n15312;
  assign n17372 = n15312 & ~n15553;
  assign n17373 = ~n17371 & ~n17372;
  assign n17374 = n15326 & ~n17373;
  assign n17375 = ~pi0862 & ~n15326;
  assign po1050 = n17374 | n17375;
  assign n17377 = ~pi0863 & ~n15312;
  assign n17378 = n15312 & ~n15700;
  assign n17379 = ~n17377 & ~n17378;
  assign n17380 = n15326 & ~n17379;
  assign n17381 = ~pi0863 & ~n15326;
  assign po1051 = n17380 | n17381;
  assign n17383 = ~pi0864 & ~n15312;
  assign n17384 = n15312 & ~n15562;
  assign n17385 = ~n17383 & ~n17384;
  assign n17386 = n15326 & ~n17385;
  assign n17387 = ~pi0864 & ~n15326;
  assign po1052 = n17386 | n17387;
  assign n17389 = ~pi0865 & ~n15312;
  assign n17390 = n15312 & ~n15571;
  assign n17391 = ~n17389 & ~n17390;
  assign n17392 = n15326 & ~n17391;
  assign n17393 = ~pi0865 & ~n15326;
  assign po1053 = n17392 | n17393;
  assign n17395 = ~pi0866 & ~n15312;
  assign n17396 = n15312 & ~n15580;
  assign n17397 = ~n17395 & ~n17396;
  assign n17398 = n15326 & ~n17397;
  assign n17399 = ~pi0866 & ~n15326;
  assign po1054 = n17398 | n17399;
  assign n17401 = ~pi0867 & ~n15312;
  assign n17402 = n15312 & ~n15589;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = n15326 & ~n17403;
  assign n17405 = ~pi0867 & ~n15326;
  assign po1055 = n17404 | n17405;
  assign n17407 = ~pi0868 & ~n15312;
  assign n17408 = n15312 & n15377;
  assign n17409 = ~n17407 & ~n17408;
  assign n17410 = n15326 & ~n17409;
  assign n17411 = ~pi0868 & ~n15326;
  assign po1056 = n17410 | n17411;
  assign n17413 = ~pi0869 & ~n15312;
  assign n17414 = n15312 & ~n15598;
  assign n17415 = ~n17413 & ~n17414;
  assign n17416 = n15326 & ~n17415;
  assign n17417 = ~pi0869 & ~n15326;
  assign po1057 = n17416 | n17417;
  assign n17419 = ~pi0870 & ~n15312;
  assign n17420 = n15312 & ~n15607;
  assign n17421 = ~n17419 & ~n17420;
  assign n17422 = n15326 & ~n17421;
  assign n17423 = ~pi0870 & ~n15326;
  assign po1058 = n17422 | n17423;
  assign n17425 = ~pi0871 & ~n15312;
  assign n17426 = n15312 & ~n15616;
  assign n17427 = ~n17425 & ~n17426;
  assign n17428 = n15326 & ~n17427;
  assign n17429 = ~pi0871 & ~n15326;
  assign po1059 = n17428 | n17429;
  assign n17431 = ~pi0872 & ~n15312;
  assign n17432 = n15312 & ~n15625;
  assign n17433 = ~n17431 & ~n17432;
  assign n17434 = n15326 & ~n17433;
  assign n17435 = ~pi0872 & ~n15326;
  assign po1060 = n17434 | n17435;
  assign n17437 = n15310 & n15334;
  assign n17438 = ~pi0873 & ~n17437;
  assign n17439 = ~n15442 & n17437;
  assign n17440 = ~n17438 & ~n17439;
  assign n17441 = n15326 & ~n17440;
  assign n17442 = ~pi0873 & ~n15326;
  assign po1061 = n17441 | n17442;
  assign n17444 = ~pi0874 & ~n17437;
  assign n17445 = ~n15451 & n17437;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = n15326 & ~n17446;
  assign n17448 = ~pi0874 & ~n15326;
  assign po1062 = n17447 | n17448;
  assign n17450 = ~pi0875 & ~n17437;
  assign n17451 = ~n15316 & n17437;
  assign n17452 = ~n17450 & ~n17451;
  assign n17453 = n15326 & ~n17452;
  assign n17454 = ~pi0875 & ~n15326;
  assign po1063 = n17453 | n17454;
  assign n17456 = ~pi0876 & ~n17437;
  assign n17457 = ~n15466 & n17437;
  assign n17458 = ~n17456 & ~n17457;
  assign n17459 = n15326 & ~n17458;
  assign n17460 = ~pi0876 & ~n15326;
  assign po1064 = n17459 | n17460;
  assign po1065 = ~n15362 & ~po0719;
  assign n17463 = ~pi0878 & ~n17437;
  assign n17464 = ~n15475 & n17437;
  assign n17465 = ~n17463 & ~n17464;
  assign n17466 = n15326 & ~n17465;
  assign n17467 = ~pi0878 & ~n15326;
  assign po1066 = n17466 | n17467;
  assign n17469 = ~pi0879 & ~n17437;
  assign n17470 = ~n15484 & n17437;
  assign n17471 = ~n17469 & ~n17470;
  assign n17472 = n15326 & ~n17471;
  assign n17473 = ~pi0879 & ~n15326;
  assign po1067 = n17472 | n17473;
  assign n17475 = ~pi0880 & ~n17437;
  assign n17476 = ~n15493 & n17437;
  assign n17477 = ~n17475 & ~n17476;
  assign n17478 = n15326 & ~n17477;
  assign n17479 = ~pi0880 & ~n15326;
  assign po1068 = n17478 | n17479;
  assign n17481 = ~pi0881 & ~n17437;
  assign n17482 = ~n15332 & n17437;
  assign n17483 = ~n17481 & ~n17482;
  assign n17484 = n15326 & ~n17483;
  assign n17485 = ~pi0881 & ~n15326;
  assign po1069 = n17484 | n17485;
  assign n17487 = ~pi0882 & ~n17437;
  assign n17488 = ~n15709 & n17437;
  assign n17489 = ~n17487 & ~n17488;
  assign n17490 = n15326 & ~n17489;
  assign n17491 = ~pi0882 & ~n15326;
  assign po1070 = n17490 | n17491;
  assign n17493 = ~pi0883 & ~n17437;
  assign n17494 = ~n15517 & n17437;
  assign n17495 = ~n17493 & ~n17494;
  assign n17496 = n15326 & ~n17495;
  assign n17497 = ~pi0883 & ~n15326;
  assign po1071 = n17496 | n17497;
  assign n17499 = ~pi0884 & ~n17437;
  assign n17500 = ~n15535 & n17437;
  assign n17501 = ~n17499 & ~n17500;
  assign n17502 = n15326 & ~n17501;
  assign n17503 = ~pi0884 & ~n15326;
  assign po1072 = n17502 | n17503;
  assign n17505 = ~pi0885 & ~n17437;
  assign n17506 = ~n15544 & n17437;
  assign n17507 = ~n17505 & ~n17506;
  assign n17508 = n15326 & ~n17507;
  assign n17509 = ~pi0885 & ~n15326;
  assign po1073 = n17508 | n17509;
  assign n17511 = ~pi0886 & ~n17437;
  assign n17512 = ~n15553 & n17437;
  assign n17513 = ~n17511 & ~n17512;
  assign n17514 = n15326 & ~n17513;
  assign n17515 = ~pi0886 & ~n15326;
  assign po1074 = n17514 | n17515;
  assign n17517 = ~pi0887 & ~n17437;
  assign n17518 = ~n15700 & n17437;
  assign n17519 = ~n17517 & ~n17518;
  assign n17520 = n15326 & ~n17519;
  assign n17521 = ~pi0887 & ~n15326;
  assign po1075 = n17520 | n17521;
  assign n17523 = ~pi0888 & ~n17437;
  assign n17524 = ~n15562 & n17437;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = n15326 & ~n17525;
  assign n17527 = ~pi0888 & ~n15326;
  assign po1076 = n17526 | n17527;
  assign n17529 = ~pi0889 & ~n17437;
  assign n17530 = ~n15580 & n17437;
  assign n17531 = ~n17529 & ~n17530;
  assign n17532 = n15326 & ~n17531;
  assign n17533 = ~pi0889 & ~n15326;
  assign po1077 = n17532 | n17533;
  assign n17535 = ~pi0890 & ~n17437;
  assign n17536 = ~n15589 & n17437;
  assign n17537 = ~n17535 & ~n17536;
  assign n17538 = n15326 & ~n17537;
  assign n17539 = ~pi0890 & ~n15326;
  assign po1078 = n17538 | n17539;
  assign n17541 = ~pi0891 & ~n17437;
  assign n17542 = n15377 & n17437;
  assign n17543 = ~n17541 & ~n17542;
  assign n17544 = n15326 & ~n17543;
  assign n17545 = ~pi0891 & ~n15326;
  assign po1079 = n17544 | n17545;
  assign n17547 = ~pi0892 & ~n17437;
  assign n17548 = ~n15598 & n17437;
  assign n17549 = ~n17547 & ~n17548;
  assign n17550 = n15326 & ~n17549;
  assign n17551 = ~pi0892 & ~n15326;
  assign po1080 = n17550 | n17551;
  assign n17553 = ~pi0893 & ~n17437;
  assign n17554 = ~n15607 & n17437;
  assign n17555 = ~n17553 & ~n17554;
  assign n17556 = n15326 & ~n17555;
  assign n17557 = ~pi0893 & ~n15326;
  assign po1081 = n17556 | n17557;
  assign n17559 = ~pi0894 & ~n17437;
  assign n17560 = ~n15616 & n17437;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = n15326 & ~n17561;
  assign n17563 = ~pi0894 & ~n15326;
  assign po1082 = n17562 | n17563;
  assign n17565 = ~pi0895 & ~n17437;
  assign n17566 = ~n15625 & n17437;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = n15326 & ~n17567;
  assign n17569 = ~pi0895 & ~n15326;
  assign po1083 = n17568 | n17569;
  assign n17571 = n15348 & n15352;
  assign po1084 = ~po0719 & ~n17571;
  assign n17573 = n15414 & ~n15451;
  assign n17574 = ~pi0897 & ~n15414;
  assign n17575 = ~n17573 & ~n17574;
  assign n17576 = n15326 & ~n17575;
  assign n17577 = ~pi0897 & ~n15326;
  assign po1085 = n17576 | n17577;
  assign n17579 = ~pi0898 & ~n17154;
  assign n17580 = ~n15332 & n17154;
  assign n17581 = ~n17579 & ~n17580;
  assign n17582 = n15326 & ~n17581;
  assign n17583 = ~pi0898 & ~n15326;
  assign po1086 = n17582 | n17583;
  assign n17585 = ~n15316 & n15335;
  assign n17586 = ~pi0899 & ~n15335;
  assign n17587 = ~n17585 & ~n17586;
  assign n17588 = n15326 & ~n17587;
  assign n17589 = ~pi0899 & ~n15326;
  assign po1087 = n17588 | n17589;
  assign n17591 = n15414 & ~n15571;
  assign n17592 = ~pi0900 & ~n15414;
  assign n17593 = ~n17591 & ~n17592;
  assign n17594 = n15326 & ~n17593;
  assign n17595 = ~pi0900 & ~n15326;
  assign po1088 = n17594 | n17595;
  assign n17597 = n15414 & ~n15526;
  assign n17598 = ~pi0901 & ~n15414;
  assign n17599 = ~n17597 & ~n17598;
  assign n17600 = n15326 & ~n17599;
  assign n17601 = ~pi0901 & ~n15326;
  assign po1089 = n17600 | n17601;
  assign n17603 = ~pi0902 & ~n17015;
  assign n17604 = ~n15332 & n17015;
  assign n17605 = ~n17603 & ~n17604;
  assign n17606 = n15326 & ~n17605;
  assign n17607 = ~pi0902 & ~n15326;
  assign po1090 = n17606 | n17607;
  assign n17609 = ~pi0903 & ~n17015;
  assign n17610 = ~n15316 & n17015;
  assign n17611 = ~n17609 & ~n17610;
  assign n17612 = n15326 & ~n17611;
  assign n17613 = ~pi0903 & ~n15326;
  assign po1091 = n17612 | n17613;
  assign n17615 = n15393 & ~n15562;
  assign n17616 = ~pi0904 & ~n15393;
  assign n17617 = ~n17615 & ~n17616;
  assign n17618 = n15326 & ~n17617;
  assign n17619 = ~pi0904 & ~n15326;
  assign po1092 = n17618 | n17619;
  assign n17621 = n15393 & ~n15571;
  assign n17622 = ~pi0905 & ~n15393;
  assign n17623 = ~n17621 & ~n17622;
  assign n17624 = n15326 & ~n17623;
  assign n17625 = ~pi0905 & ~n15326;
  assign po1093 = n17624 | n17625;
  assign n17627 = n15393 & ~n15526;
  assign n17628 = ~pi0906 & ~n15393;
  assign n17629 = ~n17627 & ~n17628;
  assign n17630 = n15326 & ~n17629;
  assign n17631 = ~pi0906 & ~n15326;
  assign po1094 = n17630 | n17631;
  assign n17633 = n15393 & ~n15493;
  assign n17634 = ~pi0907 & ~n15393;
  assign n17635 = ~n17633 & ~n17634;
  assign n17636 = n15326 & ~n17635;
  assign n17637 = ~pi0907 & ~n15326;
  assign po1095 = n17636 | n17637;
  assign n17639 = ~pi0908 & ~n16870;
  assign n17640 = ~n15332 & n16870;
  assign n17641 = ~n17639 & ~n17640;
  assign n17642 = n15326 & ~n17641;
  assign n17643 = ~pi0908 & ~n15326;
  assign po1096 = n17642 | n17643;
  assign n17645 = n15393 & ~n15442;
  assign n17646 = ~pi0909 & ~n15393;
  assign n17647 = ~n17645 & ~n17646;
  assign n17648 = n15326 & ~n17647;
  assign n17649 = ~pi0909 & ~n15326;
  assign po1097 = n17648 | n17649;
  assign n17651 = n15434 & ~n15571;
  assign n17652 = ~pi0910 & ~n15434;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = n15326 & ~n17653;
  assign n17655 = ~pi0910 & ~n15326;
  assign po1098 = n17654 | n17655;
  assign n17657 = n15434 & ~n15598;
  assign n17658 = ~pi0911 & ~n15434;
  assign n17659 = ~n17657 & ~n17658;
  assign n17660 = n15326 & ~n17659;
  assign n17661 = ~pi0911 & ~n15326;
  assign po1099 = n17660 | n17661;
  assign n17663 = ~n15562 & n16136;
  assign n17664 = ~pi0912 & ~n16136;
  assign n17665 = ~n17663 & ~n17664;
  assign n17666 = n15326 & ~n17665;
  assign n17667 = ~pi0912 & ~n15326;
  assign po1100 = n17666 | n17667;
  assign n17669 = n15386 & ~n15700;
  assign n17670 = ~pi0913 & ~n15386;
  assign n17671 = ~n17669 & ~n17670;
  assign n17672 = n15326 & ~n17671;
  assign n17673 = ~pi0913 & ~n15326;
  assign po1101 = n17672 | n17673;
  assign n17675 = n15434 & ~n15451;
  assign n17676 = ~pi0914 & ~n15434;
  assign n17677 = ~n17675 & ~n17676;
  assign n17678 = n15326 & ~n17677;
  assign n17679 = ~pi0914 & ~n15326;
  assign po1102 = n17678 | n17679;
  assign n17681 = n15434 & ~n15502;
  assign n17682 = ~pi0915 & ~n15434;
  assign n17683 = ~n17681 & ~n17682;
  assign n17684 = n15326 & ~n17683;
  assign n17685 = ~pi0915 & ~n15326;
  assign po1103 = n17684 | n17685;
  assign n17687 = n15386 & ~n15709;
  assign n17688 = ~pi0916 & ~n15386;
  assign n17689 = ~n17687 & ~n17688;
  assign n17690 = n15326 & ~n17689;
  assign n17691 = ~pi0916 & ~n15326;
  assign po1104 = n17690 | n17691;
  assign n17693 = ~n15598 & n16635;
  assign n17694 = ~pi0917 & ~n16635;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = n15326 & ~n17695;
  assign n17697 = ~pi0917 & ~n15326;
  assign po1105 = n17696 | n17697;
  assign n17699 = ~n15526 & n16635;
  assign n17700 = ~pi0918 & ~n16635;
  assign n17701 = ~n17699 & ~n17700;
  assign n17702 = n15326 & ~n17701;
  assign n17703 = ~pi0918 & ~n15326;
  assign po1106 = n17702 | n17703;
  assign n17705 = ~n15571 & n16635;
  assign n17706 = ~pi0919 & ~n16635;
  assign n17707 = ~n17705 & ~n17706;
  assign n17708 = n15326 & ~n17707;
  assign n17709 = ~pi0919 & ~n15326;
  assign po1107 = n17708 | n17709;
  assign n17711 = ~pi0920 & ~n15326;
  assign n17712 = n15377 & n16136;
  assign n17713 = ~pi0920 & ~n16136;
  assign n17714 = ~n17712 & ~n17713;
  assign n17715 = n15326 & ~n17714;
  assign po1108 = n17711 | n17715;
  assign n17717 = ~n15502 & n16635;
  assign n17718 = ~pi0921 & ~n16635;
  assign n17719 = ~n17717 & ~n17718;
  assign n17720 = n15326 & ~n17719;
  assign n17721 = ~pi0921 & ~n15326;
  assign po1109 = n17720 | n17721;
  assign n17723 = n15407 & ~n15451;
  assign n17724 = ~pi0922 & ~n15407;
  assign n17725 = ~n17723 & ~n17724;
  assign n17726 = n15326 & ~n17725;
  assign n17727 = ~pi0922 & ~n15326;
  assign po1110 = n17726 | n17727;
  assign n17729 = ~pi0923 & ~n15326;
  assign n17730 = n15377 & n16635;
  assign n17731 = ~pi0923 & ~n16635;
  assign n17732 = ~n17730 & ~n17731;
  assign n17733 = n15326 & ~n17732;
  assign po1111 = n17729 | n17733;
  assign n17735 = ~n15451 & n16635;
  assign n17736 = ~pi0924 & ~n16635;
  assign n17737 = ~n17735 & ~n17736;
  assign n17738 = n15326 & ~n17737;
  assign n17739 = ~pi0924 & ~n15326;
  assign po1112 = n17738 | n17739;
  assign n17741 = ~n15332 & n15407;
  assign n17742 = ~pi0925 & ~n15407;
  assign n17743 = ~n17741 & ~n17742;
  assign n17744 = n15326 & ~n17743;
  assign n17745 = ~pi0925 & ~n15326;
  assign po1113 = n17744 | n17745;
  assign n17747 = n15374 & ~n15571;
  assign n17748 = ~pi0926 & ~n15374;
  assign n17749 = ~n17747 & ~n17748;
  assign n17750 = n15326 & ~n17749;
  assign n17751 = ~pi0926 & ~n15326;
  assign po1114 = n17750 | n17751;
  assign n17753 = n15400 & ~n15598;
  assign n17754 = ~pi0927 & ~n15400;
  assign n17755 = ~n17753 & ~n17754;
  assign n17756 = n15326 & ~n17755;
  assign n17757 = ~pi0927 & ~n15326;
  assign po1115 = n17756 | n17757;
  assign n17759 = n15400 & ~n15571;
  assign n17760 = ~pi0929 & ~n15400;
  assign n17761 = ~n17759 & ~n17760;
  assign n17762 = n15326 & ~n17761;
  assign n17763 = ~pi0929 & ~n15326;
  assign po1116 = n17762 | n17763;
  assign n17765 = n15400 & ~n15502;
  assign n17766 = ~pi0932 & ~n15400;
  assign n17767 = ~n17765 & ~n17766;
  assign n17768 = n15326 & ~n17767;
  assign n17769 = ~pi0932 & ~n15326;
  assign po1117 = n17768 | n17769;
  assign n17771 = n15400 & ~n15451;
  assign n17772 = ~pi0936 & ~n15400;
  assign n17773 = ~n17771 & ~n17772;
  assign n17774 = n15326 & ~n17773;
  assign n17775 = ~pi0936 & ~n15326;
  assign po1118 = n17774 | n17775;
  assign n17777 = n15374 & ~n15598;
  assign n17778 = ~pi0937 & ~n15374;
  assign n17779 = ~n17777 & ~n17778;
  assign n17780 = n15326 & ~n17779;
  assign n17781 = ~pi0937 & ~n15326;
  assign po1119 = n17780 | n17781;
  assign n17783 = n15374 & ~n15502;
  assign n17784 = ~pi0940 & ~n15374;
  assign n17785 = ~n17783 & ~n17784;
  assign n17786 = n15326 & ~n17785;
  assign n17787 = ~pi0940 & ~n15326;
  assign po1120 = n17786 | n17787;
  assign n17789 = n15374 & ~n15451;
  assign n17790 = ~pi0941 & ~n15374;
  assign n17791 = ~n17789 & ~n17790;
  assign n17792 = n15326 & ~n17791;
  assign n17793 = ~pi0941 & ~n15326;
  assign po1121 = n17792 | n17793;
  assign n17795 = ~n15517 & n16136;
  assign n17796 = ~pi0942 & ~n16136;
  assign n17797 = ~n17795 & ~n17796;
  assign n17798 = n15326 & ~n17797;
  assign n17799 = ~pi0942 & ~n15326;
  assign po1122 = n17798 | n17799;
  assign n17801 = ~n15442 & n16136;
  assign n17802 = ~pi0943 & ~n16136;
  assign n17803 = ~n17801 & ~n17802;
  assign n17804 = n15326 & ~n17803;
  assign n17805 = ~pi0943 & ~n15326;
  assign po1123 = n17804 | n17805;
  assign n17807 = n15427 & ~n15709;
  assign n17808 = ~pi0944 & ~n15427;
  assign n17809 = ~n17807 & ~n17808;
  assign n17810 = n15326 & ~n17809;
  assign n17811 = ~pi0944 & ~n15326;
  assign po1124 = n17810 | n17811;
  assign n17813 = n15427 & ~n15484;
  assign n17814 = ~pi0945 & ~n15427;
  assign n17815 = ~n17813 & ~n17814;
  assign n17816 = n15326 & ~n17815;
  assign n17817 = ~pi0945 & ~n15326;
  assign po1125 = n17816 | n17817;
  assign n17819 = n15335 & ~n15625;
  assign n17820 = ~pi0946 & ~n15335;
  assign n17821 = ~n17819 & ~n17820;
  assign n17822 = n15326 & ~n17821;
  assign n17823 = ~pi0946 & ~n15326;
  assign po1126 = n17822 | n17823;
  assign n17825 = ~pi0947 & ~n17437;
  assign n17826 = ~n15571 & n17437;
  assign n17827 = ~n17825 & ~n17826;
  assign n17828 = n15326 & ~n17827;
  assign n17829 = ~pi0947 & ~n15326;
  assign po1127 = n17828 | n17829;
  assign n17831 = ~pi0948 & ~n17437;
  assign n17832 = ~n15526 & n17437;
  assign n17833 = ~n17831 & ~n17832;
  assign n17834 = n15326 & ~n17833;
  assign n17835 = ~pi0948 & ~n15326;
  assign po1128 = n17834 | n17835;
  assign n17837 = ~pi0949 & ~n17437;
  assign n17838 = ~n15502 & n17437;
  assign n17839 = ~n17837 & ~n17838;
  assign n17840 = n15326 & ~n17839;
  assign n17841 = ~pi0949 & ~n15326;
  assign po1129 = n17840 | n17841;
  assign n17843 = ~pi0950 & ~n15312;
  assign n17844 = pi1345 & ~n15376;
  assign n17845 = ~pi1290 & n17844;
  assign n17846 = n15312 & ~n17845;
  assign n17847 = ~n17843 & ~n17846;
  assign n17848 = n15326 & ~n17847;
  assign n17849 = ~pi0950 & ~n15326;
  assign po1130 = n17848 | n17849;
  assign n17851 = ~pi1289 & n17844;
  assign n17852 = n15386 & ~n17851;
  assign n17853 = ~pi0951 & ~n15386;
  assign n17854 = ~n17852 & ~n17853;
  assign n17855 = n15326 & ~n17854;
  assign n17856 = ~pi0951 & ~n15326;
  assign po1131 = n17855 | n17856;
  assign n17858 = n15386 & ~n17845;
  assign n17859 = ~pi0952 & ~n15386;
  assign n17860 = ~n17858 & ~n17859;
  assign n17861 = n15326 & ~n17860;
  assign n17862 = ~pi0952 & ~n15326;
  assign po1132 = n17861 | n17862;
  assign n17864 = n15393 & ~n17845;
  assign n17865 = ~pi0953 & ~n15393;
  assign n17866 = ~n17864 & ~n17865;
  assign n17867 = n15326 & ~n17866;
  assign n17868 = ~pi0953 & ~n15326;
  assign po1133 = n17867 | n17868;
  assign n17870 = n15393 & ~n17851;
  assign n17871 = ~pi0954 & ~n15393;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = n15326 & ~n17872;
  assign n17874 = ~pi0954 & ~n15326;
  assign po1134 = n17873 | n17874;
  assign n17876 = n15414 & ~n17851;
  assign n17877 = ~pi0955 & ~n15414;
  assign n17878 = ~n17876 & ~n17877;
  assign n17879 = n15326 & ~n17878;
  assign n17880 = ~pi0955 & ~n15326;
  assign po1135 = n17879 | n17880;
  assign n17882 = n15414 & ~n17845;
  assign n17883 = ~pi0956 & ~n15414;
  assign n17884 = ~n17882 & ~n17883;
  assign n17885 = n15326 & ~n17884;
  assign n17886 = ~pi0956 & ~n15326;
  assign po1136 = n17885 | n17886;
  assign n17888 = n15335 & ~n17851;
  assign n17889 = ~pi0957 & ~n15335;
  assign n17890 = ~n17888 & ~n17889;
  assign n17891 = n15326 & ~n17890;
  assign n17892 = ~pi0957 & ~n15326;
  assign po1137 = n17891 | n17892;
  assign n17894 = n15427 & ~n17851;
  assign n17895 = ~pi0958 & ~n15427;
  assign n17896 = ~n17894 & ~n17895;
  assign n17897 = n15326 & ~n17896;
  assign n17898 = ~pi0958 & ~n15326;
  assign po1138 = n17897 | n17898;
  assign n17900 = n15427 & ~n17845;
  assign n17901 = ~pi0959 & ~n15427;
  assign n17902 = ~n17900 & ~n17901;
  assign n17903 = n15326 & ~n17902;
  assign n17904 = ~pi0959 & ~n15326;
  assign po1139 = n17903 | n17904;
  assign n17906 = n16136 & ~n17845;
  assign n17907 = ~pi0960 & ~n16136;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = n15326 & ~n17908;
  assign n17910 = ~pi0960 & ~n15326;
  assign po1140 = n17909 | n17910;
  assign n17912 = n16136 & ~n17851;
  assign n17913 = ~pi0961 & ~n16136;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = n15326 & ~n17914;
  assign n17916 = ~pi0961 & ~n15326;
  assign po1141 = n17915 | n17916;
  assign n17918 = n15374 & ~n17851;
  assign n17919 = ~pi0962 & ~n15374;
  assign n17920 = ~n17918 & ~n17919;
  assign n17921 = n15326 & ~n17920;
  assign n17922 = ~pi0962 & ~n15326;
  assign po1142 = n17921 | n17922;
  assign n17924 = ~pi0963 & ~n16870;
  assign n17925 = n16870 & ~n17851;
  assign n17926 = ~n17924 & ~n17925;
  assign n17927 = n15326 & ~n17926;
  assign n17928 = ~pi0963 & ~n15326;
  assign po1143 = n17927 | n17928;
  assign n17930 = ~pi0964 & ~n17015;
  assign n17931 = n17015 & ~n17851;
  assign n17932 = ~n17930 & ~n17931;
  assign n17933 = n15326 & ~n17932;
  assign n17934 = ~pi0964 & ~n15326;
  assign po1144 = n17933 | n17934;
  assign n17936 = ~pi0965 & ~n17154;
  assign n17937 = n17154 & ~n17851;
  assign n17938 = ~n17936 & ~n17937;
  assign n17939 = n15326 & ~n17938;
  assign n17940 = ~pi0965 & ~n15326;
  assign po1145 = n17939 | n17940;
  assign n17942 = ~pi0966 & ~n15312;
  assign n17943 = n15312 & ~n17851;
  assign n17944 = ~n17942 & ~n17943;
  assign n17945 = n15326 & ~n17944;
  assign n17946 = ~pi0966 & ~n15326;
  assign po1146 = n17945 | n17946;
  assign n17948 = n15400 & ~n17851;
  assign n17949 = ~pi0967 & ~n15400;
  assign n17950 = ~n17948 & ~n17949;
  assign n17951 = n15326 & ~n17950;
  assign n17952 = ~pi0967 & ~n15326;
  assign po1147 = n17951 | n17952;
  assign n17954 = n15400 & ~n17845;
  assign n17955 = ~pi0968 & ~n15400;
  assign n17956 = ~n17954 & ~n17955;
  assign n17957 = n15326 & ~n17956;
  assign n17958 = ~pi0968 & ~n15326;
  assign po1148 = n17957 | n17958;
  assign n17960 = n15407 & ~n17851;
  assign n17961 = ~pi0969 & ~n15407;
  assign n17962 = ~n17960 & ~n17961;
  assign n17963 = n15326 & ~n17962;
  assign n17964 = ~pi0969 & ~n15326;
  assign po1149 = n17963 | n17964;
  assign n17966 = n15407 & ~n17845;
  assign n17967 = ~pi0970 & ~n15407;
  assign n17968 = ~n17966 & ~n17967;
  assign n17969 = n15326 & ~n17968;
  assign n17970 = ~pi0970 & ~n15326;
  assign po1150 = n17969 | n17970;
  assign n17972 = n16635 & ~n17851;
  assign n17973 = ~pi0971 & ~n16635;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = n15326 & ~n17974;
  assign n17976 = ~pi0971 & ~n15326;
  assign po1151 = n17975 | n17976;
  assign n17978 = n16635 & ~n17845;
  assign n17979 = ~pi0972 & ~n16635;
  assign n17980 = ~n17978 & ~n17979;
  assign n17981 = n15326 & ~n17980;
  assign n17982 = ~pi0972 & ~n15326;
  assign po1152 = n17981 | n17982;
  assign n17984 = ~pi0973 & ~n17437;
  assign n17985 = n17437 & ~n17851;
  assign n17986 = ~n17984 & ~n17985;
  assign n17987 = n15326 & ~n17986;
  assign n17988 = ~pi0973 & ~n15326;
  assign po1153 = n17987 | n17988;
  assign n17990 = n15434 & ~n17851;
  assign n17991 = ~pi0974 & ~n15434;
  assign n17992 = ~n17990 & ~n17991;
  assign n17993 = n15326 & ~n17992;
  assign n17994 = ~pi0974 & ~n15326;
  assign po1154 = n17993 | n17994;
  assign n17996 = n7066 & n7078;
  assign n17997 = ~pi1686 & n7124;
  assign po3086 = n7101 & ~n7117;
  assign n17999 = pi1687 & ~n7109;
  assign n18000 = ~po3086 & ~n17999;
  assign n18001 = ~n17997 & n18000;
  assign n18002 = ~n17996 & n18001;
  assign n18003 = ~n7121 & n18002;
  assign n18004 = ~n7063 & n18003;
  assign po1155 = ~n7166 & n18004;
  assign n18006 = ~pi0976 & ~n17154;
  assign n18007 = n17154 & ~n17845;
  assign n18008 = ~n18006 & ~n18007;
  assign n18009 = n15326 & ~n18008;
  assign n18010 = ~pi0976 & ~n15326;
  assign po1156 = n18009 | n18010;
  assign n18012 = ~pi0977 & ~n17015;
  assign n18013 = n17015 & ~n17845;
  assign n18014 = ~n18012 & ~n18013;
  assign n18015 = n15326 & ~n18014;
  assign n18016 = ~pi0977 & ~n15326;
  assign po1157 = n18015 | n18016;
  assign n18018 = ~pi0978 & ~n16870;
  assign n18019 = n16870 & ~n17845;
  assign n18020 = ~n18018 & ~n18019;
  assign n18021 = n15326 & ~n18020;
  assign n18022 = ~pi0978 & ~n15326;
  assign po1158 = n18021 | n18022;
  assign n18024 = n15374 & ~n17845;
  assign n18025 = ~pi0979 & ~n15374;
  assign n18026 = ~n18024 & ~n18025;
  assign n18027 = n15326 & ~n18026;
  assign n18028 = ~pi0979 & ~n15326;
  assign po1159 = n18027 | n18028;
  assign n18030 = n15434 & ~n17845;
  assign n18031 = ~pi0980 & ~n15434;
  assign n18032 = ~n18030 & ~n18031;
  assign n18033 = n15326 & ~n18032;
  assign n18034 = ~pi0980 & ~n15326;
  assign po1160 = n18033 | n18034;
  assign n18036 = ~pi0981 & ~n17437;
  assign n18037 = n17437 & ~n17845;
  assign n18038 = ~n18036 & ~n18037;
  assign n18039 = n15326 & ~n18038;
  assign n18040 = ~pi0981 & ~n15326;
  assign po1161 = n18039 | n18040;
  assign n18042 = n15335 & ~n17845;
  assign n18043 = ~pi0982 & ~n15335;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = n15326 & ~n18044;
  assign n18046 = ~pi0982 & ~n15326;
  assign po1162 = n18045 | n18046;
  assign n18048 = ~pi1291 & pi1345;
  assign n18049 = ~n15376 & ~n18048;
  assign n18050 = n15400 & n18049;
  assign n18051 = ~pi0983 & ~n15400;
  assign n18052 = ~n18050 & ~n18051;
  assign n18053 = n15326 & ~n18052;
  assign n18054 = ~pi0983 & ~n15326;
  assign po1163 = n18053 | n18054;
  assign n18056 = ~pi0984 & ~n15312;
  assign n18057 = pi0504 & ~pi1345;
  assign n18058 = ~pi1293 & pi1345;
  assign n18059 = ~n18057 & ~n18058;
  assign n18060 = n15312 & ~n18059;
  assign n18061 = ~n18056 & ~n18060;
  assign n18062 = n15326 & ~n18061;
  assign n18063 = ~pi0984 & ~n15326;
  assign po1164 = n18062 | n18063;
  assign n18065 = ~pi0985 & ~n15312;
  assign n18066 = pi0514 & ~pi1345;
  assign n18067 = ~pi1320 & pi1345;
  assign n18068 = ~n18066 & ~n18067;
  assign n18069 = n15312 & ~n18068;
  assign n18070 = ~n18065 & ~n18069;
  assign n18071 = n15326 & ~n18070;
  assign n18072 = ~pi0985 & ~n15326;
  assign po1165 = n18071 | n18072;
  assign n18074 = ~pi0986 & ~n15312;
  assign n18075 = pi0515 & ~pi1345;
  assign n18076 = ~pi1287 & pi1345;
  assign n18077 = ~n18075 & ~n18076;
  assign n18078 = n15312 & ~n18077;
  assign n18079 = ~n18074 & ~n18078;
  assign n18080 = n15326 & ~n18079;
  assign n18081 = ~pi0986 & ~n15326;
  assign po1166 = n18080 | n18081;
  assign n18083 = ~pi0987 & ~n15312;
  assign n18084 = pi0497 & ~pi1345;
  assign n18085 = ~pi1283 & pi1345;
  assign n18086 = ~n18084 & ~n18085;
  assign n18087 = n15312 & ~n18086;
  assign n18088 = ~n18083 & ~n18087;
  assign n18089 = n15326 & ~n18088;
  assign n18090 = ~pi0987 & ~n15326;
  assign po1167 = n18089 | n18090;
  assign n18092 = pi0988 & ~pi3362;
  assign po1168 = ~n11017 | n18092;
  assign n18094 = ~pi0989 & ~n15312;
  assign n18095 = pi0488 & ~pi1345;
  assign n18096 = ~pi1276 & pi1345;
  assign n18097 = ~n18095 & ~n18096;
  assign n18098 = n15312 & ~n18097;
  assign n18099 = ~n18094 & ~n18098;
  assign n18100 = n15326 & ~n18099;
  assign n18101 = ~pi0989 & ~n15326;
  assign po1169 = n18100 | n18101;
  assign n18103 = pi0510 & ~pi1345;
  assign n18104 = ~pi1323 & pi1345;
  assign n18105 = ~n18103 & ~n18104;
  assign n18106 = n15386 & ~n18105;
  assign n18107 = ~pi0990 & ~n15386;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = n15326 & ~n18108;
  assign n18110 = ~pi0990 & ~n15326;
  assign po1170 = n18109 | n18110;
  assign n18112 = n15386 & ~n18086;
  assign n18113 = ~pi0991 & ~n15386;
  assign n18114 = ~n18112 & ~n18113;
  assign n18115 = n15326 & ~n18114;
  assign n18116 = ~pi0991 & ~n15326;
  assign po1171 = n18115 | n18116;
  assign n18118 = n15386 & ~n18068;
  assign n18119 = ~pi0992 & ~n15386;
  assign n18120 = ~n18118 & ~n18119;
  assign n18121 = n15326 & ~n18120;
  assign n18122 = ~pi0992 & ~n15326;
  assign po1172 = n18121 | n18122;
  assign n18124 = n15386 & ~n18059;
  assign n18125 = ~pi0993 & ~n15386;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = n15326 & ~n18126;
  assign n18128 = ~pi0993 & ~n15326;
  assign po1173 = n18127 | n18128;
  assign n18130 = n15393 & ~n18097;
  assign n18131 = ~pi0994 & ~n15393;
  assign n18132 = ~n18130 & ~n18131;
  assign n18133 = n15326 & ~n18132;
  assign n18134 = ~pi0994 & ~n15326;
  assign po1174 = n18133 | n18134;
  assign n18136 = n15393 & ~n18105;
  assign n18137 = ~pi0995 & ~n15393;
  assign n18138 = ~n18136 & ~n18137;
  assign n18139 = n15326 & ~n18138;
  assign n18140 = ~pi0995 & ~n15326;
  assign po1175 = n18139 | n18140;
  assign n18142 = n15393 & ~n18077;
  assign n18143 = ~pi0996 & ~n15393;
  assign n18144 = ~n18142 & ~n18143;
  assign n18145 = n15326 & ~n18144;
  assign n18146 = ~pi0996 & ~n15326;
  assign po1176 = n18145 | n18146;
  assign n18148 = n15393 & ~n18059;
  assign n18149 = ~pi0997 & ~n15393;
  assign n18150 = ~n18148 & ~n18149;
  assign n18151 = n15326 & ~n18150;
  assign n18152 = ~pi0997 & ~n15326;
  assign po1177 = n18151 | n18152;
  assign n18154 = n15393 & ~n18068;
  assign n18155 = ~pi0998 & ~n15393;
  assign n18156 = ~n18154 & ~n18155;
  assign n18157 = n15326 & ~n18156;
  assign n18158 = ~pi0998 & ~n15326;
  assign po1178 = n18157 | n18158;
  assign n18160 = pi0499 & ~pi1345;
  assign n18161 = ~pi1328 & pi1345;
  assign n18162 = ~n18160 & ~n18161;
  assign n18163 = n15414 & ~n18162;
  assign n18164 = ~pi0999 & ~n15414;
  assign n18165 = ~n18163 & ~n18164;
  assign n18166 = n15326 & ~n18165;
  assign n18167 = ~pi0999 & ~n15326;
  assign po1179 = n18166 | n18167;
  assign n18169 = n15414 & ~n18105;
  assign n18170 = ~pi1000 & ~n15414;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = n15326 & ~n18171;
  assign n18173 = ~pi1000 & ~n15326;
  assign po1180 = n18172 | n18173;
  assign n18175 = n15414 & ~n18077;
  assign n18176 = ~pi1001 & ~n15414;
  assign n18177 = ~n18175 & ~n18176;
  assign n18178 = n15326 & ~n18177;
  assign n18179 = ~pi1001 & ~n15326;
  assign po1181 = n18178 | n18179;
  assign n18181 = n15414 & n18049;
  assign n18182 = ~pi1002 & ~n15414;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = n15326 & ~n18183;
  assign n18185 = ~pi1002 & ~n15326;
  assign po1182 = n18184 | n18185;
  assign n18187 = n15414 & ~n18059;
  assign n18188 = ~pi1003 & ~n15414;
  assign n18189 = ~n18187 & ~n18188;
  assign n18190 = n15326 & ~n18189;
  assign n18191 = ~pi1003 & ~n15326;
  assign po1183 = n18190 | n18191;
  assign n18193 = n15335 & ~n18162;
  assign n18194 = ~pi1004 & ~n15335;
  assign n18195 = ~n18193 & ~n18194;
  assign n18196 = n15326 & ~n18195;
  assign n18197 = ~pi1004 & ~n15326;
  assign po1184 = n18196 | n18197;
  assign n18199 = n15335 & n18049;
  assign n18200 = ~pi1005 & ~n15335;
  assign n18201 = ~n18199 & ~n18200;
  assign n18202 = n15326 & ~n18201;
  assign n18203 = ~pi1005 & ~n15326;
  assign po1185 = n18202 | n18203;
  assign n18205 = n15335 & ~n18068;
  assign n18206 = ~pi1006 & ~n15335;
  assign n18207 = ~n18205 & ~n18206;
  assign n18208 = n15326 & ~n18207;
  assign n18209 = ~pi1006 & ~n15326;
  assign po1186 = n18208 | n18209;
  assign n18211 = pi0505 & ~pi1345;
  assign n18212 = ~pi1308 & pi1345;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = n15335 & ~n18213;
  assign n18215 = ~pi1007 & ~n15335;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = n15326 & ~n18216;
  assign n18218 = ~pi1007 & ~n15326;
  assign po1187 = n18217 | n18218;
  assign n18220 = n15427 & ~n18162;
  assign n18221 = ~pi1008 & ~n15427;
  assign n18222 = ~n18220 & ~n18221;
  assign n18223 = n15326 & ~n18222;
  assign n18224 = ~pi1008 & ~n15326;
  assign po1188 = n18223 | n18224;
  assign n18226 = n15427 & ~n18097;
  assign n18227 = ~pi1009 & ~n15427;
  assign n18228 = ~n18226 & ~n18227;
  assign n18229 = n15326 & ~n18228;
  assign n18230 = ~pi1009 & ~n15326;
  assign po1189 = n18229 | n18230;
  assign n18232 = n15427 & ~n18068;
  assign n18233 = ~pi1010 & ~n15427;
  assign n18234 = ~n18232 & ~n18233;
  assign n18235 = n15326 & ~n18234;
  assign n18236 = ~pi1010 & ~n15326;
  assign po1190 = n18235 | n18236;
  assign n18238 = n15427 & ~n18059;
  assign n18239 = ~pi1011 & ~n15427;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = n15326 & ~n18240;
  assign n18242 = ~pi1011 & ~n15326;
  assign po1191 = n18241 | n18242;
  assign n18244 = n16136 & ~n18105;
  assign n18245 = ~pi1012 & ~n16136;
  assign n18246 = ~n18244 & ~n18245;
  assign n18247 = n15326 & ~n18246;
  assign n18248 = ~pi1012 & ~n15326;
  assign po1192 = n18247 | n18248;
  assign n18250 = n16136 & ~n18086;
  assign n18251 = ~pi1013 & ~n16136;
  assign n18252 = ~n18250 & ~n18251;
  assign n18253 = n15326 & ~n18252;
  assign n18254 = ~pi1013 & ~n15326;
  assign po1193 = n18253 | n18254;
  assign n18256 = n16136 & ~n18068;
  assign n18257 = ~pi1014 & ~n16136;
  assign n18258 = ~n18256 & ~n18257;
  assign n18259 = n15326 & ~n18258;
  assign n18260 = ~pi1014 & ~n15326;
  assign po1194 = n18259 | n18260;
  assign n18262 = n16136 & ~n18059;
  assign n18263 = ~pi1015 & ~n16136;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = n15326 & ~n18264;
  assign n18266 = ~pi1015 & ~n15326;
  assign po1195 = n18265 | n18266;
  assign n18268 = n15374 & ~n18162;
  assign n18269 = ~pi1016 & ~n15374;
  assign n18270 = ~n18268 & ~n18269;
  assign n18271 = n15326 & ~n18270;
  assign n18272 = ~pi1016 & ~n15326;
  assign po1196 = n18271 | n18272;
  assign n18274 = n15374 & ~n18097;
  assign n18275 = ~pi1017 & ~n15374;
  assign n18276 = ~n18274 & ~n18275;
  assign n18277 = n15326 & ~n18276;
  assign n18278 = ~pi1017 & ~n15326;
  assign po1197 = n18277 | n18278;
  assign n18280 = n15374 & ~n18105;
  assign n18281 = ~pi1018 & ~n15374;
  assign n18282 = ~n18280 & ~n18281;
  assign n18283 = n15326 & ~n18282;
  assign n18284 = ~pi1018 & ~n15326;
  assign po1198 = n18283 | n18284;
  assign n18286 = n15374 & ~n18077;
  assign n18287 = ~pi1019 & ~n15374;
  assign n18288 = ~n18286 & ~n18287;
  assign n18289 = n15326 & ~n18288;
  assign n18290 = ~pi1019 & ~n15326;
  assign po1199 = n18289 | n18290;
  assign n18292 = n15374 & ~n18068;
  assign n18293 = ~pi1020 & ~n15374;
  assign n18294 = ~n18292 & ~n18293;
  assign n18295 = n15326 & ~n18294;
  assign n18296 = ~pi1020 & ~n15326;
  assign po1200 = n18295 | n18296;
  assign n18298 = n15374 & ~n18213;
  assign n18299 = ~pi1021 & ~n15374;
  assign n18300 = ~n18298 & ~n18299;
  assign n18301 = n15326 & ~n18300;
  assign n18302 = ~pi1021 & ~n15326;
  assign po1201 = n18301 | n18302;
  assign n18304 = n15374 & ~n18059;
  assign n18305 = ~pi1022 & ~n15374;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = n15326 & ~n18306;
  assign n18308 = ~pi1022 & ~n15326;
  assign po1202 = n18307 | n18308;
  assign n18310 = n15400 & ~n18162;
  assign n18311 = ~pi1023 & ~n15400;
  assign n18312 = ~n18310 & ~n18311;
  assign n18313 = n15326 & ~n18312;
  assign n18314 = ~pi1023 & ~n15326;
  assign po1203 = n18313 | n18314;
  assign n18316 = n15400 & ~n18105;
  assign n18317 = ~pi1024 & ~n15400;
  assign n18318 = ~n18316 & ~n18317;
  assign n18319 = n15326 & ~n18318;
  assign n18320 = ~pi1024 & ~n15326;
  assign po1204 = n18319 | n18320;
  assign n18322 = n15400 & ~n18077;
  assign n18323 = ~pi1025 & ~n15400;
  assign n18324 = ~n18322 & ~n18323;
  assign n18325 = n15326 & ~n18324;
  assign n18326 = ~pi1025 & ~n15326;
  assign po1205 = n18325 | n18326;
  assign n18328 = n15400 & ~n18068;
  assign n18329 = ~pi1026 & ~n15400;
  assign n18330 = ~n18328 & ~n18329;
  assign n18331 = n15326 & ~n18330;
  assign n18332 = ~pi1026 & ~n15326;
  assign po1206 = n18331 | n18332;
  assign n18334 = n15400 & ~n18059;
  assign n18335 = ~pi1027 & ~n15400;
  assign n18336 = ~n18334 & ~n18335;
  assign n18337 = n15326 & ~n18336;
  assign n18338 = ~pi1027 & ~n15326;
  assign po1207 = n18337 | n18338;
  assign n18340 = n15407 & ~n18162;
  assign n18341 = ~pi1028 & ~n15407;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = n15326 & ~n18342;
  assign n18344 = ~pi1028 & ~n15326;
  assign po1208 = n18343 | n18344;
  assign n18346 = n15407 & ~n18059;
  assign n18347 = ~pi1029 & ~n15407;
  assign n18348 = ~n18346 & ~n18347;
  assign n18349 = n15326 & ~n18348;
  assign n18350 = ~pi1029 & ~n15326;
  assign po1209 = n18349 | n18350;
  assign n18352 = n16635 & ~n18162;
  assign n18353 = ~pi1030 & ~n16635;
  assign n18354 = ~n18352 & ~n18353;
  assign n18355 = n15326 & ~n18354;
  assign n18356 = ~pi1030 & ~n15326;
  assign po1210 = n18355 | n18356;
  assign n18358 = n16635 & ~n18105;
  assign n18359 = ~pi1031 & ~n16635;
  assign n18360 = ~n18358 & ~n18359;
  assign n18361 = n15326 & ~n18360;
  assign n18362 = ~pi1031 & ~n15326;
  assign po1211 = n18361 | n18362;
  assign n18364 = n16635 & ~n18077;
  assign n18365 = ~pi1032 & ~n16635;
  assign n18366 = ~n18364 & ~n18365;
  assign n18367 = n15326 & ~n18366;
  assign n18368 = ~pi1032 & ~n15326;
  assign po1212 = n18367 | n18368;
  assign n18370 = n16635 & ~n18068;
  assign n18371 = ~pi1033 & ~n16635;
  assign n18372 = ~n18370 & ~n18371;
  assign n18373 = n15326 & ~n18372;
  assign n18374 = ~pi1033 & ~n15326;
  assign po1213 = n18373 | n18374;
  assign n18376 = n16635 & ~n18059;
  assign n18377 = ~pi1034 & ~n16635;
  assign n18378 = ~n18376 & ~n18377;
  assign n18379 = n15326 & ~n18378;
  assign n18380 = ~pi1034 & ~n15326;
  assign po1214 = n18379 | n18380;
  assign n18382 = n15434 & ~n18162;
  assign n18383 = ~pi1035 & ~n15434;
  assign n18384 = ~n18382 & ~n18383;
  assign n18385 = n15326 & ~n18384;
  assign n18386 = ~pi1035 & ~n15326;
  assign po1215 = n18385 | n18386;
  assign n18388 = n15434 & ~n18105;
  assign n18389 = ~pi1036 & ~n15434;
  assign n18390 = ~n18388 & ~n18389;
  assign n18391 = n15326 & ~n18390;
  assign n18392 = ~pi1036 & ~n15326;
  assign po1216 = n18391 | n18392;
  assign n18394 = n15434 & ~n18077;
  assign n18395 = ~pi1037 & ~n15434;
  assign n18396 = ~n18394 & ~n18395;
  assign n18397 = n15326 & ~n18396;
  assign n18398 = ~pi1037 & ~n15326;
  assign po1217 = n18397 | n18398;
  assign n18400 = n15434 & ~n18068;
  assign n18401 = ~pi1038 & ~n15434;
  assign n18402 = ~n18400 & ~n18401;
  assign n18403 = n15326 & ~n18402;
  assign n18404 = ~pi1038 & ~n15326;
  assign po1218 = n18403 | n18404;
  assign n18406 = n15434 & ~n18059;
  assign n18407 = ~pi1039 & ~n15434;
  assign n18408 = ~n18406 & ~n18407;
  assign n18409 = n15326 & ~n18408;
  assign n18410 = ~pi1039 & ~n15326;
  assign po1219 = n18409 | n18410;
  assign n18412 = ~pi1040 & ~n16870;
  assign n18413 = n16870 & ~n18162;
  assign n18414 = ~n18412 & ~n18413;
  assign n18415 = n15326 & ~n18414;
  assign n18416 = ~pi1040 & ~n15326;
  assign po1220 = n18415 | n18416;
  assign n18418 = ~pi1041 & ~n16870;
  assign n18419 = n16870 & ~n18059;
  assign n18420 = ~n18418 & ~n18419;
  assign n18421 = n15326 & ~n18420;
  assign n18422 = ~pi1041 & ~n15326;
  assign po1221 = n18421 | n18422;
  assign n18424 = ~pi1042 & ~n17015;
  assign n18425 = n17015 & ~n18162;
  assign n18426 = ~n18424 & ~n18425;
  assign n18427 = n15326 & ~n18426;
  assign n18428 = ~pi1042 & ~n15326;
  assign po1222 = n18427 | n18428;
  assign n18430 = ~pi1043 & ~n17015;
  assign n18431 = n17015 & n18049;
  assign n18432 = ~n18430 & ~n18431;
  assign n18433 = n15326 & ~n18432;
  assign n18434 = ~pi1043 & ~n15326;
  assign po1223 = n18433 | n18434;
  assign n18436 = ~pi1044 & ~n17015;
  assign n18437 = n17015 & ~n18213;
  assign n18438 = ~n18436 & ~n18437;
  assign n18439 = n15326 & ~n18438;
  assign n18440 = ~pi1044 & ~n15326;
  assign po1224 = n18439 | n18440;
  assign n18442 = ~pi1045 & ~n17154;
  assign n18443 = n17154 & ~n18162;
  assign n18444 = ~n18442 & ~n18443;
  assign n18445 = n15326 & ~n18444;
  assign n18446 = ~pi1045 & ~n15326;
  assign po1225 = n18445 | n18446;
  assign n18448 = ~pi1046 & ~n17154;
  assign n18449 = n17154 & ~n18059;
  assign n18450 = ~n18448 & ~n18449;
  assign n18451 = n15326 & ~n18450;
  assign n18452 = ~pi1046 & ~n15326;
  assign po1226 = n18451 | n18452;
  assign n18454 = ~pi1047 & ~n17154;
  assign n18455 = n17154 & ~n18213;
  assign n18456 = ~n18454 & ~n18455;
  assign n18457 = n15326 & ~n18456;
  assign n18458 = ~pi1047 & ~n15326;
  assign po1227 = n18457 | n18458;
  assign n18460 = ~pi1048 & ~n15312;
  assign n18461 = n15312 & ~n18162;
  assign n18462 = ~n18460 & ~n18461;
  assign n18463 = n15326 & ~n18462;
  assign n18464 = ~pi1048 & ~n15326;
  assign po1228 = n18463 | n18464;
  assign n18466 = ~pi1049 & ~n15312;
  assign n18467 = n15312 & ~n18105;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = n15326 & ~n18468;
  assign n18470 = ~pi1049 & ~n15326;
  assign po1229 = n18469 | n18470;
  assign n18472 = ~pi1050 & ~n15312;
  assign n18473 = n15312 & n18049;
  assign n18474 = ~n18472 & ~n18473;
  assign n18475 = n15326 & ~n18474;
  assign n18476 = ~pi1050 & ~n15326;
  assign po1230 = n18475 | n18476;
  assign n18478 = ~pi1051 & ~n15312;
  assign n18479 = n15312 & ~n18213;
  assign n18480 = ~n18478 & ~n18479;
  assign n18481 = n15326 & ~n18480;
  assign n18482 = ~pi1051 & ~n15326;
  assign po1231 = n18481 | n18482;
  assign n18484 = n16635 & n18049;
  assign n18485 = ~pi1052 & ~n16635;
  assign n18486 = ~n18484 & ~n18485;
  assign n18487 = n15326 & ~n18486;
  assign n18488 = ~pi1052 & ~n15326;
  assign po1232 = n18487 | n18488;
  assign n18490 = ~pi1053 & ~n17437;
  assign n18491 = n17437 & ~n18162;
  assign n18492 = ~n18490 & ~n18491;
  assign n18493 = n15326 & ~n18492;
  assign n18494 = ~pi1053 & ~n15326;
  assign po1233 = n18493 | n18494;
  assign n18496 = ~pi1054 & ~n17437;
  assign n18497 = n17437 & ~n18105;
  assign n18498 = ~n18496 & ~n18497;
  assign n18499 = n15326 & ~n18498;
  assign n18500 = ~pi1054 & ~n15326;
  assign po1234 = n18499 | n18500;
  assign n18502 = ~pi1055 & ~n17437;
  assign n18503 = n17437 & n18049;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = n15326 & ~n18504;
  assign n18506 = ~pi1055 & ~n15326;
  assign po1235 = n18505 | n18506;
  assign n18508 = ~pi1056 & ~n17437;
  assign n18509 = n17437 & ~n18068;
  assign n18510 = ~n18508 & ~n18509;
  assign n18511 = n15326 & ~n18510;
  assign n18512 = ~pi1056 & ~n15326;
  assign po1236 = n18511 | n18512;
  assign n18514 = ~pi1057 & ~n17437;
  assign n18515 = n17437 & ~n18059;
  assign n18516 = ~n18514 & ~n18515;
  assign n18517 = n15326 & ~n18516;
  assign n18518 = ~pi1057 & ~n15326;
  assign po1237 = n18517 | n18518;
  assign n18520 = n15434 & n18049;
  assign n18521 = ~pi1058 & ~n15434;
  assign n18522 = ~n18520 & ~n18521;
  assign n18523 = n15326 & ~n18522;
  assign n18524 = ~pi1058 & ~n15326;
  assign po1238 = n18523 | n18524;
  assign n18526 = ~pi1059 & ~n17154;
  assign n18527 = n17154 & n18049;
  assign n18528 = ~n18526 & ~n18527;
  assign n18529 = n15326 & ~n18528;
  assign n18530 = ~pi1059 & ~n15326;
  assign po1239 = n18529 | n18530;
  assign n18532 = ~pi1060 & ~n17154;
  assign n18533 = n17154 & ~n18068;
  assign n18534 = ~n18532 & ~n18533;
  assign n18535 = n15326 & ~n18534;
  assign n18536 = ~pi1060 & ~n15326;
  assign po1240 = n18535 | n18536;
  assign n18538 = n15335 & ~n18097;
  assign n18539 = ~pi1061 & ~n15335;
  assign n18540 = ~n18538 & ~n18539;
  assign n18541 = n15326 & ~n18540;
  assign n18542 = ~pi1061 & ~n15326;
  assign po1241 = n18541 | n18542;
  assign n18544 = n15414 & ~n18213;
  assign n18545 = ~pi1062 & ~n15414;
  assign n18546 = ~n18544 & ~n18545;
  assign n18547 = n15326 & ~n18546;
  assign n18548 = ~pi1062 & ~n15326;
  assign po1242 = n18547 | n18548;
  assign n18550 = ~pi1063 & ~n17154;
  assign n18551 = n17154 & ~n18077;
  assign n18552 = ~n18550 & ~n18551;
  assign n18553 = n15326 & ~n18552;
  assign n18554 = ~pi1063 & ~n15326;
  assign po1243 = n18553 | n18554;
  assign n18556 = ~pi1064 & ~n17154;
  assign n18557 = n17154 & ~n18086;
  assign n18558 = ~n18556 & ~n18557;
  assign n18559 = n15326 & ~n18558;
  assign n18560 = ~pi1064 & ~n15326;
  assign po1244 = n18559 | n18560;
  assign n18562 = n15414 & ~n18068;
  assign n18563 = ~pi1065 & ~n15414;
  assign n18564 = ~n18562 & ~n18563;
  assign n18565 = n15326 & ~n18564;
  assign n18566 = ~pi1065 & ~n15326;
  assign po1245 = n18565 | n18566;
  assign n18568 = ~pi1066 & ~n17154;
  assign n18569 = n17154 & ~n18105;
  assign n18570 = ~n18568 & ~n18569;
  assign n18571 = n15326 & ~n18570;
  assign n18572 = ~pi1066 & ~n15326;
  assign po1246 = n18571 | n18572;
  assign n18574 = ~pi1067 & ~n17015;
  assign n18575 = n17015 & ~n18068;
  assign n18576 = ~n18574 & ~n18575;
  assign n18577 = n15326 & ~n18576;
  assign n18578 = ~pi1067 & ~n15326;
  assign po1247 = n18577 | n18578;
  assign n18580 = ~pi1068 & ~n17154;
  assign n18581 = n17154 & ~n18097;
  assign n18582 = ~n18580 & ~n18581;
  assign n18583 = n15326 & ~n18582;
  assign n18584 = ~pi1068 & ~n15326;
  assign po1248 = n18583 | n18584;
  assign n18586 = n15414 & ~n18086;
  assign n18587 = ~pi1069 & ~n15414;
  assign n18588 = ~n18586 & ~n18587;
  assign n18589 = n15326 & ~n18588;
  assign n18590 = ~pi1069 & ~n15326;
  assign po1249 = n18589 | n18590;
  assign n18592 = ~pi1070 & ~n17015;
  assign n18593 = n17015 & ~n18059;
  assign n18594 = ~n18592 & ~n18593;
  assign n18595 = n15326 & ~n18594;
  assign n18596 = ~pi1070 & ~n15326;
  assign po1250 = n18595 | n18596;
  assign n18598 = ~pi1071 & ~n17015;
  assign n18599 = n17015 & ~n18105;
  assign n18600 = ~n18598 & ~n18599;
  assign n18601 = n15326 & ~n18600;
  assign n18602 = ~pi1071 & ~n15326;
  assign po1251 = n18601 | n18602;
  assign n18604 = ~pi1072 & ~n17015;
  assign n18605 = n17015 & ~n18077;
  assign n18606 = ~n18604 & ~n18605;
  assign n18607 = n15326 & ~n18606;
  assign n18608 = ~pi1072 & ~n15326;
  assign po1252 = n18607 | n18608;
  assign n18610 = n15414 & ~n18097;
  assign n18611 = ~pi1073 & ~n15414;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = n15326 & ~n18612;
  assign n18614 = ~pi1073 & ~n15326;
  assign po1253 = n18613 | n18614;
  assign n18616 = ~pi1074 & ~n17015;
  assign n18617 = n17015 & ~n18086;
  assign n18618 = ~n18616 & ~n18617;
  assign n18619 = n15326 & ~n18618;
  assign n18620 = ~pi1074 & ~n15326;
  assign po1254 = n18619 | n18620;
  assign n18622 = n15434 & ~n18086;
  assign n18623 = ~pi1075 & ~n15434;
  assign n18624 = ~n18622 & ~n18623;
  assign n18625 = n15326 & ~n18624;
  assign n18626 = ~pi1075 & ~n15326;
  assign po1255 = n18625 | n18626;
  assign n18628 = n15393 & ~n18213;
  assign n18629 = ~pi1076 & ~n15393;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = n15326 & ~n18630;
  assign n18632 = ~pi1076 & ~n15326;
  assign po1256 = n18631 | n18632;
  assign n18634 = ~pi1077 & ~n16870;
  assign n18635 = n16870 & ~n18213;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = n15326 & ~n18636;
  assign n18638 = ~pi1077 & ~n15326;
  assign po1257 = n18637 | n18638;
  assign n18640 = n15386 & ~n18077;
  assign n18641 = ~pi1078 & ~n15386;
  assign n18642 = ~n18640 & ~n18641;
  assign n18643 = n15326 & ~n18642;
  assign n18644 = ~pi1078 & ~n15326;
  assign po1258 = n18643 | n18644;
  assign n18646 = ~pi1079 & ~n17015;
  assign n18647 = n17015 & ~n18097;
  assign n18648 = ~n18646 & ~n18647;
  assign n18649 = n15326 & ~n18648;
  assign n18650 = ~pi1079 & ~n15326;
  assign po1259 = n18649 | n18650;
  assign n18652 = n15393 & n18049;
  assign n18653 = ~pi1080 & ~n15393;
  assign n18654 = ~n18652 & ~n18653;
  assign n18655 = n15326 & ~n18654;
  assign n18656 = ~pi1080 & ~n15326;
  assign po1260 = n18655 | n18656;
  assign n18658 = ~pi1081 & ~n16870;
  assign n18659 = n16870 & ~n18086;
  assign n18660 = ~n18658 & ~n18659;
  assign n18661 = n15326 & ~n18660;
  assign n18662 = ~pi1081 & ~n15326;
  assign po1261 = n18661 | n18662;
  assign n18664 = ~pi1082 & ~n16870;
  assign n18665 = n16870 & n18049;
  assign n18666 = ~n18664 & ~n18665;
  assign n18667 = n15326 & ~n18666;
  assign n18668 = ~pi1082 & ~n15326;
  assign po1262 = n18667 | n18668;
  assign n18670 = ~pi1083 & ~n16870;
  assign n18671 = n16870 & ~n18068;
  assign n18672 = ~n18670 & ~n18671;
  assign n18673 = n15326 & ~n18672;
  assign n18674 = ~pi1083 & ~n15326;
  assign po1263 = n18673 | n18674;
  assign n18676 = n15393 & ~n18086;
  assign n18677 = ~pi1084 & ~n15393;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 = n15326 & ~n18678;
  assign n18680 = ~pi1084 & ~n15326;
  assign po1264 = n18679 | n18680;
  assign n18682 = ~pi1085 & ~n16870;
  assign n18683 = n16870 & ~n18077;
  assign n18684 = ~n18682 & ~n18683;
  assign n18685 = n15326 & ~n18684;
  assign n18686 = ~pi1085 & ~n15326;
  assign po1265 = n18685 | n18686;
  assign n18688 = n15374 & n18049;
  assign n18689 = ~pi1086 & ~n15374;
  assign n18690 = ~n18688 & ~n18689;
  assign n18691 = n15326 & ~n18690;
  assign n18692 = ~pi1086 & ~n15326;
  assign po1266 = n18691 | n18692;
  assign n18694 = ~pi1087 & ~n16870;
  assign n18695 = n16870 & ~n18105;
  assign n18696 = ~n18694 & ~n18695;
  assign n18697 = n15326 & ~n18696;
  assign n18698 = ~pi1087 & ~n15326;
  assign po1267 = n18697 | n18698;
  assign n18700 = n15393 & ~n18162;
  assign n18701 = ~pi1088 & ~n15393;
  assign n18702 = ~n18700 & ~n18701;
  assign n18703 = n15326 & ~n18702;
  assign n18704 = ~pi1088 & ~n15326;
  assign po1268 = n18703 | n18704;
  assign n18706 = ~pi1089 & ~n16870;
  assign n18707 = n16870 & ~n18097;
  assign n18708 = ~n18706 & ~n18707;
  assign n18709 = n15326 & ~n18708;
  assign n18710 = ~pi1089 & ~n15326;
  assign po1269 = n18709 | n18710;
  assign n18712 = n15386 & ~n18213;
  assign n18713 = ~pi1090 & ~n15386;
  assign n18714 = ~n18712 & ~n18713;
  assign n18715 = n15326 & ~n18714;
  assign n18716 = ~pi1090 & ~n15326;
  assign po1270 = n18715 | n18716;
  assign n18718 = n15434 & ~n18213;
  assign n18719 = ~pi1091 & ~n15434;
  assign n18720 = ~n18718 & ~n18719;
  assign n18721 = n15326 & ~n18720;
  assign n18722 = ~pi1091 & ~n15326;
  assign po1271 = n18721 | n18722;
  assign n18724 = n15386 & n18049;
  assign n18725 = ~pi1092 & ~n15386;
  assign n18726 = ~n18724 & ~n18725;
  assign n18727 = n15326 & ~n18726;
  assign n18728 = ~pi1092 & ~n15326;
  assign po1272 = n18727 | n18728;
  assign n18730 = n15434 & ~n18097;
  assign n18731 = ~pi1093 & ~n15434;
  assign n18732 = ~n18730 & ~n18731;
  assign n18733 = n15326 & ~n18732;
  assign n18734 = ~pi1093 & ~n15326;
  assign po1273 = n18733 | n18734;
  assign n18736 = n16635 & ~n18213;
  assign n18737 = ~pi1094 & ~n16635;
  assign n18738 = ~n18736 & ~n18737;
  assign n18739 = n15326 & ~n18738;
  assign n18740 = ~pi1094 & ~n15326;
  assign po1274 = n18739 | n18740;
  assign n18742 = n15386 & ~n18097;
  assign n18743 = ~pi1095 & ~n15386;
  assign n18744 = ~n18742 & ~n18743;
  assign n18745 = n15326 & ~n18744;
  assign n18746 = ~pi1095 & ~n15326;
  assign po1275 = n18745 | n18746;
  assign n18748 = n15386 & ~n18162;
  assign n18749 = ~pi1096 & ~n15386;
  assign n18750 = ~n18748 & ~n18749;
  assign n18751 = n15326 & ~n18750;
  assign n18752 = ~pi1096 & ~n15326;
  assign po1276 = n18751 | n18752;
  assign n18754 = n16635 & ~n18086;
  assign n18755 = ~pi1097 & ~n16635;
  assign n18756 = ~n18754 & ~n18755;
  assign n18757 = n15326 & ~n18756;
  assign n18758 = ~pi1097 & ~n15326;
  assign po1277 = n18757 | n18758;
  assign n18760 = n16635 & ~n18097;
  assign n18761 = ~pi1098 & ~n16635;
  assign n18762 = ~n18760 & ~n18761;
  assign n18763 = n15326 & ~n18762;
  assign n18764 = ~pi1098 & ~n15326;
  assign po1278 = n18763 | n18764;
  assign n18766 = n15407 & ~n18068;
  assign n18767 = ~pi1099 & ~n15407;
  assign n18768 = ~n18766 & ~n18767;
  assign n18769 = n15326 & ~n18768;
  assign n18770 = ~pi1099 & ~n15326;
  assign po1279 = n18769 | n18770;
  assign n18772 = n15407 & ~n18213;
  assign n18773 = ~pi1100 & ~n15407;
  assign n18774 = ~n18772 & ~n18773;
  assign n18775 = n15326 & ~n18774;
  assign n18776 = ~pi1100 & ~n15326;
  assign po1280 = n18775 | n18776;
  assign n18778 = n15407 & ~n18077;
  assign n18779 = ~pi1101 & ~n15407;
  assign n18780 = ~n18778 & ~n18779;
  assign n18781 = n15326 & ~n18780;
  assign n18782 = ~pi1101 & ~n15326;
  assign po1281 = n18781 | n18782;
  assign n18784 = n15407 & ~n18086;
  assign n18785 = ~pi1102 & ~n15407;
  assign n18786 = ~n18784 & ~n18785;
  assign n18787 = n15326 & ~n18786;
  assign n18788 = ~pi1102 & ~n15326;
  assign po1282 = n18787 | n18788;
  assign n18790 = n15407 & ~n18105;
  assign n18791 = ~pi1103 & ~n15407;
  assign n18792 = ~n18790 & ~n18791;
  assign n18793 = n15326 & ~n18792;
  assign n18794 = ~pi1103 & ~n15326;
  assign po1283 = n18793 | n18794;
  assign n18796 = n15407 & ~n18097;
  assign n18797 = ~pi1104 & ~n15407;
  assign n18798 = ~n18796 & ~n18797;
  assign n18799 = n15326 & ~n18798;
  assign n18800 = ~pi1104 & ~n15326;
  assign po1284 = n18799 | n18800;
  assign n18802 = n15400 & ~n18213;
  assign n18803 = ~pi1105 & ~n15400;
  assign n18804 = ~n18802 & ~n18803;
  assign n18805 = n15326 & ~n18804;
  assign n18806 = ~pi1105 & ~n15326;
  assign po1285 = n18805 | n18806;
  assign n18808 = n15400 & ~n18086;
  assign n18809 = ~pi1106 & ~n15400;
  assign n18810 = ~n18808 & ~n18809;
  assign n18811 = n15326 & ~n18810;
  assign n18812 = ~pi1106 & ~n15326;
  assign po1286 = n18811 | n18812;
  assign n18814 = n15400 & ~n18097;
  assign n18815 = ~pi1107 & ~n15400;
  assign n18816 = ~n18814 & ~n18815;
  assign n18817 = n15326 & ~n18816;
  assign n18818 = ~pi1107 & ~n15326;
  assign po1287 = n18817 | n18818;
  assign n18820 = n15374 & ~n18086;
  assign n18821 = ~pi1108 & ~n15374;
  assign n18822 = ~n18820 & ~n18821;
  assign n18823 = n15326 & ~n18822;
  assign n18824 = ~pi1108 & ~n15326;
  assign po1288 = n18823 | n18824;
  assign n18826 = n16136 & ~n18213;
  assign n18827 = ~pi1109 & ~n16136;
  assign n18828 = ~n18826 & ~n18827;
  assign n18829 = n15326 & ~n18828;
  assign n18830 = ~pi1109 & ~n15326;
  assign po1289 = n18829 | n18830;
  assign n18832 = n16136 & n18049;
  assign n18833 = ~pi1110 & ~n16136;
  assign n18834 = ~n18832 & ~n18833;
  assign n18835 = n15326 & ~n18834;
  assign n18836 = ~pi1110 & ~n15326;
  assign po1290 = n18835 | n18836;
  assign n18838 = n16136 & ~n18077;
  assign n18839 = ~pi1111 & ~n16136;
  assign n18840 = ~n18838 & ~n18839;
  assign n18841 = n15326 & ~n18840;
  assign n18842 = ~pi1111 & ~n15326;
  assign po1291 = n18841 | n18842;
  assign n18844 = n15335 & ~n18105;
  assign n18845 = ~pi1112 & ~n15335;
  assign n18846 = ~n18844 & ~n18845;
  assign n18847 = n15326 & ~n18846;
  assign n18848 = ~pi1112 & ~n15326;
  assign po1292 = n18847 | n18848;
  assign n18850 = n15427 & ~n18086;
  assign n18851 = ~pi1113 & ~n15427;
  assign n18852 = ~n18850 & ~n18851;
  assign n18853 = n15326 & ~n18852;
  assign n18854 = ~pi1113 & ~n15326;
  assign po1293 = n18853 | n18854;
  assign n18856 = n16136 & ~n18097;
  assign n18857 = ~pi1114 & ~n16136;
  assign n18858 = ~n18856 & ~n18857;
  assign n18859 = n15326 & ~n18858;
  assign n18860 = ~pi1114 & ~n15326;
  assign po1294 = n18859 | n18860;
  assign n18862 = n16136 & ~n18162;
  assign n18863 = ~pi1115 & ~n16136;
  assign n18864 = ~n18862 & ~n18863;
  assign n18865 = n15326 & ~n18864;
  assign n18866 = ~pi1115 & ~n15326;
  assign po1295 = n18865 | n18866;
  assign n18868 = n15427 & n18049;
  assign n18869 = ~pi1116 & ~n15427;
  assign n18870 = ~n18868 & ~n18869;
  assign n18871 = n15326 & ~n18870;
  assign n18872 = ~pi1116 & ~n15326;
  assign po1296 = n18871 | n18872;
  assign n18874 = n15427 & ~n18213;
  assign n18875 = ~pi1117 & ~n15427;
  assign n18876 = ~n18874 & ~n18875;
  assign n18877 = n15326 & ~n18876;
  assign n18878 = ~pi1117 & ~n15326;
  assign po1297 = n18877 | n18878;
  assign n18880 = n15427 & ~n18077;
  assign n18881 = ~pi1118 & ~n15427;
  assign n18882 = ~n18880 & ~n18881;
  assign n18883 = n15326 & ~n18882;
  assign n18884 = ~pi1118 & ~n15326;
  assign po1298 = n18883 | n18884;
  assign n18886 = n15427 & ~n18105;
  assign n18887 = ~pi1119 & ~n15427;
  assign n18888 = ~n18886 & ~n18887;
  assign n18889 = n15326 & ~n18888;
  assign n18890 = ~pi1119 & ~n15326;
  assign po1299 = n18889 | n18890;
  assign n18892 = ~pi1120 & ~n17437;
  assign n18893 = n17437 & ~n18077;
  assign n18894 = ~n18892 & ~n18893;
  assign n18895 = n15326 & ~n18894;
  assign n18896 = ~pi1120 & ~n15326;
  assign po1300 = n18895 | n18896;
  assign n18898 = ~pi1121 & ~n17437;
  assign n18899 = n17437 & ~n18213;
  assign n18900 = ~n18898 & ~n18899;
  assign n18901 = n15326 & ~n18900;
  assign n18902 = ~pi1121 & ~n15326;
  assign po1301 = n18901 | n18902;
  assign n18904 = n15335 & ~n18059;
  assign n18905 = ~pi1122 & ~n15335;
  assign n18906 = ~n18904 & ~n18905;
  assign n18907 = n15326 & ~n18906;
  assign n18908 = ~pi1122 & ~n15326;
  assign po1302 = n18907 | n18908;
  assign n18910 = n15407 & n18049;
  assign n18911 = ~pi1123 & ~n15407;
  assign n18912 = ~n18910 & ~n18911;
  assign n18913 = n15326 & ~n18912;
  assign n18914 = ~pi1123 & ~n15326;
  assign po1303 = n18913 | n18914;
  assign n18916 = ~pi1124 & ~n17437;
  assign n18917 = n17437 & ~n18086;
  assign n18918 = ~n18916 & ~n18917;
  assign n18919 = n15326 & ~n18918;
  assign n18920 = ~pi1124 & ~n15326;
  assign po1304 = n18919 | n18920;
  assign n18922 = ~pi1125 & ~n17437;
  assign n18923 = n17437 & ~n18097;
  assign n18924 = ~n18922 & ~n18923;
  assign n18925 = n15326 & ~n18924;
  assign n18926 = ~pi1125 & ~n15326;
  assign po1305 = n18925 | n18926;
  assign n18928 = n15335 & ~n18086;
  assign n18929 = ~pi1126 & ~n15335;
  assign n18930 = ~n18928 & ~n18929;
  assign n18931 = n15326 & ~n18930;
  assign n18932 = ~pi1126 & ~n15326;
  assign po1306 = n18931 | n18932;
  assign n18934 = n15335 & ~n18077;
  assign n18935 = ~pi1127 & ~n15335;
  assign n18936 = ~n18934 & ~n18935;
  assign n18937 = n15326 & ~n18936;
  assign n18938 = ~pi1127 & ~n15326;
  assign po1307 = n18937 | n18938;
  assign n18940 = pi0134 & ~pi3206;
  assign n18941 = pi1984 & ~n18940;
  assign n18942 = n11945 & n18940;
  assign po1308 = n18941 | n18942;
  assign n18944 = ~pi1129 & ~n11939;
  assign n18945 = ~n11943 & ~n18944;
  assign n18946 = n18940 & ~n18945;
  assign n18947 = ~pi1984 & ~n18940;
  assign po1309 = n18946 | n18947;
  assign n18949 = pi1828 & ~n18940;
  assign n18950 = ~n11955 & n18940;
  assign po1310 = n18949 | n18950;
  assign n18952 = pi1985 & ~n18940;
  assign n18953 = n11971 & n18940;
  assign po1311 = n18952 | n18953;
  assign n18955 = pi1679 & n8187;
  assign n18956 = ~n8206 & n15319;
  assign n18957 = n8198 & n18956;
  assign n18958 = n18955 & n18957;
  assign n18959 = pi0081 & ~pi1353;
  assign n18960 = n18958 & ~n18959;
  assign n18961 = ~pi1353 & n18960;
  assign n18962 = ~pi1132 & ~n18961;
  assign n18963 = ~n15442 & n18961;
  assign po1312 = n18962 | n18963;
  assign n18965 = ~pi1133 & ~n18961;
  assign n18966 = ~n15451 & n18961;
  assign po1313 = n18965 | n18966;
  assign n18968 = ~pi1134 & ~n18961;
  assign n18969 = ~n15316 & n18961;
  assign po1314 = n18968 | n18969;
  assign n18971 = ~pi1135 & ~n18961;
  assign n18972 = ~n15466 & n18961;
  assign po1315 = n18971 | n18972;
  assign n18974 = ~pi1136 & ~n18961;
  assign n18975 = ~n15475 & n18961;
  assign po1316 = n18974 | n18975;
  assign n18977 = ~pi1137 & ~n18961;
  assign n18978 = ~n15484 & n18961;
  assign po1317 = n18977 | n18978;
  assign n18980 = ~pi1138 & ~n18961;
  assign n18981 = ~n15493 & n18961;
  assign po1318 = n18980 | n18981;
  assign n18983 = ~pi1139 & ~n18961;
  assign n18984 = ~n15332 & n18961;
  assign po1319 = n18983 | n18984;
  assign n18986 = ~pi1140 & ~n18961;
  assign n18987 = ~n15709 & n18961;
  assign po1320 = n18986 | n18987;
  assign n18989 = ~pi1141 & ~n18961;
  assign n18990 = ~n15517 & n18961;
  assign po1321 = n18989 | n18990;
  assign n18992 = ~pi1142 & ~n18961;
  assign n18993 = ~n15535 & n18961;
  assign po1322 = n18992 | n18993;
  assign n18995 = ~pi1143 & ~n18961;
  assign n18996 = ~n15544 & n18961;
  assign po1323 = n18995 | n18996;
  assign n18998 = ~pi1144 & ~n18961;
  assign n18999 = ~n15553 & n18961;
  assign po1324 = n18998 | n18999;
  assign n19001 = ~pi1145 & ~n18961;
  assign n19002 = ~n15700 & n18961;
  assign po1325 = n19001 | n19002;
  assign n19004 = ~pi1146 & ~n18961;
  assign n19005 = ~n15562 & n18961;
  assign po1326 = n19004 | n19005;
  assign n19007 = ~pi1147 & ~n18961;
  assign n19008 = ~n15580 & n18961;
  assign po1327 = n19007 | n19008;
  assign n19010 = ~pi1148 & ~n18961;
  assign n19011 = ~n15589 & n18961;
  assign po1328 = n19010 | n19011;
  assign n19013 = ~pi1149 & ~n18961;
  assign n19014 = ~n15607 & n18961;
  assign po1329 = n19013 | n19014;
  assign n19016 = ~pi1150 & ~n18961;
  assign n19017 = ~n15616 & n18961;
  assign po1330 = n19016 | n19017;
  assign n19019 = ~pi1151 & ~n18961;
  assign n19020 = ~n15625 & n18961;
  assign po1331 = n19019 | n19020;
  assign n19022 = pi1152 & ~n15326;
  assign n19023 = pi1152 & pi1154;
  assign n19024 = ~pi1152 & ~pi1154;
  assign n19025 = ~n19023 & ~n19024;
  assign n19026 = n15326 & n19025;
  assign po1332 = n19022 | n19026;
  assign n19028 = pi1153 & ~n15326;
  assign po1333 = n19026 | n19028;
  assign n19030 = pi1154 & ~n15326;
  assign n19031 = ~pi1154 & n15326;
  assign po1334 = n19030 | n19031;
  assign n19033 = ~pi1155 & ~n18961;
  assign n19034 = ~n15598 & n18961;
  assign po1335 = n19033 | n19034;
  assign n19036 = ~pi1156 & ~n18961;
  assign n19037 = ~n15571 & n18961;
  assign po1336 = n19036 | n19037;
  assign n19039 = ~pi1157 & ~n18961;
  assign n19040 = ~n15502 & n18961;
  assign po1337 = n19039 | n19040;
  assign n19042 = ~pi1158 & ~n18961;
  assign n19043 = ~n15526 & n18961;
  assign po1338 = n19042 | n19043;
  assign n19045 = ~pi1161 & n8074;
  assign n19046 = pi1160 & pi1161;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = pi1159 & pi1161;
  assign n19049 = n19047 & ~n19048;
  assign n19050 = pi1159 & pi1160;
  assign n19051 = ~n8046 & n9242;
  assign n19052 = n8075 & ~n8078;
  assign n19053 = n19051 & ~n19052;
  assign n19054 = ~n19050 & n19053;
  assign n19055 = n19049 & n19054;
  assign n19056 = pi1159 & n19055;
  assign n19057 = ~pi1161 & ~n8074;
  assign n19058 = ~n19050 & n19057;
  assign n19059 = ~n19055 & ~n19058;
  assign po1339 = n19056 | n19059;
  assign n19061 = pi1160 & n19055;
  assign n19062 = n8044 & ~n19055;
  assign po1340 = n19061 | n19062;
  assign n19064 = pi1161 & n19055;
  assign n19065 = n8046 & ~n19055;
  assign po1341 = n19064 | n19065;
  assign n19067 = pi1828 & pi1984;
  assign n19068 = ~pi1985 & ~n19067;
  assign n19069 = pi1984 & pi1985;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = ~pi1828 & pi1985;
  assign n19072 = ~n19070 & ~n19071;
  assign n19073 = ~n18940 & ~n19072;
  assign n19074 = ~pi1162 & ~n11939;
  assign n19075 = ~pi1129 & ~pi1177;
  assign n19076 = pi1162 & n19075;
  assign n19077 = ~pi1162 & ~n19075;
  assign n19078 = ~n19076 & ~n19077;
  assign n19079 = n11939 & ~n19078;
  assign n19080 = ~n19074 & ~n19079;
  assign n19081 = n18940 & ~n19080;
  assign po1342 = n19073 | n19081;
  assign n19083 = ~pi1877 & ~n18940;
  assign n19084 = pi1163 & ~n11939;
  assign n19085 = ~pi1128 & pi1130;
  assign n19086 = pi1128 & ~pi1130;
  assign n19087 = ~n19085 & ~n19086;
  assign n19088 = n11939 & ~n19087;
  assign n19089 = ~n19084 & ~n19088;
  assign n19090 = n18940 & ~n19089;
  assign po1343 = n19083 | n19090;
  assign n19092 = ~pi2384 & ~n18940;
  assign n19093 = pi1164 & ~n11939;
  assign n19094 = ~pi1130 & pi1131;
  assign n19095 = pi1130 & ~pi1131;
  assign n19096 = ~n19094 & ~n19095;
  assign n19097 = n11939 & ~n19096;
  assign n19098 = ~n19093 & ~n19097;
  assign n19099 = n18940 & ~n19098;
  assign po1344 = n19092 | n19099;
  assign n19101 = ~pi1986 & ~n18940;
  assign n19102 = pi1165 & ~n11939;
  assign n19103 = ~pi1181 & n11939;
  assign n19104 = ~n19102 & ~n19103;
  assign n19105 = n18940 & ~n19104;
  assign po1345 = n19101 | n19105;
  assign n19107 = ~n15333 & ~n15384;
  assign n19108 = n15326 & ~n19107;
  assign n19109 = pi1166 & ~n15326;
  assign po1346 = n19108 | n19109;
  assign n19111 = pi1154 & n15310;
  assign n19112 = pi1167 & ~n19111;
  assign n19113 = ~pi1167 & n19111;
  assign n19114 = ~n19112 & ~n19113;
  assign n19115 = n15326 & ~n19114;
  assign n19116 = pi1167 & ~n15326;
  assign po1347 = n19115 | n19116;
  assign n19118 = pi1153 & n15326;
  assign n19119 = pi1168 & ~n15326;
  assign po1348 = n19118 | n19119;
  assign n19121 = pi1166 & n15326;
  assign n19122 = pi1169 & ~n15326;
  assign po1349 = n19121 | n19122;
  assign n19124 = pi1172 & n15326;
  assign n19125 = pi1170 & ~n15326;
  assign po1350 = n19124 | n19125;
  assign n19127 = pi1175 & n15326;
  assign n19128 = pi1171 & ~n15326;
  assign po1351 = n19127 | n19128;
  assign n19130 = pi1167 & ~pi1176;
  assign n19131 = ~pi1167 & pi1176;
  assign n19132 = ~n19130 & ~n19131;
  assign n19133 = n15326 & ~n19132;
  assign n19134 = pi1172 & ~n15326;
  assign po1352 = n19133 | n19134;
  assign n19136 = ~pi1173 & ~n16136;
  assign n19137 = n15323 & n16136;
  assign n19138 = ~n19136 & ~n19137;
  assign n19139 = n15326 & ~n19138;
  assign n19140 = ~pi1173 & ~n15326;
  assign po1353 = n19139 | n19140;
  assign n19142 = n15323 & n17437;
  assign n19143 = ~pi1174 & ~n17437;
  assign n19144 = ~n19142 & ~n19143;
  assign n19145 = n15326 & ~n19144;
  assign n19146 = ~pi1174 & ~n15326;
  assign po1354 = n19145 | n19146;
  assign n19148 = pi1167 & n15326;
  assign n19149 = pi1175 & ~n15326;
  assign po1355 = n19148 | n19149;
  assign n19151 = ~pi1176 & ~n19023;
  assign n19152 = pi1154 & pi1176;
  assign n19153 = ~n19151 & ~n19152;
  assign n19154 = ~n15333 & ~n19153;
  assign n19155 = n15326 & ~n19154;
  assign n19156 = pi1176 & ~n15326;
  assign po1356 = n19155 | n19156;
  assign n19158 = pi1828 & ~pi1984;
  assign n19159 = ~pi1828 & pi1984;
  assign n19160 = ~n19158 & ~n19159;
  assign n19161 = ~n18940 & ~n19160;
  assign n19162 = ~pi1177 & ~n11939;
  assign n19163 = ~pi1129 & pi1177;
  assign n19164 = pi1129 & ~pi1177;
  assign n19165 = ~n19163 & ~n19164;
  assign n19166 = n11939 & ~n19165;
  assign n19167 = ~n19162 & ~n19166;
  assign n19168 = n18940 & ~n19167;
  assign po1357 = n19161 | n19168;
  assign n19170 = ~pi2358 & ~n18940;
  assign n19171 = pi1178 & ~n11939;
  assign n19172 = pi1131 & ~pi1181;
  assign n19173 = ~pi1131 & pi1181;
  assign n19174 = ~n19172 & ~n19173;
  assign n19175 = n11939 & ~n19174;
  assign n19176 = ~n19171 & ~n19175;
  assign n19177 = n18940 & ~n19176;
  assign po1358 = n19170 | n19177;
  assign n19179 = pi1828 & pi1985;
  assign n19180 = pi1984 & n19179;
  assign n19181 = pi1983 & ~n19180;
  assign n19182 = ~pi1983 & n19180;
  assign n19183 = ~n19181 & ~n19182;
  assign n19184 = ~n18940 & ~n19183;
  assign n19185 = ~pi1179 & ~n11939;
  assign n19186 = ~pi1162 & n19075;
  assign n19187 = pi1179 & n19186;
  assign n19188 = ~pi1179 & ~n19186;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = n11939 & ~n19189;
  assign n19191 = ~n19185 & ~n19190;
  assign n19192 = n18940 & ~n19191;
  assign po1359 = n19184 | n19192;
  assign n19194 = ~pi1180 & ~n14364;
  assign n19195 = pi1180 & n14364;
  assign n19196 = ~n19194 & ~n19195;
  assign n19197 = pi2913 & ~n19196;
  assign n19198 = ~pi1371 & ~pi2913;
  assign po1360 = n19197 | n19198;
  assign n19200 = pi1983 & ~n18940;
  assign n19201 = ~n11958 & n18940;
  assign po1361 = n19200 | n19201;
  assign n19203 = n15323 & n15326;
  assign n19204 = pi1182 & pi1209;
  assign n19205 = ~pi1182 & ~pi1209;
  assign n19206 = ~n19204 & ~n19205;
  assign n19207 = n19203 & n19206;
  assign n19208 = ~pi1182 & ~n19203;
  assign po1362 = n19207 | n19208;
  assign n19210 = ~pi1183 & ~n18961;
  assign n19211 = ~n18162 & n18961;
  assign po1363 = n19210 | n19211;
  assign n19213 = ~pi1184 & ~n18961;
  assign n19214 = ~n18105 & n18961;
  assign po1364 = n19213 | n19214;
  assign n19216 = ~pi1185 & ~n18961;
  assign n19217 = ~n18077 & n18961;
  assign po1365 = n19216 | n19217;
  assign n19219 = ~pi1186 & ~n18961;
  assign n19220 = ~n18059 & n18961;
  assign po1366 = n19219 | n19220;
  assign n19222 = ~pi1187 & ~n18961;
  assign n19223 = ~n18068 & n18961;
  assign po1367 = n19222 | n19223;
  assign n19225 = ~pi1188 & ~n15374;
  assign n19226 = n15323 & n15374;
  assign n19227 = ~n19225 & ~n19226;
  assign n19228 = n15326 & ~n19227;
  assign n19229 = ~pi1188 & ~n15326;
  assign po1368 = n19228 | n19229;
  assign n19231 = ~pi1189 & ~n15434;
  assign n19232 = n15323 & n15434;
  assign n19233 = ~n19231 & ~n19232;
  assign n19234 = n15326 & ~n19233;
  assign n19235 = ~pi1189 & ~n15326;
  assign po1369 = n19234 | n19235;
  assign n19237 = n15323 & n16870;
  assign n19238 = ~pi1190 & ~n16870;
  assign n19239 = ~n19237 & ~n19238;
  assign n19240 = n15326 & ~n19239;
  assign n19241 = ~pi1190 & ~n15326;
  assign po1370 = n19240 | n19241;
  assign n19243 = ~pi1191 & ~n18961;
  assign n19244 = ~n18086 & n18961;
  assign po1371 = n19243 | n19244;
  assign n19246 = ~pi1192 & ~n18961;
  assign n19247 = ~n18213 & n18961;
  assign po1372 = n19246 | n19247;
  assign n19249 = ~pi1193 & ~n18961;
  assign n19250 = ~n18097 & n18961;
  assign po1373 = n19249 | n19250;
  assign n19252 = ~pi1194 & ~n19203;
  assign po1374 = n19207 | n19252;
  assign n19254 = ~pi1195 & ~n19203;
  assign n19255 = pi1195 & ~pi1209;
  assign n19256 = ~pi1182 & n19255;
  assign n19257 = ~pi1195 & pi1209;
  assign n19258 = ~n19256 & ~n19257;
  assign n19259 = pi1182 & ~pi1195;
  assign n19260 = n19258 & ~n19259;
  assign n19261 = n19203 & ~n19260;
  assign po1375 = n19254 | n19261;
  assign n19263 = ~pi1196 & ~n19203;
  assign n19264 = ~pi1182 & pi1195;
  assign n19265 = ~n19259 & ~n19264;
  assign n19266 = n19203 & ~n19265;
  assign po1376 = n19263 | n19266;
  assign n19268 = ~pi1197 & ~n15386;
  assign n19269 = n15323 & n15386;
  assign n19270 = ~n19268 & ~n19269;
  assign n19271 = n15326 & ~n19270;
  assign n19272 = ~pi1197 & ~n15326;
  assign po1377 = n19271 | n19272;
  assign n19274 = ~pi1198 & ~n15400;
  assign n19275 = n15323 & n15400;
  assign n19276 = ~n19274 & ~n19275;
  assign n19277 = n15326 & ~n19276;
  assign n19278 = ~pi1198 & ~n15326;
  assign po1378 = n19277 | n19278;
  assign n19280 = ~pi1199 & ~n15407;
  assign n19281 = n15323 & n15407;
  assign n19282 = ~n19280 & ~n19281;
  assign n19283 = n15326 & ~n19282;
  assign n19284 = ~pi1199 & ~n15326;
  assign po1379 = n19283 | n19284;
  assign n19286 = ~pi1200 & ~n15414;
  assign n19287 = n15323 & n15414;
  assign n19288 = ~n19286 & ~n19287;
  assign n19289 = n15326 & ~n19288;
  assign n19290 = ~pi1200 & ~n15326;
  assign po1380 = n19289 | n19290;
  assign n19292 = ~pi1201 & ~n15427;
  assign n19293 = n15323 & n15427;
  assign n19294 = ~n19292 & ~n19293;
  assign n19295 = n15326 & ~n19294;
  assign n19296 = ~pi1201 & ~n15326;
  assign po1381 = n19295 | n19296;
  assign n19298 = n15323 & n17015;
  assign n19299 = ~pi1202 & ~n17015;
  assign n19300 = ~n19298 & ~n19299;
  assign n19301 = n15326 & ~n19300;
  assign n19302 = ~pi1202 & ~n15326;
  assign po1382 = n19301 | n19302;
  assign n19304 = n15323 & n17154;
  assign n19305 = ~pi1203 & ~n17154;
  assign n19306 = ~n19304 & ~n19305;
  assign n19307 = n15326 & ~n19306;
  assign n19308 = ~pi1203 & ~n15326;
  assign po1383 = n19307 | n19308;
  assign n19310 = ~pi1204 & ~n15393;
  assign n19311 = n15323 & n15393;
  assign n19312 = ~n19310 & ~n19311;
  assign n19313 = n15326 & ~n19312;
  assign n19314 = ~pi1204 & ~n15326;
  assign po1384 = n19313 | n19314;
  assign n19316 = n15312 & n15323;
  assign n19317 = ~pi1205 & ~n15312;
  assign n19318 = ~n19316 & ~n19317;
  assign n19319 = n15326 & ~n19318;
  assign n19320 = ~pi1205 & ~n15326;
  assign po1385 = n19319 | n19320;
  assign n19322 = ~pi1206 & ~n15335;
  assign n19323 = n15323 & n15335;
  assign n19324 = ~n19322 & ~n19323;
  assign n19325 = n15326 & ~n19324;
  assign n19326 = ~pi1206 & ~n15326;
  assign po1386 = n19325 | n19326;
  assign n19328 = ~pi1207 & ~n16635;
  assign n19329 = n15323 & n16635;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = n15326 & ~n19330;
  assign n19332 = ~pi1207 & ~n15326;
  assign po1387 = n19331 | n19332;
  assign n19334 = ~pi1208 & ~n19203;
  assign n19335 = ~pi1195 & n19203;
  assign po1388 = n19334 | n19335;
  assign n19337 = ~pi1209 & ~n19203;
  assign n19338 = pi1209 & n19203;
  assign po1389 = n19337 | n19338;
  assign n19340 = ~pi1210 & ~n14907;
  assign n19341 = pi1210 & ~pi3362;
  assign po1390 = n19340 | n19341;
  assign n19343 = ~pi1367 & pi1407;
  assign n19344 = ~pi1371 & pi1407;
  assign n19345 = ~n19343 & ~n19344;
  assign n19346 = pi1367 & pi1371;
  assign n19347 = ~pi1407 & n19346;
  assign n19348 = n19345 & ~n19347;
  assign n19349 = ~pi2913 & ~n19348;
  assign n19350 = ~pi1180 & pi1224;
  assign n19351 = pi1211 & n19350;
  assign n19352 = ~pi1211 & ~n19350;
  assign n19353 = ~n19351 & ~n19352;
  assign n19354 = n14364 & ~n19353;
  assign n19355 = ~pi1211 & ~n14364;
  assign n19356 = ~n19354 & ~n19355;
  assign n19357 = pi2913 & ~n19356;
  assign po1391 = n19349 | n19357;
  assign n19359 = pi1367 & ~pi2913;
  assign n19360 = pi2913 & ~n14373;
  assign po1392 = n19359 | n19360;
  assign n19362 = pi1407 & ~pi2913;
  assign n19363 = pi2913 & ~n14370;
  assign po1393 = n19362 | n19363;
  assign n19365 = ~pi1408 & ~pi2913;
  assign n19366 = ~pi1216 & n14364;
  assign n19367 = pi1214 & ~n14364;
  assign n19368 = ~n19366 & ~n19367;
  assign n19369 = pi2913 & ~n19368;
  assign po1394 = n19365 | n19369;
  assign n19371 = ~pi1383 & ~pi2913;
  assign n19372 = ~pi1217 & n14364;
  assign n19373 = pi1215 & ~n14364;
  assign n19374 = ~n19372 & ~n19373;
  assign n19375 = pi2913 & ~n19374;
  assign po1395 = n19371 | n19375;
  assign n19377 = pi1375 & ~pi2913;
  assign n19378 = pi1212 & ~pi1221;
  assign n19379 = ~pi1212 & pi1221;
  assign n19380 = ~n19378 & ~n19379;
  assign n19381 = n14364 & ~n19380;
  assign n19382 = ~pi1216 & ~n14364;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = pi2913 & ~n19383;
  assign po1396 = n19377 | n19384;
  assign n19386 = pi1369 & ~pi2913;
  assign n19387 = pi1212 & ~pi1213;
  assign n19388 = ~pi1212 & pi1213;
  assign n19389 = ~n19387 & ~n19388;
  assign n19390 = n14364 & ~n19389;
  assign n19391 = ~pi1217 & ~n14364;
  assign n19392 = ~n19390 & ~n19391;
  assign n19393 = pi2913 & ~n19392;
  assign po1397 = n19386 | n19393;
  assign n19395 = pi1218 & ~n18961;
  assign n19396 = pi1680 & pi1681;
  assign n19397 = n18961 & ~n19396;
  assign n19398 = pi2465 & ~pi2960;
  assign n19399 = pi3125 & n19398;
  assign n19400 = n19397 & n19399;
  assign po1398 = n19395 | n19400;
  assign n19402 = pi3117 & ~pi3120;
  assign n19403 = pi3042 & pi3124;
  assign n19404 = n19402 & ~n19403;
  assign n19405 = ~po3257 & ~po3302;
  assign n19406 = ~n19404 & ~n19405;
  assign po1405 = n19051 & ~n19406;
  assign n19408 = pi1371 & ~pi2913;
  assign n19409 = pi2913 & ~n14367;
  assign po1401 = n19408 | n19409;
  assign n19411 = ~pi1409 & ~pi2913;
  assign n19412 = ~pi1223 & n14364;
  assign n19413 = pi1222 & ~n14364;
  assign n19414 = ~n19412 & ~n19413;
  assign n19415 = pi2913 & ~n19414;
  assign po1402 = n19411 | n19415;
  assign n19417 = pi1410 & ~pi2913;
  assign n19418 = ~pi1213 & n14364;
  assign n19419 = ~pi1223 & ~n14364;
  assign n19420 = ~n19418 & ~n19419;
  assign n19421 = pi2913 & ~n19420;
  assign po1403 = n19417 | n19421;
  assign n19423 = ~pi1367 & pi1371;
  assign n19424 = pi1367 & ~pi1371;
  assign n19425 = ~n19423 & ~n19424;
  assign n19426 = ~pi2913 & ~n19425;
  assign n19427 = pi1180 & pi1224;
  assign n19428 = ~pi1180 & ~pi1224;
  assign n19429 = ~n19427 & ~n19428;
  assign n19430 = n14364 & ~n19429;
  assign n19431 = pi1224 & ~n14364;
  assign n19432 = ~n19430 & ~n19431;
  assign n19433 = pi2913 & ~n19432;
  assign po1404 = n19426 | n19433;
  assign n19435 = pi1228 & pi1376;
  assign n19436 = ~pi3365 & n19435;
  assign n19437 = pi1376 & ~n7075;
  assign n19438 = pi3365 & n19437;
  assign n19439 = ~pi1228 & n19438;
  assign po1406 = n19436 | n19439;
  assign n19441 = pi1229 & ~n13171;
  assign n19442 = ~pi1229 & n13171;
  assign po1407 = n19441 | n19442;
  assign n19444 = ~pi1762 & n18961;
  assign n19445 = ~pi1680 & n19444;
  assign n19446 = pi2465 & n19445;
  assign n19447 = ~pi1230 & ~n18961;
  assign po1408 = n19446 | n19447;
  assign n19449 = n9391 & ~n15368;
  assign n19450 = ~n9382 & ~n19449;
  assign n19451 = ~pi3027 & n19450;
  assign n19452 = ~n9380 & n19451;
  assign n19453 = ~pi0444 & n9404;
  assign n19454 = pi1692 & ~n9404;
  assign n19455 = ~n19453 & ~n19454;
  assign n19456 = pi1858 & ~n19455;
  assign n19457 = ~pi1218 & pi1337;
  assign n19458 = ~n19456 & ~n19457;
  assign n19459 = pi1337 & pi2519;
  assign n19460 = n19458 & ~n19459;
  assign n19461 = ~pi2911 & n19460;
  assign n19462 = n9391 & ~n19461;
  assign n19463 = ~n15367 & ~n19462;
  assign n19464 = ~pi2461 & ~pi2526;
  assign n19465 = ~pi1971 & n19464;
  assign n19466 = ~pi1972 & ~pi2252;
  assign n19467 = ~pi2463 & n19466;
  assign n19468 = ~pi2757 & n19467;
  assign n19469 = n19465 & n19468;
  assign n19470 = pi3369 & n19469;
  assign n19471 = ~pi3027 & ~n19470;
  assign n19472 = ~pi1805 & n19471;
  assign n19473 = n19463 & n19472;
  assign n19474 = ~n19452 & ~n19473;
  assign n19475 = ~n9382 & n19474;
  assign n19476 = pi1232 & n19452;
  assign po1410 = n19475 | n19476;
  assign n19478 = pi3365 & n7075;
  assign n19479 = pi1238 & pi1257;
  assign n19480 = pi1237 & n19479;
  assign n19481 = pi1228 & pi1236;
  assign n19482 = n19480 & n19481;
  assign n19483 = pi1233 & ~n19482;
  assign n19484 = ~pi1233 & n19482;
  assign n19485 = ~n19483 & ~n19484;
  assign n19486 = pi3365 & ~n19485;
  assign n19487 = ~n19478 & ~n19486;
  assign n19488 = pi1233 & ~pi3365;
  assign n19489 = n19487 & ~n19488;
  assign po1411 = pi1376 & ~n19489;
  assign n19491 = n7071 & n19481;
  assign n19492 = pi1238 & n19491;
  assign n19493 = pi1233 & n19492;
  assign n19494 = pi1234 & ~n19493;
  assign n19495 = ~pi1234 & n19493;
  assign n19496 = ~n19494 & ~n19495;
  assign n19497 = pi3365 & ~n19496;
  assign n19498 = ~n19478 & ~n19497;
  assign n19499 = pi1234 & ~pi3365;
  assign n19500 = n19498 & ~n19499;
  assign po1412 = pi1376 & ~n19500;
  assign n19502 = ~pi1235 & ~n18961;
  assign po1413 = n19444 | n19502;
  assign n19504 = pi1228 & ~pi1236;
  assign n19505 = ~n7072 & ~n19504;
  assign n19506 = pi3365 & ~n19505;
  assign n19507 = pi1236 & ~pi3365;
  assign n19508 = ~n19506 & ~n19507;
  assign n19509 = ~n19478 & n19508;
  assign po1414 = pi1376 & ~n19509;
  assign n19511 = pi1237 & ~pi3365;
  assign n19512 = pi1237 & ~n19481;
  assign n19513 = ~pi1237 & n19481;
  assign n19514 = ~n19512 & ~n19513;
  assign n19515 = pi3365 & ~n19514;
  assign n19516 = ~n19478 & ~n19515;
  assign n19517 = ~n19511 & n19516;
  assign po1415 = pi1376 & ~n19517;
  assign n19519 = pi1238 & ~pi3365;
  assign n19520 = pi1237 & n19481;
  assign n19521 = pi1257 & n19520;
  assign n19522 = pi1238 & ~n19521;
  assign n19523 = ~pi1238 & n19521;
  assign n19524 = ~n19522 & ~n19523;
  assign n19525 = pi3365 & ~n19524;
  assign n19526 = ~n19478 & ~n19525;
  assign n19527 = ~n19519 & n19526;
  assign po1416 = pi1376 & ~n19527;
  assign n19529 = ~n11155 & n13169;
  assign n19530 = ~pi0444 & ~n19529;
  assign n19531 = pi1239 & ~n19530;
  assign n19532 = pi1266 & pi1305;
  assign n19533 = ~pi1266 & ~pi1305;
  assign n19534 = ~n19532 & ~n19533;
  assign n19535 = n19530 & n19534;
  assign po1417 = n19531 | n19535;
  assign n19537 = pi1229 & pi1242;
  assign n19538 = pi1240 & ~n19537;
  assign n19539 = ~pi1240 & n19537;
  assign n19540 = ~n19538 & ~n19539;
  assign n19541 = n13171 & ~n19540;
  assign n19542 = pi1240 & ~n13171;
  assign po1418 = n19541 | n19542;
  assign n19544 = pi1240 & n19537;
  assign n19545 = pi1241 & ~n19544;
  assign n19546 = ~pi1241 & n19544;
  assign n19547 = ~n19545 & ~n19546;
  assign n19548 = n13171 & ~n19547;
  assign n19549 = pi1241 & ~n13171;
  assign po1419 = n19548 | n19549;
  assign n19551 = pi1229 & ~pi1242;
  assign n19552 = ~pi1229 & pi1242;
  assign n19553 = ~n19551 & ~n19552;
  assign n19554 = n13171 & ~n19553;
  assign n19555 = pi1242 & ~n13171;
  assign po1420 = n19554 | n19555;
  assign n19557 = pi1250 & n13171;
  assign n19558 = ~pi1244 & ~n13171;
  assign po1422 = n19557 | n19558;
  assign n19560 = pi1254 & n13171;
  assign n19561 = ~pi1245 & ~n13171;
  assign po1423 = n19560 | n19561;
  assign n19563 = pi1251 & n13171;
  assign n19564 = ~pi1246 & ~n13171;
  assign po1424 = n19563 | n19564;
  assign n19566 = ~pi1244 & n13171;
  assign n19567 = ~pi1247 & ~n13171;
  assign po1425 = n19566 | n19567;
  assign n19569 = ~pi1245 & n13171;
  assign n19570 = ~pi1248 & ~n13171;
  assign po1426 = n19569 | n19570;
  assign n19572 = ~pi1246 & n13171;
  assign n19573 = ~pi1249 & ~n13171;
  assign po1427 = n19572 | n19573;
  assign n19575 = pi1231 & ~pi1267;
  assign n19576 = ~pi1231 & pi1267;
  assign n19577 = ~n19575 & ~n19576;
  assign n19578 = n13171 & ~n19577;
  assign n19579 = pi1250 & ~n13171;
  assign po1428 = n19578 | n19579;
  assign n19581 = ~pi1243 & pi1256;
  assign n19582 = pi1243 & ~pi1256;
  assign n19583 = ~n19581 & ~n19582;
  assign n19584 = n13171 & ~n19583;
  assign n19585 = pi1251 & ~n13171;
  assign po1429 = n19584 | n19585;
  assign n19587 = pi1256 & n13171;
  assign n19588 = pi1252 & ~n13171;
  assign po1430 = n19587 | n19588;
  assign n19590 = ~pi1255 & n13171;
  assign n19591 = ~pi1253 & ~n13171;
  assign po1431 = n19590 | n19591;
  assign n19593 = pi1243 & ~pi1267;
  assign n19594 = ~pi1243 & pi1267;
  assign n19595 = ~n19593 & ~n19594;
  assign n19596 = n13171 & ~n19595;
  assign n19597 = pi1254 & ~n13171;
  assign po1432 = n19596 | n19597;
  assign n19599 = pi1252 & n13171;
  assign n19600 = ~pi1255 & ~n13171;
  assign po1433 = n19599 | n19600;
  assign n19602 = pi1257 & ~pi3365;
  assign n19603 = pi1257 & ~n19520;
  assign n19604 = ~pi1257 & n19520;
  assign n19605 = ~n19603 & ~n19604;
  assign n19606 = pi3365 & ~n19605;
  assign n19607 = ~n19478 & ~n19606;
  assign n19608 = ~n19602 & n19607;
  assign po1435 = pi1376 & ~n19608;
  assign n19610 = n19479 & n19520;
  assign n19611 = pi1233 & n19610;
  assign n19612 = pi1234 & n19611;
  assign n19613 = pi1258 & ~n19612;
  assign n19614 = ~pi1258 & n19612;
  assign n19615 = ~n19613 & ~n19614;
  assign n19616 = pi3365 & ~n19615;
  assign n19617 = ~n19478 & ~n19616;
  assign n19618 = pi1258 & ~pi3365;
  assign n19619 = n19617 & ~n19618;
  assign po1436 = pi1376 & ~n19619;
  assign n19621 = pi1259 & n19452;
  assign po1437 = n19475 | n19621;
  assign n19623 = ~pi3123 & n8009;
  assign n19624 = ~n9089 & n19623;
  assign n19625 = ~po3339 & n19624;
  assign n19626 = ~pi1260 & ~n8009;
  assign po1438 = n19625 | n19626;
  assign n19628 = pi1261 & ~n8009;
  assign n19629 = n9089 & ~po3339;
  assign n19630 = n8009 & n19629;
  assign n19631 = ~n19628 & ~n19630;
  assign n19632 = n11154 & po3339;
  assign n19633 = n8009 & n19632;
  assign n19634 = ~pi1858 & n19633;
  assign po1439 = ~n19631 | n19634;
  assign n19636 = pi1262 & ~n18961;
  assign n19637 = pi2955 & n18961;
  assign po1440 = n19636 | n19637;
  assign n19639 = pi1263 & ~n18961;
  assign n19640 = pi2958 & n18961;
  assign po1441 = n19639 | n19640;
  assign n19642 = pi1264 & ~n18961;
  assign n19643 = pi2952 & n18961;
  assign po1442 = n19642 | n19643;
  assign n19645 = ~pi1265 & ~n18961;
  assign n19646 = pi2960 & n18961;
  assign po1443 = n19645 | n19646;
  assign n19648 = ~pi1266 & ~n19530;
  assign po1444 = n19535 | n19648;
  assign n19650 = pi1268 & ~n18961;
  assign n19651 = pi2959 & n18961;
  assign po1446 = n19650 | n19651;
  assign n19653 = ~pi1269 & ~n18961;
  assign n19654 = ~pi1680 & ~pi1762;
  assign n19655 = pi2465 & n19654;
  assign n19656 = ~pi1681 & n19655;
  assign n19657 = n18961 & ~n19656;
  assign po1447 = n19653 | n19657;
  assign n19659 = ~pi1303 & ~pi1330;
  assign n19660 = pi1302 & pi1313;
  assign n19661 = pi1296 & pi1300;
  assign n19662 = pi1316 & n19661;
  assign n19663 = pi1301 & n19662;
  assign n19664 = pi1314 & n19663;
  assign n19665 = pi1304 & n19664;
  assign n19666 = n19660 & n19665;
  assign n19667 = ~pi1297 & n19666;
  assign n19668 = ~pi1298 & n19667;
  assign n19669 = n19659 & n19668;
  assign n19670 = ~pi1270 & n19669;
  assign n19671 = pi1270 & ~n19669;
  assign n19672 = ~n19670 & ~n19671;
  assign n19673 = pi1318 & n18959;
  assign n19674 = ~n11950 & n19673;
  assign n19675 = ~n8229 & n19674;
  assign po1448 = n19672 & n19675;
  assign n19677 = pi1271 & ~n8009;
  assign n19678 = pi1338 & ~n9089;
  assign n19679 = n8009 & n19678;
  assign po1449 = n19677 | n19679;
  assign n19681 = ~n10999 & ~n15322;
  assign n19682 = ~pi1272 & n19681;
  assign n19683 = ~pi1899 & ~n19681;
  assign po1450 = n19682 | n19683;
  assign n19685 = ~pi1273 & n19681;
  assign n19686 = ~pi1900 & ~n19681;
  assign po1451 = n19685 | n19686;
  assign n19688 = ~pi1274 & n19681;
  assign n19689 = ~pi1898 & ~n19681;
  assign po1452 = n19688 | n19689;
  assign n19691 = ~pi1275 & n19681;
  assign n19692 = ~pi1885 & ~n19681;
  assign po1453 = n19691 | n19692;
  assign n19694 = ~pi1276 & n19681;
  assign n19695 = ~pi1876 & ~n19681;
  assign po1454 = n19694 | n19695;
  assign n19697 = ~pi1277 & n19681;
  assign n19698 = ~pi1886 & ~n19681;
  assign po1455 = n19697 | n19698;
  assign n19700 = ~pi1278 & n19681;
  assign n19701 = ~pi1861 & ~n19681;
  assign po1456 = n19700 | n19701;
  assign n19703 = ~pi1279 & n19681;
  assign n19704 = ~pi1893 & ~n19681;
  assign po1457 = n19703 | n19704;
  assign n19706 = ~pi1280 & n19681;
  assign n19707 = ~pi1895 & ~n19681;
  assign po1458 = n19706 | n19707;
  assign n19709 = ~pi1281 & n19681;
  assign n19710 = ~pi1894 & ~n19681;
  assign po1459 = n19709 | n19710;
  assign n19712 = ~pi1282 & n19681;
  assign n19713 = ~pi1865 & ~n19681;
  assign po1460 = n19712 | n19713;
  assign n19715 = ~pi1283 & n19681;
  assign n19716 = ~pi1897 & ~n19681;
  assign po1461 = n19715 | n19716;
  assign n19718 = ~pi1284 & n19681;
  assign n19719 = ~pi1891 & ~n19681;
  assign po1462 = n19718 | n19719;
  assign n19721 = ~pi1285 & n19681;
  assign n19722 = ~pi1860 & ~n19681;
  assign po1463 = n19721 | n19722;
  assign n19724 = ~pi1286 & n19681;
  assign n19725 = ~pi1868 & ~n19681;
  assign po1464 = n19724 | n19725;
  assign n19727 = ~pi1287 & n19681;
  assign n19728 = ~pi1869 & ~n19681;
  assign po1465 = n19727 | n19728;
  assign n19730 = ~pi1288 & n19681;
  assign n19731 = ~pi1892 & ~n19681;
  assign po1466 = n19730 | n19731;
  assign n19733 = ~pi1289 & n19681;
  assign n19734 = pi2955 & ~n19681;
  assign po1467 = n19733 | n19734;
  assign n19736 = ~pi1290 & n19681;
  assign n19737 = pi2958 & ~n19681;
  assign po1468 = n19736 | n19737;
  assign n19739 = ~pi1291 & n19681;
  assign n19740 = pi2952 & ~n19681;
  assign po1469 = n19739 | n19740;
  assign n19742 = ~pi1292 & n19681;
  assign n19743 = ~pi1871 & ~n19681;
  assign po1470 = n19742 | n19743;
  assign n19745 = ~pi1293 & n19681;
  assign n19746 = ~pi1888 & ~n19681;
  assign po1471 = n19745 | n19746;
  assign n19748 = ~pi1294 & n19681;
  assign n19749 = ~pi1874 & ~n19681;
  assign po1472 = n19748 | n19749;
  assign n19751 = ~pi1295 & n19681;
  assign n19752 = ~pi1889 & ~n19681;
  assign po1473 = n19751 | n19752;
  assign po1474 = ~pi1296 & n19675;
  assign n19755 = pi1304 & n19659;
  assign n19756 = pi1313 & n19755;
  assign n19757 = pi1301 & pi1314;
  assign n19758 = n19661 & n19757;
  assign n19759 = pi1302 & n19758;
  assign n19760 = pi1316 & n19759;
  assign n19761 = n19756 & n19760;
  assign n19762 = pi1297 & ~n19761;
  assign n19763 = ~pi1297 & n19761;
  assign n19764 = ~n19762 & ~n19763;
  assign po1475 = n19675 & n19764;
  assign n19766 = ~pi1297 & n19755;
  assign n19767 = n19660 & n19662;
  assign n19768 = n19757 & n19767;
  assign n19769 = n19766 & n19768;
  assign n19770 = ~pi1298 & n19769;
  assign n19771 = pi1298 & ~n19769;
  assign n19772 = ~n19770 & ~n19771;
  assign po1476 = n19675 & n19772;
  assign n19774 = ~pi1270 & ~pi1315;
  assign n19775 = n19763 & n19774;
  assign n19776 = ~pi1298 & n19775;
  assign n19777 = ~pi1299 & n19776;
  assign n19778 = pi1299 & ~n19776;
  assign n19779 = ~n19777 & ~n19778;
  assign po1477 = n19675 & n19779;
  assign n19781 = ~pi1296 & ~pi1300;
  assign n19782 = ~n19661 & ~n19781;
  assign po1478 = n19675 & n19782;
  assign n19784 = ~pi1301 & ~n19662;
  assign n19785 = ~n19663 & ~n19784;
  assign po1479 = n19675 & n19785;
  assign n19787 = pi1300 & n19757;
  assign n19788 = pi1296 & n19787;
  assign n19789 = pi1316 & n19788;
  assign n19790 = pi1302 & n19789;
  assign n19791 = ~pi1302 & ~n19789;
  assign n19792 = ~n19790 & ~n19791;
  assign po1480 = n19675 & n19792;
  assign n19794 = pi1304 & n19660;
  assign n19795 = ~pi1330 & n19794;
  assign n19796 = n19789 & n19795;
  assign n19797 = ~pi1303 & n19796;
  assign n19798 = pi1303 & ~n19796;
  assign n19799 = ~n19797 & ~n19798;
  assign po1481 = n19675 & n19799;
  assign n19801 = pi1304 & n19768;
  assign n19802 = ~pi1304 & ~n19768;
  assign n19803 = ~n19801 & ~n19802;
  assign po1482 = n19675 & n19803;
  assign n19805 = ~pi1305 & ~n19530;
  assign n19806 = pi1305 & n19530;
  assign po1483 = n19805 | n19806;
  assign n19808 = pi1307 & ~n19530;
  assign n19809 = ~pi1311 & n19530;
  assign po1485 = n19808 | n19809;
  assign n19811 = ~pi1308 & n19681;
  assign n19812 = ~pi1873 & ~n19681;
  assign po1486 = n19811 | n19812;
  assign n19814 = pi1309 & ~n19530;
  assign n19815 = pi1266 & ~pi1311;
  assign n19816 = ~pi1266 & pi1311;
  assign n19817 = ~n19815 & ~n19816;
  assign n19818 = n19530 & ~n19817;
  assign po1487 = n19814 | n19818;
  assign po1488 = ~pi1310 & ~n18961;
  assign n19821 = ~pi1311 & ~n19530;
  assign n19822 = ~pi1305 & pi1311;
  assign n19823 = ~pi1266 & n19822;
  assign n19824 = pi1305 & ~pi1311;
  assign n19825 = ~n19823 & ~n19824;
  assign n19826 = ~n19815 & n19825;
  assign n19827 = n19530 & ~n19826;
  assign po1489 = n19821 | n19827;
  assign n19829 = ~pi1312 & ~n14891;
  assign n19830 = pi1312 & ~pi3362;
  assign po1490 = n19829 | n19830;
  assign n19832 = pi1313 & n19760;
  assign n19833 = ~pi1313 & ~n19760;
  assign n19834 = ~n19832 & ~n19833;
  assign po1491 = n19675 & n19834;
  assign n19836 = ~pi1314 & ~n19663;
  assign n19837 = ~n19664 & ~n19836;
  assign po1492 = n19675 & n19837;
  assign n19839 = ~pi1270 & ~pi1298;
  assign n19840 = n19796 & n19839;
  assign n19841 = ~pi1303 & n19840;
  assign n19842 = ~pi1297 & n19841;
  assign n19843 = ~pi1315 & n19842;
  assign n19844 = pi1315 & ~n19842;
  assign n19845 = ~n19843 & ~n19844;
  assign po1493 = n19675 & n19845;
  assign n19847 = ~pi1316 & ~n19661;
  assign n19848 = ~n19662 & ~n19847;
  assign po1494 = n19675 & n19848;
  assign n19850 = n19769 & n19839;
  assign n19851 = ~pi1299 & n19850;
  assign n19852 = ~pi1315 & n19851;
  assign n19853 = ~pi1317 & n19852;
  assign n19854 = pi1317 & ~n19852;
  assign n19855 = ~n19853 & ~n19854;
  assign po1495 = n19675 & n19855;
  assign n19857 = n19669 & n19774;
  assign n19858 = ~pi1299 & n19857;
  assign n19859 = ~pi1317 & n19858;
  assign n19860 = ~pi1318 & n19859;
  assign n19861 = pi1318 & ~n19859;
  assign n19862 = ~n19860 & ~n19861;
  assign po1496 = n19675 & n19862;
  assign n19864 = ~pi1319 & n19681;
  assign n19865 = ~pi1887 & ~n19681;
  assign po1497 = n19864 | n19865;
  assign n19867 = ~pi1320 & n19681;
  assign n19868 = ~pi1872 & ~n19681;
  assign po1498 = n19867 | n19868;
  assign n19870 = ~pi1321 & n19681;
  assign n19871 = pi2959 & ~n19681;
  assign po1499 = n19870 | n19871;
  assign n19873 = ~pi1322 & n19681;
  assign n19874 = ~pi1870 & ~n19681;
  assign po1500 = n19873 | n19874;
  assign n19876 = ~pi1323 & n19681;
  assign n19877 = ~pi1864 & ~n19681;
  assign po1501 = n19876 | n19877;
  assign n19879 = ~pi1324 & n19681;
  assign n19880 = ~pi1867 & ~n19681;
  assign po1502 = n19879 | n19880;
  assign n19882 = ~pi1325 & n19681;
  assign n19883 = ~pi1866 & ~n19681;
  assign po1503 = n19882 | n19883;
  assign n19885 = ~pi1326 & n19681;
  assign n19886 = ~pi1875 & ~n19681;
  assign po1504 = n19885 | n19886;
  assign n19888 = ~pi1327 & n19681;
  assign n19889 = ~pi1863 & ~n19681;
  assign po1505 = n19888 | n19889;
  assign n19891 = ~pi1328 & n19681;
  assign n19892 = ~pi1896 & ~n19681;
  assign po1506 = n19891 | n19892;
  assign n19894 = ~pi1329 & n19681;
  assign n19895 = ~pi1862 & ~n19681;
  assign po1507 = n19894 | n19895;
  assign n19897 = ~pi1330 & n19666;
  assign n19898 = pi1330 & ~n19666;
  assign n19899 = ~n19897 & ~n19898;
  assign po1508 = n19675 & n19899;
  assign n19901 = pi3123 & ~po3339;
  assign n19902 = ~n8119 & ~n19901;
  assign n19903 = pi1374 & n8009;
  assign n19904 = n8143 & n19903;
  assign n19905 = ~n8090 & n19904;
  assign n19906 = n19902 & n19905;
  assign n19907 = n8009 & n9089;
  assign n19908 = pi1331 & ~n8009;
  assign n19909 = ~n19907 & ~n19908;
  assign po1509 = n19906 | ~n19909;
  assign n19911 = pi1332 & n18004;
  assign n19912 = ~n7060 & ~n8003;
  assign po1510 = n19911 | n19912;
  assign n19914 = pi2966 & pi2995;
  assign n19915 = ~pi2982 & ~pi3001;
  assign n19916 = pi2981 & ~pi2997;
  assign n19917 = pi2996 & n19916;
  assign n19918 = n19915 & n19917;
  assign n19919 = n19914 & n19918;
  assign n19920 = n7254 & n19919;
  assign n19921 = pi2920 & n19920;
  assign n19922 = ~pi3018 & n19921;
  assign n19923 = pi1333 & ~n19922;
  assign n19924 = n9530 & n19921;
  assign po1511 = n19923 | n19924;
  assign n19926 = pi2966 & ~pi2995;
  assign n19927 = n19918 & n19926;
  assign n19928 = n7254 & n19927;
  assign n19929 = pi2920 & n19928;
  assign n19930 = ~pi3018 & n19929;
  assign n19931 = pi1334 & ~n19930;
  assign n19932 = n9530 & n19929;
  assign po1512 = n19931 | n19932;
  assign n19934 = pi1335 & ~n8009;
  assign po1513 = n19907 | n19934;
  assign n19936 = ~pi0443 & n9404;
  assign n19937 = ~pi1693 & ~n9404;
  assign n19938 = ~n19936 & ~n19937;
  assign n19939 = ~pi1337 & ~n19938;
  assign n19940 = ~pi0443 & ~pi2486;
  assign n19941 = ~pi1218 & ~pi1263;
  assign n19942 = pi2486 & n19941;
  assign n19943 = ~n19940 & ~n19942;
  assign n19944 = pi1337 & ~n19943;
  assign n19945 = ~n19939 & ~n19944;
  assign n19946 = pi1676 & ~n19945;
  assign n19947 = pi1683 & n9409;
  assign n19948 = ~n19946 & ~n19947;
  assign n19949 = pi1902 & n9411;
  assign n19950 = n19948 & ~n19949;
  assign n19951 = ~n9399 & ~n19950;
  assign n19952 = pi1336 & n9399;
  assign po1514 = n19951 | n19952;
  assign n19954 = pi3118 & ~pi3124;
  assign n19955 = pi3027 & ~pi3201;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = ~n9403 & n19956;
  assign n19958 = n9402 & ~n19957;
  assign n19959 = pi2911 & n19958;
  assign n19960 = ~pi2975 & ~n19954;
  assign n19961 = pi3124 & n15360;
  assign n19962 = pi2944 & n19961;
  assign n19963 = pi2924 & n19962;
  assign n19964 = ~pi3118 & ~pi3124;
  assign n19965 = pi2944 & n19964;
  assign n19966 = ~n19955 & ~n19965;
  assign n19967 = ~n19963 & n19966;
  assign n19968 = n19960 & n19967;
  assign n19969 = n9402 & ~n19968;
  assign n19970 = pi1337 & n9402;
  assign n19971 = n19969 & n19970;
  assign n19972 = ~n19959 & ~n19971;
  assign n19973 = ~pi1750 & n11154;
  assign n19974 = ~pi1827 & n19973;
  assign n19975 = pi1265 & n19974;
  assign n19976 = n19972 & n19975;
  assign n19977 = n10977 & n19976;
  assign n19978 = pi1337 & n19960;
  assign n19979 = n19967 & n19978;
  assign n19980 = pi1337 & ~n9402;
  assign n19981 = ~n19979 & ~n19980;
  assign po1515 = n19977 | ~n19981;
  assign n19983 = ~pi2996 & n19916;
  assign n19984 = n19915 & n19983;
  assign n19985 = ~pi2966 & pi2995;
  assign n19986 = ~pi2920 & n19985;
  assign n19987 = n7254 & n19986;
  assign n19988 = n19984 & n19987;
  assign n19989 = ~pi2972 & n19988;
  assign n19990 = pi1338 & ~n19989;
  assign n19991 = ~pi2972 & pi3163;
  assign n19992 = n19988 & n19991;
  assign po1516 = n19990 | n19992;
  assign n19994 = pi1339 & ~n19989;
  assign n19995 = ~pi2972 & pi3166;
  assign n19996 = n19988 & n19995;
  assign po1517 = n19994 | n19996;
  assign n19998 = n19918 & n19985;
  assign n19999 = ~pi2920 & n19998;
  assign n20000 = n7254 & n19999;
  assign n20001 = ~pi3018 & n20000;
  assign n20002 = pi1340 & ~n20001;
  assign n20003 = n9530 & n20000;
  assign po1518 = n20002 | n20003;
  assign n20005 = pi2982 & ~pi3001;
  assign n20006 = n7246 & n19917;
  assign n20007 = pi2995 & n20006;
  assign n20008 = n20005 & n20007;
  assign n20009 = n7254 & n20008;
  assign n20010 = ~pi2972 & n20009;
  assign n20011 = pi1341 & ~n20010;
  assign n20012 = ~pi2972 & pi3136;
  assign n20013 = n20009 & n20012;
  assign po1519 = n20011 | n20013;
  assign n20015 = ~pi2920 & ~pi2966;
  assign n20016 = ~pi2982 & pi3001;
  assign n20017 = ~pi2995 & n20016;
  assign n20018 = n7254 & n20017;
  assign n20019 = n19917 & n20018;
  assign n20020 = n20015 & n20019;
  assign n20021 = ~pi3018 & n20020;
  assign n20022 = pi1342 & ~n20021;
  assign n20023 = n9530 & n20020;
  assign po1520 = n20022 | n20023;
  assign n20025 = pi1343 & n9386;
  assign n20026 = ~n9386 & ~n19950;
  assign po1521 = n20025 | n20026;
  assign n20028 = ~pi0120 & pi0126;
  assign n20029 = ~pi0128 & pi1220;
  assign n20030 = n20028 & n20029;
  assign n20031 = po3257 & ~n20030;
  assign n20032 = ~n9245 & ~n20031;
  assign n20033 = n8889 & ~n20032;
  assign n20034 = ~pi1260 & n20033;
  assign po1522 = ~pi2984 & n20034;
  assign n20036 = ~pi1969 & n8194;
  assign n20037 = n8197 & ~n20036;
  assign n20038 = ~n8197 & ~n8296;
  assign po1523 = n20037 | n20038;
  assign n20040 = ~pi1878 & pi3511;
  assign n20041 = pi1336 & pi1878;
  assign n20042 = ~n20040 & ~n20041;
  assign n20043 = ~pi1878 & pi3510;
  assign n20044 = pi0135 & pi1878;
  assign n20045 = ~n20043 & ~n20044;
  assign n20046 = ~n20042 & n20045;
  assign n20047 = n20042 & ~n20045;
  assign n20048 = ~n20046 & ~n20047;
  assign n20049 = ~pi1878 & pi3513;
  assign n20050 = pi0136 & pi1878;
  assign n20051 = ~n20049 & ~n20050;
  assign n20052 = ~pi1878 & pi3512;
  assign n20053 = pi0139 & pi1878;
  assign n20054 = ~n20052 & ~n20053;
  assign n20055 = ~n20051 & n20054;
  assign n20056 = n20051 & ~n20054;
  assign n20057 = ~n20055 & ~n20056;
  assign n20058 = pi0144 & ~pi0198;
  assign n20059 = ~pi0144 & pi0198;
  assign n20060 = ~n20058 & ~n20059;
  assign n20061 = ~pi0143 & pi0203;
  assign n20062 = pi0143 & ~pi0203;
  assign n20063 = ~n20061 & ~n20062;
  assign n20064 = ~n20060 & n20063;
  assign n20065 = n20060 & ~n20063;
  assign n20066 = ~n20064 & ~n20065;
  assign n20067 = ~pi0145 & pi0146;
  assign n20068 = pi0145 & ~pi0146;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = pi0130 & ~pi0192;
  assign n20071 = ~pi0130 & pi0192;
  assign n20072 = ~n20070 & ~n20071;
  assign n20073 = ~n20069 & n20072;
  assign n20074 = n20069 & ~n20072;
  assign n20075 = ~n20073 & ~n20074;
  assign n20076 = ~n20066 & n20075;
  assign n20077 = n20066 & ~n20075;
  assign n20078 = ~n20076 & ~n20077;
  assign n20079 = ~pi0173 & pi0174;
  assign n20080 = pi0173 & ~pi0174;
  assign n20081 = ~n20079 & ~n20080;
  assign n20082 = ~pi0175 & pi0176;
  assign n20083 = pi0175 & ~pi0176;
  assign n20084 = ~n20082 & ~n20083;
  assign n20085 = ~n20081 & n20084;
  assign n20086 = n20081 & ~n20084;
  assign n20087 = ~n20085 & ~n20086;
  assign n20088 = pi0142 & ~pi0178;
  assign n20089 = ~pi0142 & pi0178;
  assign n20090 = ~n20088 & ~n20089;
  assign n20091 = ~pi0177 & pi0195;
  assign n20092 = pi0177 & ~pi0195;
  assign n20093 = ~n20091 & ~n20092;
  assign n20094 = ~n20090 & n20093;
  assign n20095 = n20090 & ~n20093;
  assign n20096 = ~n20094 & ~n20095;
  assign n20097 = ~n20087 & n20096;
  assign n20098 = n20087 & ~n20096;
  assign n20099 = ~n20097 & ~n20098;
  assign n20100 = ~n20078 & n20099;
  assign n20101 = n20078 & ~n20099;
  assign n20102 = ~n20100 & ~n20101;
  assign n20103 = ~pi0187 & pi0189;
  assign n20104 = pi0187 & ~pi0189;
  assign n20105 = ~n20103 & ~n20104;
  assign n20106 = ~pi0153 & pi0179;
  assign n20107 = pi0153 & ~pi0179;
  assign n20108 = ~n20106 & ~n20107;
  assign n20109 = ~n20105 & n20108;
  assign n20110 = n20105 & ~n20108;
  assign n20111 = ~n20109 & ~n20110;
  assign n20112 = pi0141 & ~pi0172;
  assign n20113 = ~pi0141 & pi0172;
  assign n20114 = ~n20112 & ~n20113;
  assign n20115 = pi0171 & ~pi0190;
  assign n20116 = ~pi0171 & pi0190;
  assign n20117 = ~n20115 & ~n20116;
  assign n20118 = ~n20114 & n20117;
  assign n20119 = n20114 & ~n20117;
  assign n20120 = ~n20118 & ~n20119;
  assign n20121 = ~n20111 & n20120;
  assign n20122 = n20111 & ~n20120;
  assign n20123 = ~n20121 & ~n20122;
  assign n20124 = ~pi0147 & pi0148;
  assign n20125 = pi0147 & ~pi0148;
  assign n20126 = ~n20124 & ~n20125;
  assign n20127 = pi0191 & ~pi0201;
  assign n20128 = ~pi0191 & pi0201;
  assign n20129 = ~n20127 & ~n20128;
  assign n20130 = ~n20126 & n20129;
  assign n20131 = n20126 & ~n20129;
  assign n20132 = ~n20130 & ~n20131;
  assign n20133 = ~pi0149 & pi0150;
  assign n20134 = pi0149 & ~pi0150;
  assign n20135 = ~n20133 & ~n20134;
  assign n20136 = ~pi0151 & pi0152;
  assign n20137 = pi0151 & ~pi0152;
  assign n20138 = ~n20136 & ~n20137;
  assign n20139 = ~n20135 & n20138;
  assign n20140 = n20135 & ~n20138;
  assign n20141 = ~n20139 & ~n20140;
  assign n20142 = ~n20132 & n20141;
  assign n20143 = n20132 & ~n20141;
  assign n20144 = ~n20142 & ~n20143;
  assign n20145 = ~n20123 & n20144;
  assign n20146 = n20123 & ~n20144;
  assign n20147 = ~n20145 & ~n20146;
  assign n20148 = ~n20102 & n20147;
  assign n20149 = n20102 & ~n20147;
  assign n20150 = ~n20148 & ~n20149;
  assign n20151 = ~n20057 & n20150;
  assign n20152 = n20057 & ~n20150;
  assign n20153 = ~n20151 & ~n20152;
  assign n20154 = ~n20048 & n20153;
  assign n20155 = n20048 & ~n20153;
  assign n20156 = ~n20154 & ~n20155;
  assign n20157 = ~pi1878 & ~n20156;
  assign n20158 = pi0139 & ~pi1336;
  assign n20159 = ~pi0139 & pi1336;
  assign n20160 = ~n20158 & ~n20159;
  assign n20161 = pi0136 & n20150;
  assign n20162 = ~pi0136 & ~n20150;
  assign n20163 = ~n20161 & ~n20162;
  assign n20164 = pi0135 & n20163;
  assign n20165 = ~pi0135 & ~n20163;
  assign n20166 = ~n20164 & ~n20165;
  assign n20167 = ~n20160 & n20166;
  assign n20168 = n20160 & ~n20166;
  assign n20169 = ~n20167 & ~n20168;
  assign n20170 = pi1878 & ~n20169;
  assign po1524 = n20157 | n20170;
  assign n20172 = ~pi2966 & ~pi2995;
  assign n20173 = pi2982 & pi3001;
  assign n20174 = n19983 & n20173;
  assign n20175 = ~pi2920 & n20174;
  assign n20176 = n20172 & n20175;
  assign n20177 = n7254 & n20176;
  assign n20178 = ~pi2972 & n20177;
  assign n20179 = pi1348 & ~n20178;
  assign n20180 = n20012 & n20177;
  assign po1525 = n20179 | n20180;
  assign n20182 = n7254 & n20172;
  assign n20183 = pi2920 & n20182;
  assign n20184 = n19918 & n20183;
  assign n20185 = ~pi2972 & n20184;
  assign n20186 = pi1349 & ~n20185;
  assign n20187 = n19995 & n20184;
  assign po1526 = n20186 | n20187;
  assign n20189 = pi2920 & n7244;
  assign n20190 = pi2966 & n20189;
  assign n20191 = pi3001 & n20190;
  assign n20192 = pi2995 & n20191;
  assign n20193 = n7254 & n20192;
  assign n20194 = ~pi2972 & n20193;
  assign n20195 = pi1350 & ~n20194;
  assign n20196 = ~pi2972 & pi3159;
  assign n20197 = n20193 & n20196;
  assign po1527 = n20195 | n20197;
  assign n20199 = pi2920 & n19998;
  assign n20200 = n7254 & n20199;
  assign n20201 = ~pi2972 & n20200;
  assign n20202 = pi1351 & ~n20201;
  assign n20203 = n19991 & n20200;
  assign po1528 = n20202 | n20203;
  assign n20205 = pi1352 & ~n20194;
  assign n20206 = n19995 & n20193;
  assign po1529 = n20205 | n20206;
  assign n20208 = pi3156 & pi3249;
  assign n20209 = ~pi0081 & ~n20208;
  assign n20210 = ~pi1353 & ~n18958;
  assign po1530 = n20209 & ~n20210;
  assign n20212 = pi1354 & ~n20185;
  assign n20213 = n20012 & n20184;
  assign po1531 = n20212 | n20213;
  assign n20215 = pi1355 & ~n20185;
  assign n20216 = n19991 & n20184;
  assign po1532 = n20215 | n20216;
  assign n20218 = pi1356 & ~n20194;
  assign n20219 = n20012 & n20193;
  assign po1533 = n20218 | n20219;
  assign n20221 = pi1357 & ~n20194;
  assign n20222 = n19991 & n20193;
  assign po1534 = n20221 | n20222;
  assign n20224 = pi1358 & ~n20201;
  assign n20225 = n20012 & n20200;
  assign po1535 = n20224 | n20225;
  assign n20227 = pi1359 & ~n20201;
  assign n20228 = n19995 & n20200;
  assign po1536 = n20227 | n20228;
  assign n20230 = n7247 & n7254;
  assign n20231 = ~pi2972 & n20230;
  assign n20232 = pi1360 & ~n20231;
  assign n20233 = n20012 & n20230;
  assign po1537 = n20232 | n20233;
  assign n20235 = pi1361 & ~n20231;
  assign n20236 = n19991 & n20230;
  assign po1538 = n20235 | n20236;
  assign n20238 = pi1362 & ~n20231;
  assign n20239 = n19995 & n20230;
  assign po1539 = n20238 | n20239;
  assign n20241 = ~pi2920 & n19928;
  assign n20242 = ~pi2972 & n20241;
  assign n20243 = pi1363 & ~n20242;
  assign n20244 = n20012 & n20241;
  assign po1540 = n20243 | n20244;
  assign n20246 = ~pi2920 & n19920;
  assign n20247 = ~pi2972 & n20246;
  assign n20248 = pi1364 & ~n20247;
  assign n20249 = n20012 & n20246;
  assign po1541 = n20248 | n20249;
  assign n20251 = ~pi3057 & n20230;
  assign n20252 = pi1365 & ~n20251;
  assign n20253 = ~pi3057 & pi3170;
  assign n20254 = n20230 & n20253;
  assign po1542 = n20252 | n20254;
  assign n20256 = n20008 & n20253;
  assign n20257 = n7254 & n20256;
  assign n20258 = pi1366 & ~n20257;
  assign po3245 = n9402 & n19954;
  assign n20260 = n9402 & n19955;
  assign n20261 = ~po3245 & ~n20260;
  assign n20262 = pi1858 & ~n20261;
  assign n20263 = pi1341 & n20262;
  assign po1543 = n20258 | n20263;
  assign n20265 = ~pi1369 & pi3233;
  assign n20266 = pi1369 & ~pi3233;
  assign n20267 = ~n20265 & ~n20266;
  assign n20268 = ~pi1410 & pi3240;
  assign n20269 = pi1410 & ~pi3240;
  assign n20270 = ~n20268 & ~n20269;
  assign n20271 = n20267 & n20270;
  assign n20272 = pi2968 & ~n20271;
  assign n20273 = ~pi1375 & pi3224;
  assign n20274 = pi1375 & ~pi3224;
  assign n20275 = ~n20273 & ~n20274;
  assign n20276 = pi2968 & ~n20275;
  assign n20277 = ~n20272 & ~n20276;
  assign n20278 = pi1367 & n20277;
  assign n20279 = ~n19425 & ~n20277;
  assign po1544 = n20278 | n20279;
  assign n20281 = ~pi3018 & pi3172;
  assign n20282 = n7247 & n20281;
  assign n20283 = n7254 & n20282;
  assign n20284 = pi1368 & ~n20283;
  assign po1545 = n20030 | n20284;
  assign n20286 = pi1369 & n20277;
  assign n20287 = pi1367 & ~pi1407;
  assign n20288 = ~n19343 & ~n20287;
  assign n20289 = ~n20277 & ~n20288;
  assign po1546 = n20286 | n20289;
  assign n20291 = ~pi3018 & pi3135;
  assign n20292 = n7247 & n20291;
  assign n20293 = n7254 & n20292;
  assign n20294 = pi1370 & ~n20293;
  assign po1547 = ~pi3071 | n20294;
  assign n20296 = pi1371 & n20277;
  assign n20297 = ~pi1371 & ~n20277;
  assign po1548 = n20296 | n20297;
  assign n20299 = ~pi3018 & pi3150;
  assign n20300 = n7247 & n20299;
  assign n20301 = n7254 & n20300;
  assign n20302 = pi1372 & ~n20301;
  assign po1549 = n19955 | n20302;
  assign n20304 = n19917 & n20173;
  assign n20305 = n19986 & n20304;
  assign n20306 = n19991 & n20305;
  assign n20307 = n7254 & n20306;
  assign n20308 = pi1373 & ~n20307;
  assign n20309 = pi1341 & pi1396;
  assign n20310 = n20262 & n20309;
  assign po1550 = n20308 | n20310;
  assign n20312 = ~pi1750 & ~n19972;
  assign n20313 = pi1374 & ~n20312;
  assign n20314 = pi3174 & pi3348;
  assign po1551 = ~n20313 & ~n20314;
  assign n20316 = pi1375 & n20277;
  assign po1552 = n20279 | n20316;
  assign po1553 = ~n7067 | ~n18004;
  assign n20319 = ~pi3018 & n20246;
  assign n20320 = pi1377 & ~n20319;
  assign n20321 = n9530 & n20246;
  assign po1554 = n20320 | n20321;
  assign n20323 = ~pi3018 & n20241;
  assign n20324 = pi1378 & ~n20323;
  assign n20325 = n9530 & n20241;
  assign po1555 = n20324 | n20325;
  assign n20327 = pi1379 & ~n20231;
  assign n20328 = n20196 & n20230;
  assign po1556 = n20327 | n20328;
  assign n20330 = pi1407 & n19346;
  assign n20331 = pi3316 & n20330;
  assign n20332 = ~pi1380 & ~n20330;
  assign n20333 = ~n20331 & ~n20332;
  assign n20334 = ~n20277 & ~n20333;
  assign n20335 = ~pi1380 & n20277;
  assign po1557 = n20334 | n20335;
  assign n20337 = ~pi1407 & n19424;
  assign n20338 = ~pi1381 & ~n20337;
  assign n20339 = pi3293 & n20337;
  assign n20340 = ~n20338 & ~n20339;
  assign n20341 = ~n20277 & ~n20340;
  assign n20342 = ~pi1381 & n20277;
  assign po1558 = n20341 | n20342;
  assign n20344 = ~pi1382 & ~n19347;
  assign n20345 = pi3346 & n19347;
  assign n20346 = ~n20344 & ~n20345;
  assign n20347 = ~n20277 & ~n20346;
  assign n20348 = ~pi1382 & n20277;
  assign po1559 = n20347 | n20348;
  assign n20350 = pi1369 & ~n20277;
  assign n20351 = ~pi1383 & n20277;
  assign po1560 = n20350 | n20351;
  assign n20353 = ~pi1384 & ~n19347;
  assign n20354 = pi3318 & n19347;
  assign n20355 = ~n20353 & ~n20354;
  assign n20356 = ~n20277 & ~n20355;
  assign n20357 = ~pi1384 & n20277;
  assign po1561 = n20356 | n20357;
  assign n20359 = ~pi1385 & ~n19347;
  assign n20360 = pi3341 & n19347;
  assign n20361 = ~n20359 & ~n20360;
  assign n20362 = ~n20277 & ~n20361;
  assign n20363 = ~pi1385 & n20277;
  assign po1562 = n20362 | n20363;
  assign n20365 = ~pi1386 & ~n19347;
  assign n20366 = pi3355 & n19347;
  assign n20367 = ~n20365 & ~n20366;
  assign n20368 = ~n20277 & ~n20367;
  assign n20369 = ~pi1386 & n20277;
  assign po1563 = n20368 | n20369;
  assign n20371 = ~pi1387 & ~n19347;
  assign n20372 = pi3321 & n19347;
  assign n20373 = ~n20371 & ~n20372;
  assign n20374 = ~n20277 & ~n20373;
  assign n20375 = ~pi1387 & n20277;
  assign po1564 = n20374 | n20375;
  assign n20377 = ~pi1388 & ~n19347;
  assign n20378 = pi3336 & n19347;
  assign n20379 = ~n20377 & ~n20378;
  assign n20380 = ~n20277 & ~n20379;
  assign n20381 = ~pi1388 & n20277;
  assign po1565 = n20380 | n20381;
  assign n20383 = ~pi1389 & ~n19347;
  assign n20384 = pi3298 & n19347;
  assign n20385 = ~n20383 & ~n20384;
  assign n20386 = ~n20277 & ~n20385;
  assign n20387 = ~pi1389 & n20277;
  assign po1566 = n20386 | n20387;
  assign n20389 = ~pi1390 & ~n19347;
  assign n20390 = pi3333 & n19347;
  assign n20391 = ~n20389 & ~n20390;
  assign n20392 = ~n20277 & ~n20391;
  assign n20393 = ~pi1390 & n20277;
  assign po1567 = n20392 | n20393;
  assign n20395 = ~pi1391 & ~n19347;
  assign n20396 = pi3287 & n19347;
  assign n20397 = ~n20395 & ~n20396;
  assign n20398 = ~n20277 & ~n20397;
  assign n20399 = ~pi1391 & n20277;
  assign po1568 = n20398 | n20399;
  assign n20401 = ~pi1392 & ~n19347;
  assign n20402 = pi3343 & n19347;
  assign n20403 = ~n20401 & ~n20402;
  assign n20404 = ~n20277 & ~n20403;
  assign n20405 = ~pi1392 & n20277;
  assign po1569 = n20404 | n20405;
  assign n20407 = ~pi1393 & ~n20337;
  assign n20408 = pi3313 & n20337;
  assign n20409 = ~n20407 & ~n20408;
  assign n20410 = ~n20277 & ~n20409;
  assign n20411 = ~pi1393 & n20277;
  assign po1570 = n20410 | n20411;
  assign n20413 = ~pi1394 & ~n19347;
  assign n20414 = pi3290 & n19347;
  assign n20415 = ~n20413 & ~n20414;
  assign n20416 = ~n20277 & ~n20415;
  assign n20417 = ~pi1394 & n20277;
  assign po1571 = n20416 | n20417;
  assign n20419 = n7254 & n20304;
  assign n20420 = pi2920 & n20419;
  assign n20421 = n19926 & n20420;
  assign n20422 = ~pi2972 & n20421;
  assign n20423 = pi1395 & ~n20422;
  assign n20424 = n20012 & n20421;
  assign po1572 = n20423 | n20424;
  assign n20426 = pi1396 & ~n20422;
  assign n20427 = n19991 & n20421;
  assign po1573 = n20426 | n20427;
  assign n20429 = pi1397 & ~n20422;
  assign n20430 = n19995 & n20421;
  assign po1574 = n20429 | n20430;
  assign n20432 = ~pi1398 & ~n20337;
  assign n20433 = pi3311 & n20337;
  assign n20434 = ~n20432 & ~n20433;
  assign n20435 = ~n20277 & ~n20434;
  assign n20436 = ~pi1398 & n20277;
  assign po1575 = n20435 | n20436;
  assign n20438 = pi1399 & ~n7254;
  assign n20439 = ~pi2972 & pi3142;
  assign n20440 = n20192 & n20439;
  assign n20441 = ~pi2972 & n20192;
  assign n20442 = pi1399 & ~n20441;
  assign n20443 = ~n20440 & ~n20442;
  assign n20444 = n7254 & ~n20443;
  assign po1576 = n20438 | n20444;
  assign n20446 = pi1400 & ~n7254;
  assign n20447 = pi2920 & n7245;
  assign n20448 = pi2966 & n20447;
  assign n20449 = n20439 & n20448;
  assign n20450 = ~pi2972 & n20448;
  assign n20451 = pi1400 & ~n20450;
  assign n20452 = ~n20449 & ~n20451;
  assign n20453 = n7254 & ~n20452;
  assign po1577 = n20446 | n20453;
  assign n20455 = pi1401 & ~n7254;
  assign n20456 = ~pi2972 & pi3169;
  assign n20457 = n20192 & n20456;
  assign n20458 = pi1401 & ~n20441;
  assign n20459 = ~n20457 & ~n20458;
  assign n20460 = n7254 & ~n20459;
  assign po1578 = n20455 | n20460;
  assign n20462 = pi1402 & ~n7254;
  assign n20463 = ~pi2972 & pi3145;
  assign n20464 = n20192 & n20463;
  assign n20465 = pi1402 & ~n20441;
  assign n20466 = ~n20464 & ~n20465;
  assign n20467 = n7254 & ~n20466;
  assign po1579 = n20462 | n20467;
  assign n20469 = pi1403 & ~n7254;
  assign n20470 = n20448 & n20456;
  assign n20471 = pi1403 & ~n20450;
  assign n20472 = ~n20470 & ~n20471;
  assign n20473 = n7254 & ~n20472;
  assign po1580 = n20469 | n20473;
  assign n20475 = pi1404 & ~n7254;
  assign n20476 = n20448 & n20463;
  assign n20477 = pi1404 & ~n20450;
  assign n20478 = ~n20476 & ~n20477;
  assign n20479 = n7254 & ~n20478;
  assign po1581 = n20475 | n20479;
  assign n20481 = n19995 & n20305;
  assign n20482 = n7254 & n20481;
  assign n20483 = pi1405 & ~n20482;
  assign n20484 = pi3186 & pi3248;
  assign po1582 = ~n20483 & ~n20484;
  assign n20486 = n20176 & n20253;
  assign n20487 = n7254 & n20486;
  assign n20488 = pi1406 & ~n20487;
  assign n20489 = pi3185 & pi3250;
  assign po1583 = ~n20488 & ~n20489;
  assign n20491 = ~n19348 & ~n20277;
  assign n20492 = pi1407 & n20277;
  assign po1584 = n20491 | n20492;
  assign n20494 = pi1375 & ~n20277;
  assign n20495 = ~pi1408 & n20277;
  assign po1585 = n20494 | n20495;
  assign n20497 = pi1410 & ~n20277;
  assign n20498 = ~pi1409 & n20277;
  assign po1586 = n20497 | n20498;
  assign n20500 = pi1407 & ~n20277;
  assign n20501 = pi1410 & n20277;
  assign po1587 = n20500 | n20501;
  assign n20503 = ~pi1367 & ~pi1371;
  assign n20504 = pi1407 & n20503;
  assign n20505 = pi3343 & n20504;
  assign n20506 = ~pi1411 & ~n20504;
  assign n20507 = ~n20505 & ~n20506;
  assign n20508 = ~n20277 & ~n20507;
  assign n20509 = ~pi1411 & n20277;
  assign po1588 = n20508 | n20509;
  assign n20511 = pi3288 & n20504;
  assign n20512 = ~pi1412 & ~n20504;
  assign n20513 = ~n20511 & ~n20512;
  assign n20514 = ~n20277 & ~n20513;
  assign n20515 = ~pi1412 & n20277;
  assign po1589 = n20514 | n20515;
  assign n20517 = pi3328 & n20504;
  assign n20518 = ~pi1413 & ~n20504;
  assign n20519 = ~n20517 & ~n20518;
  assign n20520 = ~n20277 & ~n20519;
  assign n20521 = ~pi1413 & n20277;
  assign po1590 = n20520 | n20521;
  assign n20523 = pi3340 & n20504;
  assign n20524 = ~pi1414 & ~n20504;
  assign n20525 = ~n20523 & ~n20524;
  assign n20526 = ~n20277 & ~n20525;
  assign n20527 = ~pi1414 & n20277;
  assign po1591 = n20526 | n20527;
  assign n20529 = pi3314 & n20504;
  assign n20530 = ~pi1415 & ~n20504;
  assign n20531 = ~n20529 & ~n20530;
  assign n20532 = ~n20277 & ~n20531;
  assign n20533 = ~pi1415 & n20277;
  assign po1592 = n20532 | n20533;
  assign n20535 = pi3347 & n20504;
  assign n20536 = ~pi1416 & ~n20504;
  assign n20537 = ~n20535 & ~n20536;
  assign n20538 = ~n20277 & ~n20537;
  assign n20539 = ~pi1416 & n20277;
  assign po1593 = n20538 | n20539;
  assign n20541 = pi3316 & n20504;
  assign n20542 = ~pi1417 & ~n20504;
  assign n20543 = ~n20541 & ~n20542;
  assign n20544 = ~n20277 & ~n20543;
  assign n20545 = ~pi1417 & n20277;
  assign po1594 = n20544 | n20545;
  assign n20547 = pi3333 & n20504;
  assign n20548 = ~pi1418 & ~n20504;
  assign n20549 = ~n20547 & ~n20548;
  assign n20550 = ~n20277 & ~n20549;
  assign n20551 = ~pi1418 & n20277;
  assign po1595 = n20550 | n20551;
  assign n20553 = pi3330 & n20504;
  assign n20554 = ~pi1419 & ~n20504;
  assign n20555 = ~n20553 & ~n20554;
  assign n20556 = ~n20277 & ~n20555;
  assign n20557 = ~pi1419 & n20277;
  assign po1596 = n20556 | n20557;
  assign n20559 = pi3326 & n20504;
  assign n20560 = ~pi1420 & ~n20504;
  assign n20561 = ~n20559 & ~n20560;
  assign n20562 = ~n20277 & ~n20561;
  assign n20563 = ~pi1420 & n20277;
  assign po1597 = n20562 | n20563;
  assign n20565 = pi3295 & n20504;
  assign n20566 = ~pi1421 & ~n20504;
  assign n20567 = ~n20565 & ~n20566;
  assign n20568 = ~n20277 & ~n20567;
  assign n20569 = ~pi1421 & n20277;
  assign po1598 = n20568 | n20569;
  assign n20571 = pi3349 & n20504;
  assign n20572 = ~pi1422 & ~n20504;
  assign n20573 = ~n20571 & ~n20572;
  assign n20574 = ~n20277 & ~n20573;
  assign n20575 = ~pi1422 & n20277;
  assign po1599 = n20574 | n20575;
  assign n20577 = pi3354 & n20504;
  assign n20578 = ~pi1423 & ~n20504;
  assign n20579 = ~n20577 & ~n20578;
  assign n20580 = ~n20277 & ~n20579;
  assign n20581 = ~pi1423 & n20277;
  assign po1600 = n20580 | n20581;
  assign n20583 = pi3299 & n20504;
  assign n20584 = ~pi1424 & ~n20504;
  assign n20585 = ~n20583 & ~n20584;
  assign n20586 = ~n20277 & ~n20585;
  assign n20587 = ~pi1424 & n20277;
  assign po1601 = n20586 | n20587;
  assign n20589 = pi2994 & n20504;
  assign n20590 = ~pi1425 & ~n20504;
  assign n20591 = ~n20589 & ~n20590;
  assign n20592 = ~n20277 & ~n20591;
  assign n20593 = ~pi1425 & n20277;
  assign po1602 = n20592 | n20593;
  assign n20595 = pi3311 & n20504;
  assign n20596 = ~pi1426 & ~n20504;
  assign n20597 = ~n20595 & ~n20596;
  assign n20598 = ~n20277 & ~n20597;
  assign n20599 = ~pi1426 & n20277;
  assign po1603 = n20598 | n20599;
  assign n20601 = pi3353 & n20504;
  assign n20602 = ~pi1427 & ~n20504;
  assign n20603 = ~n20601 & ~n20602;
  assign n20604 = ~n20277 & ~n20603;
  assign n20605 = ~pi1427 & n20277;
  assign po1604 = n20604 | n20605;
  assign n20607 = pi3293 & n20504;
  assign n20608 = ~pi1428 & ~n20504;
  assign n20609 = ~n20607 & ~n20608;
  assign n20610 = ~n20277 & ~n20609;
  assign n20611 = ~pi1428 & n20277;
  assign po1605 = n20610 | n20611;
  assign n20613 = pi3313 & n20504;
  assign n20614 = ~pi1429 & ~n20504;
  assign n20615 = ~n20613 & ~n20614;
  assign n20616 = ~n20277 & ~n20615;
  assign n20617 = ~pi1429 & n20277;
  assign po1606 = n20616 | n20617;
  assign n20619 = pi1407 & n19423;
  assign n20620 = pi3343 & n20619;
  assign n20621 = ~pi1430 & ~n20619;
  assign n20622 = ~n20620 & ~n20621;
  assign n20623 = ~n20277 & ~n20622;
  assign n20624 = ~pi1430 & n20277;
  assign po1607 = n20623 | n20624;
  assign n20626 = pi3287 & n20619;
  assign n20627 = ~pi1431 & ~n20619;
  assign n20628 = ~n20626 & ~n20627;
  assign n20629 = ~n20277 & ~n20628;
  assign n20630 = ~pi1431 & n20277;
  assign po1608 = n20629 | n20630;
  assign n20632 = pi3328 & n20619;
  assign n20633 = ~pi1432 & ~n20619;
  assign n20634 = ~n20632 & ~n20633;
  assign n20635 = ~n20277 & ~n20634;
  assign n20636 = ~pi1432 & n20277;
  assign po1609 = n20635 | n20636;
  assign n20638 = pi3286 & n20619;
  assign n20639 = ~pi1433 & ~n20619;
  assign n20640 = ~n20638 & ~n20639;
  assign n20641 = ~n20277 & ~n20640;
  assign n20642 = ~pi1433 & n20277;
  assign po1610 = n20641 | n20642;
  assign n20644 = pi3290 & n20619;
  assign n20645 = ~pi1434 & ~n20619;
  assign n20646 = ~n20644 & ~n20645;
  assign n20647 = ~n20277 & ~n20646;
  assign n20648 = ~pi1434 & n20277;
  assign po1611 = n20647 | n20648;
  assign n20650 = pi3314 & n20619;
  assign n20651 = ~pi1435 & ~n20619;
  assign n20652 = ~n20650 & ~n20651;
  assign n20653 = ~n20277 & ~n20652;
  assign n20654 = ~pi1435 & n20277;
  assign po1612 = n20653 | n20654;
  assign n20656 = pi3315 & n20619;
  assign n20657 = ~pi1436 & ~n20619;
  assign n20658 = ~n20656 & ~n20657;
  assign n20659 = ~n20277 & ~n20658;
  assign n20660 = ~pi1436 & n20277;
  assign po1613 = n20659 | n20660;
  assign n20662 = pi3298 & n20619;
  assign n20663 = ~pi1437 & ~n20619;
  assign n20664 = ~n20662 & ~n20663;
  assign n20665 = ~n20277 & ~n20664;
  assign n20666 = ~pi1437 & n20277;
  assign po1614 = n20665 | n20666;
  assign n20668 = pi3316 & n20619;
  assign n20669 = ~pi1438 & ~n20619;
  assign n20670 = ~n20668 & ~n20669;
  assign n20671 = ~n20277 & ~n20670;
  assign n20672 = ~pi1438 & n20277;
  assign po1615 = n20671 | n20672;
  assign n20674 = pi3333 & n20619;
  assign n20675 = ~pi1439 & ~n20619;
  assign n20676 = ~n20674 & ~n20675;
  assign n20677 = ~n20277 & ~n20676;
  assign n20678 = ~pi1439 & n20277;
  assign po1616 = n20677 | n20678;
  assign n20680 = pi3321 & n20619;
  assign n20681 = ~pi1440 & ~n20619;
  assign n20682 = ~n20680 & ~n20681;
  assign n20683 = ~n20277 & ~n20682;
  assign n20684 = ~pi1440 & n20277;
  assign po1617 = n20683 | n20684;
  assign n20686 = pi3336 & n20619;
  assign n20687 = ~pi1441 & ~n20619;
  assign n20688 = ~n20686 & ~n20687;
  assign n20689 = ~n20277 & ~n20688;
  assign n20690 = ~pi1441 & n20277;
  assign po1618 = n20689 | n20690;
  assign n20692 = pi3318 & n20619;
  assign n20693 = ~pi1442 & ~n20619;
  assign n20694 = ~n20692 & ~n20693;
  assign n20695 = ~n20277 & ~n20694;
  assign n20696 = ~pi1442 & n20277;
  assign po1619 = n20695 | n20696;
  assign n20698 = pi3350 & n20619;
  assign n20699 = ~pi1443 & ~n20619;
  assign n20700 = ~n20698 & ~n20699;
  assign n20701 = ~n20277 & ~n20700;
  assign n20702 = ~pi1443 & n20277;
  assign po1620 = n20701 | n20702;
  assign n20704 = pi3355 & n20619;
  assign n20705 = ~pi1444 & ~n20619;
  assign n20706 = ~n20704 & ~n20705;
  assign n20707 = ~n20277 & ~n20706;
  assign n20708 = ~pi1444 & n20277;
  assign po1621 = n20707 | n20708;
  assign n20710 = pi3341 & n20619;
  assign n20711 = ~pi1445 & ~n20619;
  assign n20712 = ~n20710 & ~n20711;
  assign n20713 = ~n20277 & ~n20712;
  assign n20714 = ~pi1445 & n20277;
  assign po1622 = n20713 | n20714;
  assign n20716 = pi3346 & n20619;
  assign n20717 = ~pi1446 & ~n20619;
  assign n20718 = ~n20716 & ~n20717;
  assign n20719 = ~n20277 & ~n20718;
  assign n20720 = ~pi1446 & n20277;
  assign po1623 = n20719 | n20720;
  assign n20722 = pi3311 & n20619;
  assign n20723 = ~pi1447 & ~n20619;
  assign n20724 = ~n20722 & ~n20723;
  assign n20725 = ~n20277 & ~n20724;
  assign n20726 = ~pi1447 & n20277;
  assign po1624 = n20725 | n20726;
  assign n20728 = pi3353 & n20619;
  assign n20729 = ~pi1448 & ~n20619;
  assign n20730 = ~n20728 & ~n20729;
  assign n20731 = ~n20277 & ~n20730;
  assign n20732 = ~pi1448 & n20277;
  assign po1625 = n20731 | n20732;
  assign n20734 = pi3337 & n20619;
  assign n20735 = ~pi1449 & ~n20619;
  assign n20736 = ~n20734 & ~n20735;
  assign n20737 = ~n20277 & ~n20736;
  assign n20738 = ~pi1449 & n20277;
  assign po1626 = n20737 | n20738;
  assign n20740 = pi3313 & n20619;
  assign n20741 = ~pi1450 & ~n20619;
  assign n20742 = ~n20740 & ~n20741;
  assign n20743 = ~n20277 & ~n20742;
  assign n20744 = ~pi1450 & n20277;
  assign po1627 = n20743 | n20744;
  assign n20746 = pi3335 & n20619;
  assign n20747 = ~pi1451 & ~n20619;
  assign n20748 = ~n20746 & ~n20747;
  assign n20749 = ~n20277 & ~n20748;
  assign n20750 = ~pi1451 & n20277;
  assign po1628 = n20749 | n20750;
  assign n20752 = pi1407 & n19424;
  assign n20753 = pi3288 & n20752;
  assign n20754 = ~pi1452 & ~n20752;
  assign n20755 = ~n20753 & ~n20754;
  assign n20756 = ~n20277 & ~n20755;
  assign n20757 = ~pi1452 & n20277;
  assign po1629 = n20756 | n20757;
  assign n20759 = pi3287 & n20752;
  assign n20760 = ~pi1453 & ~n20752;
  assign n20761 = ~n20759 & ~n20760;
  assign n20762 = ~n20277 & ~n20761;
  assign n20763 = ~pi1453 & n20277;
  assign po1630 = n20762 | n20763;
  assign n20765 = pi3328 & n20752;
  assign n20766 = ~pi1454 & ~n20752;
  assign n20767 = ~n20765 & ~n20766;
  assign n20768 = ~n20277 & ~n20767;
  assign n20769 = ~pi1454 & n20277;
  assign po1631 = n20768 | n20769;
  assign n20771 = pi3340 & n20752;
  assign n20772 = ~pi1455 & ~n20752;
  assign n20773 = ~n20771 & ~n20772;
  assign n20774 = ~n20277 & ~n20773;
  assign n20775 = ~pi1455 & n20277;
  assign po1632 = n20774 | n20775;
  assign n20777 = pi3314 & n20752;
  assign n20778 = ~pi1456 & ~n20752;
  assign n20779 = ~n20777 & ~n20778;
  assign n20780 = ~n20277 & ~n20779;
  assign n20781 = ~pi1456 & n20277;
  assign po1633 = n20780 | n20781;
  assign n20783 = pi3347 & n20752;
  assign n20784 = ~pi1457 & ~n20752;
  assign n20785 = ~n20783 & ~n20784;
  assign n20786 = ~n20277 & ~n20785;
  assign n20787 = ~pi1457 & n20277;
  assign po1634 = n20786 | n20787;
  assign n20789 = pi3298 & n20752;
  assign n20790 = ~pi1458 & ~n20752;
  assign n20791 = ~n20789 & ~n20790;
  assign n20792 = ~n20277 & ~n20791;
  assign n20793 = ~pi1458 & n20277;
  assign po1635 = n20792 | n20793;
  assign n20795 = pi3316 & n20752;
  assign n20796 = ~pi1459 & ~n20752;
  assign n20797 = ~n20795 & ~n20796;
  assign n20798 = ~n20277 & ~n20797;
  assign n20799 = ~pi1459 & n20277;
  assign po1636 = n20798 | n20799;
  assign n20801 = pi3330 & n20752;
  assign n20802 = ~pi1460 & ~n20752;
  assign n20803 = ~n20801 & ~n20802;
  assign n20804 = ~n20277 & ~n20803;
  assign n20805 = ~pi1460 & n20277;
  assign po1637 = n20804 | n20805;
  assign n20807 = pi3326 & n20752;
  assign n20808 = ~pi1461 & ~n20752;
  assign n20809 = ~n20807 & ~n20808;
  assign n20810 = ~n20277 & ~n20809;
  assign n20811 = ~pi1461 & n20277;
  assign po1638 = n20810 | n20811;
  assign n20813 = pi3295 & n20752;
  assign n20814 = ~pi1462 & ~n20752;
  assign n20815 = ~n20813 & ~n20814;
  assign n20816 = ~n20277 & ~n20815;
  assign n20817 = ~pi1462 & n20277;
  assign po1639 = n20816 | n20817;
  assign n20819 = pi3318 & n20752;
  assign n20820 = ~pi1463 & ~n20752;
  assign n20821 = ~n20819 & ~n20820;
  assign n20822 = ~n20277 & ~n20821;
  assign n20823 = ~pi1463 & n20277;
  assign po1640 = n20822 | n20823;
  assign n20825 = pi3349 & n20752;
  assign n20826 = ~pi1464 & ~n20752;
  assign n20827 = ~n20825 & ~n20826;
  assign n20828 = ~n20277 & ~n20827;
  assign n20829 = ~pi1464 & n20277;
  assign po1641 = n20828 | n20829;
  assign n20831 = pi3354 & n20752;
  assign n20832 = ~pi1465 & ~n20752;
  assign n20833 = ~n20831 & ~n20832;
  assign n20834 = ~n20277 & ~n20833;
  assign n20835 = ~pi1465 & n20277;
  assign po1642 = n20834 | n20835;
  assign n20837 = pi3299 & n20752;
  assign n20838 = ~pi1466 & ~n20752;
  assign n20839 = ~n20837 & ~n20838;
  assign n20840 = ~n20277 & ~n20839;
  assign n20841 = ~pi1466 & n20277;
  assign po1643 = n20840 | n20841;
  assign n20843 = pi2994 & n20752;
  assign n20844 = ~pi1467 & ~n20752;
  assign n20845 = ~n20843 & ~n20844;
  assign n20846 = ~n20277 & ~n20845;
  assign n20847 = ~pi1467 & n20277;
  assign po1644 = n20846 | n20847;
  assign n20849 = pi3346 & n20752;
  assign n20850 = ~pi1468 & ~n20752;
  assign n20851 = ~n20849 & ~n20850;
  assign n20852 = ~n20277 & ~n20851;
  assign n20853 = ~pi1468 & n20277;
  assign po1645 = n20852 | n20853;
  assign n20855 = pi3311 & n20752;
  assign n20856 = ~pi1469 & ~n20752;
  assign n20857 = ~n20855 & ~n20856;
  assign n20858 = ~n20277 & ~n20857;
  assign n20859 = ~pi1469 & n20277;
  assign po1646 = n20858 | n20859;
  assign n20861 = pi3293 & n20752;
  assign n20862 = ~pi1470 & ~n20752;
  assign n20863 = ~n20861 & ~n20862;
  assign n20864 = ~n20277 & ~n20863;
  assign n20865 = ~pi1470 & n20277;
  assign po1647 = n20864 | n20865;
  assign n20867 = pi3337 & n20752;
  assign n20868 = ~pi1471 & ~n20752;
  assign n20869 = ~n20867 & ~n20868;
  assign n20870 = ~n20277 & ~n20869;
  assign n20871 = ~pi1471 & n20277;
  assign po1648 = n20870 | n20871;
  assign n20873 = pi3313 & n20752;
  assign n20874 = ~pi1472 & ~n20752;
  assign n20875 = ~n20873 & ~n20874;
  assign n20876 = ~n20277 & ~n20875;
  assign n20877 = ~pi1472 & n20277;
  assign po1649 = n20876 | n20877;
  assign n20879 = pi3343 & n20330;
  assign n20880 = ~pi1473 & ~n20330;
  assign n20881 = ~n20879 & ~n20880;
  assign n20882 = ~n20277 & ~n20881;
  assign n20883 = ~pi1473 & n20277;
  assign po1650 = n20882 | n20883;
  assign n20885 = pi3288 & n20330;
  assign n20886 = ~pi1474 & ~n20330;
  assign n20887 = ~n20885 & ~n20886;
  assign n20888 = ~n20277 & ~n20887;
  assign n20889 = ~pi1474 & n20277;
  assign po1651 = n20888 | n20889;
  assign n20891 = pi3287 & n20330;
  assign n20892 = ~pi1475 & ~n20330;
  assign n20893 = ~n20891 & ~n20892;
  assign n20894 = ~n20277 & ~n20893;
  assign n20895 = ~pi1475 & n20277;
  assign po1652 = n20894 | n20895;
  assign n20897 = pi3286 & n20330;
  assign n20898 = ~pi1476 & ~n20330;
  assign n20899 = ~n20897 & ~n20898;
  assign n20900 = ~n20277 & ~n20899;
  assign n20901 = ~pi1476 & n20277;
  assign po1653 = n20900 | n20901;
  assign n20903 = pi3290 & n20330;
  assign n20904 = ~pi1477 & ~n20330;
  assign n20905 = ~n20903 & ~n20904;
  assign n20906 = ~n20277 & ~n20905;
  assign n20907 = ~pi1477 & n20277;
  assign po1654 = n20906 | n20907;
  assign n20909 = pi3315 & n20330;
  assign n20910 = ~pi1478 & ~n20330;
  assign n20911 = ~n20909 & ~n20910;
  assign n20912 = ~n20277 & ~n20911;
  assign n20913 = ~pi1478 & n20277;
  assign po1655 = n20912 | n20913;
  assign n20915 = pi3347 & n20330;
  assign n20916 = ~pi1479 & ~n20330;
  assign n20917 = ~n20915 & ~n20916;
  assign n20918 = ~n20277 & ~n20917;
  assign n20919 = ~pi1479 & n20277;
  assign po1656 = n20918 | n20919;
  assign n20921 = pi3298 & n20330;
  assign n20922 = ~pi1480 & ~n20330;
  assign n20923 = ~n20921 & ~n20922;
  assign n20924 = ~n20277 & ~n20923;
  assign n20925 = ~pi1480 & n20277;
  assign po1657 = n20924 | n20925;
  assign n20927 = pi3333 & n20330;
  assign n20928 = ~pi1481 & ~n20330;
  assign n20929 = ~n20927 & ~n20928;
  assign n20930 = ~n20277 & ~n20929;
  assign n20931 = ~pi1481 & n20277;
  assign po1658 = n20930 | n20931;
  assign n20933 = pi3321 & n20330;
  assign n20934 = ~pi1482 & ~n20330;
  assign n20935 = ~n20933 & ~n20934;
  assign n20936 = ~n20277 & ~n20935;
  assign n20937 = ~pi1482 & n20277;
  assign po1659 = n20936 | n20937;
  assign n20939 = pi3336 & n20330;
  assign n20940 = ~pi1483 & ~n20330;
  assign n20941 = ~n20939 & ~n20940;
  assign n20942 = ~n20277 & ~n20941;
  assign n20943 = ~pi1483 & n20277;
  assign po1660 = n20942 | n20943;
  assign n20945 = pi3295 & n20330;
  assign n20946 = ~pi1484 & ~n20330;
  assign n20947 = ~n20945 & ~n20946;
  assign n20948 = ~n20277 & ~n20947;
  assign n20949 = ~pi1484 & n20277;
  assign po1661 = n20948 | n20949;
  assign n20951 = pi3318 & n20330;
  assign n20952 = ~pi1485 & ~n20330;
  assign n20953 = ~n20951 & ~n20952;
  assign n20954 = ~n20277 & ~n20953;
  assign n20955 = ~pi1485 & n20277;
  assign po1662 = n20954 | n20955;
  assign n20957 = pi3350 & n20330;
  assign n20958 = ~pi1486 & ~n20330;
  assign n20959 = ~n20957 & ~n20958;
  assign n20960 = ~n20277 & ~n20959;
  assign n20961 = ~pi1486 & n20277;
  assign po1663 = n20960 | n20961;
  assign n20963 = pi3354 & n20330;
  assign n20964 = ~pi1487 & ~n20330;
  assign n20965 = ~n20963 & ~n20964;
  assign n20966 = ~n20277 & ~n20965;
  assign n20967 = ~pi1487 & n20277;
  assign po1664 = n20966 | n20967;
  assign n20969 = pi3355 & n20330;
  assign n20970 = ~pi1488 & ~n20330;
  assign n20971 = ~n20969 & ~n20970;
  assign n20972 = ~n20277 & ~n20971;
  assign n20973 = ~pi1488 & n20277;
  assign po1665 = n20972 | n20973;
  assign n20975 = pi3341 & n20330;
  assign n20976 = ~pi1489 & ~n20330;
  assign n20977 = ~n20975 & ~n20976;
  assign n20978 = ~n20277 & ~n20977;
  assign n20979 = ~pi1489 & n20277;
  assign po1666 = n20978 | n20979;
  assign n20981 = pi2994 & n20330;
  assign n20982 = ~pi1490 & ~n20330;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = ~n20277 & ~n20983;
  assign n20985 = ~pi1490 & n20277;
  assign po1667 = n20984 | n20985;
  assign n20987 = pi3346 & n20330;
  assign n20988 = ~pi1491 & ~n20330;
  assign n20989 = ~n20987 & ~n20988;
  assign n20990 = ~n20277 & ~n20989;
  assign n20991 = ~pi1491 & n20277;
  assign po1668 = n20990 | n20991;
  assign n20993 = pi3353 & n20330;
  assign n20994 = ~pi1492 & ~n20330;
  assign n20995 = ~n20993 & ~n20994;
  assign n20996 = ~n20277 & ~n20995;
  assign n20997 = ~pi1492 & n20277;
  assign po1669 = n20996 | n20997;
  assign n20999 = pi3337 & n20330;
  assign n21000 = ~pi1493 & ~n20330;
  assign n21001 = ~n20999 & ~n21000;
  assign n21002 = ~n20277 & ~n21001;
  assign n21003 = ~pi1493 & n20277;
  assign po1670 = n21002 | n21003;
  assign n21005 = pi3335 & n20330;
  assign n21006 = ~pi1494 & ~n20330;
  assign n21007 = ~n21005 & ~n21006;
  assign n21008 = ~n20277 & ~n21007;
  assign n21009 = ~pi1494 & n20277;
  assign po1671 = n21008 | n21009;
  assign n21011 = ~pi1407 & n19423;
  assign n21012 = ~pi1495 & ~n21011;
  assign n21013 = pi3340 & n21011;
  assign n21014 = ~n21012 & ~n21013;
  assign n21015 = ~n20277 & ~n21014;
  assign n21016 = ~pi1495 & n20277;
  assign po1672 = n21015 | n21016;
  assign n21018 = ~pi1496 & ~n21011;
  assign n21019 = pi3290 & n21011;
  assign n21020 = ~n21018 & ~n21019;
  assign n21021 = ~n20277 & ~n21020;
  assign n21022 = ~pi1496 & n20277;
  assign po1673 = n21021 | n21022;
  assign n21024 = ~pi1497 & ~n21011;
  assign n21025 = pi3314 & n21011;
  assign n21026 = ~n21024 & ~n21025;
  assign n21027 = ~n20277 & ~n21026;
  assign n21028 = ~pi1497 & n20277;
  assign po1674 = n21027 | n21028;
  assign n21030 = ~pi1498 & ~n21011;
  assign n21031 = pi3347 & n21011;
  assign n21032 = ~n21030 & ~n21031;
  assign n21033 = ~n20277 & ~n21032;
  assign n21034 = ~pi1498 & n20277;
  assign po1675 = n21033 | n21034;
  assign n21036 = ~pi1499 & ~n21011;
  assign n21037 = pi3316 & n21011;
  assign n21038 = ~n21036 & ~n21037;
  assign n21039 = ~n20277 & ~n21038;
  assign n21040 = ~pi1499 & n20277;
  assign po1676 = n21039 | n21040;
  assign n21042 = ~pi1500 & ~n21011;
  assign n21043 = pi3330 & n21011;
  assign n21044 = ~n21042 & ~n21043;
  assign n21045 = ~n20277 & ~n21044;
  assign n21046 = ~pi1500 & n20277;
  assign po1677 = n21045 | n21046;
  assign n21048 = ~pi1501 & ~n21011;
  assign n21049 = pi3321 & n21011;
  assign n21050 = ~n21048 & ~n21049;
  assign n21051 = ~n20277 & ~n21050;
  assign n21052 = ~pi1501 & n20277;
  assign po1678 = n21051 | n21052;
  assign n21054 = ~pi1502 & ~n21011;
  assign n21055 = pi3326 & n21011;
  assign n21056 = ~n21054 & ~n21055;
  assign n21057 = ~n20277 & ~n21056;
  assign n21058 = ~pi1502 & n20277;
  assign po1679 = n21057 | n21058;
  assign n21060 = ~pi1503 & ~n21011;
  assign n21061 = pi3295 & n21011;
  assign n21062 = ~n21060 & ~n21061;
  assign n21063 = ~n20277 & ~n21062;
  assign n21064 = ~pi1503 & n20277;
  assign po1680 = n21063 | n21064;
  assign n21066 = ~pi1504 & ~n21011;
  assign n21067 = pi3349 & n21011;
  assign n21068 = ~n21066 & ~n21067;
  assign n21069 = ~n20277 & ~n21068;
  assign n21070 = ~pi1504 & n20277;
  assign po1681 = n21069 | n21070;
  assign n21072 = ~pi1505 & ~n21011;
  assign n21073 = pi3354 & n21011;
  assign n21074 = ~n21072 & ~n21073;
  assign n21075 = ~n20277 & ~n21074;
  assign n21076 = ~pi1505 & n20277;
  assign po1682 = n21075 | n21076;
  assign n21078 = ~pi1506 & ~n21011;
  assign n21079 = pi3355 & n21011;
  assign n21080 = ~n21078 & ~n21079;
  assign n21081 = ~n20277 & ~n21080;
  assign n21082 = ~pi1506 & n20277;
  assign po1683 = n21081 | n21082;
  assign n21084 = ~pi1507 & ~n21011;
  assign n21085 = pi3299 & n21011;
  assign n21086 = ~n21084 & ~n21085;
  assign n21087 = ~n20277 & ~n21086;
  assign n21088 = ~pi1507 & n20277;
  assign po1684 = n21087 | n21088;
  assign n21090 = ~pi1508 & ~n21011;
  assign n21091 = pi2994 & n21011;
  assign n21092 = ~n21090 & ~n21091;
  assign n21093 = ~n20277 & ~n21092;
  assign n21094 = ~pi1508 & n20277;
  assign po1685 = n21093 | n21094;
  assign n21096 = ~pi1509 & ~n21011;
  assign n21097 = pi3311 & n21011;
  assign n21098 = ~n21096 & ~n21097;
  assign n21099 = ~n20277 & ~n21098;
  assign n21100 = ~pi1509 & n20277;
  assign po1686 = n21099 | n21100;
  assign n21102 = ~pi1510 & ~n21011;
  assign n21103 = pi3293 & n21011;
  assign n21104 = ~n21102 & ~n21103;
  assign n21105 = ~n20277 & ~n21104;
  assign n21106 = ~pi1510 & n20277;
  assign po1687 = n21105 | n21106;
  assign n21108 = ~pi1511 & ~n21011;
  assign n21109 = pi3337 & n21011;
  assign n21110 = ~n21108 & ~n21109;
  assign n21111 = ~n20277 & ~n21110;
  assign n21112 = ~pi1511 & n20277;
  assign po1688 = n21111 | n21112;
  assign n21114 = ~pi1512 & ~n21011;
  assign n21115 = pi3313 & n21011;
  assign n21116 = ~n21114 & ~n21115;
  assign n21117 = ~n20277 & ~n21116;
  assign n21118 = ~pi1512 & n20277;
  assign po1689 = n21117 | n21118;
  assign n21120 = ~pi1513 & ~n20337;
  assign n21121 = pi3343 & n20337;
  assign n21122 = ~n21120 & ~n21121;
  assign n21123 = ~n20277 & ~n21122;
  assign n21124 = ~pi1513 & n20277;
  assign po1690 = n21123 | n21124;
  assign n21126 = ~pi1514 & ~n20337;
  assign n21127 = pi3287 & n20337;
  assign n21128 = ~n21126 & ~n21127;
  assign n21129 = ~n20277 & ~n21128;
  assign n21130 = ~pi1514 & n20277;
  assign po1691 = n21129 | n21130;
  assign n21132 = ~pi1515 & ~n20337;
  assign n21133 = pi3286 & n20337;
  assign n21134 = ~n21132 & ~n21133;
  assign n21135 = ~n20277 & ~n21134;
  assign n21136 = ~pi1515 & n20277;
  assign po1692 = n21135 | n21136;
  assign n21138 = ~pi1516 & ~n20337;
  assign n21139 = pi3340 & n20337;
  assign n21140 = ~n21138 & ~n21139;
  assign n21141 = ~n20277 & ~n21140;
  assign n21142 = ~pi1516 & n20277;
  assign po1693 = n21141 | n21142;
  assign n21144 = ~pi1517 & ~n20337;
  assign n21145 = pi3290 & n20337;
  assign n21146 = ~n21144 & ~n21145;
  assign n21147 = ~n20277 & ~n21146;
  assign n21148 = ~pi1517 & n20277;
  assign po1694 = n21147 | n21148;
  assign n21150 = ~pi1518 & ~n20337;
  assign n21151 = pi3315 & n20337;
  assign n21152 = ~n21150 & ~n21151;
  assign n21153 = ~n20277 & ~n21152;
  assign n21154 = ~pi1518 & n20277;
  assign po1695 = n21153 | n21154;
  assign n21156 = ~pi1519 & ~n20337;
  assign n21157 = pi3347 & n20337;
  assign n21158 = ~n21156 & ~n21157;
  assign n21159 = ~n20277 & ~n21158;
  assign n21160 = ~pi1519 & n20277;
  assign po1696 = n21159 | n21160;
  assign n21162 = ~pi1520 & ~n20337;
  assign n21163 = pi3298 & n20337;
  assign n21164 = ~n21162 & ~n21163;
  assign n21165 = ~n20277 & ~n21164;
  assign n21166 = ~pi1520 & n20277;
  assign po1697 = n21165 | n21166;
  assign n21168 = ~pi1521 & ~n20337;
  assign n21169 = pi3333 & n20337;
  assign n21170 = ~n21168 & ~n21169;
  assign n21171 = ~n20277 & ~n21170;
  assign n21172 = ~pi1521 & n20277;
  assign po1698 = n21171 | n21172;
  assign n21174 = ~pi1522 & ~n20337;
  assign n21175 = pi3321 & n20337;
  assign n21176 = ~n21174 & ~n21175;
  assign n21177 = ~n20277 & ~n21176;
  assign n21178 = ~pi1522 & n20277;
  assign po1699 = n21177 | n21178;
  assign n21180 = ~pi1523 & ~n20337;
  assign n21181 = pi3336 & n20337;
  assign n21182 = ~n21180 & ~n21181;
  assign n21183 = ~n20277 & ~n21182;
  assign n21184 = ~pi1523 & n20277;
  assign po1700 = n21183 | n21184;
  assign n21186 = ~pi1524 & ~n20337;
  assign n21187 = pi3318 & n20337;
  assign n21188 = ~n21186 & ~n21187;
  assign n21189 = ~n20277 & ~n21188;
  assign n21190 = ~pi1524 & n20277;
  assign po1701 = n21189 | n21190;
  assign n21192 = ~pi1525 & ~n20337;
  assign n21193 = pi3350 & n20337;
  assign n21194 = ~n21192 & ~n21193;
  assign n21195 = ~n20277 & ~n21194;
  assign n21196 = ~pi1525 & n20277;
  assign po1702 = n21195 | n21196;
  assign n21198 = ~pi1526 & ~n20337;
  assign n21199 = pi3354 & n20337;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 = ~n20277 & ~n21200;
  assign n21202 = ~pi1526 & n20277;
  assign po1703 = n21201 | n21202;
  assign n21204 = ~pi1527 & ~n20337;
  assign n21205 = pi3355 & n20337;
  assign n21206 = ~n21204 & ~n21205;
  assign n21207 = ~n20277 & ~n21206;
  assign n21208 = ~pi1527 & n20277;
  assign po1704 = n21207 | n21208;
  assign n21210 = ~pi1528 & ~n20337;
  assign n21211 = pi3341 & n20337;
  assign n21212 = ~n21210 & ~n21211;
  assign n21213 = ~n20277 & ~n21212;
  assign n21214 = ~pi1528 & n20277;
  assign po1705 = n21213 | n21214;
  assign n21216 = ~pi1529 & ~n20337;
  assign n21217 = pi3346 & n20337;
  assign n21218 = ~n21216 & ~n21217;
  assign n21219 = ~n20277 & ~n21218;
  assign n21220 = ~pi1529 & n20277;
  assign po1706 = n21219 | n21220;
  assign n21222 = ~pi1530 & ~n20337;
  assign n21223 = pi3353 & n20337;
  assign n21224 = ~n21222 & ~n21223;
  assign n21225 = ~n20277 & ~n21224;
  assign n21226 = ~pi1530 & n20277;
  assign po1707 = n21225 | n21226;
  assign n21228 = ~pi1531 & ~n20337;
  assign n21229 = pi3337 & n20337;
  assign n21230 = ~n21228 & ~n21229;
  assign n21231 = ~n20277 & ~n21230;
  assign n21232 = ~pi1531 & n20277;
  assign po1708 = n21231 | n21232;
  assign n21234 = ~pi1532 & ~n20337;
  assign n21235 = pi3335 & n20337;
  assign n21236 = ~n21234 & ~n21235;
  assign n21237 = ~n20277 & ~n21236;
  assign n21238 = ~pi1532 & n20277;
  assign po1709 = n21237 | n21238;
  assign n21240 = ~pi1533 & ~n19347;
  assign n21241 = pi3288 & n19347;
  assign n21242 = ~n21240 & ~n21241;
  assign n21243 = ~n20277 & ~n21242;
  assign n21244 = ~pi1533 & n20277;
  assign po1710 = n21243 | n21244;
  assign n21246 = ~pi1534 & ~n19347;
  assign n21247 = pi3328 & n19347;
  assign n21248 = ~n21246 & ~n21247;
  assign n21249 = ~n20277 & ~n21248;
  assign n21250 = ~pi1534 & n20277;
  assign po1711 = n21249 | n21250;
  assign n21252 = ~pi1535 & ~n19347;
  assign n21253 = pi3286 & n19347;
  assign n21254 = ~n21252 & ~n21253;
  assign n21255 = ~n20277 & ~n21254;
  assign n21256 = ~pi1535 & n20277;
  assign po1712 = n21255 | n21256;
  assign n21258 = ~pi1536 & ~n19347;
  assign n21259 = pi3340 & n19347;
  assign n21260 = ~n21258 & ~n21259;
  assign n21261 = ~n20277 & ~n21260;
  assign n21262 = ~pi1536 & n20277;
  assign po1713 = n21261 | n21262;
  assign n21264 = ~pi1537 & ~n19347;
  assign n21265 = pi3314 & n19347;
  assign n21266 = ~n21264 & ~n21265;
  assign n21267 = ~n20277 & ~n21266;
  assign n21268 = ~pi1537 & n20277;
  assign po1714 = n21267 | n21268;
  assign n21270 = ~pi1538 & ~n19347;
  assign n21271 = pi3315 & n19347;
  assign n21272 = ~n21270 & ~n21271;
  assign n21273 = ~n20277 & ~n21272;
  assign n21274 = ~pi1538 & n20277;
  assign po1715 = n21273 | n21274;
  assign n21276 = ~pi1539 & ~n19347;
  assign n21277 = pi3347 & n19347;
  assign n21278 = ~n21276 & ~n21277;
  assign n21279 = ~n20277 & ~n21278;
  assign n21280 = ~pi1539 & n20277;
  assign po1716 = n21279 | n21280;
  assign n21282 = ~pi1540 & ~n19347;
  assign n21283 = pi3316 & n19347;
  assign n21284 = ~n21282 & ~n21283;
  assign n21285 = ~n20277 & ~n21284;
  assign n21286 = ~pi1540 & n20277;
  assign po1717 = n21285 | n21286;
  assign n21288 = ~pi1541 & ~n19347;
  assign n21289 = pi3330 & n19347;
  assign n21290 = ~n21288 & ~n21289;
  assign n21291 = ~n20277 & ~n21290;
  assign n21292 = ~pi1541 & n20277;
  assign po1718 = n21291 | n21292;
  assign n21294 = ~pi1542 & ~n19347;
  assign n21295 = pi3326 & n19347;
  assign n21296 = ~n21294 & ~n21295;
  assign n21297 = ~n20277 & ~n21296;
  assign n21298 = ~pi1542 & n20277;
  assign po1719 = n21297 | n21298;
  assign n21300 = ~pi1543 & ~n19347;
  assign n21301 = pi3295 & n19347;
  assign n21302 = ~n21300 & ~n21301;
  assign n21303 = ~n20277 & ~n21302;
  assign n21304 = ~pi1543 & n20277;
  assign po1720 = n21303 | n21304;
  assign n21306 = ~pi1544 & ~n19347;
  assign n21307 = pi3349 & n19347;
  assign n21308 = ~n21306 & ~n21307;
  assign n21309 = ~n20277 & ~n21308;
  assign n21310 = ~pi1544 & n20277;
  assign po1721 = n21309 | n21310;
  assign n21312 = ~pi1545 & ~n19347;
  assign n21313 = pi3350 & n19347;
  assign n21314 = ~n21312 & ~n21313;
  assign n21315 = ~n20277 & ~n21314;
  assign n21316 = ~pi1545 & n20277;
  assign po1722 = n21315 | n21316;
  assign n21318 = ~pi1546 & ~n19347;
  assign n21319 = pi3354 & n19347;
  assign n21320 = ~n21318 & ~n21319;
  assign n21321 = ~n20277 & ~n21320;
  assign n21322 = ~pi1546 & n20277;
  assign po1723 = n21321 | n21322;
  assign n21324 = ~pi1547 & ~n19347;
  assign n21325 = pi3299 & n19347;
  assign n21326 = ~n21324 & ~n21325;
  assign n21327 = ~n20277 & ~n21326;
  assign n21328 = ~pi1547 & n20277;
  assign po1724 = n21327 | n21328;
  assign n21330 = ~pi1548 & ~n19347;
  assign n21331 = pi2994 & n19347;
  assign n21332 = ~n21330 & ~n21331;
  assign n21333 = ~n20277 & ~n21332;
  assign n21334 = ~pi1548 & n20277;
  assign po1725 = n21333 | n21334;
  assign n21336 = ~pi1549 & ~n19347;
  assign n21337 = pi3311 & n19347;
  assign n21338 = ~n21336 & ~n21337;
  assign n21339 = ~n20277 & ~n21338;
  assign n21340 = ~pi1549 & n20277;
  assign po1726 = n21339 | n21340;
  assign n21342 = ~pi1550 & ~n19347;
  assign n21343 = pi3353 & n19347;
  assign n21344 = ~n21342 & ~n21343;
  assign n21345 = ~n20277 & ~n21344;
  assign n21346 = ~pi1550 & n20277;
  assign po1727 = n21345 | n21346;
  assign n21348 = ~pi1551 & ~n19347;
  assign n21349 = pi3293 & n19347;
  assign n21350 = ~n21348 & ~n21349;
  assign n21351 = ~n20277 & ~n21350;
  assign n21352 = ~pi1551 & n20277;
  assign po1728 = n21351 | n21352;
  assign n21354 = ~pi1552 & ~n19347;
  assign n21355 = pi3313 & n19347;
  assign n21356 = ~n21354 & ~n21355;
  assign n21357 = ~n20277 & ~n21356;
  assign n21358 = ~pi1552 & n20277;
  assign po1729 = n21357 | n21358;
  assign n21360 = ~pi1553 & ~n19347;
  assign n21361 = pi3335 & n19347;
  assign n21362 = ~n21360 & ~n21361;
  assign n21363 = ~n20277 & ~n21362;
  assign n21364 = ~pi1553 & n20277;
  assign po1730 = n21363 | n21364;
  assign n21366 = ~pi1407 & n20503;
  assign n21367 = ~pi1554 & ~n21366;
  assign n21368 = pi3343 & n21366;
  assign n21369 = ~n21367 & ~n21368;
  assign n21370 = ~n20277 & ~n21369;
  assign n21371 = ~pi1554 & n20277;
  assign po1731 = n21370 | n21371;
  assign n21373 = ~pi1555 & ~n21366;
  assign n21374 = pi3287 & n21366;
  assign n21375 = ~n21373 & ~n21374;
  assign n21376 = ~n20277 & ~n21375;
  assign n21377 = ~pi1555 & n20277;
  assign po1732 = n21376 | n21377;
  assign n21379 = ~pi1556 & ~n21366;
  assign n21380 = pi3286 & n21366;
  assign n21381 = ~n21379 & ~n21380;
  assign n21382 = ~n20277 & ~n21381;
  assign n21383 = ~pi1556 & n20277;
  assign po1733 = n21382 | n21383;
  assign n21385 = ~pi1557 & ~n21366;
  assign n21386 = pi3290 & n21366;
  assign n21387 = ~n21385 & ~n21386;
  assign n21388 = ~n20277 & ~n21387;
  assign n21389 = ~pi1557 & n20277;
  assign po1734 = n21388 | n21389;
  assign n21391 = ~pi1558 & ~n21366;
  assign n21392 = pi3315 & n21366;
  assign n21393 = ~n21391 & ~n21392;
  assign n21394 = ~n20277 & ~n21393;
  assign n21395 = ~pi1558 & n20277;
  assign po1735 = n21394 | n21395;
  assign n21397 = ~pi1559 & ~n21366;
  assign n21398 = pi3298 & n21366;
  assign n21399 = ~n21397 & ~n21398;
  assign n21400 = ~n20277 & ~n21399;
  assign n21401 = ~pi1559 & n20277;
  assign po1736 = n21400 | n21401;
  assign n21403 = ~pi1560 & ~n21366;
  assign n21404 = pi3316 & n21366;
  assign n21405 = ~n21403 & ~n21404;
  assign n21406 = ~n20277 & ~n21405;
  assign n21407 = ~pi1560 & n20277;
  assign po1737 = n21406 | n21407;
  assign n21409 = ~pi1561 & ~n21366;
  assign n21410 = pi3333 & n21366;
  assign n21411 = ~n21409 & ~n21410;
  assign n21412 = ~n20277 & ~n21411;
  assign n21413 = ~pi1561 & n20277;
  assign po1738 = n21412 | n21413;
  assign n21415 = ~pi1562 & ~n21366;
  assign n21416 = pi3321 & n21366;
  assign n21417 = ~n21415 & ~n21416;
  assign n21418 = ~n20277 & ~n21417;
  assign n21419 = ~pi1562 & n20277;
  assign po1739 = n21418 | n21419;
  assign n21421 = ~pi1563 & ~n21366;
  assign n21422 = pi3336 & n21366;
  assign n21423 = ~n21421 & ~n21422;
  assign n21424 = ~n20277 & ~n21423;
  assign n21425 = ~pi1563 & n20277;
  assign po1740 = n21424 | n21425;
  assign n21427 = ~pi1564 & ~n21366;
  assign n21428 = pi3318 & n21366;
  assign n21429 = ~n21427 & ~n21428;
  assign n21430 = ~n20277 & ~n21429;
  assign n21431 = ~pi1564 & n20277;
  assign po1741 = n21430 | n21431;
  assign n21433 = ~pi1565 & ~n21366;
  assign n21434 = pi3349 & n21366;
  assign n21435 = ~n21433 & ~n21434;
  assign n21436 = ~n20277 & ~n21435;
  assign n21437 = ~pi1565 & n20277;
  assign po1742 = n21436 | n21437;
  assign n21439 = ~pi1566 & ~n21366;
  assign n21440 = pi3350 & n21366;
  assign n21441 = ~n21439 & ~n21440;
  assign n21442 = ~n20277 & ~n21441;
  assign n21443 = ~pi1566 & n20277;
  assign po1743 = n21442 | n21443;
  assign n21445 = ~pi1567 & ~n21366;
  assign n21446 = pi3355 & n21366;
  assign n21447 = ~n21445 & ~n21446;
  assign n21448 = ~n20277 & ~n21447;
  assign n21449 = ~pi1567 & n20277;
  assign po1744 = n21448 | n21449;
  assign n21451 = ~pi1568 & ~n21366;
  assign n21452 = pi3341 & n21366;
  assign n21453 = ~n21451 & ~n21452;
  assign n21454 = ~n20277 & ~n21453;
  assign n21455 = ~pi1568 & n20277;
  assign po1745 = n21454 | n21455;
  assign n21457 = ~pi1569 & ~n21366;
  assign n21458 = pi3346 & n21366;
  assign n21459 = ~n21457 & ~n21458;
  assign n21460 = ~n20277 & ~n21459;
  assign n21461 = ~pi1569 & n20277;
  assign po1746 = n21460 | n21461;
  assign n21463 = ~pi1570 & ~n21366;
  assign n21464 = pi3311 & n21366;
  assign n21465 = ~n21463 & ~n21464;
  assign n21466 = ~n20277 & ~n21465;
  assign n21467 = ~pi1570 & n20277;
  assign po1747 = n21466 | n21467;
  assign n21469 = ~pi1571 & ~n21366;
  assign n21470 = pi3353 & n21366;
  assign n21471 = ~n21469 & ~n21470;
  assign n21472 = ~n20277 & ~n21471;
  assign n21473 = ~pi1571 & n20277;
  assign po1748 = n21472 | n21473;
  assign n21475 = ~pi1572 & ~n21366;
  assign n21476 = pi3337 & n21366;
  assign n21477 = ~n21475 & ~n21476;
  assign n21478 = ~n20277 & ~n21477;
  assign n21479 = ~pi1572 & n20277;
  assign po1749 = n21478 | n21479;
  assign n21481 = ~pi1573 & ~n21366;
  assign n21482 = pi3335 & n21366;
  assign n21483 = ~n21481 & ~n21482;
  assign n21484 = ~n20277 & ~n21483;
  assign n21485 = ~pi1573 & n20277;
  assign po1750 = n21484 | n21485;
  assign n21487 = ~pi1574 & ~n21011;
  assign n21488 = pi3288 & n21011;
  assign n21489 = ~n21487 & ~n21488;
  assign n21490 = ~n20277 & ~n21489;
  assign n21491 = ~pi1574 & n20277;
  assign po1751 = n21490 | n21491;
  assign n21493 = ~pi1575 & ~n21011;
  assign n21494 = pi3328 & n21011;
  assign n21495 = ~n21493 & ~n21494;
  assign n21496 = ~n20277 & ~n21495;
  assign n21497 = ~pi1575 & n20277;
  assign po1752 = n21496 | n21497;
  assign n21499 = ~pi1576 & ~n20337;
  assign n21500 = pi3299 & n20337;
  assign n21501 = ~n21499 & ~n21500;
  assign n21502 = ~n20277 & ~n21501;
  assign n21503 = ~pi1576 & n20277;
  assign po1753 = n21502 | n21503;
  assign n21505 = ~pi1577 & ~n20337;
  assign n21506 = pi2994 & n20337;
  assign n21507 = ~n21505 & ~n21506;
  assign n21508 = ~n20277 & ~n21507;
  assign n21509 = ~pi1577 & n20277;
  assign po1754 = n21508 | n21509;
  assign n21511 = ~pi1578 & ~n20337;
  assign n21512 = pi3295 & n20337;
  assign n21513 = ~n21511 & ~n21512;
  assign n21514 = ~n20277 & ~n21513;
  assign n21515 = ~pi1578 & n20277;
  assign po1755 = n21514 | n21515;
  assign n21517 = ~pi1579 & ~n20337;
  assign n21518 = pi3349 & n20337;
  assign n21519 = ~n21517 & ~n21518;
  assign n21520 = ~n20277 & ~n21519;
  assign n21521 = ~pi1579 & n20277;
  assign po1756 = n21520 | n21521;
  assign n21523 = ~pi1580 & ~n20337;
  assign n21524 = pi3326 & n20337;
  assign n21525 = ~n21523 & ~n21524;
  assign n21526 = ~n20277 & ~n21525;
  assign n21527 = ~pi1580 & n20277;
  assign po1757 = n21526 | n21527;
  assign n21529 = ~pi1581 & ~n20337;
  assign n21530 = pi3330 & n20337;
  assign n21531 = ~n21529 & ~n21530;
  assign n21532 = ~n20277 & ~n21531;
  assign n21533 = ~pi1581 & n20277;
  assign po1758 = n21532 | n21533;
  assign n21535 = ~pi1582 & ~n20337;
  assign n21536 = pi3316 & n20337;
  assign n21537 = ~n21535 & ~n21536;
  assign n21538 = ~n20277 & ~n21537;
  assign n21539 = ~pi1582 & n20277;
  assign po1759 = n21538 | n21539;
  assign n21541 = ~pi1583 & ~n20337;
  assign n21542 = pi3314 & n20337;
  assign n21543 = ~n21541 & ~n21542;
  assign n21544 = ~n20277 & ~n21543;
  assign n21545 = ~pi1583 & n20277;
  assign po1760 = n21544 | n21545;
  assign n21547 = ~pi1584 & ~n21011;
  assign n21548 = pi3335 & n21011;
  assign n21549 = ~n21547 & ~n21548;
  assign n21550 = ~n20277 & ~n21549;
  assign n21551 = ~pi1584 & n20277;
  assign po1761 = n21550 | n21551;
  assign n21553 = ~pi1585 & ~n20337;
  assign n21554 = pi3288 & n20337;
  assign n21555 = ~n21553 & ~n21554;
  assign n21556 = ~n20277 & ~n21555;
  assign n21557 = ~pi1585 & n20277;
  assign po1762 = n21556 | n21557;
  assign n21559 = ~pi1586 & ~n20337;
  assign n21560 = pi3328 & n20337;
  assign n21561 = ~n21559 & ~n21560;
  assign n21562 = ~n20277 & ~n21561;
  assign n21563 = ~pi1586 & n20277;
  assign po1763 = n21562 | n21563;
  assign n21565 = ~pi1587 & ~n21011;
  assign n21566 = pi3318 & n21011;
  assign n21567 = ~n21565 & ~n21566;
  assign n21568 = ~n20277 & ~n21567;
  assign n21569 = ~pi1587 & n20277;
  assign po1764 = n21568 | n21569;
  assign n21571 = pi3330 & n20330;
  assign n21572 = ~pi1588 & ~n20330;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = ~n20277 & ~n21573;
  assign n21575 = ~pi1588 & n20277;
  assign po1765 = n21574 | n21575;
  assign n21577 = pi1589 & ~n7254;
  assign n21578 = ~pi2972 & pi3131;
  assign n21579 = n20448 & n21578;
  assign n21580 = pi1589 & ~n20450;
  assign n21581 = ~n21579 & ~n21580;
  assign n21582 = n7254 & ~n21581;
  assign po1766 = n21577 | n21582;
  assign n21584 = ~pi1590 & ~n21011;
  assign n21585 = pi3346 & n21011;
  assign n21586 = ~n21584 & ~n21585;
  assign n21587 = ~n20277 & ~n21586;
  assign n21588 = ~pi1590 & n20277;
  assign po1767 = n21587 | n21588;
  assign n21590 = ~pi1591 & ~n21011;
  assign n21591 = pi3353 & n21011;
  assign n21592 = ~n21590 & ~n21591;
  assign n21593 = ~n20277 & ~n21592;
  assign n21594 = ~pi1591 & n20277;
  assign po1768 = n21593 | n21594;
  assign n21596 = ~pi1592 & ~n21011;
  assign n21597 = pi3341 & n21011;
  assign n21598 = ~n21596 & ~n21597;
  assign n21599 = ~n20277 & ~n21598;
  assign n21600 = ~pi1592 & n20277;
  assign po1769 = n21599 | n21600;
  assign n21602 = ~pi1593 & ~n21011;
  assign n21603 = pi3350 & n21011;
  assign n21604 = ~n21602 & ~n21603;
  assign n21605 = ~n20277 & ~n21604;
  assign n21606 = ~pi1593 & n20277;
  assign po1770 = n21605 | n21606;
  assign n21608 = ~pi1594 & ~n21011;
  assign n21609 = pi3336 & n21011;
  assign n21610 = ~n21608 & ~n21609;
  assign n21611 = ~n20277 & ~n21610;
  assign n21612 = ~pi1594 & n20277;
  assign po1771 = n21611 | n21612;
  assign n21614 = pi1595 & ~n7254;
  assign n21615 = n20192 & n21578;
  assign n21616 = pi1595 & ~n20441;
  assign n21617 = ~n21615 & ~n21616;
  assign n21618 = n7254 & ~n21617;
  assign po1772 = n21614 | n21618;
  assign n21620 = ~pi1596 & ~n21011;
  assign n21621 = pi3298 & n21011;
  assign n21622 = ~n21620 & ~n21621;
  assign n21623 = ~n20277 & ~n21622;
  assign n21624 = ~pi1596 & n20277;
  assign po1773 = n21623 | n21624;
  assign n21626 = ~pi1597 & ~n21011;
  assign n21627 = pi3333 & n21011;
  assign n21628 = ~n21626 & ~n21627;
  assign n21629 = ~n20277 & ~n21628;
  assign n21630 = ~pi1597 & n20277;
  assign po1774 = n21629 | n21630;
  assign n21632 = ~pi1598 & ~n21011;
  assign n21633 = pi3315 & n21011;
  assign n21634 = ~n21632 & ~n21633;
  assign n21635 = ~n20277 & ~n21634;
  assign n21636 = ~pi1598 & n20277;
  assign po1775 = n21635 | n21636;
  assign n21638 = pi3311 & n20330;
  assign n21639 = ~pi1599 & ~n20330;
  assign n21640 = ~n21638 & ~n21639;
  assign n21641 = ~n20277 & ~n21640;
  assign n21642 = ~pi1599 & n20277;
  assign po1776 = n21641 | n21642;
  assign n21644 = pi3313 & n20330;
  assign n21645 = ~pi1600 & ~n20330;
  assign n21646 = ~n21644 & ~n21645;
  assign n21647 = ~n20277 & ~n21646;
  assign n21648 = ~pi1600 & n20277;
  assign po1777 = n21647 | n21648;
  assign n21650 = pi3293 & n20330;
  assign n21651 = ~pi1601 & ~n20330;
  assign n21652 = ~n21650 & ~n21651;
  assign n21653 = ~n20277 & ~n21652;
  assign n21654 = ~pi1601 & n20277;
  assign po1778 = n21653 | n21654;
  assign n21656 = pi3299 & n20330;
  assign n21657 = ~pi1602 & ~n20330;
  assign n21658 = ~n21656 & ~n21657;
  assign n21659 = ~n20277 & ~n21658;
  assign n21660 = ~pi1602 & n20277;
  assign po1779 = n21659 | n21660;
  assign n21662 = pi3349 & n20330;
  assign n21663 = ~pi1603 & ~n20330;
  assign n21664 = ~n21662 & ~n21663;
  assign n21665 = ~n20277 & ~n21664;
  assign n21666 = ~pi1603 & n20277;
  assign po1780 = n21665 | n21666;
  assign n21668 = pi3326 & n20330;
  assign n21669 = ~pi1604 & ~n20330;
  assign n21670 = ~n21668 & ~n21669;
  assign n21671 = ~n20277 & ~n21670;
  assign n21672 = ~pi1604 & n20277;
  assign po1781 = n21671 | n21672;
  assign n21674 = ~pi1605 & ~n21366;
  assign n21675 = pi3313 & n21366;
  assign n21676 = ~n21674 & ~n21675;
  assign n21677 = ~n20277 & ~n21676;
  assign n21678 = ~pi1605 & n20277;
  assign po1782 = n21677 | n21678;
  assign n21680 = pi3335 & n20752;
  assign n21681 = ~pi1606 & ~n20752;
  assign n21682 = ~n21680 & ~n21681;
  assign n21683 = ~n20277 & ~n21682;
  assign n21684 = ~pi1606 & n20277;
  assign po1783 = n21683 | n21684;
  assign n21686 = pi3350 & n20752;
  assign n21687 = ~pi1607 & ~n20752;
  assign n21688 = ~n21686 & ~n21687;
  assign n21689 = ~n20277 & ~n21688;
  assign n21690 = ~pi1607 & n20277;
  assign po1784 = n21689 | n21690;
  assign n21692 = pi3340 & n20330;
  assign n21693 = ~pi1608 & ~n20330;
  assign n21694 = ~n21692 & ~n21693;
  assign n21695 = ~n20277 & ~n21694;
  assign n21696 = ~pi1608 & n20277;
  assign po1785 = n21695 | n21696;
  assign n21698 = pi3314 & n20330;
  assign n21699 = ~pi1609 & ~n20330;
  assign n21700 = ~n21698 & ~n21699;
  assign n21701 = ~n20277 & ~n21700;
  assign n21702 = ~pi1609 & n20277;
  assign po1786 = n21701 | n21702;
  assign n21704 = pi3328 & n20330;
  assign n21705 = ~pi1610 & ~n20330;
  assign n21706 = ~n21704 & ~n21705;
  assign n21707 = ~n20277 & ~n21706;
  assign n21708 = ~pi1610 & n20277;
  assign po1787 = n21707 | n21708;
  assign n21710 = pi3353 & n20752;
  assign n21711 = ~pi1611 & ~n20752;
  assign n21712 = ~n21710 & ~n21711;
  assign n21713 = ~n20277 & ~n21712;
  assign n21714 = ~pi1611 & n20277;
  assign po1788 = n21713 | n21714;
  assign n21716 = pi3355 & n20752;
  assign n21717 = ~pi1612 & ~n20752;
  assign n21718 = ~n21716 & ~n21717;
  assign n21719 = ~n20277 & ~n21718;
  assign n21720 = ~pi1612 & n20277;
  assign po1789 = n21719 | n21720;
  assign n21722 = pi3341 & n20752;
  assign n21723 = ~pi1613 & ~n20752;
  assign n21724 = ~n21722 & ~n21723;
  assign n21725 = ~n20277 & ~n21724;
  assign n21726 = ~pi1613 & n20277;
  assign po1790 = n21725 | n21726;
  assign n21728 = pi3336 & n20752;
  assign n21729 = ~pi1614 & ~n20752;
  assign n21730 = ~n21728 & ~n21729;
  assign n21731 = ~n20277 & ~n21730;
  assign n21732 = ~pi1614 & n20277;
  assign po1791 = n21731 | n21732;
  assign n21734 = pi3321 & n20752;
  assign n21735 = ~pi1615 & ~n20752;
  assign n21736 = ~n21734 & ~n21735;
  assign n21737 = ~n20277 & ~n21736;
  assign n21738 = ~pi1615 & n20277;
  assign po1792 = n21737 | n21738;
  assign n21740 = pi3343 & n20752;
  assign n21741 = ~pi1616 & ~n20752;
  assign n21742 = ~n21740 & ~n21741;
  assign n21743 = ~n20277 & ~n21742;
  assign n21744 = ~pi1616 & n20277;
  assign po1793 = n21743 | n21744;
  assign n21746 = ~pi1617 & ~n21011;
  assign n21747 = pi3343 & n21011;
  assign n21748 = ~n21746 & ~n21747;
  assign n21749 = ~n20277 & ~n21748;
  assign n21750 = ~pi1617 & n20277;
  assign po1794 = n21749 | n21750;
  assign n21752 = pi3333 & n20752;
  assign n21753 = ~pi1618 & ~n20752;
  assign n21754 = ~n21752 & ~n21753;
  assign n21755 = ~n20277 & ~n21754;
  assign n21756 = ~pi1618 & n20277;
  assign po1795 = n21755 | n21756;
  assign n21758 = ~pi1619 & ~n21011;
  assign n21759 = pi3287 & n21011;
  assign n21760 = ~n21758 & ~n21759;
  assign n21761 = ~n20277 & ~n21760;
  assign n21762 = ~pi1619 & n20277;
  assign po1796 = n21761 | n21762;
  assign n21764 = pi3286 & n20752;
  assign n21765 = ~pi1620 & ~n20752;
  assign n21766 = ~n21764 & ~n21765;
  assign n21767 = ~n20277 & ~n21766;
  assign n21768 = ~pi1620 & n20277;
  assign po1797 = n21767 | n21768;
  assign n21770 = pi3315 & n20752;
  assign n21771 = ~pi1621 & ~n20752;
  assign n21772 = ~n21770 & ~n21771;
  assign n21773 = ~n20277 & ~n21772;
  assign n21774 = ~pi1621 & n20277;
  assign po1798 = n21773 | n21774;
  assign n21776 = ~pi1622 & ~n21011;
  assign n21777 = pi3286 & n21011;
  assign n21778 = ~n21776 & ~n21777;
  assign n21779 = ~n20277 & ~n21778;
  assign n21780 = ~pi1622 & n20277;
  assign po1799 = n21779 | n21780;
  assign n21782 = pi3290 & n20752;
  assign n21783 = ~pi1623 & ~n20752;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = ~n20277 & ~n21784;
  assign n21786 = ~pi1623 & n20277;
  assign po1800 = n21785 | n21786;
  assign n21788 = pi3354 & n20619;
  assign n21789 = ~pi1624 & ~n20619;
  assign n21790 = ~n21788 & ~n21789;
  assign n21791 = ~n20277 & ~n21790;
  assign n21792 = ~pi1624 & n20277;
  assign po1801 = n21791 | n21792;
  assign n21794 = ~pi1625 & ~n21366;
  assign n21795 = pi3293 & n21366;
  assign n21796 = ~n21794 & ~n21795;
  assign n21797 = ~n20277 & ~n21796;
  assign n21798 = ~pi1625 & n20277;
  assign po1802 = n21797 | n21798;
  assign n21800 = pi3293 & n20619;
  assign n21801 = ~pi1626 & ~n20619;
  assign n21802 = ~n21800 & ~n21801;
  assign n21803 = ~n20277 & ~n21802;
  assign n21804 = ~pi1626 & n20277;
  assign po1803 = n21803 | n21804;
  assign n21806 = ~pi1627 & ~n21366;
  assign n21807 = pi2994 & n21366;
  assign n21808 = ~n21806 & ~n21807;
  assign n21809 = ~n20277 & ~n21808;
  assign n21810 = ~pi1627 & n20277;
  assign po1804 = n21809 | n21810;
  assign n21812 = ~pi1628 & ~n21366;
  assign n21813 = pi3330 & n21366;
  assign n21814 = ~n21812 & ~n21813;
  assign n21815 = ~n20277 & ~n21814;
  assign n21816 = ~pi1628 & n20277;
  assign po1805 = n21815 | n21816;
  assign n21818 = ~pi1629 & ~n21366;
  assign n21819 = pi3299 & n21366;
  assign n21820 = ~n21818 & ~n21819;
  assign n21821 = ~n20277 & ~n21820;
  assign n21822 = ~pi1629 & n20277;
  assign po1806 = n21821 | n21822;
  assign n21824 = ~pi1630 & ~n21366;
  assign n21825 = pi3354 & n21366;
  assign n21826 = ~n21824 & ~n21825;
  assign n21827 = ~n20277 & ~n21826;
  assign n21828 = ~pi1630 & n20277;
  assign po1807 = n21827 | n21828;
  assign n21830 = pi3299 & n20619;
  assign n21831 = ~pi1631 & ~n20619;
  assign n21832 = ~n21830 & ~n21831;
  assign n21833 = ~n20277 & ~n21832;
  assign n21834 = ~pi1631 & n20277;
  assign po1808 = n21833 | n21834;
  assign n21836 = pi2994 & n20619;
  assign n21837 = ~pi1632 & ~n20619;
  assign n21838 = ~n21836 & ~n21837;
  assign n21839 = ~n20277 & ~n21838;
  assign n21840 = ~pi1632 & n20277;
  assign po1809 = n21839 | n21840;
  assign n21842 = ~pi1633 & ~n21366;
  assign n21843 = pi3295 & n21366;
  assign n21844 = ~n21842 & ~n21843;
  assign n21845 = ~n20277 & ~n21844;
  assign n21846 = ~pi1633 & n20277;
  assign po1810 = n21845 | n21846;
  assign n21848 = ~pi1634 & ~n21366;
  assign n21849 = pi3326 & n21366;
  assign n21850 = ~n21848 & ~n21849;
  assign n21851 = ~n20277 & ~n21850;
  assign n21852 = ~pi1634 & n20277;
  assign po1811 = n21851 | n21852;
  assign n21854 = pi3295 & n20619;
  assign n21855 = ~pi1635 & ~n20619;
  assign n21856 = ~n21854 & ~n21855;
  assign n21857 = ~n20277 & ~n21856;
  assign n21858 = ~pi1635 & n20277;
  assign po1812 = n21857 | n21858;
  assign n21860 = ~pi1636 & ~n21366;
  assign n21861 = pi3288 & n21366;
  assign n21862 = ~n21860 & ~n21861;
  assign n21863 = ~n20277 & ~n21862;
  assign n21864 = ~pi1636 & n20277;
  assign po1813 = n21863 | n21864;
  assign n21866 = ~pi1637 & ~n21366;
  assign n21867 = pi3347 & n21366;
  assign n21868 = ~n21866 & ~n21867;
  assign n21869 = ~n20277 & ~n21868;
  assign n21870 = ~pi1637 & n20277;
  assign po1814 = n21869 | n21870;
  assign n21872 = pi3349 & n20619;
  assign n21873 = ~pi1638 & ~n20619;
  assign n21874 = ~n21872 & ~n21873;
  assign n21875 = ~n20277 & ~n21874;
  assign n21876 = ~pi1638 & n20277;
  assign po1815 = n21875 | n21876;
  assign n21878 = ~pi1639 & ~n21366;
  assign n21879 = pi3314 & n21366;
  assign n21880 = ~n21878 & ~n21879;
  assign n21881 = ~n20277 & ~n21880;
  assign n21882 = ~pi1639 & n20277;
  assign po1816 = n21881 | n21882;
  assign n21884 = pi3347 & n20619;
  assign n21885 = ~pi1640 & ~n20619;
  assign n21886 = ~n21884 & ~n21885;
  assign n21887 = ~n20277 & ~n21886;
  assign n21888 = ~pi1640 & n20277;
  assign po1817 = n21887 | n21888;
  assign n21890 = pi3326 & n20619;
  assign n21891 = ~pi1641 & ~n20619;
  assign n21892 = ~n21890 & ~n21891;
  assign n21893 = ~n20277 & ~n21892;
  assign n21894 = ~pi1641 & n20277;
  assign po1818 = n21893 | n21894;
  assign n21896 = ~pi1642 & ~n21366;
  assign n21897 = pi3328 & n21366;
  assign n21898 = ~n21896 & ~n21897;
  assign n21899 = ~n20277 & ~n21898;
  assign n21900 = ~pi1642 & n20277;
  assign po1819 = n21899 | n21900;
  assign n21902 = ~pi1643 & ~n21366;
  assign n21903 = pi3340 & n21366;
  assign n21904 = ~n21902 & ~n21903;
  assign n21905 = ~n20277 & ~n21904;
  assign n21906 = ~pi1643 & n20277;
  assign po1820 = n21905 | n21906;
  assign n21908 = pi3330 & n20619;
  assign n21909 = ~pi1644 & ~n20619;
  assign n21910 = ~n21908 & ~n21909;
  assign n21911 = ~n20277 & ~n21910;
  assign n21912 = ~pi1644 & n20277;
  assign po1821 = n21911 | n21912;
  assign n21914 = pi3340 & n20619;
  assign n21915 = ~pi1645 & ~n20619;
  assign n21916 = ~n21914 & ~n21915;
  assign n21917 = ~n20277 & ~n21916;
  assign n21918 = ~pi1645 & n20277;
  assign po1822 = n21917 | n21918;
  assign n21920 = pi3288 & n20619;
  assign n21921 = ~pi1646 & ~n20619;
  assign n21922 = ~n21920 & ~n21921;
  assign n21923 = ~n20277 & ~n21922;
  assign n21924 = ~pi1646 & n20277;
  assign po1823 = n21923 | n21924;
  assign n21926 = pi3335 & n20504;
  assign n21927 = ~pi1647 & ~n20504;
  assign n21928 = ~n21926 & ~n21927;
  assign n21929 = ~n20277 & ~n21928;
  assign n21930 = ~pi1647 & n20277;
  assign po1824 = n21929 | n21930;
  assign n21932 = ~pi1648 & ~n19347;
  assign n21933 = pi3337 & n19347;
  assign n21934 = ~n21932 & ~n21933;
  assign n21935 = ~n20277 & ~n21934;
  assign n21936 = ~pi1648 & n20277;
  assign po1825 = n21935 | n21936;
  assign n21938 = pi3337 & n20504;
  assign n21939 = ~pi1649 & ~n20504;
  assign n21940 = ~n21938 & ~n21939;
  assign n21941 = ~n20277 & ~n21940;
  assign n21942 = ~pi1649 & n20277;
  assign po1826 = n21941 | n21942;
  assign n21944 = pi3350 & n20504;
  assign n21945 = ~pi1650 & ~n20504;
  assign n21946 = ~n21944 & ~n21945;
  assign n21947 = ~n20277 & ~n21946;
  assign n21948 = ~pi1650 & n20277;
  assign po1827 = n21947 | n21948;
  assign n21950 = pi3355 & n20504;
  assign n21951 = ~pi1651 & ~n20504;
  assign n21952 = ~n21950 & ~n21951;
  assign n21953 = ~n20277 & ~n21952;
  assign n21954 = ~pi1651 & n20277;
  assign po1828 = n21953 | n21954;
  assign n21956 = pi3346 & n20504;
  assign n21957 = ~pi1652 & ~n20504;
  assign n21958 = ~n21956 & ~n21957;
  assign n21959 = ~n20277 & ~n21958;
  assign n21960 = ~pi1652 & n20277;
  assign po1829 = n21959 | n21960;
  assign n21962 = pi3341 & n20504;
  assign n21963 = ~pi1653 & ~n20504;
  assign n21964 = ~n21962 & ~n21963;
  assign n21965 = ~n20277 & ~n21964;
  assign n21966 = ~pi1653 & n20277;
  assign po1830 = n21965 | n21966;
  assign n21968 = pi3318 & n20504;
  assign n21969 = ~pi1654 & ~n20504;
  assign n21970 = ~n21968 & ~n21969;
  assign n21971 = ~n20277 & ~n21970;
  assign n21972 = ~pi1654 & n20277;
  assign po1831 = n21971 | n21972;
  assign n21974 = pi3321 & n20504;
  assign n21975 = ~pi1655 & ~n20504;
  assign n21976 = ~n21974 & ~n21975;
  assign n21977 = ~n20277 & ~n21976;
  assign n21978 = ~pi1655 & n20277;
  assign po1832 = n21977 | n21978;
  assign n21980 = pi3336 & n20504;
  assign n21981 = ~pi1656 & ~n20504;
  assign n21982 = ~n21980 & ~n21981;
  assign n21983 = ~n20277 & ~n21982;
  assign n21984 = ~pi1656 & n20277;
  assign po1833 = n21983 | n21984;
  assign n21986 = pi3286 & n20504;
  assign n21987 = ~pi1657 & ~n20504;
  assign n21988 = ~n21986 & ~n21987;
  assign n21989 = ~n20277 & ~n21988;
  assign n21990 = ~pi1657 & n20277;
  assign po1834 = n21989 | n21990;
  assign n21992 = pi3298 & n20504;
  assign n21993 = ~pi1658 & ~n20504;
  assign n21994 = ~n21992 & ~n21993;
  assign n21995 = ~n20277 & ~n21994;
  assign n21996 = ~pi1658 & n20277;
  assign po1835 = n21995 | n21996;
  assign n21998 = pi3315 & n20504;
  assign n21999 = ~pi1659 & ~n20504;
  assign n22000 = ~n21998 & ~n21999;
  assign n22001 = ~n20277 & ~n22000;
  assign n22002 = ~pi1659 & n20277;
  assign po1836 = n22001 | n22002;
  assign n22004 = pi3290 & n20504;
  assign n22005 = ~pi1660 & ~n20504;
  assign n22006 = ~n22004 & ~n22005;
  assign n22007 = ~n20277 & ~n22006;
  assign n22008 = ~pi1660 & n20277;
  assign po1837 = n22007 | n22008;
  assign n22010 = pi3287 & n20504;
  assign n22011 = ~pi1661 & ~n20504;
  assign n22012 = ~n22010 & ~n22011;
  assign n22013 = ~n20277 & ~n22012;
  assign n22014 = ~pi1661 & n20277;
  assign po1838 = n22013 | n22014;
  assign n22016 = ~pi0327 & n11459;
  assign n22017 = pi1662 & ~n11459;
  assign po1839 = n22016 | n22017;
  assign n22019 = ~pi0296 & n11459;
  assign n22020 = pi1663 & ~n11459;
  assign po1840 = n22019 | n22020;
  assign n22022 = ~pi0297 & n11459;
  assign n22023 = pi1664 & ~n11459;
  assign po1841 = n22022 | n22023;
  assign n22025 = ~pi0330 & n11459;
  assign n22026 = pi1665 & ~n11459;
  assign po1842 = n22025 | n22026;
  assign n22028 = ~pi0294 & n11459;
  assign n22029 = pi1666 & ~n11459;
  assign po1843 = n22028 | n22029;
  assign n22031 = ~pi0292 & n11459;
  assign n22032 = pi1667 & ~n11459;
  assign po1844 = n22031 | n22032;
  assign n22034 = pi2920 & n19984;
  assign n22035 = n20172 & n22034;
  assign n22036 = ~pi2966 & ~pi3001;
  assign n22037 = n7244 & n22036;
  assign n22038 = ~pi2920 & n22037;
  assign n22039 = pi2995 & n22038;
  assign n22040 = ~n22035 & ~n22039;
  assign n22041 = n7254 & ~n22040;
  assign n22042 = ~pi3057 & n22041;
  assign n22043 = pi1668 & ~n22042;
  assign n22044 = ~pi3057 & pi3141;
  assign n22045 = n22041 & n22044;
  assign po1845 = n22043 | n22045;
  assign n22047 = ~pi0288 & n11459;
  assign n22048 = pi1669 & ~n11459;
  assign po1846 = n22047 | n22048;
  assign n22050 = n7254 & n20448;
  assign n22051 = ~pi3057 & n22050;
  assign n22052 = pi1670 & ~n22051;
  assign n22053 = ~pi3057 & pi3146;
  assign n22054 = n22050 & n22053;
  assign po1847 = n22052 | n22054;
  assign n22056 = ~pi0278 & n11459;
  assign n22057 = pi1671 & ~n11459;
  assign po1848 = n22056 | n22057;
  assign n22059 = ~pi0329 & n11459;
  assign n22060 = pi1672 & ~n11459;
  assign po1849 = n22059 | n22060;
  assign n22062 = ~pi0333 & n11459;
  assign n22063 = pi1673 & ~n11459;
  assign po1850 = n22062 | n22063;
  assign n22065 = ~pi0280 & n11459;
  assign n22066 = pi1674 & ~n11459;
  assign po1851 = n22065 | n22066;
  assign n22068 = ~pi0331 & n11459;
  assign n22069 = pi1675 & ~n11459;
  assign po1852 = n22068 | n22069;
  assign n22071 = n9391 & ~n15354;
  assign n22072 = ~n19449 & ~n22071;
  assign po3300 = ~n9382 | n10977;
  assign n22074 = pi2989 & n9384;
  assign n22075 = ~po3300 & n22074;
  assign n22076 = ~n9380 & ~n15360;
  assign n22077 = ~n22075 & n22076;
  assign n22078 = n22072 & n22077;
  assign n22079 = pi1676 & n22078;
  assign n22080 = ~n9380 & ~n9391;
  assign n22081 = ~n22078 & ~n22080;
  assign po1853 = n22079 | n22081;
  assign n22083 = ~pi3018 & n20421;
  assign n22084 = pi1677 & ~n22083;
  assign n22085 = n9530 & n20421;
  assign po1854 = n22084 | n22085;
  assign n22087 = pi1678 & ~n8238;
  assign n22088 = ~n8276 & ~n8293;
  assign n22089 = ~pi1685 & n22088;
  assign n22090 = ~pi1353 & n22089;
  assign n22091 = n8238 & n22090;
  assign n22092 = pi3246 & n22091;
  assign n22093 = pi3149 & n22092;
  assign po1855 = n22087 | n22093;
  assign n22095 = pi1679 & ~n8238;
  assign n22096 = n8238 & ~n18959;
  assign n22097 = pi3246 & n22096;
  assign n22098 = pi3149 & n22097;
  assign n22099 = ~pi1353 & n22098;
  assign po1856 = n22095 | n22099;
  assign n22101 = ~pi1680 & ~n8238;
  assign n22102 = ~pi0502 & pi1334;
  assign n22103 = n9489 & n22102;
  assign n22104 = ~n9489 & ~n22102;
  assign n22105 = ~n22103 & ~n22104;
  assign n22106 = pi1334 & ~n22105;
  assign n22107 = pi1354 & n22106;
  assign n22108 = ~pi0502 & pi1333;
  assign n22109 = n9464 & n22108;
  assign n22110 = ~n9464 & ~n22108;
  assign n22111 = ~n22109 & ~n22110;
  assign n22112 = pi1333 & ~n22111;
  assign n22113 = pi1358 & n22112;
  assign n22114 = ~n22107 & ~n22113;
  assign n22115 = pi3125 & n8238;
  assign n22116 = ~n22114 & n22115;
  assign po1857 = n22101 | n22116;
  assign n22118 = ~pi1681 & ~n8238;
  assign n22119 = pi1355 & n22106;
  assign n22120 = pi1351 & n22112;
  assign n22121 = ~n22119 & ~n22120;
  assign n22122 = n22115 & ~n22121;
  assign po1858 = n22118 | n22122;
  assign n22124 = pi1682 & ~n8238;
  assign n22125 = pi1264 & ~pi2952;
  assign n22126 = ~pi1264 & pi2952;
  assign n22127 = ~n22125 & ~n22126;
  assign n22128 = pi1268 & ~pi2959;
  assign n22129 = ~pi1268 & pi2959;
  assign n22130 = ~n22128 & ~n22129;
  assign n22131 = n22127 & n22130;
  assign n22132 = pi1263 & ~pi2958;
  assign n22133 = ~pi1263 & pi2958;
  assign n22134 = ~n22132 & ~n22133;
  assign n22135 = pi1262 & ~pi2955;
  assign n22136 = ~pi1262 & pi2955;
  assign n22137 = ~n22135 & ~n22136;
  assign n22138 = n22134 & n22137;
  assign n22139 = ~pi0504 & ~pi1186;
  assign n22140 = pi0504 & pi1186;
  assign n22141 = ~n22139 & ~n22140;
  assign n22142 = ~pi0514 & ~pi1187;
  assign n22143 = pi0514 & pi1187;
  assign n22144 = ~n22142 & ~n22143;
  assign n22145 = n22141 & n22144;
  assign n22146 = ~pi0505 & ~pi1192;
  assign n22147 = pi0505 & pi1192;
  assign n22148 = ~n22146 & ~n22147;
  assign n22149 = ~pi0506 & ~pi1149;
  assign n22150 = pi0506 & pi1149;
  assign n22151 = ~n22149 & ~n22150;
  assign n22152 = n22148 & n22151;
  assign n22153 = ~pi0515 & ~pi1185;
  assign n22154 = pi0515 & pi1185;
  assign n22155 = ~n22153 & ~n22154;
  assign n22156 = ~pi0503 & ~pi1155;
  assign n22157 = pi0503 & pi1155;
  assign n22158 = ~n22156 & ~n22157;
  assign n22159 = n22155 & n22158;
  assign n22160 = pi1132 & pi2938;
  assign n22161 = ~pi1132 & ~pi2938;
  assign n22162 = ~n22160 & ~n22161;
  assign n22163 = pi1140 & pi2941;
  assign n22164 = ~pi1140 & ~pi2941;
  assign n22165 = ~n22163 & ~n22164;
  assign n22166 = n22162 & n22165;
  assign n22167 = n22159 & n22166;
  assign n22168 = n22152 & n22167;
  assign n22169 = n22145 & n22168;
  assign n22170 = ~pi0485 & ~pi1134;
  assign n22171 = pi0485 & pi1134;
  assign n22172 = ~n22170 & ~n22171;
  assign n22173 = ~pi0507 & ~pi1151;
  assign n22174 = pi0507 & pi1151;
  assign n22175 = ~n22173 & ~n22174;
  assign n22176 = n22172 & n22175;
  assign n22177 = ~pi0486 & ~pi1133;
  assign n22178 = pi0486 & pi1133;
  assign n22179 = ~n22177 & ~n22178;
  assign n22180 = ~pi0512 & ~pi1150;
  assign n22181 = pi0512 & pi1150;
  assign n22182 = ~n22180 & ~n22181;
  assign n22183 = n22179 & n22182;
  assign n22184 = ~pi0487 & ~pi1135;
  assign n22185 = pi0487 & pi1135;
  assign n22186 = ~n22184 & ~n22185;
  assign n22187 = ~pi0488 & ~pi1193;
  assign n22188 = pi0488 & pi1193;
  assign n22189 = ~n22187 & ~n22188;
  assign n22190 = n22186 & n22189;
  assign n22191 = ~pi0489 & ~pi1136;
  assign n22192 = pi0489 & pi1136;
  assign n22193 = ~n22191 & ~n22192;
  assign n22194 = ~pi0499 & ~pi1183;
  assign n22195 = pi0499 & pi1183;
  assign n22196 = ~n22194 & ~n22195;
  assign n22197 = n22193 & n22196;
  assign n22198 = n22190 & n22197;
  assign n22199 = n22183 & n22198;
  assign n22200 = n22176 & n22199;
  assign n22201 = n22169 & n22200;
  assign n22202 = n8238 & n22201;
  assign n22203 = ~pi0495 & ~pi1142;
  assign n22204 = pi0495 & pi1142;
  assign n22205 = ~n22203 & ~n22204;
  assign n22206 = ~pi0494 & ~pi1158;
  assign n22207 = pi0494 & pi1158;
  assign n22208 = ~n22206 & ~n22207;
  assign n22209 = n22205 & n22208;
  assign n22210 = ~pi0510 & ~pi1184;
  assign n22211 = pi0510 & pi1184;
  assign n22212 = ~n22210 & ~n22211;
  assign n22213 = ~pi0493 & ~pi1141;
  assign n22214 = pi0493 & pi1141;
  assign n22215 = ~n22213 & ~n22214;
  assign n22216 = n22212 & n22215;
  assign n22217 = ~pi0511 & ~pi1157;
  assign n22218 = pi0511 & pi1157;
  assign n22219 = ~n22217 & ~n22218;
  assign n22220 = ~pi0490 & ~pi1137;
  assign n22221 = pi0490 & pi1137;
  assign n22222 = ~n22220 & ~n22221;
  assign n22223 = n22219 & n22222;
  assign n22224 = ~pi0492 & ~pi1139;
  assign n22225 = pi0492 & pi1139;
  assign n22226 = ~n22224 & ~n22225;
  assign n22227 = ~pi0491 & ~pi1138;
  assign n22228 = pi0491 & pi1138;
  assign n22229 = ~n22227 & ~n22228;
  assign n22230 = n22226 & n22229;
  assign n22231 = n22223 & n22230;
  assign n22232 = n22216 & n22231;
  assign n22233 = n22209 & n22232;
  assign n22234 = pi0502 & ~pi1148;
  assign n22235 = ~pi0502 & pi1148;
  assign n22236 = ~n22234 & ~n22235;
  assign n22237 = ~pi0508 & ~pi1146;
  assign n22238 = pi0508 & pi1146;
  assign n22239 = ~n22237 & ~n22238;
  assign n22240 = n22236 & n22239;
  assign n22241 = pi0500 & ~pi1156;
  assign n22242 = ~pi0500 & pi1156;
  assign n22243 = ~n22241 & ~n22242;
  assign n22244 = ~pi0501 & ~pi1147;
  assign n22245 = pi0501 & pi1147;
  assign n22246 = ~n22244 & ~n22245;
  assign n22247 = n22243 & n22246;
  assign n22248 = ~pi0498 & ~pi1145;
  assign n22249 = pi0498 & pi1145;
  assign n22250 = ~n22248 & ~n22249;
  assign n22251 = ~pi0513 & ~pi1144;
  assign n22252 = pi0513 & pi1144;
  assign n22253 = ~n22251 & ~n22252;
  assign n22254 = n22250 & n22253;
  assign n22255 = ~pi0496 & ~pi1143;
  assign n22256 = pi0496 & pi1143;
  assign n22257 = ~n22255 & ~n22256;
  assign n22258 = ~pi0497 & ~pi1191;
  assign n22259 = pi0497 & pi1191;
  assign n22260 = ~n22258 & ~n22259;
  assign n22261 = n22257 & n22260;
  assign n22262 = n22254 & n22261;
  assign n22263 = n22247 & n22262;
  assign n22264 = n22240 & n22263;
  assign n22265 = n22233 & n22264;
  assign n22266 = n22202 & n22265;
  assign n22267 = n22138 & n22266;
  assign n22268 = n22131 & n22267;
  assign po1859 = n22124 | n22268;
  assign n22270 = pi1683 & ~n10977;
  assign n22271 = ~pi0443 & n11155;
  assign n22272 = ~pi1269 & ~n11155;
  assign n22273 = ~n22271 & ~n22272;
  assign n22274 = n10977 & ~n22273;
  assign po1860 = n22270 | n22274;
  assign n22276 = pi2960 & n18959;
  assign n22277 = ~pi1265 & n22276;
  assign n22278 = pi1265 & n18959;
  assign n22279 = ~pi2960 & n22278;
  assign n22280 = ~pi1332 & ~n8224;
  assign n22281 = n22279 & n22280;
  assign n22282 = ~n22277 & ~n22281;
  assign n22283 = n8238 & ~n22282;
  assign n22284 = pi1684 & ~n8238;
  assign po1861 = n22283 | n22284;
  assign n22286 = pi1686 & pi2912;
  assign n22287 = ~pi1685 & ~n22286;
  assign n22288 = pi3148 & ~pi3191;
  assign po1862 = ~n22287 & ~n22288;
  assign n22290 = ~pi2908 & pi3191;
  assign n22291 = ~pi1685 & n22290;
  assign n22292 = ~pi3190 & n22291;
  assign n22293 = pi1686 & ~n22291;
  assign n22294 = ~n22292 & ~n22293;
  assign n22295 = pi0222 & n7068;
  assign n22296 = n7101 & n22295;
  assign n22297 = n7075 & n22296;
  assign n22298 = ~pi2912 & ~n22297;
  assign n22299 = pi1686 & ~n22298;
  assign po1863 = ~n22294 & ~n22299;
  assign n22301 = ~pi2922 & ~pi2923;
  assign n22302 = pi2949 & n22301;
  assign n22303 = pi2946 & n22302;
  assign n22304 = ~pi1688 & ~n22302;
  assign n22305 = ~n22303 & ~n22304;
  assign n22306 = pi1306 & ~n8131;
  assign n22307 = ~n22305 & n22306;
  assign n22308 = ~pi1688 & ~n22306;
  assign po1865 = n22307 | n22308;
  assign n22310 = ~pi2922 & pi2923;
  assign n22311 = pi2949 & n22310;
  assign n22312 = pi2946 & n22311;
  assign n22313 = ~pi1689 & ~n22311;
  assign n22314 = ~n22312 & ~n22313;
  assign n22315 = n22306 & ~n22314;
  assign n22316 = ~pi1689 & ~n22306;
  assign po1866 = n22315 | n22316;
  assign n22318 = ~pi2949 & n22301;
  assign n22319 = ~pi1690 & ~n22318;
  assign n22320 = pi2946 & n22318;
  assign n22321 = ~n22319 & ~n22320;
  assign n22322 = n22306 & ~n22321;
  assign n22323 = ~pi1690 & ~n22306;
  assign po1867 = n22322 | n22323;
  assign n22325 = pi2922 & pi2923;
  assign n22326 = ~pi2949 & n22325;
  assign n22327 = ~pi1691 & ~n22326;
  assign n22328 = pi2946 & n22326;
  assign n22329 = ~n22327 & ~n22328;
  assign n22330 = n22306 & ~n22329;
  assign n22331 = ~pi1691 & ~n22306;
  assign po1868 = n22330 | n22331;
  assign n22333 = pi1692 & n11462;
  assign n22334 = ~pi0444 & pi1858;
  assign n22335 = ~pi2911 & ~n22334;
  assign n22336 = ~n11462 & ~n22335;
  assign po1869 = n22333 | n22336;
  assign n22338 = ~pi1693 & n11462;
  assign n22339 = ~n11462 & ~n19943;
  assign po1870 = n22338 | n22339;
  assign n22341 = pi1694 & n22078;
  assign n22342 = n9382 & ~n9391;
  assign n22343 = ~n22078 & n22342;
  assign po1871 = n22341 | n22343;
  assign n22345 = pi1695 & n22078;
  assign n22346 = ~pi1696 & ~n9389;
  assign n22347 = pi1694 & pi1695;
  assign n22348 = ~pi1697 & ~n22347;
  assign n22349 = n22346 & n22348;
  assign n22350 = ~n9391 & ~n22349;
  assign n22351 = ~n22078 & n22350;
  assign po1872 = n22345 | n22351;
  assign n22353 = pi1696 & n22078;
  assign n22354 = ~pi1232 & n9391;
  assign n22355 = n9380 & ~n9391;
  assign n22356 = ~n22354 & ~n22355;
  assign n22357 = ~n22078 & ~n22356;
  assign po1873 = n22353 | n22357;
  assign n22359 = pi1697 & n22078;
  assign n22360 = pi1232 & n9391;
  assign n22361 = ~n22078 & n22360;
  assign po1874 = n22359 | n22361;
  assign n22363 = pi1698 & n22078;
  assign n22364 = ~pi1694 & ~pi1697;
  assign n22365 = ~pi1696 & n22364;
  assign n22366 = pi1695 & n22365;
  assign n22367 = ~n22078 & ~n22366;
  assign po1875 = n22363 | n22367;
  assign n22369 = pi1699 & ~n22051;
  assign n22370 = n20253 & n22050;
  assign po1876 = n22369 | n22370;
  assign n22372 = pi1700 & ~n22051;
  assign n22373 = ~pi3057 & pi3139;
  assign n22374 = n22050 & n22373;
  assign po1877 = n22372 | n22374;
  assign n22376 = pi1701 & ~n22051;
  assign n22377 = ~pi3057 & pi3168;
  assign n22378 = n22050 & n22377;
  assign po1878 = n22376 | n22378;
  assign n22380 = pi1702 & ~n22051;
  assign n22381 = n22044 & n22050;
  assign po1879 = n22380 | n22381;
  assign n22383 = pi1703 & ~n22051;
  assign n22384 = ~pi3057 & pi3143;
  assign n22385 = n22050 & n22384;
  assign po1880 = n22383 | n22385;
  assign n22387 = pi1704 & ~n22051;
  assign n22388 = ~pi3057 & pi3147;
  assign n22389 = n22050 & n22388;
  assign po1881 = n22387 | n22389;
  assign n22391 = pi1705 & ~n22051;
  assign n22392 = ~pi3057 & pi3153;
  assign n22393 = n22050 & n22392;
  assign po1882 = n22391 | n22393;
  assign n22395 = ~pi2972 & n22050;
  assign n22396 = pi1706 & ~n22395;
  assign n22397 = n20012 & n22050;
  assign po1883 = n22396 | n22397;
  assign n22399 = pi1707 & ~n22042;
  assign n22400 = n22041 & n22388;
  assign po1884 = n22399 | n22400;
  assign n22402 = pi1708 & ~n22395;
  assign n22403 = n19991 & n22050;
  assign po1885 = n22402 | n22403;
  assign n22405 = pi1709 & ~n22395;
  assign n22406 = n19995 & n22050;
  assign po1886 = n22405 | n22406;
  assign n22408 = pi1710 & ~n22042;
  assign n22409 = n22041 & n22384;
  assign po1887 = n22408 | n22409;
  assign n22411 = ~pi3020 & n22041;
  assign n22412 = pi1711 & ~n22411;
  assign n22413 = ~pi3020 & pi3132;
  assign n22414 = n22041 & n22413;
  assign po1888 = n22412 | n22414;
  assign n22416 = pi1712 & ~n22395;
  assign n22417 = n20196 & n22050;
  assign po1889 = n22416 | n22417;
  assign n22419 = pi1713 & ~n22411;
  assign n22420 = ~pi3020 & pi3134;
  assign n22421 = n22041 & n22420;
  assign po1890 = n22419 | n22421;
  assign n22423 = pi1714 & ~n22411;
  assign n22424 = ~pi3020 & pi3155;
  assign n22425 = n22041 & n22424;
  assign po1891 = n22423 | n22425;
  assign n22427 = pi1715 & ~n22411;
  assign n22428 = ~pi3020 & pi3154;
  assign n22429 = n22041 & n22428;
  assign po1892 = n22427 | n22429;
  assign n22431 = pi1716 & ~n22411;
  assign n22432 = ~pi3020 & pi3164;
  assign n22433 = n22041 & n22432;
  assign po1893 = n22431 | n22433;
  assign n22435 = pi1717 & ~n22042;
  assign n22436 = n22041 & n22392;
  assign po1894 = n22435 | n22436;
  assign n22438 = pi1718 & ~n22411;
  assign n22439 = ~pi3020 & pi3171;
  assign n22440 = n22041 & n22439;
  assign po1895 = n22438 | n22440;
  assign n22442 = ~pi3018 & n22041;
  assign n22443 = pi1719 & ~n22442;
  assign n22444 = ~pi3018 & pi3151;
  assign n22445 = n22041 & n22444;
  assign po1896 = n22443 | n22445;
  assign n22447 = pi1720 & ~n22442;
  assign n22448 = n20281 & n22041;
  assign po1897 = n22447 | n22448;
  assign n22450 = pi1721 & ~n22442;
  assign n22451 = n20291 & n22041;
  assign po1898 = n22450 | n22451;
  assign n22453 = pi1722 & ~n22442;
  assign n22454 = n10806 & n22041;
  assign po1899 = n22453 | n22454;
  assign n22456 = pi1723 & ~n22442;
  assign n22457 = n20299 & n22041;
  assign po1900 = n22456 | n22457;
  assign n22459 = ~pi2967 & n7111;
  assign n22460 = n7161 & n22459;
  assign n22461 = ~pi1724 & ~pi1796;
  assign n22462 = pi1724 & pi1796;
  assign n22463 = ~n22461 & ~n22462;
  assign n22464 = n7496 & ~n22463;
  assign n22465 = pi1724 & ~n7496;
  assign n22466 = ~n22464 & ~n22465;
  assign n22467 = ~n22459 & ~n22466;
  assign po1901 = n22460 | n22467;
  assign n22469 = ~n7153 & ~n7161;
  assign n22470 = n22459 & ~n22469;
  assign n22471 = ~pi1725 & ~n22461;
  assign n22472 = pi1725 & n22461;
  assign n22473 = ~n22471 & ~n22472;
  assign n22474 = n7496 & ~n22473;
  assign n22475 = ~pi1725 & ~n7496;
  assign n22476 = ~n22474 & ~n22475;
  assign n22477 = ~n22459 & ~n22476;
  assign po1902 = n22470 | n22477;
  assign n22479 = ~pi0275 & n11459;
  assign n22480 = pi1726 & ~n11459;
  assign po1903 = n22479 | n22480;
  assign n22482 = ~pi0276 & n11459;
  assign n22483 = pi1727 & ~n11459;
  assign po1904 = n22482 | n22483;
  assign n22485 = ~pi0277 & n11459;
  assign n22486 = pi1728 & ~n11459;
  assign po1905 = n22485 | n22486;
  assign n22488 = ~pi0279 & n11459;
  assign n22489 = pi1729 & ~n11459;
  assign po1906 = n22488 | n22489;
  assign n22491 = ~pi0281 & n11459;
  assign n22492 = pi1730 & ~n11459;
  assign po1907 = n22491 | n22492;
  assign n22494 = ~pi0282 & n11459;
  assign n22495 = pi1731 & ~n11459;
  assign po1908 = n22494 | n22495;
  assign n22497 = ~pi0283 & n11459;
  assign n22498 = pi1732 & ~n11459;
  assign po1909 = n22497 | n22498;
  assign n22500 = ~pi0284 & n11459;
  assign n22501 = pi1733 & ~n11459;
  assign po1910 = n22500 | n22501;
  assign n22503 = ~pi0285 & n11459;
  assign n22504 = pi1734 & ~n11459;
  assign po1911 = n22503 | n22504;
  assign n22506 = ~pi0286 & n11459;
  assign n22507 = pi1735 & ~n11459;
  assign po1912 = n22506 | n22507;
  assign n22509 = ~pi0287 & n11459;
  assign n22510 = pi1736 & ~n11459;
  assign po1913 = n22509 | n22510;
  assign n22512 = ~pi0334 & n11459;
  assign n22513 = pi1737 & ~n11459;
  assign po1914 = n22512 | n22513;
  assign n22515 = ~pi0264 & n11459;
  assign n22516 = pi1738 & ~n11459;
  assign po1915 = n22515 | n22516;
  assign n22518 = ~pi0289 & n11459;
  assign n22519 = pi1739 & ~n11459;
  assign po1916 = n22518 | n22519;
  assign n22521 = ~pi0290 & n11459;
  assign n22522 = pi1740 & ~n11459;
  assign po1917 = n22521 | n22522;
  assign n22524 = ~pi0291 & n11459;
  assign n22525 = pi1741 & ~n11459;
  assign po1918 = n22524 | n22525;
  assign n22527 = ~pi0293 & n11459;
  assign n22528 = pi1742 & ~n11459;
  assign po1919 = n22527 | n22528;
  assign n22530 = ~pi0295 & n11459;
  assign n22531 = pi1743 & ~n11459;
  assign po1920 = n22530 | n22531;
  assign n22533 = ~pi0328 & n11459;
  assign n22534 = pi1744 & ~n11459;
  assign po1921 = n22533 | n22534;
  assign n22536 = ~pi0352 & n11459;
  assign n22537 = pi1745 & ~n11459;
  assign po1922 = n22536 | n22537;
  assign n22539 = ~pi2949 & n22310;
  assign n22540 = ~pi1746 & ~n22539;
  assign n22541 = pi2946 & n22539;
  assign n22542 = ~n22540 & ~n22541;
  assign n22543 = n22306 & ~n22542;
  assign n22544 = ~pi1746 & ~n22306;
  assign po1923 = n22543 | n22544;
  assign n22546 = pi2922 & ~pi2923;
  assign n22547 = ~pi2949 & n22546;
  assign n22548 = ~pi1747 & ~n22547;
  assign n22549 = pi2946 & n22547;
  assign n22550 = ~n22548 & ~n22549;
  assign n22551 = n22306 & ~n22550;
  assign n22552 = ~pi1747 & ~n22306;
  assign po1924 = n22551 | n22552;
  assign n22554 = pi2949 & n22325;
  assign n22555 = pi2946 & n22554;
  assign n22556 = ~pi1748 & ~n22554;
  assign n22557 = ~n22555 & ~n22556;
  assign n22558 = n22306 & ~n22557;
  assign n22559 = ~pi1748 & ~n22306;
  assign po1925 = n22558 | n22559;
  assign n22561 = pi2949 & n22546;
  assign n22562 = pi2946 & n22561;
  assign n22563 = ~pi1749 & ~n22561;
  assign n22564 = ~n22562 & ~n22563;
  assign n22565 = n22306 & ~n22564;
  assign n22566 = ~pi1749 & ~n22306;
  assign po1926 = n22565 | n22566;
  assign n22568 = pi1374 & ~pi2948;
  assign n22569 = ~pi3174 & n22568;
  assign n22570 = pi1750 & pi3200;
  assign n22571 = n22569 & n22570;
  assign n22572 = pi1750 & ~n22569;
  assign n22573 = ~pi3200 & n22569;
  assign n22574 = ~n22572 & ~n22573;
  assign n22575 = n19972 & n22574;
  assign po1927 = n22571 | n22575;
  assign n22577 = pi1751 & ~n22442;
  assign n22578 = n9530 & n22041;
  assign po1928 = n22577 | n22578;
  assign n22580 = pi1752 & ~n22442;
  assign n22581 = ~pi3018 & pi3157;
  assign n22582 = n22041 & n22581;
  assign po1929 = n22580 | n22582;
  assign n22584 = pi1753 & ~n22442;
  assign n22585 = n7248 & n22041;
  assign po1930 = n22584 | n22585;
  assign n22587 = pi1754 & ~n22411;
  assign n22588 = ~pi3020 & pi3162;
  assign n22589 = n22041 & n22588;
  assign po1931 = n22587 | n22589;
  assign n22591 = pi1755 & ~n22411;
  assign n22592 = ~pi3020 & pi3165;
  assign n22593 = n22041 & n22592;
  assign po1932 = n22591 | n22593;
  assign n22595 = n19914 & n19984;
  assign n22596 = ~pi2920 & n22595;
  assign n22597 = n7254 & n22596;
  assign n22598 = ~pi3020 & n22597;
  assign n22599 = pi1756 & ~n22598;
  assign n22600 = n22420 & n22597;
  assign po1933 = n22599 | n22600;
  assign n22602 = ~pi3057 & n22597;
  assign n22603 = pi1757 & ~n22602;
  assign n22604 = n22392 & n22597;
  assign po1934 = n22603 | n22604;
  assign n22606 = ~pi3018 & n22597;
  assign n22607 = pi1758 & ~n22606;
  assign n22608 = n7248 & n22597;
  assign po1935 = n22607 | n22608;
  assign n22610 = n7254 & n22036;
  assign n22611 = n7242 & n22610;
  assign n22612 = n9425 & n22611;
  assign n22613 = ~pi3057 & n22612;
  assign n22614 = pi1759 & ~n22613;
  assign n22615 = n22377 & n22612;
  assign po1936 = n22614 | n22615;
  assign n22617 = pi1760 & ~n22613;
  assign n22618 = n22392 & n22612;
  assign po1937 = n22617 | n22618;
  assign n22620 = n9396 & n19970;
  assign n22621 = pi1218 & n22620;
  assign n22622 = pi1337 & ~n22621;
  assign n22623 = pi1269 & pi1310;
  assign n22624 = ~pi1589 & ~pi1712;
  assign n22625 = ~pi1403 & ~pi1404;
  assign n22626 = n22624 & n22625;
  assign n22627 = ~n22623 & n22626;
  assign n22628 = ~pi1337 & ~n22627;
  assign n22629 = ~pi1337 & pi1400;
  assign n22630 = ~n22628 & ~n22629;
  assign n22631 = ~n22622 & ~n22630;
  assign n22632 = ~pi2525 & ~pi2874;
  assign n22633 = ~pi1816 & n22632;
  assign n22634 = ~pi1761 & ~n22633;
  assign n22635 = pi1761 & n22633;
  assign n22636 = ~n22634 & ~n22635;
  assign n22637 = pi1337 & ~n22622;
  assign n22638 = ~n22636 & n22637;
  assign n22639 = ~n22631 & ~n22638;
  assign n22640 = ~pi1761 & n22622;
  assign po1938 = ~n22639 | n22640;
  assign n22642 = pi1762 & ~n8238;
  assign n22643 = pi1363 & n22106;
  assign n22644 = pi1364 & n22112;
  assign n22645 = ~n22643 & ~n22644;
  assign n22646 = n8238 & ~n22645;
  assign po1939 = n22642 | n22646;
  assign n22648 = ~pi3020 & n22612;
  assign n22649 = pi1763 & ~n22648;
  assign n22650 = n22432 & n22612;
  assign po1940 = n22649 | n22650;
  assign n22652 = pi1764 & ~n22648;
  assign n22653 = n22439 & n22612;
  assign po1941 = n22652 | n22653;
  assign n22655 = pi1765 & ~n22648;
  assign n22656 = n22424 & n22612;
  assign po1942 = n22655 | n22656;
  assign n22658 = pi1766 & ~n22648;
  assign n22659 = n22588 & n22612;
  assign po1943 = n22658 | n22659;
  assign n22661 = pi1767 & ~n22648;
  assign n22662 = n22428 & n22612;
  assign po1944 = n22661 | n22662;
  assign n22664 = ~pi3018 & n22612;
  assign n22665 = pi1768 & ~n22664;
  assign n22666 = n22444 & n22612;
  assign po1945 = n22665 | n22666;
  assign n22668 = pi1769 & ~n22664;
  assign n22669 = n22581 & n22612;
  assign po1946 = n22668 | n22669;
  assign n22671 = pi1770 & ~n22664;
  assign n22672 = n20281 & n22612;
  assign po1947 = n22671 | n22672;
  assign n22674 = pi1771 & ~n22664;
  assign n22675 = n20299 & n22612;
  assign po1948 = n22674 | n22675;
  assign n22677 = pi1772 & ~n22664;
  assign n22678 = n10806 & n22612;
  assign po1949 = n22677 | n22678;
  assign n22680 = pi1773 & ~n22613;
  assign n22681 = n22373 & n22612;
  assign po1950 = n22680 | n22681;
  assign n22683 = pi1774 & ~n22613;
  assign n22684 = n22044 & n22612;
  assign po1951 = n22683 | n22684;
  assign n22686 = pi1775 & ~n22613;
  assign n22687 = n22384 & n22612;
  assign po1952 = n22686 | n22687;
  assign n22689 = pi1776 & ~n22613;
  assign n22690 = n22388 & n22612;
  assign po1953 = n22689 | n22690;
  assign n22692 = pi1777 & ~n22648;
  assign n22693 = n22420 & n22612;
  assign po1954 = n22692 | n22693;
  assign n22695 = pi1779 & ~n22598;
  assign n22696 = n22588 & n22597;
  assign po1956 = n22695 | n22696;
  assign n22698 = pi1780 & ~n22602;
  assign n22699 = n22373 & n22597;
  assign po1957 = n22698 | n22699;
  assign n22701 = pi1781 & ~n22602;
  assign n22702 = n22044 & n22597;
  assign po1958 = n22701 | n22702;
  assign n22704 = pi1782 & ~n22602;
  assign n22705 = n22377 & n22597;
  assign po1959 = n22704 | n22705;
  assign n22707 = pi1783 & ~n22602;
  assign n22708 = n22384 & n22597;
  assign po1960 = n22707 | n22708;
  assign n22710 = pi1784 & ~n22598;
  assign n22711 = n22432 & n22597;
  assign po1961 = n22710 | n22711;
  assign n22713 = pi1785 & ~n22598;
  assign n22714 = n22413 & n22597;
  assign po1962 = n22713 | n22714;
  assign n22716 = pi1786 & ~n22598;
  assign n22717 = n22424 & n22597;
  assign po1963 = n22716 | n22717;
  assign n22719 = pi1787 & ~n22602;
  assign n22720 = n22388 & n22597;
  assign po1964 = n22719 | n22720;
  assign n22722 = pi1788 & ~n22598;
  assign n22723 = n22592 & n22597;
  assign po1965 = n22722 | n22723;
  assign n22725 = pi1789 & ~n22598;
  assign n22726 = n22428 & n22597;
  assign po1966 = n22725 | n22726;
  assign n22728 = pi1790 & ~n22606;
  assign n22729 = n22444 & n22597;
  assign po1967 = n22728 | n22729;
  assign n22731 = pi1791 & ~n22598;
  assign n22732 = n22439 & n22597;
  assign po1968 = n22731 | n22732;
  assign n22734 = pi1792 & ~n22606;
  assign n22735 = n20299 & n22597;
  assign po1969 = n22734 | n22735;
  assign n22737 = pi1793 & ~n22606;
  assign n22738 = n9530 & n22597;
  assign po1970 = n22737 | n22738;
  assign n22740 = pi1794 & ~n22606;
  assign n22741 = n10806 & n22597;
  assign po1971 = n22740 | n22741;
  assign n22743 = pi1795 & ~n22606;
  assign n22744 = n20291 & n22597;
  assign po1972 = n22743 | n22744;
  assign n22746 = pi1796 & ~n7496;
  assign n22747 = ~pi1796 & n7496;
  assign n22748 = ~n22746 & ~n22747;
  assign n22749 = ~n22459 & ~n22748;
  assign n22750 = ~n7159 & n22459;
  assign po1973 = n22749 | n22750;
  assign n22752 = pi1797 & ~n22664;
  assign n22753 = n9530 & n22612;
  assign po1974 = n22752 | n22753;
  assign n22755 = n8238 & n22112;
  assign n22756 = pi1798 & ~n8238;
  assign po1975 = n22755 | n22756;
  assign n22758 = pi1799 & ~n22613;
  assign n22759 = n20253 & n22612;
  assign po1976 = n22758 | n22759;
  assign n22761 = pi1800 & ~n22613;
  assign n22762 = n22053 & n22612;
  assign po1977 = n22761 | n22762;
  assign n22764 = pi1801 & ~n22648;
  assign n22765 = n22592 & n22612;
  assign po1978 = n22764 | n22765;
  assign n22767 = pi1802 & ~n22664;
  assign n22768 = n20291 & n22612;
  assign po1979 = n22767 | n22768;
  assign n22770 = pi1803 & ~n22664;
  assign n22771 = n7248 & n22612;
  assign po1980 = n22770 | n22771;
  assign n22773 = pi1804 & ~n22648;
  assign n22774 = n22413 & n22612;
  assign po1981 = n22773 | n22774;
  assign n22776 = n9396 & ~n10977;
  assign n22777 = n9402 & n22776;
  assign n22778 = ~n10978 & ~n22777;
  assign n22779 = ~n19461 & ~n22778;
  assign n22780 = pi1805 & n22778;
  assign po1982 = n22779 | n22780;
  assign n22782 = n8238 & n22106;
  assign n22783 = pi1806 & ~n8238;
  assign po1983 = n22782 | n22783;
  assign n22785 = pi1807 & ~n22606;
  assign n22786 = n22581 & n22597;
  assign po1984 = n22785 | n22786;
  assign n22788 = pi1808 & ~n22602;
  assign n22789 = n20253 & n22597;
  assign po1985 = n22788 | n22789;
  assign n22791 = pi1809 & ~n22602;
  assign n22792 = n22053 & n22597;
  assign po1986 = n22791 | n22792;
  assign n22794 = pi1810 & ~n22606;
  assign n22795 = n20281 & n22597;
  assign po1987 = n22794 | n22795;
  assign po1988 = n8238 | n8305;
  assign n22798 = pi2920 & n7254;
  assign n22799 = n22595 & n22798;
  assign n22800 = ~pi3057 & n22799;
  assign n22801 = pi1812 & ~n22800;
  assign n22802 = n22373 & n22799;
  assign po1989 = n22801 | n22802;
  assign n22804 = pi1813 & ~n7496;
  assign n22805 = n7184 & n7496;
  assign n22806 = ~n22804 & ~n22805;
  assign po1990 = ~n22459 & ~n22806;
  assign n22808 = ~pi3018 & n22799;
  assign n22809 = pi1814 & ~n22808;
  assign n22810 = n20299 & n22799;
  assign po1991 = n22809 | n22810;
  assign n22812 = ~pi3020 & n22799;
  assign n22813 = pi1815 & ~n22812;
  assign n22814 = n22420 & n22799;
  assign po1992 = n22813 | n22814;
  assign n22816 = ~pi1816 & n22622;
  assign n22817 = ~pi1337 & pi1709;
  assign n22818 = ~n22628 & ~n22817;
  assign n22819 = ~n22622 & n22818;
  assign n22820 = ~n22816 & ~n22819;
  assign n22821 = pi1816 & ~n22632;
  assign n22822 = ~n22633 & ~n22821;
  assign n22823 = n22637 & ~n22822;
  assign po1993 = n22820 | n22823;
  assign n22825 = pi1817 & ~n22812;
  assign n22826 = n22413 & n22799;
  assign po1994 = n22825 | n22826;
  assign n22828 = pi1818 & ~n22812;
  assign n22829 = n22432 & n22799;
  assign po1995 = n22828 | n22829;
  assign n22831 = pi1819 & ~n22812;
  assign n22832 = n22424 & n22799;
  assign po1996 = n22831 | n22832;
  assign n22834 = pi1820 & ~n22812;
  assign n22835 = n22588 & n22799;
  assign po1997 = n22834 | n22835;
  assign n22837 = pi1821 & ~n22808;
  assign n22838 = n7248 & n22799;
  assign po1998 = n22837 | n22838;
  assign n22840 = pi1822 & ~n22812;
  assign n22841 = n22428 & n22799;
  assign po1999 = n22840 | n22841;
  assign n22843 = pi1823 & ~n22808;
  assign n22844 = n10806 & n22799;
  assign po2000 = n22843 | n22844;
  assign n22846 = pi1824 & ~n22808;
  assign n22847 = n20291 & n22799;
  assign po2001 = n22846 | n22847;
  assign n22849 = pi1825 & ~n22808;
  assign n22850 = n9530 & n22799;
  assign po2002 = n22849 | n22850;
  assign n22852 = pi1826 & ~n22800;
  assign n22853 = n22388 & n22799;
  assign po2003 = n22852 | n22853;
  assign n22855 = ~pi1692 & n20262;
  assign n22856 = ~pi1805 & n22855;
  assign n22857 = ~pi1827 & n22856;
  assign n22858 = pi0444 & pi1827;
  assign po2004 = n22857 | n22858;
  assign n22860 = ~n19957 & n19970;
  assign n22861 = pi1828 & ~n22860;
  assign n22862 = ~n19160 & n22860;
  assign po2005 = n22861 | n22862;
  assign n22864 = ~pi1829 & ~n22860;
  assign n22865 = pi1828 & ~pi1985;
  assign n22866 = pi1983 & ~pi1984;
  assign n22867 = n22865 & n22866;
  assign n22868 = ~pi1829 & ~n22867;
  assign n22869 = ~pi0305 & pi0306;
  assign n22870 = pi1683 & n22869;
  assign n22871 = n19955 & ~n22870;
  assign n22872 = ~n19954 & ~n22871;
  assign n22873 = n22867 & ~n22872;
  assign n22874 = ~n22868 & ~n22873;
  assign n22875 = n22860 & ~n22874;
  assign po2006 = n22864 | n22875;
  assign n22877 = ~pi1830 & ~n22860;
  assign n22878 = pi1983 & pi1984;
  assign n22879 = n22865 & n22878;
  assign n22880 = ~n22872 & n22879;
  assign n22881 = ~pi1830 & ~n22879;
  assign n22882 = ~n22880 & ~n22881;
  assign n22883 = n22860 & ~n22882;
  assign po2007 = n22877 | n22883;
  assign n22885 = ~pi1831 & ~n22860;
  assign n22886 = n19071 & n22866;
  assign n22887 = ~pi1831 & ~n22886;
  assign n22888 = ~n22872 & n22886;
  assign n22889 = ~n22887 & ~n22888;
  assign n22890 = n22860 & ~n22889;
  assign po2008 = n22885 | n22890;
  assign n22892 = ~pi1832 & ~n22860;
  assign n22893 = n19071 & n22878;
  assign n22894 = ~n22872 & n22893;
  assign n22895 = ~pi1832 & ~n22893;
  assign n22896 = ~n22894 & ~n22895;
  assign n22897 = n22860 & ~n22896;
  assign po2009 = n22892 | n22897;
  assign n22899 = ~pi1833 & ~n22860;
  assign n22900 = n19179 & n22866;
  assign n22901 = ~n22872 & n22900;
  assign n22902 = ~pi1833 & ~n22900;
  assign n22903 = ~n22901 & ~n22902;
  assign n22904 = n22860 & ~n22903;
  assign po2010 = n22899 | n22904;
  assign n22906 = ~pi1834 & ~n22860;
  assign n22907 = ~pi1983 & pi1984;
  assign n22908 = ~pi1828 & ~pi1985;
  assign n22909 = n22907 & n22908;
  assign n22910 = ~pi1834 & ~n22909;
  assign n22911 = ~n22872 & n22909;
  assign n22912 = ~n22910 & ~n22911;
  assign n22913 = n22860 & ~n22912;
  assign po2011 = n22906 | n22913;
  assign n22915 = ~pi1835 & ~n22860;
  assign n22916 = ~pi1983 & ~pi1984;
  assign n22917 = n22865 & n22916;
  assign n22918 = ~pi1835 & ~n22917;
  assign n22919 = ~n22872 & n22917;
  assign n22920 = ~n22918 & ~n22919;
  assign n22921 = n22860 & ~n22920;
  assign po2012 = n22915 | n22921;
  assign n22923 = ~pi1836 & ~n22860;
  assign n22924 = n22865 & n22907;
  assign n22925 = ~pi1836 & ~n22924;
  assign n22926 = ~n22872 & n22924;
  assign n22927 = ~n22925 & ~n22926;
  assign n22928 = n22860 & ~n22927;
  assign po2013 = n22923 | n22928;
  assign n22930 = ~pi1837 & ~n22860;
  assign n22931 = n19071 & n22916;
  assign n22932 = ~pi1837 & ~n22931;
  assign n22933 = ~n22872 & n22931;
  assign n22934 = ~n22932 & ~n22933;
  assign n22935 = n22860 & ~n22934;
  assign po2014 = n22930 | n22935;
  assign n22937 = ~pi1838 & ~n22860;
  assign n22938 = n19179 & n22907;
  assign n22939 = ~n22872 & n22938;
  assign n22940 = ~pi1838 & ~n22938;
  assign n22941 = ~n22939 & ~n22940;
  assign n22942 = n22860 & ~n22941;
  assign po2015 = n22937 | n22942;
  assign n22944 = ~pi1839 & ~n22860;
  assign n22945 = n22866 & n22908;
  assign n22946 = ~pi1839 & ~n22945;
  assign n22947 = ~n22872 & n22945;
  assign n22948 = ~n22946 & ~n22947;
  assign n22949 = n22860 & ~n22948;
  assign po2016 = n22944 | n22949;
  assign n22951 = ~pi1840 & ~n22860;
  assign n22952 = n22878 & n22908;
  assign n22953 = ~pi1840 & ~n22952;
  assign n22954 = ~n22872 & n22952;
  assign n22955 = ~n22953 & ~n22954;
  assign n22956 = n22860 & ~n22955;
  assign po2017 = n22951 | n22956;
  assign n22958 = ~pi1841 & ~n22860;
  assign n22959 = n22908 & n22916;
  assign n22960 = ~pi1841 & ~n22959;
  assign n22961 = ~n22872 & n22959;
  assign n22962 = ~n22960 & ~n22961;
  assign n22963 = n22860 & ~n22962;
  assign po2018 = n22958 | n22963;
  assign n22965 = ~pi1842 & ~n22860;
  assign n22966 = n19071 & n22907;
  assign n22967 = ~pi1842 & ~n22966;
  assign n22968 = ~n22872 & n22966;
  assign n22969 = ~n22967 & ~n22968;
  assign n22970 = n22860 & ~n22969;
  assign po2019 = n22965 | n22970;
  assign n22972 = ~pi1843 & ~n22860;
  assign n22973 = n19179 & n22916;
  assign n22974 = ~pi1843 & ~n22973;
  assign n22975 = ~n22872 & n22973;
  assign n22976 = ~n22974 & ~n22975;
  assign n22977 = n22860 & ~n22976;
  assign po2020 = n22972 | n22977;
  assign n22979 = ~pi1844 & ~n22860;
  assign n22980 = n19179 & n22878;
  assign n22981 = ~n22872 & n22980;
  assign n22982 = ~pi1844 & ~n22980;
  assign n22983 = ~n22981 & ~n22982;
  assign n22984 = n22860 & ~n22983;
  assign po2021 = n22979 | n22984;
  assign n22986 = pi1845 & ~n22800;
  assign n22987 = n22377 & n22799;
  assign po2022 = n22986 | n22987;
  assign n22989 = pi1846 & ~n22800;
  assign n22990 = n22384 & n22799;
  assign po2023 = n22989 | n22990;
  assign n22992 = pi1847 & ~n22800;
  assign n22993 = n22392 & n22799;
  assign po2024 = n22992 | n22993;
  assign n22995 = pi1848 & ~n22800;
  assign n22996 = n22044 & n22799;
  assign po2025 = n22995 | n22996;
  assign n22998 = pi1849 & ~n22800;
  assign n22999 = n20253 & n22799;
  assign po2026 = n22998 | n22999;
  assign n23001 = pi1850 & ~n22800;
  assign n23002 = n22053 & n22799;
  assign po2027 = n23001 | n23002;
  assign n23004 = pi1851 & ~n22808;
  assign n23005 = n20281 & n22799;
  assign po2028 = n23004 | n23005;
  assign n23007 = pi1852 & ~n22808;
  assign n23008 = n22581 & n22799;
  assign po2029 = n23007 | n23008;
  assign n23010 = pi1853 & ~n22808;
  assign n23011 = n22444 & n22799;
  assign po2030 = n23010 | n23011;
  assign n23013 = pi1854 & ~n22812;
  assign n23014 = n22592 & n22799;
  assign po2031 = n23013 | n23014;
  assign n23016 = pi1855 & ~n22812;
  assign n23017 = n22439 & n22799;
  assign po2032 = n23016 | n23017;
  assign n23019 = pi2976 & n22554;
  assign n23020 = ~pi1856 & ~n22554;
  assign n23021 = ~n23019 & ~n23020;
  assign n23022 = n22306 & ~n23021;
  assign n23023 = ~pi1856 & ~n22306;
  assign po2033 = n23022 | n23023;
  assign n23025 = pi2976 & n22311;
  assign n23026 = ~pi1857 & ~n22311;
  assign n23027 = ~n23025 & ~n23026;
  assign n23028 = n22306 & ~n23027;
  assign n23029 = ~pi1857 & ~n22306;
  assign po2034 = n23028 | n23029;
  assign n23031 = ~n19955 & n19960;
  assign n23032 = n9402 & ~n23031;
  assign n23033 = pi1858 & ~n23032;
  assign po2035 = n11155 | n23033;
  assign n23035 = n15368 & n22360;
  assign n23036 = ~pi3027 & n23035;
  assign n23037 = ~pi3201 & n23036;
  assign n23038 = ~n22075 & ~n23037;
  assign n23039 = ~n22354 & n23038;
  assign po2036 = ~n9380 & n23039;
  assign n23041 = pi3437 & n15250;
  assign n23042 = ~pi1860 & ~n15250;
  assign n23043 = ~n23041 & ~n23042;
  assign n23044 = ~pi0509 & ~n23043;
  assign n23045 = pi0509 & ~pi1860;
  assign po2037 = n23044 | n23045;
  assign n23047 = pi3427 & n15250;
  assign n23048 = ~pi1861 & ~n15250;
  assign n23049 = ~n23047 & ~n23048;
  assign n23050 = ~pi0509 & ~n23049;
  assign n23051 = pi0509 & ~pi1861;
  assign po2038 = n23050 | n23051;
  assign n23053 = pi3429 & n15250;
  assign n23054 = ~pi1862 & ~n15250;
  assign n23055 = ~n23053 & ~n23054;
  assign n23056 = ~pi0509 & ~n23055;
  assign n23057 = pi0509 & ~pi1862;
  assign po2039 = n23056 | n23057;
  assign n23059 = pi3430 & n15250;
  assign n23060 = ~pi1863 & ~n15250;
  assign n23061 = ~n23059 & ~n23060;
  assign n23062 = ~pi0509 & ~n23061;
  assign n23063 = pi0509 & ~pi1863;
  assign po2040 = n23062 | n23063;
  assign n23065 = pi3432 & n15250;
  assign n23066 = ~pi1864 & ~n15250;
  assign n23067 = ~n23065 & ~n23066;
  assign n23068 = ~pi0509 & ~n23067;
  assign n23069 = pi0509 & ~pi1864;
  assign po2041 = n23068 | n23069;
  assign n23071 = pi3433 & n15250;
  assign n23072 = ~pi1865 & ~n15250;
  assign n23073 = ~n23071 & ~n23072;
  assign n23074 = ~pi0509 & ~n23073;
  assign n23075 = pi0509 & ~pi1865;
  assign po2042 = n23074 | n23075;
  assign n23077 = pi3434 & n15250;
  assign n23078 = ~pi1866 & ~n15250;
  assign n23079 = ~n23077 & ~n23078;
  assign n23080 = ~pi0509 & ~n23079;
  assign n23081 = pi0509 & ~pi1866;
  assign po2043 = n23080 | n23081;
  assign n23083 = pi3438 & n15250;
  assign n23084 = ~pi1867 & ~n15250;
  assign n23085 = ~n23083 & ~n23084;
  assign n23086 = ~pi0509 & ~n23085;
  assign n23087 = pi0509 & ~pi1867;
  assign po2044 = n23086 | n23087;
  assign n23089 = pi3439 & n15250;
  assign n23090 = ~pi1868 & ~n15250;
  assign n23091 = ~n23089 & ~n23090;
  assign n23092 = ~pi0509 & ~n23091;
  assign n23093 = pi0509 & ~pi1868;
  assign po2045 = n23092 | n23093;
  assign n23095 = pi3412 & n15250;
  assign n23096 = ~pi1869 & ~n15250;
  assign n23097 = ~n23095 & ~n23096;
  assign n23098 = ~pi0509 & ~n23097;
  assign n23099 = pi0509 & ~pi1869;
  assign po2046 = n23098 | n23099;
  assign n23101 = pi3441 & n15250;
  assign n23102 = ~pi1870 & ~n15250;
  assign n23103 = ~n23101 & ~n23102;
  assign n23104 = ~pi0509 & ~n23103;
  assign n23105 = pi0509 & ~pi1870;
  assign po2047 = n23104 | n23105;
  assign n23107 = pi3413 & n15250;
  assign n23108 = ~pi1871 & ~n15250;
  assign n23109 = ~n23107 & ~n23108;
  assign n23110 = ~pi0509 & ~n23109;
  assign n23111 = pi0509 & ~pi1871;
  assign po2048 = n23110 | n23111;
  assign n23113 = pi3414 & n15250;
  assign n23114 = ~pi1872 & ~n15250;
  assign n23115 = ~n23113 & ~n23114;
  assign n23116 = ~pi0509 & ~n23115;
  assign n23117 = pi0509 & ~pi1872;
  assign po2049 = n23116 | n23117;
  assign n23119 = pi3416 & n15250;
  assign n23120 = ~pi1873 & ~n15250;
  assign n23121 = ~n23119 & ~n23120;
  assign n23122 = ~pi0509 & ~n23121;
  assign n23123 = pi0509 & ~pi1873;
  assign po2050 = n23122 | n23123;
  assign n23125 = pi3418 & n15250;
  assign n23126 = ~pi1874 & ~n15250;
  assign n23127 = ~n23125 & ~n23126;
  assign n23128 = ~pi0509 & ~n23127;
  assign n23129 = pi0509 & ~pi1874;
  assign po2051 = n23128 | n23129;
  assign n23131 = pi3426 & n15250;
  assign n23132 = ~pi1875 & ~n15250;
  assign n23133 = ~n23131 & ~n23132;
  assign n23134 = ~pi0509 & ~n23133;
  assign n23135 = pi0509 & ~pi1875;
  assign po2052 = n23134 | n23135;
  assign n23137 = pi3424 & n15250;
  assign n23138 = ~pi1876 & ~n15250;
  assign n23139 = ~n23137 & ~n23138;
  assign n23140 = ~pi0509 & ~n23139;
  assign n23141 = pi0509 & ~pi1876;
  assign po2053 = n23140 | n23141;
  assign n23143 = ~pi1877 & ~n22860;
  assign po2054 = n22862 | n23143;
  assign n23145 = n9386 & ~n23037;
  assign n23146 = ~n15361 & ~n22354;
  assign po2158 = n23145 & n23146;
  assign n23148 = pi2976 & n22561;
  assign n23149 = ~pi1879 & ~n22561;
  assign n23150 = ~n23148 & ~n23149;
  assign n23151 = n22306 & ~n23150;
  assign n23152 = ~pi1879 & ~n22306;
  assign po2056 = n23151 | n23152;
  assign n23154 = pi2976 & n22302;
  assign n23155 = ~pi1880 & ~n22302;
  assign n23156 = ~n23154 & ~n23155;
  assign n23157 = n22306 & ~n23156;
  assign n23158 = ~pi1880 & ~n22306;
  assign po2057 = n23157 | n23158;
  assign n23160 = ~pi1881 & ~n22318;
  assign n23161 = pi2976 & n22318;
  assign n23162 = ~n23160 & ~n23161;
  assign n23163 = n22306 & ~n23162;
  assign n23164 = ~pi1881 & ~n22306;
  assign po2058 = n23163 | n23164;
  assign n23166 = ~pi1882 & ~n22547;
  assign n23167 = pi2976 & n22547;
  assign n23168 = ~n23166 & ~n23167;
  assign n23169 = n22306 & ~n23168;
  assign n23170 = ~pi1882 & ~n22306;
  assign po2059 = n23169 | n23170;
  assign n23172 = ~pi3082 & n22539;
  assign n23173 = ~pi1883 & ~n22539;
  assign n23174 = ~n23172 & ~n23173;
  assign n23175 = n22306 & ~n23174;
  assign n23176 = ~pi1883 & ~n22306;
  assign po2060 = n23175 | n23176;
  assign n23178 = ~pi1884 & ~n22326;
  assign n23179 = pi2976 & n22326;
  assign n23180 = ~n23178 & ~n23179;
  assign n23181 = n22306 & ~n23180;
  assign n23182 = ~pi1884 & ~n22306;
  assign po2061 = n23181 | n23182;
  assign n23184 = pi3423 & n15250;
  assign n23185 = ~pi1885 & ~n15250;
  assign n23186 = ~n23184 & ~n23185;
  assign n23187 = ~pi0509 & ~n23186;
  assign n23188 = pi0509 & ~pi1885;
  assign po2062 = n23187 | n23188;
  assign n23190 = pi3425 & n15250;
  assign n23191 = ~pi1886 & ~n15250;
  assign n23192 = ~n23190 & ~n23191;
  assign n23193 = ~pi0509 & ~n23192;
  assign n23194 = pi0509 & ~pi1886;
  assign po2063 = n23193 | n23194;
  assign n23196 = pi3419 & n15250;
  assign n23197 = ~pi1887 & ~n15250;
  assign n23198 = ~n23196 & ~n23197;
  assign n23199 = ~pi0509 & ~n23198;
  assign n23200 = pi0509 & ~pi1887;
  assign po2064 = n23199 | n23200;
  assign n23202 = pi3415 & n15250;
  assign n23203 = ~pi1888 & ~n15250;
  assign n23204 = ~n23202 & ~n23203;
  assign n23205 = ~pi0509 & ~n23204;
  assign n23206 = pi0509 & ~pi1888;
  assign po2065 = n23205 | n23206;
  assign n23208 = pi3417 & n15250;
  assign n23209 = ~pi1889 & ~n15250;
  assign n23210 = ~n23208 & ~n23209;
  assign n23211 = ~pi0509 & ~n23210;
  assign n23212 = pi0509 & ~pi1889;
  assign po2066 = n23211 | n23212;
  assign n23214 = ~pi3082 & n22547;
  assign n23215 = ~pi1890 & ~n22547;
  assign n23216 = ~n23214 & ~n23215;
  assign n23217 = n22306 & ~n23216;
  assign n23218 = ~pi1890 & ~n22306;
  assign po2067 = n23217 | n23218;
  assign n23220 = pi3436 & n15250;
  assign n23221 = ~pi1891 & ~n15250;
  assign n23222 = ~n23220 & ~n23221;
  assign n23223 = ~pi0509 & ~n23222;
  assign n23224 = pi0509 & ~pi1891;
  assign po2068 = n23223 | n23224;
  assign n23226 = pi3440 & n15250;
  assign n23227 = ~pi1892 & ~n15250;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = ~pi0509 & ~n23228;
  assign n23230 = pi0509 & ~pi1892;
  assign po2069 = n23229 | n23230;
  assign n23232 = pi3428 & n15250;
  assign n23233 = ~pi1893 & ~n15250;
  assign n23234 = ~n23232 & ~n23233;
  assign n23235 = ~pi0509 & ~n23234;
  assign n23236 = pi0509 & ~pi1893;
  assign po2070 = n23235 | n23236;
  assign n23238 = pi3431 & n15250;
  assign n23239 = ~pi1894 & ~n15250;
  assign n23240 = ~n23238 & ~n23239;
  assign n23241 = ~pi0509 & ~n23240;
  assign n23242 = pi0509 & ~pi1894;
  assign po2071 = n23241 | n23242;
  assign n23244 = pi3411 & n15250;
  assign n23245 = ~pi1895 & ~n15250;
  assign n23246 = ~n23244 & ~n23245;
  assign n23247 = ~pi0509 & ~n23246;
  assign n23248 = pi0509 & ~pi1895;
  assign po2072 = n23247 | n23248;
  assign n23250 = pi3422 & n15250;
  assign n23251 = ~pi1896 & ~n15250;
  assign n23252 = ~n23250 & ~n23251;
  assign n23253 = ~pi0509 & ~n23252;
  assign n23254 = pi0509 & ~pi1896;
  assign po2073 = n23253 | n23254;
  assign n23256 = pi3435 & n15250;
  assign n23257 = ~pi1897 & ~n15250;
  assign n23258 = ~n23256 & ~n23257;
  assign n23259 = ~pi0509 & ~n23258;
  assign n23260 = pi0509 & ~pi1897;
  assign po2074 = n23259 | n23260;
  assign n23262 = pi3421 & n15250;
  assign n23263 = ~pi1898 & ~n15250;
  assign n23264 = ~n23262 & ~n23263;
  assign n23265 = ~pi0509 & ~n23264;
  assign n23266 = pi0509 & ~pi1898;
  assign po2075 = n23265 | n23266;
  assign n23268 = pi3410 & n15250;
  assign n23269 = ~pi1899 & ~n15250;
  assign n23270 = ~n23268 & ~n23269;
  assign n23271 = ~pi0509 & ~n23270;
  assign n23272 = pi0509 & ~pi1899;
  assign po2076 = n23271 | n23272;
  assign n23274 = pi3420 & n15250;
  assign n23275 = ~pi1900 & ~n15250;
  assign n23276 = ~n23274 & ~n23275;
  assign n23277 = ~pi0509 & ~n23276;
  assign n23278 = pi0509 & ~pi1900;
  assign po2077 = n23277 | n23278;
  assign n23280 = ~pi3082 & n22326;
  assign n23281 = ~pi1901 & ~n22326;
  assign n23282 = ~n23280 & ~n23281;
  assign n23283 = n22306 & ~n23282;
  assign n23284 = ~pi1901 & ~n22306;
  assign po2078 = n23283 | n23284;
  assign n23286 = ~pi1693 & pi1858;
  assign n23287 = ~pi1858 & ~n19943;
  assign n23288 = ~n23286 & ~n23287;
  assign n23289 = ~n10979 & ~n23288;
  assign n23290 = pi1902 & n10979;
  assign po2079 = n23289 | n23290;
  assign n23292 = ~pi1903 & ~n22539;
  assign n23293 = pi2976 & n22539;
  assign n23294 = ~n23292 & ~n23293;
  assign n23295 = n22306 & ~n23294;
  assign n23296 = ~pi1903 & ~n22306;
  assign po2080 = n23295 | n23296;
  assign n23298 = ~pi3082 & n22318;
  assign n23299 = ~pi1904 & ~n22318;
  assign n23300 = ~n23298 & ~n23299;
  assign n23301 = n22306 & ~n23300;
  assign n23302 = ~pi1904 & ~n22306;
  assign po2081 = n23301 | n23302;
  assign n23304 = ~pi1905 & ~n22860;
  assign n23305 = ~pi1905 & ~n22900;
  assign n23306 = ~pi3159 & ~n19955;
  assign n23307 = n22900 & ~n23306;
  assign n23308 = ~n23305 & ~n23307;
  assign n23309 = n22860 & ~n23308;
  assign po2082 = n23304 | n23309;
  assign n23311 = ~pi1906 & ~n22860;
  assign n23312 = ~pi1906 & ~n22879;
  assign n23313 = ~pi3145 & ~n19955;
  assign n23314 = n22879 & ~n23313;
  assign n23315 = ~n23312 & ~n23314;
  assign n23316 = n22860 & ~n23315;
  assign po2083 = n23311 | n23316;
  assign n23318 = ~pi1907 & ~n22860;
  assign n23319 = ~pi1907 & ~n22980;
  assign n23320 = ~pi3143 & ~n19955;
  assign n23321 = n22980 & ~n23320;
  assign n23322 = ~n23319 & ~n23321;
  assign n23323 = n22860 & ~n23322;
  assign po2084 = n23318 | n23323;
  assign n23325 = ~pi1908 & ~n22860;
  assign n23326 = ~pi1908 & ~n22938;
  assign n23327 = ~pi3142 & ~n19955;
  assign n23328 = n22938 & ~n23327;
  assign n23329 = ~n23326 & ~n23328;
  assign n23330 = n22860 & ~n23329;
  assign po2085 = n23325 | n23330;
  assign n23332 = ~pi1909 & ~n22860;
  assign n23333 = ~pi1909 & ~n22893;
  assign n23334 = ~pi3131 & ~n19955;
  assign n23335 = n22893 & ~n23334;
  assign n23336 = ~n23333 & ~n23335;
  assign n23337 = n22860 & ~n23336;
  assign po2086 = n23332 | n23337;
  assign n23339 = ~pi1910 & ~n22860;
  assign n23340 = ~pi1910 & ~n22893;
  assign n23341 = ~pi3146 & ~n19955;
  assign n23342 = n22893 & ~n23341;
  assign n23343 = ~n23340 & ~n23342;
  assign n23344 = n22860 & ~n23343;
  assign po2087 = n23339 | n23344;
  assign n23346 = ~pi1911 & ~n22860;
  assign n23347 = ~pi1911 & ~n22893;
  assign n23348 = ~pi3136 & ~n19955;
  assign n23349 = n22893 & ~n23348;
  assign n23350 = ~n23347 & ~n23349;
  assign n23351 = n22860 & ~n23350;
  assign po2088 = n23346 | n23351;
  assign n23353 = ~pi1912 & ~n22860;
  assign n23354 = ~pi1912 & ~n22980;
  assign n23355 = ~pi3171 & ~n19955;
  assign n23356 = n22980 & ~n23355;
  assign n23357 = ~n23354 & ~n23356;
  assign n23358 = n22860 & ~n23357;
  assign po2089 = n23353 | n23358;
  assign n23360 = ~pi1913 & ~n22860;
  assign n23361 = ~pi1913 & ~n22879;
  assign n23362 = n22879 & ~n23306;
  assign n23363 = ~n23361 & ~n23362;
  assign n23364 = n22860 & ~n23363;
  assign po2090 = n23360 | n23364;
  assign n23366 = ~pi1914 & ~n22860;
  assign n23367 = ~pi1914 & ~n22980;
  assign n23368 = ~pi3153 & ~n19955;
  assign n23369 = n22980 & ~n23368;
  assign n23370 = ~n23367 & ~n23369;
  assign n23371 = n22860 & ~n23370;
  assign po2091 = n23366 | n23371;
  assign n23373 = ~pi1915 & ~n22860;
  assign n23374 = ~pi1915 & ~n22879;
  assign n23375 = n22879 & ~n23334;
  assign n23376 = ~n23374 & ~n23375;
  assign n23377 = n22860 & ~n23376;
  assign po2092 = n23373 | n23377;
  assign n23379 = ~pi1916 & ~n22860;
  assign n23380 = ~pi1916 & ~n22980;
  assign n23381 = ~pi3134 & ~n19955;
  assign n23382 = n22980 & ~n23381;
  assign n23383 = ~n23380 & ~n23382;
  assign n23384 = n22860 & ~n23383;
  assign po2093 = n23379 | n23384;
  assign n23386 = ~pi1917 & ~n22860;
  assign n23387 = ~pi1917 & ~n22879;
  assign n23388 = ~pi3170 & ~n19955;
  assign n23389 = n22879 & ~n23388;
  assign n23390 = ~n23387 & ~n23389;
  assign n23391 = n22860 & ~n23390;
  assign po2094 = n23386 | n23391;
  assign n23393 = ~pi1918 & ~n22860;
  assign n23394 = ~pi1918 & ~n22980;
  assign n23395 = ~pi3132 & ~n19955;
  assign n23396 = n22980 & ~n23395;
  assign n23397 = ~n23394 & ~n23396;
  assign n23398 = n22860 & ~n23397;
  assign po2095 = n23393 | n23398;
  assign n23400 = ~pi1919 & ~n22860;
  assign n23401 = ~pi1919 & ~n22900;
  assign n23402 = n22900 & ~n23334;
  assign n23403 = ~n23401 & ~n23402;
  assign n23404 = n22860 & ~n23403;
  assign po2096 = n23400 | n23404;
  assign n23406 = ~pi1920 & ~n22860;
  assign n23407 = ~pi1920 & ~n22879;
  assign n23408 = ~pi3133 & ~n19955;
  assign n23409 = n22879 & ~n23408;
  assign n23410 = ~n23407 & ~n23409;
  assign n23411 = n22860 & ~n23410;
  assign po2097 = n23406 | n23411;
  assign n23413 = ~pi1921 & ~n22860;
  assign n23414 = ~pi1921 & ~n22879;
  assign n23415 = ~pi3151 & ~n19955;
  assign n23416 = n22879 & ~n23415;
  assign n23417 = ~n23414 & ~n23416;
  assign n23418 = n22860 & ~n23417;
  assign po2098 = n23413 | n23418;
  assign n23420 = ~pi1922 & ~n22860;
  assign n23421 = ~pi1922 & ~n22980;
  assign n23422 = n22980 & ~n23348;
  assign n23423 = ~n23421 & ~n23422;
  assign n23424 = n22860 & ~n23423;
  assign po2099 = n23420 | n23424;
  assign po2100 = pi1923 & ~n8238;
  assign n23427 = ~pi1924 & ~n22860;
  assign n23428 = ~pi3141 & ~n19955;
  assign n23429 = n22867 & ~n23428;
  assign n23430 = ~pi1924 & ~n22867;
  assign n23431 = ~n23429 & ~n23430;
  assign n23432 = n22860 & ~n23431;
  assign po2101 = n23427 | n23432;
  assign n23434 = ~pi1925 & ~n22860;
  assign n23435 = ~pi1925 & ~n22879;
  assign n23436 = n22879 & ~n23327;
  assign n23437 = ~n23435 & ~n23436;
  assign n23438 = n22860 & ~n23437;
  assign po2102 = n23434 | n23438;
  assign n23440 = ~pi1926 & ~n22860;
  assign n23441 = ~pi1926 & ~n22980;
  assign n23442 = n22980 & ~n23428;
  assign n23443 = ~n23441 & ~n23442;
  assign n23444 = n22860 & ~n23443;
  assign po2103 = n23440 | n23444;
  assign n23446 = ~pi1927 & ~n22860;
  assign n23447 = ~pi1927 & ~n22980;
  assign n23448 = ~pi3139 & ~n19955;
  assign n23449 = n22980 & ~n23448;
  assign n23450 = ~n23447 & ~n23449;
  assign n23451 = n22860 & ~n23450;
  assign po2104 = n23446 | n23451;
  assign n23453 = ~pi1928 & ~n22860;
  assign n23454 = ~pi1928 & ~n22879;
  assign n23455 = pi2975 & n22879;
  assign n23456 = ~n23454 & ~n23455;
  assign n23457 = n22860 & ~n23456;
  assign po2105 = n23453 | n23457;
  assign n23459 = ~pi1929 & ~n22860;
  assign n23460 = ~pi1929 & ~n22980;
  assign n23461 = ~pi3168 & ~n19955;
  assign n23462 = n22980 & ~n23461;
  assign n23463 = ~n23460 & ~n23462;
  assign n23464 = n22860 & ~n23463;
  assign po2106 = n23459 | n23464;
  assign n23466 = ~pi1930 & ~n22860;
  assign n23467 = ~pi1930 & ~n22900;
  assign n23468 = n22900 & ~n23341;
  assign n23469 = ~n23467 & ~n23468;
  assign n23470 = n22860 & ~n23469;
  assign po2107 = n23466 | n23470;
  assign n23472 = ~pi1931 & ~n22860;
  assign n23473 = ~pi1931 & ~n22879;
  assign n23474 = ~pi3166 & ~n19955;
  assign n23475 = n22879 & ~n23474;
  assign n23476 = ~n23473 & ~n23475;
  assign n23477 = n22860 & ~n23476;
  assign po2108 = n23472 | n23477;
  assign n23479 = ~pi1932 & ~n22860;
  assign n23480 = ~pi1932 & ~n22879;
  assign n23481 = ~pi3150 & ~n19955;
  assign n23482 = n22879 & ~n23481;
  assign n23483 = ~n23480 & ~n23482;
  assign n23484 = n22860 & ~n23483;
  assign po2109 = n23479 | n23484;
  assign n23486 = ~pi1933 & ~n22860;
  assign n23487 = ~pi1933 & ~n22900;
  assign n23488 = n22900 & ~n23388;
  assign n23489 = ~n23487 & ~n23488;
  assign n23490 = n22860 & ~n23489;
  assign po2110 = n23486 | n23490;
  assign n23492 = ~pi1934 & ~n22860;
  assign n23493 = n22931 & ~n23334;
  assign n23494 = ~pi1934 & ~n22931;
  assign n23495 = ~n23493 & ~n23494;
  assign n23496 = n22860 & ~n23495;
  assign po2111 = n23492 | n23496;
  assign n23498 = ~pi1935 & ~n22860;
  assign n23499 = n22966 & ~n23388;
  assign n23500 = ~pi1935 & ~n22966;
  assign n23501 = ~n23499 & ~n23500;
  assign n23502 = n22860 & ~n23501;
  assign po2112 = n23498 | n23502;
  assign n23504 = ~pi1936 & ~n22860;
  assign n23505 = n22973 & ~n23415;
  assign n23506 = ~pi1936 & ~n22973;
  assign n23507 = ~n23505 & ~n23506;
  assign n23508 = n22860 & ~n23507;
  assign po2113 = n23504 | n23508;
  assign n23510 = ~pi1937 & ~n22860;
  assign n23511 = ~pi3154 & ~n19955;
  assign n23512 = n22973 & ~n23511;
  assign n23513 = ~pi1937 & ~n22973;
  assign n23514 = ~n23512 & ~n23513;
  assign n23515 = n22860 & ~n23514;
  assign po2114 = n23510 | n23515;
  assign n23517 = ~pi1938 & ~n22860;
  assign n23518 = ~pi3147 & ~n19955;
  assign n23519 = n22867 & ~n23518;
  assign n23520 = ~pi1938 & ~n22867;
  assign n23521 = ~n23519 & ~n23520;
  assign n23522 = n22860 & ~n23521;
  assign po2115 = n23517 | n23522;
  assign n23524 = ~pi1939 & ~n22860;
  assign n23525 = n22867 & ~n23306;
  assign n23526 = ~pi1939 & ~n22867;
  assign n23527 = ~n23525 & ~n23526;
  assign n23528 = n22860 & ~n23527;
  assign po2116 = n23524 | n23528;
  assign n23530 = ~pi1940 & ~n22860;
  assign n23531 = n22924 & ~n23381;
  assign n23532 = ~pi1940 & ~n22924;
  assign n23533 = ~n23531 & ~n23532;
  assign n23534 = n22860 & ~n23533;
  assign po2117 = n23530 | n23534;
  assign n23536 = ~pi1941 & ~n22860;
  assign n23537 = ~pi3172 & ~n19955;
  assign n23538 = n22886 & ~n23537;
  assign n23539 = ~pi1941 & ~n22886;
  assign n23540 = ~n23538 & ~n23539;
  assign n23541 = n22860 & ~n23540;
  assign po2118 = n23536 | n23541;
  assign n23543 = ~pi1942 & ~n22860;
  assign n23544 = n22924 & ~n23320;
  assign n23545 = ~pi1942 & ~n22924;
  assign n23546 = ~n23544 & ~n23545;
  assign n23547 = n22860 & ~n23546;
  assign po2119 = n23543 | n23547;
  assign n23549 = ~pi1943 & ~n22860;
  assign n23550 = ~pi3135 & ~n19955;
  assign n23551 = n22886 & ~n23550;
  assign n23552 = ~pi1943 & ~n22886;
  assign n23553 = ~n23551 & ~n23552;
  assign n23554 = n22860 & ~n23553;
  assign po2120 = n23549 | n23554;
  assign n23556 = ~pi1944 & ~n22860;
  assign n23557 = ~pi3163 & ~n19955;
  assign n23558 = n22886 & ~n23557;
  assign n23559 = ~pi1944 & ~n22886;
  assign n23560 = ~n23558 & ~n23559;
  assign n23561 = n22860 & ~n23560;
  assign po2121 = n23556 | n23561;
  assign n23563 = ~pi1945 & ~n22860;
  assign n23564 = n22886 & ~n23415;
  assign n23565 = ~pi1945 & ~n22886;
  assign n23566 = ~n23564 & ~n23565;
  assign n23567 = n22860 & ~n23566;
  assign po2122 = n23563 | n23567;
  assign n23569 = ~pi1946 & ~n22860;
  assign n23570 = ~pi3157 & ~n19955;
  assign n23571 = n22886 & ~n23570;
  assign n23572 = ~pi1946 & ~n22886;
  assign n23573 = ~n23571 & ~n23572;
  assign n23574 = n22860 & ~n23573;
  assign po2123 = n23569 | n23574;
  assign n23576 = ~pi1947 & ~n22860;
  assign n23577 = n22886 & ~n23511;
  assign n23578 = ~pi1947 & ~n22886;
  assign n23579 = ~n23577 & ~n23578;
  assign n23580 = n22860 & ~n23579;
  assign po2124 = n23576 | n23580;
  assign n23582 = ~pi1948 & ~n22860;
  assign n23583 = n22867 & ~n23381;
  assign n23584 = ~pi1948 & ~n22867;
  assign n23585 = ~n23583 & ~n23584;
  assign n23586 = n22860 & ~n23585;
  assign po2125 = n23582 | n23586;
  assign n23588 = ~pi1949 & ~n22860;
  assign n23589 = n22886 & ~n23381;
  assign n23590 = ~pi1949 & ~n22886;
  assign n23591 = ~n23589 & ~n23590;
  assign n23592 = n22860 & ~n23591;
  assign po2126 = n23588 | n23592;
  assign n23594 = ~pi1950 & ~n22860;
  assign n23595 = n22867 & ~n23388;
  assign n23596 = ~pi1950 & ~n22867;
  assign n23597 = ~n23595 & ~n23596;
  assign n23598 = n22860 & ~n23597;
  assign po2127 = n23594 | n23598;
  assign n23600 = ~pi1951 & ~n22860;
  assign n23601 = n22886 & ~n23428;
  assign n23602 = ~pi1951 & ~n22886;
  assign n23603 = ~n23601 & ~n23602;
  assign n23604 = n22860 & ~n23603;
  assign po2128 = n23600 | n23604;
  assign n23606 = ~pi1952 & ~n22860;
  assign n23607 = n22886 & ~n23448;
  assign n23608 = ~pi1952 & ~n22886;
  assign n23609 = ~n23607 & ~n23608;
  assign n23610 = n22860 & ~n23609;
  assign po2129 = n23606 | n23610;
  assign n23612 = ~pi1953 & ~n22860;
  assign n23613 = n22867 & ~n23341;
  assign n23614 = ~pi1953 & ~n22867;
  assign n23615 = ~n23613 & ~n23614;
  assign n23616 = n22860 & ~n23615;
  assign po2130 = n23612 | n23616;
  assign n23618 = ~pi1954 & ~n22860;
  assign n23619 = n22867 & ~n23415;
  assign n23620 = ~pi1954 & ~n22867;
  assign n23621 = ~n23619 & ~n23620;
  assign n23622 = n22860 & ~n23621;
  assign po2131 = n23618 | n23622;
  assign n23624 = ~pi1955 & ~n22860;
  assign n23625 = ~pi3158 & ~n19955;
  assign n23626 = n22867 & ~n23625;
  assign n23627 = ~pi1955 & ~n22867;
  assign n23628 = ~n23626 & ~n23627;
  assign n23629 = n22860 & ~n23628;
  assign po2132 = n23624 | n23629;
  assign n23631 = ~pi1956 & ~n22860;
  assign n23632 = n22867 & ~n23313;
  assign n23633 = ~pi1956 & ~n22867;
  assign n23634 = ~n23632 & ~n23633;
  assign n23635 = n22860 & ~n23634;
  assign po2133 = n23631 | n23635;
  assign n23637 = ~pi1957 & ~n22860;
  assign n23638 = ~pi3165 & ~n19955;
  assign n23639 = n22945 & ~n23638;
  assign n23640 = ~pi1957 & ~n22945;
  assign n23641 = ~n23639 & ~n23640;
  assign n23642 = n22860 & ~n23641;
  assign po2134 = n23637 | n23642;
  assign n23644 = ~pi1958 & ~n22860;
  assign n23645 = ~pi3164 & ~n19955;
  assign n23646 = n22867 & ~n23645;
  assign n23647 = ~pi1958 & ~n22867;
  assign n23648 = ~n23646 & ~n23647;
  assign n23649 = n22860 & ~n23648;
  assign po2135 = n23644 | n23649;
  assign n23651 = ~pi1959 & ~n22860;
  assign n23652 = n22867 & ~n23537;
  assign n23653 = ~pi1959 & ~n22867;
  assign n23654 = ~n23652 & ~n23653;
  assign n23655 = n22860 & ~n23654;
  assign po2136 = n23651 | n23655;
  assign n23657 = ~pi1960 & ~n22860;
  assign n23658 = n22867 & ~n23481;
  assign n23659 = ~pi1960 & ~n22867;
  assign n23660 = ~n23658 & ~n23659;
  assign n23661 = n22860 & ~n23660;
  assign po2137 = n23657 | n23661;
  assign n23663 = ~pi1961 & ~n22860;
  assign n23664 = ~pi3162 & ~n19955;
  assign n23665 = n22867 & ~n23664;
  assign n23666 = ~pi1961 & ~n22867;
  assign n23667 = ~n23665 & ~n23666;
  assign n23668 = n22860 & ~n23667;
  assign po2138 = n23663 | n23668;
  assign n23670 = ~pi1962 & ~n22860;
  assign n23671 = ~pi1962 & ~n22879;
  assign n23672 = n22879 & ~n23537;
  assign n23673 = ~n23671 & ~n23672;
  assign n23674 = n22860 & ~n23673;
  assign po2139 = n23670 | n23674;
  assign n23676 = ~pi1963 & ~n22860;
  assign n23677 = n22867 & ~n23511;
  assign n23678 = ~pi1963 & ~n22867;
  assign n23679 = ~n23677 & ~n23678;
  assign n23680 = n22860 & ~n23679;
  assign po2140 = n23676 | n23680;
  assign n23682 = ~pi1964 & ~n22860;
  assign n23683 = n22867 & ~n23557;
  assign n23684 = ~pi1964 & ~n22867;
  assign n23685 = ~n23683 & ~n23684;
  assign n23686 = n22860 & ~n23685;
  assign po2141 = n23682 | n23686;
  assign n23688 = pi2973 & pi2978;
  assign n23689 = pi2983 & pi2998;
  assign n23690 = pi2999 & pi3002;
  assign n23691 = pi2991 & n23690;
  assign n23692 = pi2986 & n23691;
  assign n23693 = pi2979 & n23692;
  assign n23694 = pi2977 & n23693;
  assign n23695 = n23689 & n23694;
  assign n23696 = pi2970 & n23695;
  assign n23697 = pi2962 & n23696;
  assign n23698 = n23688 & n23697;
  assign n23699 = pi2957 & pi2974;
  assign n23700 = n23698 & n23699;
  assign n23701 = pi2947 & n23700;
  assign n23702 = pi2939 & n23701;
  assign n23703 = ~pi1965 & n23702;
  assign n23704 = pi1965 & ~n23702;
  assign n23705 = ~n23703 & ~n23704;
  assign n23706 = pi0120 & n7250;
  assign n23707 = pi2758 & n23706;
  assign n23708 = pi1965 & ~n23707;
  assign n23709 = po3339 & n23708;
  assign po2142 = n23705 & n23709;
  assign n23711 = pi3182 & pi3320;
  assign n23712 = ~pi1966 & ~n23711;
  assign n23713 = n7066 & n7068;
  assign n23714 = n7075 & n23713;
  assign n23715 = ~n17996 & ~n23714;
  assign n23716 = pi1348 & ~n23715;
  assign n23717 = pi1397 & n23716;
  assign po2143 = n23712 | n23717;
  assign po2144 = pi1967 & ~n8238;
  assign po2145 = pi1968 & ~n8238;
  assign po2146 = pi1969 & ~n8238;
  assign n23722 = pi1970 & ~n20262;
  assign n23723 = ~n10917 & n20262;
  assign po2147 = n23722 | n23723;
  assign n23725 = pi1704 & n22080;
  assign n23726 = ~n19469 & ~n22080;
  assign n23727 = pi1971 & ~n23726;
  assign n23728 = ~pi2294 & ~pi2463;
  assign n23729 = n19466 & n23728;
  assign n23730 = n19464 & n23729;
  assign n23731 = pi1971 & n23730;
  assign n23732 = ~pi1971 & ~n23730;
  assign n23733 = ~n23731 & ~n23732;
  assign n23734 = n23726 & n23733;
  assign n23735 = ~n23727 & ~n23734;
  assign n23736 = ~n22080 & ~n23735;
  assign po2148 = n23725 | n23736;
  assign n23738 = pi1700 & n22080;
  assign n23739 = pi1972 & ~n23726;
  assign n23740 = ~pi1972 & n23728;
  assign n23741 = pi1972 & ~n23728;
  assign n23742 = ~n23740 & ~n23741;
  assign n23743 = n23726 & ~n23742;
  assign n23744 = ~n23739 & ~n23743;
  assign n23745 = ~n22080 & ~n23744;
  assign po2149 = n23738 | n23745;
  assign n23747 = pi2987 & n22561;
  assign n23748 = ~pi1974 & ~n22561;
  assign n23749 = ~n23747 & ~n23748;
  assign n23750 = n22306 & ~n23749;
  assign n23751 = ~pi1974 & ~n22306;
  assign po2151 = n23750 | n23751;
  assign n23753 = pi2987 & n22554;
  assign n23754 = ~pi1975 & ~n22554;
  assign n23755 = ~n23753 & ~n23754;
  assign n23756 = n22306 & ~n23755;
  assign n23757 = ~pi1975 & ~n22306;
  assign po2152 = n23756 | n23757;
  assign n23759 = ~pi1976 & ~n22318;
  assign n23760 = pi2987 & n22318;
  assign n23761 = ~n23759 & ~n23760;
  assign n23762 = n22306 & ~n23761;
  assign n23763 = ~pi1976 & ~n22306;
  assign po2153 = n23762 | n23763;
  assign n23765 = ~pi1977 & ~n22547;
  assign n23766 = pi2987 & n22547;
  assign n23767 = ~n23765 & ~n23766;
  assign n23768 = n22306 & ~n23767;
  assign n23769 = ~pi1977 & ~n22306;
  assign po2154 = n23768 | n23769;
  assign n23771 = ~pi1978 & ~n22547;
  assign n23772 = pi2988 & n22547;
  assign n23773 = ~n23771 & ~n23772;
  assign n23774 = n22306 & ~n23773;
  assign n23775 = ~pi1978 & ~n22306;
  assign po2155 = n23774 | n23775;
  assign n23777 = ~pi1979 & ~n22539;
  assign n23778 = pi2987 & n22539;
  assign n23779 = ~n23777 & ~n23778;
  assign n23780 = n22306 & ~n23779;
  assign n23781 = ~pi1979 & ~n22306;
  assign po2156 = n23780 | n23781;
  assign n23783 = ~pi1980 & ~n22326;
  assign n23784 = pi2987 & n22326;
  assign n23785 = ~n23783 & ~n23784;
  assign n23786 = n22306 & ~n23785;
  assign n23787 = ~pi1980 & ~n22306;
  assign po2157 = n23786 | n23787;
  assign n23789 = pi1983 & ~n22860;
  assign n23790 = ~n19183 & n22860;
  assign po2159 = n23789 | n23790;
  assign n23792 = pi1984 & ~n22860;
  assign n23793 = ~pi1984 & n22860;
  assign po2160 = n23792 | n23793;
  assign n23795 = pi1985 & ~n22860;
  assign n23796 = ~n19072 & n22860;
  assign po2161 = n23795 | n23796;
  assign n23798 = ~pi1986 & ~n22860;
  assign n23799 = pi1983 & n22860;
  assign po2162 = n23798 | n23799;
  assign n23801 = ~pi1987 & ~n22860;
  assign n23802 = n22959 & ~n23348;
  assign n23803 = ~pi1987 & ~n22959;
  assign n23804 = ~n23802 & ~n23803;
  assign n23805 = n22860 & ~n23804;
  assign po2163 = n23801 | n23805;
  assign n23807 = ~pi1988 & ~n22860;
  assign n23808 = n22959 & ~n23448;
  assign n23809 = ~pi1988 & ~n22959;
  assign n23810 = ~n23808 & ~n23809;
  assign n23811 = n22860 & ~n23810;
  assign po2164 = n23807 | n23811;
  assign n23813 = ~pi1989 & ~n22860;
  assign n23814 = n22959 & ~n23428;
  assign n23815 = ~pi1989 & ~n22959;
  assign n23816 = ~n23814 & ~n23815;
  assign n23817 = n22860 & ~n23816;
  assign po2165 = n23813 | n23817;
  assign n23819 = ~pi1990 & ~n22860;
  assign n23820 = n22959 & ~n23518;
  assign n23821 = ~pi1990 & ~n22959;
  assign n23822 = ~n23820 & ~n23821;
  assign n23823 = n22860 & ~n23822;
  assign po2166 = n23819 | n23823;
  assign n23825 = ~pi1991 & ~n22860;
  assign n23826 = n22867 & ~n23448;
  assign n23827 = ~pi1991 & ~n22867;
  assign n23828 = ~n23826 & ~n23827;
  assign n23829 = n22860 & ~n23828;
  assign po2167 = n23825 | n23829;
  assign n23831 = ~pi1992 & ~n22860;
  assign n23832 = n22959 & ~n23381;
  assign n23833 = ~pi1992 & ~n22959;
  assign n23834 = ~n23832 & ~n23833;
  assign n23835 = n22860 & ~n23834;
  assign po2168 = n23831 | n23835;
  assign n23837 = ~pi1993 & ~n22860;
  assign n23838 = n22959 & ~n23645;
  assign n23839 = ~pi1993 & ~n22959;
  assign n23840 = ~n23838 & ~n23839;
  assign n23841 = n22860 & ~n23840;
  assign po2169 = n23837 | n23841;
  assign n23843 = ~pi1994 & ~n22860;
  assign n23844 = n22959 & ~n23557;
  assign n23845 = ~pi1994 & ~n22959;
  assign n23846 = ~n23844 & ~n23845;
  assign n23847 = n22860 & ~n23846;
  assign po2170 = n23843 | n23847;
  assign n23849 = ~pi1995 & ~n22860;
  assign n23850 = n22959 & ~n23664;
  assign n23851 = ~pi1995 & ~n22959;
  assign n23852 = ~n23850 & ~n23851;
  assign n23853 = n22860 & ~n23852;
  assign po2171 = n23849 | n23853;
  assign n23855 = ~pi1996 & ~n22860;
  assign n23856 = n22959 & ~n23511;
  assign n23857 = ~pi1996 & ~n22959;
  assign n23858 = ~n23856 & ~n23857;
  assign n23859 = n22860 & ~n23858;
  assign po2172 = n23855 | n23859;
  assign n23861 = ~pi1997 & ~n22860;
  assign n23862 = ~pi3138 & ~n19955;
  assign n23863 = n22959 & ~n23862;
  assign n23864 = ~pi1997 & ~n22959;
  assign n23865 = ~n23863 & ~n23864;
  assign n23866 = n22860 & ~n23865;
  assign po2173 = n23861 | n23866;
  assign n23868 = ~pi1998 & ~n22860;
  assign n23869 = n22959 & ~n23415;
  assign n23870 = ~pi1998 & ~n22959;
  assign n23871 = ~n23869 & ~n23870;
  assign n23872 = n22860 & ~n23871;
  assign po2174 = n23868 | n23872;
  assign n23874 = ~pi1999 & ~n22860;
  assign n23875 = n22959 & ~n23537;
  assign n23876 = ~pi1999 & ~n22959;
  assign n23877 = ~n23875 & ~n23876;
  assign n23878 = n22860 & ~n23877;
  assign po2175 = n23874 | n23878;
  assign n23880 = ~pi2000 & ~n22860;
  assign n23881 = n22959 & ~n23550;
  assign n23882 = ~pi2000 & ~n22959;
  assign n23883 = ~n23881 & ~n23882;
  assign n23884 = n22860 & ~n23883;
  assign po2176 = n23880 | n23884;
  assign n23886 = ~pi2001 & ~n22860;
  assign n23887 = n22959 & ~n23481;
  assign n23888 = ~pi2001 & ~n22959;
  assign n23889 = ~n23887 & ~n23888;
  assign n23890 = n22860 & ~n23889;
  assign po2177 = n23886 | n23890;
  assign n23892 = ~pi2002 & ~n22860;
  assign n23893 = n22959 & ~n23408;
  assign n23894 = ~pi2002 & ~n22959;
  assign n23895 = ~n23893 & ~n23894;
  assign n23896 = n22860 & ~n23895;
  assign po2178 = n23892 | n23896;
  assign n23898 = ~pi2003 & ~n22860;
  assign n23899 = n22959 & ~n23313;
  assign n23900 = ~pi2003 & ~n22959;
  assign n23901 = ~n23899 & ~n23900;
  assign n23902 = n22860 & ~n23901;
  assign po2179 = n23898 | n23902;
  assign n23904 = ~pi2004 & ~n22860;
  assign n23905 = n22959 & ~n23306;
  assign n23906 = ~pi2004 & ~n22959;
  assign n23907 = ~n23905 & ~n23906;
  assign n23908 = n22860 & ~n23907;
  assign po2180 = n23904 | n23908;
  assign n23910 = ~pi2005 & ~n22860;
  assign n23911 = n22959 & ~n23388;
  assign n23912 = ~pi2005 & ~n22959;
  assign n23913 = ~n23911 & ~n23912;
  assign n23914 = n22860 & ~n23913;
  assign po2181 = n23910 | n23914;
  assign n23916 = ~pi2006 & ~n22860;
  assign n23917 = n22867 & ~n23348;
  assign n23918 = ~pi2006 & ~n22867;
  assign n23919 = ~n23917 & ~n23918;
  assign n23920 = n22860 & ~n23919;
  assign po2182 = n23916 | n23920;
  assign n23922 = ~pi2007 & ~n22860;
  assign n23923 = n22867 & ~n23461;
  assign n23924 = ~pi2007 & ~n22867;
  assign n23925 = ~n23923 & ~n23924;
  assign n23926 = n22860 & ~n23925;
  assign po2183 = n23922 | n23926;
  assign n23928 = ~pi2008 & ~n22860;
  assign n23929 = n22867 & ~n23320;
  assign n23930 = ~pi2008 & ~n22867;
  assign n23931 = ~n23929 & ~n23930;
  assign n23932 = n22860 & ~n23931;
  assign po2184 = n23928 | n23932;
  assign n23934 = ~pi2009 & ~n22860;
  assign n23935 = n22867 & ~n23368;
  assign n23936 = ~pi2009 & ~n22867;
  assign n23937 = ~n23935 & ~n23936;
  assign n23938 = n22860 & ~n23937;
  assign po2185 = n23934 | n23938;
  assign n23940 = ~pi2010 & ~n22860;
  assign n23941 = n22867 & ~n23395;
  assign n23942 = ~pi2010 & ~n22867;
  assign n23943 = ~n23941 & ~n23942;
  assign n23944 = n22860 & ~n23943;
  assign po2186 = n23940 | n23944;
  assign n23946 = ~pi2011 & ~n22860;
  assign n23947 = n22867 & ~n23355;
  assign n23948 = ~pi2011 & ~n22867;
  assign n23949 = ~n23947 & ~n23948;
  assign n23950 = n22860 & ~n23949;
  assign po2187 = n23946 | n23950;
  assign n23952 = ~pi2012 & ~n22860;
  assign n23953 = ~pi3155 & ~n19955;
  assign n23954 = n22867 & ~n23953;
  assign n23955 = ~pi2012 & ~n22867;
  assign n23956 = ~n23954 & ~n23955;
  assign n23957 = n22860 & ~n23956;
  assign po2188 = n23952 | n23957;
  assign n23959 = ~pi2013 & ~n22860;
  assign n23960 = n22867 & ~n23638;
  assign n23961 = ~pi2013 & ~n22867;
  assign n23962 = ~n23960 & ~n23961;
  assign n23963 = n22860 & ~n23962;
  assign po2189 = n23959 | n23963;
  assign n23965 = ~pi2014 & ~n22860;
  assign n23966 = n22867 & ~n23862;
  assign n23967 = ~pi2014 & ~n22867;
  assign n23968 = ~n23966 & ~n23967;
  assign n23969 = n22860 & ~n23968;
  assign po2190 = n23965 | n23969;
  assign n23971 = ~pi2015 & ~n22860;
  assign n23972 = n22867 & ~n23570;
  assign n23973 = ~pi2015 & ~n22867;
  assign n23974 = ~n23972 & ~n23973;
  assign n23975 = n22860 & ~n23974;
  assign po2191 = n23971 | n23975;
  assign n23977 = ~pi2016 & ~n22860;
  assign n23978 = n22867 & ~n23550;
  assign n23979 = ~pi2016 & ~n22867;
  assign n23980 = ~n23978 & ~n23979;
  assign n23981 = n22860 & ~n23980;
  assign po2192 = n23977 | n23981;
  assign n23983 = ~pi2017 & ~n22860;
  assign n23984 = n22867 & ~n23408;
  assign n23985 = ~pi2017 & ~n22867;
  assign n23986 = ~n23984 & ~n23985;
  assign n23987 = n22860 & ~n23986;
  assign po2193 = n23983 | n23987;
  assign n23989 = ~pi2018 & ~n22860;
  assign n23990 = n22867 & ~n23474;
  assign n23991 = ~pi2018 & ~n22867;
  assign n23992 = ~n23990 & ~n23991;
  assign n23993 = n22860 & ~n23992;
  assign po2194 = n23989 | n23993;
  assign n23995 = ~pi2019 & ~n22860;
  assign n23996 = n22867 & ~n23327;
  assign n23997 = ~pi2019 & ~n22867;
  assign n23998 = ~n23996 & ~n23997;
  assign n23999 = n22860 & ~n23998;
  assign po2195 = n23995 | n23999;
  assign n24001 = ~pi2020 & ~n22860;
  assign n24002 = ~pi3169 & ~n19955;
  assign n24003 = n22867 & ~n24002;
  assign n24004 = ~pi2020 & ~n22867;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = n22860 & ~n24005;
  assign po2196 = n24001 | n24006;
  assign n24008 = ~pi2021 & ~n22860;
  assign n24009 = n22867 & ~n23334;
  assign n24010 = ~pi2021 & ~n22867;
  assign n24011 = ~n24009 & ~n24010;
  assign n24012 = n22860 & ~n24011;
  assign po2197 = n24008 | n24012;
  assign n24014 = ~pi2022 & ~n22860;
  assign n24015 = n22886 & ~n23348;
  assign n24016 = ~pi2022 & ~n22886;
  assign n24017 = ~n24015 & ~n24016;
  assign n24018 = n22860 & ~n24017;
  assign po2198 = n24014 | n24018;
  assign n24020 = ~pi2023 & ~n22860;
  assign n24021 = n22886 & ~n23461;
  assign n24022 = ~pi2023 & ~n22886;
  assign n24023 = ~n24021 & ~n24022;
  assign n24024 = n22860 & ~n24023;
  assign po2199 = n24020 | n24024;
  assign n24026 = ~pi2024 & ~n22860;
  assign n24027 = n22886 & ~n23320;
  assign n24028 = ~pi2024 & ~n22886;
  assign n24029 = ~n24027 & ~n24028;
  assign n24030 = n22860 & ~n24029;
  assign po2200 = n24026 | n24030;
  assign n24032 = ~pi2025 & ~n22860;
  assign n24033 = n22886 & ~n23518;
  assign n24034 = ~pi2025 & ~n22886;
  assign n24035 = ~n24033 & ~n24034;
  assign n24036 = n22860 & ~n24035;
  assign po2201 = n24032 | n24036;
  assign n24038 = ~pi2026 & ~n22860;
  assign n24039 = n22886 & ~n23368;
  assign n24040 = ~pi2026 & ~n22886;
  assign n24041 = ~n24039 & ~n24040;
  assign n24042 = n22860 & ~n24041;
  assign po2202 = n24038 | n24042;
  assign n24044 = ~pi2027 & ~n22860;
  assign n24045 = n22886 & ~n23395;
  assign n24046 = ~pi2027 & ~n22886;
  assign n24047 = ~n24045 & ~n24046;
  assign n24048 = n22860 & ~n24047;
  assign po2203 = n24044 | n24048;
  assign n24050 = ~pi2028 & ~n22860;
  assign n24051 = n22886 & ~n23645;
  assign n24052 = ~pi2028 & ~n22886;
  assign n24053 = ~n24051 & ~n24052;
  assign n24054 = n22860 & ~n24053;
  assign po2204 = n24050 | n24054;
  assign n24056 = ~pi2029 & ~n22860;
  assign n24057 = n22886 & ~n23355;
  assign n24058 = ~pi2029 & ~n22886;
  assign n24059 = ~n24057 & ~n24058;
  assign n24060 = n22860 & ~n24059;
  assign po2205 = n24056 | n24060;
  assign n24062 = ~pi2030 & ~n22860;
  assign n24063 = n22886 & ~n23953;
  assign n24064 = ~pi2030 & ~n22886;
  assign n24065 = ~n24063 & ~n24064;
  assign n24066 = n22860 & ~n24065;
  assign po2206 = n24062 | n24066;
  assign n24068 = ~pi2031 & ~n22860;
  assign n24069 = n22886 & ~n23664;
  assign n24070 = ~pi2031 & ~n22886;
  assign n24071 = ~n24069 & ~n24070;
  assign n24072 = n22860 & ~n24071;
  assign po2207 = n24068 | n24072;
  assign n24074 = ~pi2032 & ~n22860;
  assign n24075 = n22886 & ~n23638;
  assign n24076 = ~pi2032 & ~n22886;
  assign n24077 = ~n24075 & ~n24076;
  assign n24078 = n22860 & ~n24077;
  assign po2208 = n24074 | n24078;
  assign n24080 = ~pi2033 & ~n22860;
  assign n24081 = n22886 & ~n23862;
  assign n24082 = ~pi2033 & ~n22886;
  assign n24083 = ~n24081 & ~n24082;
  assign n24084 = n22860 & ~n24083;
  assign po2209 = n24080 | n24084;
  assign n24086 = ~pi2034 & ~n22860;
  assign n24087 = n22886 & ~n23474;
  assign n24088 = ~pi2034 & ~n22886;
  assign n24089 = ~n24087 & ~n24088;
  assign n24090 = n22860 & ~n24089;
  assign po2210 = n24086 | n24090;
  assign n24092 = ~pi2035 & ~n22860;
  assign n24093 = n22886 & ~n23327;
  assign n24094 = ~pi2035 & ~n22886;
  assign n24095 = ~n24093 & ~n24094;
  assign n24096 = n22860 & ~n24095;
  assign po2211 = n24092 | n24096;
  assign n24098 = ~pi2036 & ~n22860;
  assign n24099 = n22886 & ~n24002;
  assign n24100 = ~pi2036 & ~n22886;
  assign n24101 = ~n24099 & ~n24100;
  assign n24102 = n22860 & ~n24101;
  assign po2212 = n24098 | n24102;
  assign n24104 = ~pi2037 & ~n22860;
  assign n24105 = n22886 & ~n23334;
  assign n24106 = ~pi2037 & ~n22886;
  assign n24107 = ~n24105 & ~n24106;
  assign n24108 = n22860 & ~n24107;
  assign po2213 = n24104 | n24108;
  assign n24110 = ~pi2038 & ~n22860;
  assign n24111 = n22886 & ~n23341;
  assign n24112 = ~pi2038 & ~n22886;
  assign n24113 = ~n24111 & ~n24112;
  assign n24114 = n22860 & ~n24113;
  assign po2214 = n24110 | n24114;
  assign n24116 = ~pi2039 & ~n22860;
  assign n24117 = n22909 & ~n23348;
  assign n24118 = ~pi2039 & ~n22909;
  assign n24119 = ~n24117 & ~n24118;
  assign n24120 = n22860 & ~n24119;
  assign po2215 = n24116 | n24120;
  assign n24122 = ~pi2040 & ~n22860;
  assign n24123 = n22909 & ~n23461;
  assign n24124 = ~pi2040 & ~n22909;
  assign n24125 = ~n24123 & ~n24124;
  assign n24126 = n22860 & ~n24125;
  assign po2216 = n24122 | n24126;
  assign n24128 = ~pi2041 & ~n22860;
  assign n24129 = n22909 & ~n23320;
  assign n24130 = ~pi2041 & ~n22909;
  assign n24131 = ~n24129 & ~n24130;
  assign n24132 = n22860 & ~n24131;
  assign po2217 = n24128 | n24132;
  assign n24134 = ~pi2042 & ~n22860;
  assign n24135 = n22909 & ~n23368;
  assign n24136 = ~pi2042 & ~n22909;
  assign n24137 = ~n24135 & ~n24136;
  assign n24138 = n22860 & ~n24137;
  assign po2218 = n24134 | n24138;
  assign n24140 = ~pi2043 & ~n22860;
  assign n24141 = n22909 & ~n23395;
  assign n24142 = ~pi2043 & ~n22909;
  assign n24143 = ~n24141 & ~n24142;
  assign n24144 = n22860 & ~n24143;
  assign po2219 = n24140 | n24144;
  assign n24146 = ~pi2044 & ~n22860;
  assign n24147 = n22909 & ~n23645;
  assign n24148 = ~pi2044 & ~n22909;
  assign n24149 = ~n24147 & ~n24148;
  assign n24150 = n22860 & ~n24149;
  assign po2220 = n24146 | n24150;
  assign n24152 = ~pi2045 & ~n22860;
  assign n24153 = n22909 & ~n23355;
  assign n24154 = ~pi2045 & ~n22909;
  assign n24155 = ~n24153 & ~n24154;
  assign n24156 = n22860 & ~n24155;
  assign po2221 = n24152 | n24156;
  assign n24158 = ~pi2046 & ~n22860;
  assign n24159 = n22909 & ~n23953;
  assign n24160 = ~pi2046 & ~n22909;
  assign n24161 = ~n24159 & ~n24160;
  assign n24162 = n22860 & ~n24161;
  assign po2222 = n24158 | n24162;
  assign n24164 = ~pi2047 & ~n22860;
  assign n24165 = n22909 & ~n23638;
  assign n24166 = ~pi2047 & ~n22909;
  assign n24167 = ~n24165 & ~n24166;
  assign n24168 = n22860 & ~n24167;
  assign po2223 = n24164 | n24168;
  assign n24170 = ~pi2048 & ~n22860;
  assign n24171 = n22909 & ~n23862;
  assign n24172 = ~pi2048 & ~n22909;
  assign n24173 = ~n24171 & ~n24172;
  assign n24174 = n22860 & ~n24173;
  assign po2224 = n24170 | n24174;
  assign n24176 = ~pi2049 & ~n22860;
  assign n24177 = n22909 & ~n23415;
  assign n24178 = ~pi2049 & ~n22909;
  assign n24179 = ~n24177 & ~n24178;
  assign n24180 = n22860 & ~n24179;
  assign po2225 = n24176 | n24180;
  assign n24182 = ~pi2050 & ~n22860;
  assign n24183 = n22909 & ~n23570;
  assign n24184 = ~pi2050 & ~n22909;
  assign n24185 = ~n24183 & ~n24184;
  assign n24186 = n22860 & ~n24185;
  assign po2226 = n24182 | n24186;
  assign n24188 = ~pi2051 & ~n22860;
  assign n24189 = n22909 & ~n23550;
  assign n24190 = ~pi2051 & ~n22909;
  assign n24191 = ~n24189 & ~n24190;
  assign n24192 = n22860 & ~n24191;
  assign po2227 = n24188 | n24192;
  assign n24194 = ~pi2052 & ~n22860;
  assign n24195 = n22909 & ~n23474;
  assign n24196 = ~pi2052 & ~n22909;
  assign n24197 = ~n24195 & ~n24196;
  assign n24198 = n22860 & ~n24197;
  assign po2228 = n24194 | n24198;
  assign n24200 = ~pi2053 & ~n22860;
  assign n24201 = n22909 & ~n23625;
  assign n24202 = ~pi2053 & ~n22909;
  assign n24203 = ~n24201 & ~n24202;
  assign n24204 = n22860 & ~n24203;
  assign po2229 = n24200 | n24204;
  assign n24206 = ~pi2054 & ~n22860;
  assign n24207 = n22909 & ~n23327;
  assign n24208 = ~pi2054 & ~n22909;
  assign n24209 = ~n24207 & ~n24208;
  assign n24210 = n22860 & ~n24209;
  assign po2230 = n24206 | n24210;
  assign n24212 = ~pi2055 & ~n22860;
  assign n24213 = n22909 & ~n24002;
  assign n24214 = ~pi2055 & ~n22909;
  assign n24215 = ~n24213 & ~n24214;
  assign n24216 = n22860 & ~n24215;
  assign po2231 = n24212 | n24216;
  assign n24218 = ~pi2056 & ~n22860;
  assign n24219 = n22909 & ~n23306;
  assign n24220 = ~pi2056 & ~n22909;
  assign n24221 = ~n24219 & ~n24220;
  assign n24222 = n22860 & ~n24221;
  assign po2232 = n24218 | n24222;
  assign n24224 = ~pi2057 & ~n22860;
  assign n24225 = n22909 & ~n23334;
  assign n24226 = ~pi2057 & ~n22909;
  assign n24227 = ~n24225 & ~n24226;
  assign n24228 = n22860 & ~n24227;
  assign po2233 = n24224 | n24228;
  assign n24230 = ~pi2058 & ~n22860;
  assign n24231 = n22909 & ~n23341;
  assign n24232 = ~pi2058 & ~n22909;
  assign n24233 = ~n24231 & ~n24232;
  assign n24234 = n22860 & ~n24233;
  assign po2234 = n24230 | n24234;
  assign n24236 = ~pi2059 & ~n22860;
  assign n24237 = n22917 & ~n23448;
  assign n24238 = ~pi2059 & ~n22917;
  assign n24239 = ~n24237 & ~n24238;
  assign n24240 = n22860 & ~n24239;
  assign po2235 = n24236 | n24240;
  assign n24242 = ~pi2060 & ~n22860;
  assign n24243 = n22917 & ~n23428;
  assign n24244 = ~pi2060 & ~n22917;
  assign n24245 = ~n24243 & ~n24244;
  assign n24246 = n22860 & ~n24245;
  assign po2236 = n24242 | n24246;
  assign n24248 = ~pi2061 & ~n22860;
  assign n24249 = n22917 & ~n23320;
  assign n24250 = ~pi2061 & ~n22917;
  assign n24251 = ~n24249 & ~n24250;
  assign n24252 = n22860 & ~n24251;
  assign po2237 = n24248 | n24252;
  assign n24254 = ~pi2062 & ~n22860;
  assign n24255 = n22917 & ~n23518;
  assign n24256 = ~pi2062 & ~n22917;
  assign n24257 = ~n24255 & ~n24256;
  assign n24258 = n22860 & ~n24257;
  assign po2238 = n24254 | n24258;
  assign n24260 = ~pi2063 & ~n22860;
  assign n24261 = n22917 & ~n23381;
  assign n24262 = ~pi2063 & ~n22917;
  assign n24263 = ~n24261 & ~n24262;
  assign n24264 = n22860 & ~n24263;
  assign po2239 = n24260 | n24264;
  assign n24266 = ~pi2064 & ~n22860;
  assign n24267 = n22917 & ~n23557;
  assign n24268 = ~pi2064 & ~n22917;
  assign n24269 = ~n24267 & ~n24268;
  assign n24270 = n22860 & ~n24269;
  assign po2240 = n24266 | n24270;
  assign n24272 = ~pi2065 & ~n22860;
  assign n24273 = n22917 & ~n23537;
  assign n24274 = ~pi2065 & ~n22917;
  assign n24275 = ~n24273 & ~n24274;
  assign n24276 = n22860 & ~n24275;
  assign po2241 = n24272 | n24276;
  assign n24278 = ~pi2066 & ~n22860;
  assign n24279 = n22917 & ~n23625;
  assign n24280 = ~pi2066 & ~n22917;
  assign n24281 = ~n24279 & ~n24280;
  assign n24282 = n22860 & ~n24281;
  assign po2242 = n24278 | n24282;
  assign n24284 = ~pi2067 & ~n22860;
  assign n24285 = n22917 & ~n23408;
  assign n24286 = ~pi2067 & ~n22917;
  assign n24287 = ~n24285 & ~n24286;
  assign n24288 = n22860 & ~n24287;
  assign po2243 = n24284 | n24288;
  assign n24290 = ~pi2068 & ~n22860;
  assign n24291 = n22917 & ~n23313;
  assign n24292 = ~pi2068 & ~n22917;
  assign n24293 = ~n24291 & ~n24292;
  assign n24294 = n22860 & ~n24293;
  assign po2244 = n24290 | n24294;
  assign n24296 = ~pi2069 & ~n22860;
  assign n24297 = n22917 & ~n23306;
  assign n24298 = ~pi2069 & ~n22917;
  assign n24299 = ~n24297 & ~n24298;
  assign n24300 = n22860 & ~n24299;
  assign po2245 = n24296 | n24300;
  assign n24302 = ~pi2070 & ~n22860;
  assign n24303 = n22917 & ~n23388;
  assign n24304 = ~pi2070 & ~n22917;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = n22860 & ~n24305;
  assign po2246 = n24302 | n24306;
  assign n24308 = ~pi2071 & ~n22860;
  assign n24309 = n22917 & ~n23341;
  assign n24310 = ~pi2071 & ~n22917;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = n22860 & ~n24311;
  assign po2247 = n24308 | n24312;
  assign n24314 = ~pi2072 & ~n22860;
  assign n24315 = n22924 & ~n23348;
  assign n24316 = ~pi2072 & ~n22924;
  assign n24317 = ~n24315 & ~n24316;
  assign n24318 = n22860 & ~n24317;
  assign po2248 = n24314 | n24318;
  assign n24320 = ~pi2073 & ~n22860;
  assign n24321 = n22924 & ~n23368;
  assign n24322 = ~pi2073 & ~n22924;
  assign n24323 = ~n24321 & ~n24322;
  assign n24324 = n22860 & ~n24323;
  assign po2249 = n24320 | n24324;
  assign n24326 = ~pi2074 & ~n22860;
  assign n24327 = n22924 & ~n23355;
  assign n24328 = ~pi2074 & ~n22924;
  assign n24329 = ~n24327 & ~n24328;
  assign n24330 = n22860 & ~n24329;
  assign po2250 = n24326 | n24330;
  assign n24332 = ~pi2075 & ~n22860;
  assign n24333 = n22924 & ~n23953;
  assign n24334 = ~pi2075 & ~n22924;
  assign n24335 = ~n24333 & ~n24334;
  assign n24336 = n22860 & ~n24335;
  assign po2251 = n24332 | n24336;
  assign n24338 = ~pi2076 & ~n22860;
  assign n24339 = n22924 & ~n23638;
  assign n24340 = ~pi2076 & ~n22924;
  assign n24341 = ~n24339 & ~n24340;
  assign n24342 = n22860 & ~n24341;
  assign po2252 = n24338 | n24342;
  assign n24344 = ~pi2077 & ~n22860;
  assign n24345 = n22924 & ~n23511;
  assign n24346 = ~pi2077 & ~n22924;
  assign n24347 = ~n24345 & ~n24346;
  assign n24348 = n22860 & ~n24347;
  assign po2253 = n24344 | n24348;
  assign n24350 = ~pi2078 & ~n22860;
  assign n24351 = n22924 & ~n23862;
  assign n24352 = ~pi2078 & ~n22924;
  assign n24353 = ~n24351 & ~n24352;
  assign n24354 = n22860 & ~n24353;
  assign po2254 = n24350 | n24354;
  assign n24356 = ~pi2079 & ~n22860;
  assign n24357 = n22924 & ~n23570;
  assign n24358 = ~pi2079 & ~n22924;
  assign n24359 = ~n24357 & ~n24358;
  assign n24360 = n22860 & ~n24359;
  assign po2255 = n24356 | n24360;
  assign n24362 = ~pi2080 & ~n22860;
  assign n24363 = n22924 & ~n23550;
  assign n24364 = ~pi2080 & ~n22924;
  assign n24365 = ~n24363 & ~n24364;
  assign n24366 = n22860 & ~n24365;
  assign po2256 = n24362 | n24366;
  assign n24368 = ~pi2081 & ~n22860;
  assign n24369 = n22924 & ~n23408;
  assign n24370 = ~pi2081 & ~n22924;
  assign n24371 = ~n24369 & ~n24370;
  assign n24372 = n22860 & ~n24371;
  assign po2257 = n24368 | n24372;
  assign n24374 = ~pi2082 & ~n22860;
  assign n24375 = n22924 & ~n23474;
  assign n24376 = ~pi2082 & ~n22924;
  assign n24377 = ~n24375 & ~n24376;
  assign n24378 = n22860 & ~n24377;
  assign po2258 = n24374 | n24378;
  assign n24380 = ~pi2083 & ~n22860;
  assign n24381 = n22924 & ~n23327;
  assign n24382 = ~pi2083 & ~n22924;
  assign n24383 = ~n24381 & ~n24382;
  assign n24384 = n22860 & ~n24383;
  assign po2259 = n24380 | n24384;
  assign n24386 = ~pi2084 & ~n22860;
  assign n24387 = n22924 & ~n24002;
  assign n24388 = ~pi2084 & ~n22924;
  assign n24389 = ~n24387 & ~n24388;
  assign n24390 = n22860 & ~n24389;
  assign po2260 = n24386 | n24390;
  assign n24392 = ~pi2085 & ~n22860;
  assign n24393 = n22973 & ~n23862;
  assign n24394 = ~pi2085 & ~n22973;
  assign n24395 = ~n24393 & ~n24394;
  assign n24396 = n22860 & ~n24395;
  assign po2261 = n24392 | n24396;
  assign n24398 = ~pi2086 & ~n22860;
  assign n24399 = n22924 & ~n23334;
  assign n24400 = ~pi2086 & ~n22924;
  assign n24401 = ~n24399 & ~n24400;
  assign n24402 = n22860 & ~n24401;
  assign po2262 = n24398 | n24402;
  assign n24404 = ~pi2087 & ~n22860;
  assign n24405 = n22924 & ~n23341;
  assign n24406 = ~pi2087 & ~n22924;
  assign n24407 = ~n24405 & ~n24406;
  assign n24408 = n22860 & ~n24407;
  assign po2263 = n24404 | n24408;
  assign n24410 = ~pi2088 & ~n22860;
  assign n24411 = n22931 & ~n23448;
  assign n24412 = ~pi2088 & ~n22931;
  assign n24413 = ~n24411 & ~n24412;
  assign n24414 = n22860 & ~n24413;
  assign po2264 = n24410 | n24414;
  assign n24416 = ~pi2089 & ~n22860;
  assign n24417 = n22931 & ~n23428;
  assign n24418 = ~pi2089 & ~n22931;
  assign n24419 = ~n24417 & ~n24418;
  assign n24420 = n22860 & ~n24419;
  assign po2265 = n24416 | n24420;
  assign n24422 = ~pi2090 & ~n22860;
  assign n24423 = n22931 & ~n23518;
  assign n24424 = ~pi2090 & ~n22931;
  assign n24425 = ~n24423 & ~n24424;
  assign n24426 = n22860 & ~n24425;
  assign po2266 = n24422 | n24426;
  assign n24428 = ~pi2091 & ~n22860;
  assign n24429 = n22931 & ~n23368;
  assign n24430 = ~pi2091 & ~n22931;
  assign n24431 = ~n24429 & ~n24430;
  assign n24432 = n22860 & ~n24431;
  assign po2267 = n24428 | n24432;
  assign n24434 = ~pi2092 & ~n22860;
  assign n24435 = n22931 & ~n23381;
  assign n24436 = ~pi2092 & ~n22931;
  assign n24437 = ~n24435 & ~n24436;
  assign n24438 = n22860 & ~n24437;
  assign po2268 = n24434 | n24438;
  assign n24440 = ~pi2093 & ~n22860;
  assign n24441 = n22931 & ~n23645;
  assign n24442 = ~pi2093 & ~n22931;
  assign n24443 = ~n24441 & ~n24442;
  assign n24444 = n22860 & ~n24443;
  assign po2269 = n24440 | n24444;
  assign n24446 = ~pi2094 & ~n22860;
  assign n24447 = n22931 & ~n23355;
  assign n24448 = ~pi2094 & ~n22931;
  assign n24449 = ~n24447 & ~n24448;
  assign n24450 = n22860 & ~n24449;
  assign po2270 = n24446 | n24450;
  assign n24452 = ~pi2095 & ~n22860;
  assign n24453 = n22931 & ~n23557;
  assign n24454 = ~pi2095 & ~n22931;
  assign n24455 = ~n24453 & ~n24454;
  assign n24456 = n22860 & ~n24455;
  assign po2271 = n24452 | n24456;
  assign n24458 = ~pi2096 & ~n22860;
  assign n24459 = n22931 & ~n23664;
  assign n24460 = ~pi2096 & ~n22931;
  assign n24461 = ~n24459 & ~n24460;
  assign n24462 = n22860 & ~n24461;
  assign po2272 = n24458 | n24462;
  assign n24464 = ~pi2097 & ~n22860;
  assign n24465 = n22931 & ~n23638;
  assign n24466 = ~pi2097 & ~n22931;
  assign n24467 = ~n24465 & ~n24466;
  assign n24468 = n22860 & ~n24467;
  assign po2273 = n24464 | n24468;
  assign n24470 = ~pi2098 & ~n22860;
  assign n24471 = n22931 & ~n23511;
  assign n24472 = ~pi2098 & ~n22931;
  assign n24473 = ~n24471 & ~n24472;
  assign n24474 = n22860 & ~n24473;
  assign po2274 = n24470 | n24474;
  assign n24476 = ~pi2099 & ~n22860;
  assign n24477 = n22931 & ~n23415;
  assign n24478 = ~pi2099 & ~n22931;
  assign n24479 = ~n24477 & ~n24478;
  assign n24480 = n22860 & ~n24479;
  assign po2275 = n24476 | n24480;
  assign n24482 = ~pi2100 & ~n22860;
  assign n24483 = n22931 & ~n23537;
  assign n24484 = ~pi2100 & ~n22931;
  assign n24485 = ~n24483 & ~n24484;
  assign n24486 = n22860 & ~n24485;
  assign po2276 = n24482 | n24486;
  assign n24488 = ~pi2101 & ~n22860;
  assign n24489 = n22931 & ~n23481;
  assign n24490 = ~pi2101 & ~n22931;
  assign n24491 = ~n24489 & ~n24490;
  assign n24492 = n22860 & ~n24491;
  assign po2277 = n24488 | n24492;
  assign n24494 = ~pi2102 & ~n22860;
  assign n24495 = n22931 & ~n23474;
  assign n24496 = ~pi2102 & ~n22931;
  assign n24497 = ~n24495 & ~n24496;
  assign n24498 = n22860 & ~n24497;
  assign po2278 = n24494 | n24498;
  assign n24500 = ~pi2103 & ~n22860;
  assign n24501 = n22931 & ~n23408;
  assign n24502 = ~pi2103 & ~n22931;
  assign n24503 = ~n24501 & ~n24502;
  assign n24504 = n22860 & ~n24503;
  assign po2279 = n24500 | n24504;
  assign n24506 = ~pi2104 & ~n22860;
  assign n24507 = n22931 & ~n23313;
  assign n24508 = ~pi2104 & ~n22931;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = n22860 & ~n24509;
  assign po2280 = n24506 | n24510;
  assign n24512 = ~pi2105 & ~n22860;
  assign n24513 = n22931 & ~n23306;
  assign n24514 = ~pi2105 & ~n22931;
  assign n24515 = ~n24513 & ~n24514;
  assign n24516 = n22860 & ~n24515;
  assign po2281 = n24512 | n24516;
  assign n24518 = ~pi2106 & ~n22860;
  assign n24519 = n22931 & ~n23388;
  assign n24520 = ~pi2106 & ~n22931;
  assign n24521 = ~n24519 & ~n24520;
  assign n24522 = n22860 & ~n24521;
  assign po2282 = n24518 | n24522;
  assign n24524 = ~pi2107 & ~n22860;
  assign n24525 = n22966 & ~n23348;
  assign n24526 = ~pi2107 & ~n22966;
  assign n24527 = ~n24525 & ~n24526;
  assign n24528 = n22860 & ~n24527;
  assign po2283 = n24524 | n24528;
  assign n24530 = ~pi2108 & ~n22860;
  assign n24531 = n22966 & ~n23461;
  assign n24532 = ~pi2108 & ~n22966;
  assign n24533 = ~n24531 & ~n24532;
  assign n24534 = n22860 & ~n24533;
  assign po2284 = n24530 | n24534;
  assign n24536 = ~pi2109 & ~n22860;
  assign n24537 = n22966 & ~n23320;
  assign n24538 = ~pi2109 & ~n22966;
  assign n24539 = ~n24537 & ~n24538;
  assign n24540 = n22860 & ~n24539;
  assign po2285 = n24536 | n24540;
  assign n24542 = ~pi2110 & ~n22860;
  assign n24543 = n22966 & ~n23518;
  assign n24544 = ~pi2110 & ~n22966;
  assign n24545 = ~n24543 & ~n24544;
  assign n24546 = n22860 & ~n24545;
  assign po2286 = n24542 | n24546;
  assign n24548 = ~pi2111 & ~n22860;
  assign n24549 = n22966 & ~n23368;
  assign n24550 = ~pi2111 & ~n22966;
  assign n24551 = ~n24549 & ~n24550;
  assign n24552 = n22860 & ~n24551;
  assign po2287 = n24548 | n24552;
  assign n24554 = ~pi2112 & ~n22860;
  assign n24555 = n22966 & ~n23395;
  assign n24556 = ~pi2112 & ~n22966;
  assign n24557 = ~n24555 & ~n24556;
  assign n24558 = n22860 & ~n24557;
  assign po2288 = n24554 | n24558;
  assign n24560 = ~pi2113 & ~n22860;
  assign n24561 = n22966 & ~n23645;
  assign n24562 = ~pi2113 & ~n22966;
  assign n24563 = ~n24561 & ~n24562;
  assign n24564 = n22860 & ~n24563;
  assign po2289 = n24560 | n24564;
  assign n24566 = ~pi2114 & ~n22860;
  assign n24567 = n22966 & ~n23355;
  assign n24568 = ~pi2114 & ~n22966;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = n22860 & ~n24569;
  assign po2290 = n24566 | n24570;
  assign n24572 = ~pi2115 & ~n22860;
  assign n24573 = n22966 & ~n23953;
  assign n24574 = ~pi2115 & ~n22966;
  assign n24575 = ~n24573 & ~n24574;
  assign n24576 = n22860 & ~n24575;
  assign po2291 = n24572 | n24576;
  assign n24578 = ~pi2116 & ~n22860;
  assign n24579 = n22966 & ~n23664;
  assign n24580 = ~pi2116 & ~n22966;
  assign n24581 = ~n24579 & ~n24580;
  assign n24582 = n22860 & ~n24581;
  assign po2292 = n24578 | n24582;
  assign n24584 = ~pi2117 & ~n22860;
  assign n24585 = n22966 & ~n23638;
  assign n24586 = ~pi2117 & ~n22966;
  assign n24587 = ~n24585 & ~n24586;
  assign n24588 = n22860 & ~n24587;
  assign po2293 = n24584 | n24588;
  assign n24590 = ~pi2118 & ~n22860;
  assign n24591 = n22966 & ~n23862;
  assign n24592 = ~pi2118 & ~n22966;
  assign n24593 = ~n24591 & ~n24592;
  assign n24594 = n22860 & ~n24593;
  assign po2294 = n24590 | n24594;
  assign n24596 = ~pi2119 & ~n22860;
  assign n24597 = n22966 & ~n23570;
  assign n24598 = ~pi2119 & ~n22966;
  assign n24599 = ~n24597 & ~n24598;
  assign n24600 = n22860 & ~n24599;
  assign po2295 = n24596 | n24600;
  assign n24602 = ~pi2120 & ~n22860;
  assign n24603 = n22966 & ~n23550;
  assign n24604 = ~pi2120 & ~n22966;
  assign n24605 = ~n24603 & ~n24604;
  assign n24606 = n22860 & ~n24605;
  assign po2296 = n24602 | n24606;
  assign n24608 = ~pi2121 & ~n22860;
  assign n24609 = n22966 & ~n23481;
  assign n24610 = ~pi2121 & ~n22966;
  assign n24611 = ~n24609 & ~n24610;
  assign n24612 = n22860 & ~n24611;
  assign po2297 = n24608 | n24612;
  assign n24614 = ~pi2122 & ~n22860;
  assign n24615 = n22966 & ~n23474;
  assign n24616 = ~pi2122 & ~n22966;
  assign n24617 = ~n24615 & ~n24616;
  assign n24618 = n22860 & ~n24617;
  assign po2298 = n24614 | n24618;
  assign n24620 = ~pi2123 & ~n22860;
  assign n24621 = ~pi2123 & ~n22879;
  assign n24622 = n22879 & ~n23511;
  assign n24623 = ~n24621 & ~n24622;
  assign n24624 = n22860 & ~n24623;
  assign po2299 = n24620 | n24624;
  assign n24626 = ~pi2124 & ~n22860;
  assign n24627 = n22966 & ~n23341;
  assign n24628 = ~pi2124 & ~n22966;
  assign n24629 = ~n24627 & ~n24628;
  assign n24630 = n22860 & ~n24629;
  assign po2300 = n24626 | n24630;
  assign n24632 = ~pi2125 & ~n22860;
  assign n24633 = n22973 & ~n23448;
  assign n24634 = ~pi2125 & ~n22973;
  assign n24635 = ~n24633 & ~n24634;
  assign n24636 = n22860 & ~n24635;
  assign po2301 = n24632 | n24636;
  assign n24638 = ~pi2126 & ~n22860;
  assign n24639 = n22973 & ~n23428;
  assign n24640 = ~pi2126 & ~n22973;
  assign n24641 = ~n24639 & ~n24640;
  assign n24642 = n22860 & ~n24641;
  assign po2302 = n24638 | n24642;
  assign n24644 = ~pi2127 & ~n22860;
  assign n24645 = n22973 & ~n23557;
  assign n24646 = ~pi2127 & ~n22973;
  assign n24647 = ~n24645 & ~n24646;
  assign n24648 = n22860 & ~n24647;
  assign po2303 = n24644 | n24648;
  assign n24650 = ~pi2128 & ~n22860;
  assign n24651 = n22973 & ~n23664;
  assign n24652 = ~pi2128 & ~n22973;
  assign n24653 = ~n24651 & ~n24652;
  assign n24654 = n22860 & ~n24653;
  assign po2304 = n24650 | n24654;
  assign n24656 = ~pi2129 & ~n22860;
  assign n24657 = ~pi2129 & ~n22879;
  assign n24658 = n22879 & ~n23395;
  assign n24659 = ~n24657 & ~n24658;
  assign n24660 = n22860 & ~n24659;
  assign po2305 = n24656 | n24660;
  assign n24662 = ~pi2130 & ~n22860;
  assign n24663 = n22973 & ~n23537;
  assign n24664 = ~pi2130 & ~n22973;
  assign n24665 = ~n24663 & ~n24664;
  assign n24666 = n22860 & ~n24665;
  assign po2306 = n24662 | n24666;
  assign n24668 = ~pi2131 & ~n22860;
  assign n24669 = n22973 & ~n23408;
  assign n24670 = ~pi2131 & ~n22973;
  assign n24671 = ~n24669 & ~n24670;
  assign n24672 = n22860 & ~n24671;
  assign po2307 = n24668 | n24672;
  assign n24674 = ~pi2132 & ~n22860;
  assign n24675 = n22973 & ~n23313;
  assign n24676 = ~pi2132 & ~n22973;
  assign n24677 = ~n24675 & ~n24676;
  assign n24678 = n22860 & ~n24677;
  assign po2308 = n24674 | n24678;
  assign n24680 = ~pi2133 & ~n22860;
  assign n24681 = n22945 & ~n23448;
  assign n24682 = ~pi2133 & ~n22945;
  assign n24683 = ~n24681 & ~n24682;
  assign n24684 = n22860 & ~n24683;
  assign po2309 = n24680 | n24684;
  assign n24686 = ~pi2134 & ~n22860;
  assign n24687 = n22945 & ~n23428;
  assign n24688 = ~pi2134 & ~n22945;
  assign n24689 = ~n24687 & ~n24688;
  assign n24690 = n22860 & ~n24689;
  assign po2310 = n24686 | n24690;
  assign n24692 = ~pi2135 & ~n22860;
  assign n24693 = n22945 & ~n23518;
  assign n24694 = ~pi2135 & ~n22945;
  assign n24695 = ~n24693 & ~n24694;
  assign n24696 = n22860 & ~n24695;
  assign po2311 = n24692 | n24696;
  assign n24698 = ~pi2136 & ~n22860;
  assign n24699 = n22945 & ~n23381;
  assign n24700 = ~pi2136 & ~n22945;
  assign n24701 = ~n24699 & ~n24700;
  assign n24702 = n22860 & ~n24701;
  assign po2312 = n24698 | n24702;
  assign n24704 = ~pi2137 & ~n22860;
  assign n24705 = n22945 & ~n23645;
  assign n24706 = ~pi2137 & ~n22945;
  assign n24707 = ~n24705 & ~n24706;
  assign n24708 = n22860 & ~n24707;
  assign po2313 = n24704 | n24708;
  assign n24710 = ~pi2138 & ~n22860;
  assign n24711 = n22945 & ~n23355;
  assign n24712 = ~pi2138 & ~n22945;
  assign n24713 = ~n24711 & ~n24712;
  assign n24714 = n22860 & ~n24713;
  assign po2314 = n24710 | n24714;
  assign n24716 = ~pi2139 & ~n22860;
  assign n24717 = n22945 & ~n23557;
  assign n24718 = ~pi2139 & ~n22945;
  assign n24719 = ~n24717 & ~n24718;
  assign n24720 = n22860 & ~n24719;
  assign po2315 = n24716 | n24720;
  assign n24722 = ~pi2140 & ~n22860;
  assign n24723 = n22945 & ~n23664;
  assign n24724 = ~pi2140 & ~n22945;
  assign n24725 = ~n24723 & ~n24724;
  assign n24726 = n22860 & ~n24725;
  assign po2316 = n24722 | n24726;
  assign n24728 = ~pi2141 & ~n22860;
  assign n24729 = n22945 & ~n23511;
  assign n24730 = ~pi2141 & ~n22945;
  assign n24731 = ~n24729 & ~n24730;
  assign n24732 = n22860 & ~n24731;
  assign po2317 = n24728 | n24732;
  assign n24734 = ~pi2142 & ~n22860;
  assign n24735 = n22945 & ~n23415;
  assign n24736 = ~pi2142 & ~n22945;
  assign n24737 = ~n24735 & ~n24736;
  assign n24738 = n22860 & ~n24737;
  assign po2318 = n24734 | n24738;
  assign n24740 = ~pi2143 & ~n22860;
  assign n24741 = n22945 & ~n23481;
  assign n24742 = ~pi2143 & ~n22945;
  assign n24743 = ~n24741 & ~n24742;
  assign n24744 = n22860 & ~n24743;
  assign po2319 = n24740 | n24744;
  assign n24746 = ~pi2144 & ~n22860;
  assign n24747 = n22945 & ~n23313;
  assign n24748 = ~pi2144 & ~n22945;
  assign n24749 = ~n24747 & ~n24748;
  assign n24750 = n22860 & ~n24749;
  assign po2320 = n24746 | n24750;
  assign n24752 = ~pi2145 & ~n22860;
  assign n24753 = n22952 & ~n23348;
  assign n24754 = ~pi2145 & ~n22952;
  assign n24755 = ~n24753 & ~n24754;
  assign n24756 = n22860 & ~n24755;
  assign po2321 = n24752 | n24756;
  assign n24758 = ~pi2146 & ~n22860;
  assign n24759 = n22952 & ~n23320;
  assign n24760 = ~pi2146 & ~n22952;
  assign n24761 = ~n24759 & ~n24760;
  assign n24762 = n22860 & ~n24761;
  assign po2322 = n24758 | n24762;
  assign n24764 = ~pi2147 & ~n22860;
  assign n24765 = n22952 & ~n23862;
  assign n24766 = ~pi2147 & ~n22952;
  assign n24767 = ~n24765 & ~n24766;
  assign n24768 = n22860 & ~n24767;
  assign po2323 = n24764 | n24768;
  assign n24770 = ~pi2148 & ~n22860;
  assign n24771 = n22952 & ~n23570;
  assign n24772 = ~pi2148 & ~n22952;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = n22860 & ~n24773;
  assign po2324 = n24770 | n24774;
  assign n24776 = ~pi2149 & ~n22860;
  assign n24777 = n22952 & ~n23550;
  assign n24778 = ~pi2149 & ~n22952;
  assign n24779 = ~n24777 & ~n24778;
  assign n24780 = n22860 & ~n24779;
  assign po2325 = n24776 | n24780;
  assign n24782 = ~pi2150 & ~n22860;
  assign n24783 = n22952 & ~n23481;
  assign n24784 = ~pi2150 & ~n22952;
  assign n24785 = ~n24783 & ~n24784;
  assign n24786 = n22860 & ~n24785;
  assign po2326 = n24782 | n24786;
  assign n24788 = ~pi2151 & ~n22860;
  assign n24789 = n22952 & ~n23474;
  assign n24790 = ~pi2151 & ~n22952;
  assign n24791 = ~n24789 & ~n24790;
  assign n24792 = n22860 & ~n24791;
  assign po2327 = n24788 | n24792;
  assign n24794 = ~pi2152 & ~n22860;
  assign n24795 = n22952 & ~n23327;
  assign n24796 = ~pi2152 & ~n22952;
  assign n24797 = ~n24795 & ~n24796;
  assign n24798 = n22860 & ~n24797;
  assign po2328 = n24794 | n24798;
  assign n24800 = ~pi2153 & ~n22860;
  assign n24801 = n22952 & ~n24002;
  assign n24802 = ~pi2153 & ~n22952;
  assign n24803 = ~n24801 & ~n24802;
  assign n24804 = n22860 & ~n24803;
  assign po2329 = n24800 | n24804;
  assign n24806 = ~pi2154 & ~n22860;
  assign n24807 = n22952 & ~n23306;
  assign n24808 = ~pi2154 & ~n22952;
  assign n24809 = ~n24807 & ~n24808;
  assign n24810 = n22860 & ~n24809;
  assign po2330 = n24806 | n24810;
  assign n24812 = ~pi2155 & ~n22860;
  assign n24813 = n22952 & ~n23334;
  assign n24814 = ~pi2155 & ~n22952;
  assign n24815 = ~n24813 & ~n24814;
  assign n24816 = n22860 & ~n24815;
  assign po2331 = n24812 | n24816;
  assign n24818 = ~pi2156 & ~n22860;
  assign n24819 = n22952 & ~n23341;
  assign n24820 = ~pi2156 & ~n22952;
  assign n24821 = ~n24819 & ~n24820;
  assign n24822 = n22860 & ~n24821;
  assign po2332 = n24818 | n24822;
  assign n24824 = ~pi2157 & ~n22554;
  assign n24825 = ~pi3082 & n22554;
  assign n24826 = ~n24824 & ~n24825;
  assign n24827 = n22306 & ~n24826;
  assign n24828 = ~pi2157 & ~n22306;
  assign po2333 = n24827 | n24828;
  assign n24830 = ~pi2158 & ~n22561;
  assign n24831 = ~pi3082 & n22561;
  assign n24832 = ~n24830 & ~n24831;
  assign n24833 = n22306 & ~n24832;
  assign n24834 = ~pi2158 & ~n22306;
  assign po2334 = n24833 | n24834;
  assign n24836 = ~pi2159 & ~n22860;
  assign n24837 = pi2975 & n22924;
  assign n24838 = ~pi2159 & ~n22924;
  assign n24839 = ~n24837 & ~n24838;
  assign n24840 = n22860 & ~n24839;
  assign po2335 = n24836 | n24840;
  assign n24842 = ~pi2160 & ~n22860;
  assign n24843 = pi2975 & n22966;
  assign n24844 = ~pi2160 & ~n22966;
  assign n24845 = ~n24843 & ~n24844;
  assign n24846 = n22860 & ~n24845;
  assign po2336 = n24842 | n24846;
  assign n24848 = ~pi2161 & ~n22860;
  assign n24849 = pi2975 & n22952;
  assign n24850 = ~pi2161 & ~n22952;
  assign n24851 = ~n24849 & ~n24850;
  assign n24852 = n22860 & ~n24851;
  assign po2337 = n24848 | n24852;
  assign n24854 = ~pi2162 & ~n22860;
  assign n24855 = n22952 & ~n23518;
  assign n24856 = ~pi2162 & ~n22952;
  assign n24857 = ~n24855 & ~n24856;
  assign n24858 = n22860 & ~n24857;
  assign po2338 = n24854 | n24858;
  assign n24860 = ~pi2163 & ~n22311;
  assign n24861 = ~pi3082 & n22311;
  assign n24862 = ~n24860 & ~n24861;
  assign n24863 = n22306 & ~n24862;
  assign n24864 = ~pi2163 & ~n22306;
  assign po2339 = n24863 | n24864;
  assign n24866 = ~pi2164 & ~n22302;
  assign n24867 = ~pi3082 & n22302;
  assign n24868 = ~n24866 & ~n24867;
  assign n24869 = n22306 & ~n24868;
  assign n24870 = ~pi2164 & ~n22306;
  assign po2340 = n24869 | n24870;
  assign n24872 = ~pi2165 & ~n22860;
  assign n24873 = pi2975 & n22959;
  assign n24874 = ~pi2165 & ~n22959;
  assign n24875 = ~n24873 & ~n24874;
  assign n24876 = n22860 & ~n24875;
  assign po2341 = n24872 | n24876;
  assign n24878 = ~pi2166 & ~n22860;
  assign n24879 = ~pi2166 & ~n22879;
  assign n24880 = n22879 & ~n23320;
  assign n24881 = ~n24879 & ~n24880;
  assign n24882 = n22860 & ~n24881;
  assign po2342 = n24878 | n24882;
  assign n24884 = ~pi2167 & ~n22860;
  assign n24885 = ~pi2167 & ~n22879;
  assign n24886 = n22879 & ~n23368;
  assign n24887 = ~n24885 & ~n24886;
  assign n24888 = n22860 & ~n24887;
  assign po2343 = n24884 | n24888;
  assign n24890 = ~pi2168 & ~n22860;
  assign n24891 = ~pi2168 & ~n22879;
  assign n24892 = n22879 & ~n23355;
  assign n24893 = ~n24891 & ~n24892;
  assign n24894 = n22860 & ~n24893;
  assign po2344 = n24890 | n24894;
  assign n24896 = ~pi2169 & ~n22860;
  assign n24897 = ~pi2169 & ~n22879;
  assign n24898 = n22879 & ~n23953;
  assign n24899 = ~n24897 & ~n24898;
  assign n24900 = n22860 & ~n24899;
  assign po2345 = n24896 | n24900;
  assign n24902 = ~pi2170 & ~n22860;
  assign n24903 = ~pi2170 & ~n22879;
  assign n24904 = n22879 & ~n23862;
  assign n24905 = ~n24903 & ~n24904;
  assign n24906 = n22860 & ~n24905;
  assign po2346 = n24902 | n24906;
  assign n24908 = ~pi2171 & ~n22860;
  assign n24909 = ~pi2171 & ~n22879;
  assign n24910 = n22879 & ~n23550;
  assign n24911 = ~n24909 & ~n24910;
  assign n24912 = n22860 & ~n24911;
  assign po2347 = n24908 | n24912;
  assign n24914 = ~pi2172 & ~n22860;
  assign n24915 = ~pi2172 & ~n22879;
  assign n24916 = n22879 & ~n23625;
  assign n24917 = ~n24915 & ~n24916;
  assign n24918 = n22860 & ~n24917;
  assign po2348 = n24914 | n24918;
  assign n24920 = ~pi2173 & ~n22860;
  assign n24921 = ~pi2173 & ~n22879;
  assign n24922 = n22879 & ~n24002;
  assign n24923 = ~n24921 & ~n24922;
  assign n24924 = n22860 & ~n24923;
  assign po2349 = n24920 | n24924;
  assign n24926 = ~pi2174 & ~n22860;
  assign n24927 = ~pi2174 & ~n22879;
  assign n24928 = n22879 & ~n23341;
  assign n24929 = ~n24927 & ~n24928;
  assign n24930 = n22860 & ~n24929;
  assign po2350 = n24926 | n24930;
  assign n24932 = ~pi2175 & ~n22860;
  assign n24933 = ~pi2175 & ~n22893;
  assign n24934 = n22893 & ~n23448;
  assign n24935 = ~n24933 & ~n24934;
  assign n24936 = n22860 & ~n24935;
  assign po2351 = n24932 | n24936;
  assign n24938 = ~pi2176 & ~n22860;
  assign n24939 = ~pi2176 & ~n22893;
  assign n24940 = n22893 & ~n23518;
  assign n24941 = ~n24939 & ~n24940;
  assign n24942 = n22860 & ~n24941;
  assign po2352 = n24938 | n24942;
  assign n24944 = ~pi2177 & ~n22860;
  assign n24945 = ~pi2177 & ~n22893;
  assign n24946 = n22893 & ~n23557;
  assign n24947 = ~n24945 & ~n24946;
  assign n24948 = n22860 & ~n24947;
  assign po2353 = n24944 | n24948;
  assign n24950 = ~pi2178 & ~n22860;
  assign n24951 = ~pi2178 & ~n22893;
  assign n24952 = n22893 & ~n23511;
  assign n24953 = ~n24951 & ~n24952;
  assign n24954 = n22860 & ~n24953;
  assign po2354 = n24950 | n24954;
  assign n24956 = ~pi2179 & ~n22860;
  assign n24957 = ~pi2179 & ~n22900;
  assign n24958 = n22900 & ~n23313;
  assign n24959 = ~n24957 & ~n24958;
  assign n24960 = n22860 & ~n24959;
  assign po2355 = n24956 | n24960;
  assign n24962 = ~pi2180 & ~n22860;
  assign n24963 = ~pi2180 & ~n22893;
  assign n24964 = n22893 & ~n23537;
  assign n24965 = ~n24963 & ~n24964;
  assign n24966 = n22860 & ~n24965;
  assign po2356 = n24962 | n24966;
  assign n24968 = ~pi2181 & ~n22860;
  assign n24969 = ~pi2181 & ~n22893;
  assign n24970 = n22893 & ~n23481;
  assign n24971 = ~n24969 & ~n24970;
  assign n24972 = n22860 & ~n24971;
  assign po2357 = n24968 | n24972;
  assign n24974 = ~pi2182 & ~n22860;
  assign n24975 = ~pi2182 & ~n22893;
  assign n24976 = n22893 & ~n23313;
  assign n24977 = ~n24975 & ~n24976;
  assign n24978 = n22860 & ~n24977;
  assign po2358 = n24974 | n24978;
  assign n24980 = ~pi2183 & ~n22860;
  assign n24981 = ~pi2183 & ~n22893;
  assign n24982 = n22893 & ~n23306;
  assign n24983 = ~n24981 & ~n24982;
  assign n24984 = n22860 & ~n24983;
  assign po2359 = n24980 | n24984;
  assign n24986 = ~pi2184 & ~n22860;
  assign n24987 = ~pi2184 & ~n22893;
  assign n24988 = n22893 & ~n23388;
  assign n24989 = ~n24987 & ~n24988;
  assign n24990 = n22860 & ~n24989;
  assign po2360 = n24986 | n24990;
  assign n24992 = ~pi2185 & ~n22860;
  assign n24993 = ~pi2185 & ~n22900;
  assign n24994 = n22900 & ~n23348;
  assign n24995 = ~n24993 & ~n24994;
  assign n24996 = n22860 & ~n24995;
  assign po2361 = n24992 | n24996;
  assign n24998 = ~pi2186 & ~n22860;
  assign n24999 = ~pi2186 & ~n22900;
  assign n25000 = n22900 & ~n23355;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = n22860 & ~n25001;
  assign po2362 = n24998 | n25002;
  assign n25004 = ~pi2187 & ~n22860;
  assign n25005 = ~pi2187 & ~n22900;
  assign n25006 = n22900 & ~n23953;
  assign n25007 = ~n25005 & ~n25006;
  assign n25008 = n22860 & ~n25007;
  assign po2363 = n25004 | n25008;
  assign n25010 = ~pi2188 & ~n22860;
  assign n25011 = ~pi2188 & ~n22900;
  assign n25012 = n22900 & ~n23638;
  assign n25013 = ~n25011 & ~n25012;
  assign n25014 = n22860 & ~n25013;
  assign po2364 = n25010 | n25014;
  assign n25016 = ~pi2189 & ~n22860;
  assign n25017 = ~pi2189 & ~n22900;
  assign n25018 = n22900 & ~n23474;
  assign n25019 = ~n25017 & ~n25018;
  assign n25020 = n22860 & ~n25019;
  assign po2365 = n25016 | n25020;
  assign n25022 = ~pi2190 & ~n22860;
  assign n25023 = ~pi2190 & ~n22900;
  assign n25024 = n22900 & ~n23625;
  assign n25025 = ~n25023 & ~n25024;
  assign n25026 = n22860 & ~n25025;
  assign po2366 = n25022 | n25026;
  assign n25028 = ~pi2191 & ~n22860;
  assign n25029 = ~pi2191 & ~n22900;
  assign n25030 = n22900 & ~n23327;
  assign n25031 = ~n25029 & ~n25030;
  assign n25032 = n22860 & ~n25031;
  assign po2367 = n25028 | n25032;
  assign n25034 = ~pi2192 & ~n22860;
  assign n25035 = ~pi2192 & ~n22900;
  assign n25036 = n22900 & ~n24002;
  assign n25037 = ~n25035 & ~n25036;
  assign n25038 = n22860 & ~n25037;
  assign po2368 = n25034 | n25038;
  assign n25040 = ~pi2193 & ~n22860;
  assign n25041 = ~pi2193 & ~n22980;
  assign n25042 = n22980 & ~n23518;
  assign n25043 = ~n25041 & ~n25042;
  assign n25044 = n22860 & ~n25043;
  assign po2369 = n25040 | n25044;
  assign n25046 = ~pi2194 & ~n22860;
  assign n25047 = ~pi2194 & ~n22980;
  assign n25048 = n22980 & ~n23645;
  assign n25049 = ~n25047 & ~n25048;
  assign n25050 = n22860 & ~n25049;
  assign po2370 = n25046 | n25050;
  assign n25052 = ~pi2195 & ~n22860;
  assign n25053 = ~pi2195 & ~n22980;
  assign n25054 = n22980 & ~n23557;
  assign n25055 = ~n25053 & ~n25054;
  assign n25056 = n22860 & ~n25055;
  assign po2371 = n25052 | n25056;
  assign n25058 = ~pi2196 & ~n22860;
  assign n25059 = ~pi2196 & ~n22980;
  assign n25060 = n22980 & ~n23415;
  assign n25061 = ~n25059 & ~n25060;
  assign n25062 = n22860 & ~n25061;
  assign po2372 = n25058 | n25062;
  assign n25064 = ~pi2197 & ~n22860;
  assign n25065 = ~pi2197 & ~n22980;
  assign n25066 = n22980 & ~n23537;
  assign n25067 = ~n25065 & ~n25066;
  assign n25068 = n22860 & ~n25067;
  assign po2373 = n25064 | n25068;
  assign n25070 = ~pi2198 & ~n22860;
  assign n25071 = ~pi2198 & ~n22900;
  assign n25072 = n22900 & ~n23481;
  assign n25073 = ~n25071 & ~n25072;
  assign n25074 = n22860 & ~n25073;
  assign po2374 = n25070 | n25074;
  assign n25076 = ~pi2199 & ~n22860;
  assign n25077 = ~pi2199 & ~n22980;
  assign n25078 = n22980 & ~n23481;
  assign n25079 = ~n25077 & ~n25078;
  assign n25080 = n22860 & ~n25079;
  assign po2375 = n25076 | n25080;
  assign n25082 = ~pi2200 & ~n22860;
  assign n25083 = ~pi2200 & ~n22980;
  assign n25084 = n22980 & ~n23408;
  assign n25085 = ~n25083 & ~n25084;
  assign n25086 = n22860 & ~n25085;
  assign po2376 = n25082 | n25086;
  assign n25088 = ~pi2201 & ~n22860;
  assign n25089 = ~pi2201 & ~n22980;
  assign n25090 = pi2975 & n22980;
  assign n25091 = ~n25089 & ~n25090;
  assign n25092 = n22860 & ~n25091;
  assign po2377 = n25088 | n25092;
  assign n25094 = ~pi2202 & ~n22860;
  assign n25095 = pi2975 & n22909;
  assign n25096 = ~pi2202 & ~n22909;
  assign n25097 = ~n25095 & ~n25096;
  assign n25098 = n22860 & ~n25097;
  assign po2378 = n25094 | n25098;
  assign n25100 = ~pi2203 & ~n22860;
  assign n25101 = pi2975 & n22931;
  assign n25102 = ~pi2203 & ~n22931;
  assign n25103 = ~n25101 & ~n25102;
  assign n25104 = n22860 & ~n25103;
  assign po2379 = n25100 | n25104;
  assign n25106 = ~pi2204 & ~n22860;
  assign n25107 = ~pi2204 & ~n22938;
  assign n25108 = n22938 & ~n23448;
  assign n25109 = ~n25107 & ~n25108;
  assign n25110 = n22860 & ~n25109;
  assign po2380 = n25106 | n25110;
  assign n25112 = ~pi2205 & ~n22860;
  assign n25113 = ~pi2205 & ~n22938;
  assign n25114 = n22938 & ~n23518;
  assign n25115 = ~n25113 & ~n25114;
  assign n25116 = n22860 & ~n25115;
  assign po2381 = n25112 | n25116;
  assign n25118 = ~pi2206 & ~n22860;
  assign n25119 = ~pi2206 & ~n22938;
  assign n25120 = n22938 & ~n23645;
  assign n25121 = ~n25119 & ~n25120;
  assign n25122 = n22860 & ~n25121;
  assign po2382 = n25118 | n25122;
  assign n25124 = ~pi2207 & ~n22860;
  assign n25125 = ~pi2207 & ~n22938;
  assign n25126 = n22938 & ~n23557;
  assign n25127 = ~n25125 & ~n25126;
  assign n25128 = n22860 & ~n25127;
  assign po2383 = n25124 | n25128;
  assign n25130 = ~pi2208 & ~n22860;
  assign n25131 = ~pi2208 & ~n22938;
  assign n25132 = n22938 & ~n23511;
  assign n25133 = ~n25131 & ~n25132;
  assign n25134 = n22860 & ~n25133;
  assign po2384 = n25130 | n25134;
  assign n25136 = ~pi2209 & ~n22860;
  assign n25137 = ~pi2209 & ~n22938;
  assign n25138 = n22938 & ~n23481;
  assign n25139 = ~n25137 & ~n25138;
  assign n25140 = n22860 & ~n25139;
  assign po2385 = n25136 | n25140;
  assign n25142 = ~pi2210 & ~n22860;
  assign n25143 = ~pi2210 & ~n22938;
  assign n25144 = pi2975 & n22938;
  assign n25145 = ~n25143 & ~n25144;
  assign n25146 = n22860 & ~n25145;
  assign po2386 = n25142 | n25146;
  assign n25148 = ~pi2211 & ~n22860;
  assign n25149 = ~pi2211 & ~n22938;
  assign n25150 = n22938 & ~n23306;
  assign n25151 = ~n25149 & ~n25150;
  assign n25152 = n22860 & ~n25151;
  assign po2387 = n25148 | n25152;
  assign n25154 = ~pi2212 & ~n22860;
  assign n25155 = ~pi2212 & ~n22879;
  assign n25156 = n22879 & ~n23381;
  assign n25157 = ~n25155 & ~n25156;
  assign n25158 = n22860 & ~n25157;
  assign po2388 = n25154 | n25158;
  assign n25160 = ~pi2213 & ~n22860;
  assign n25161 = ~pi2213 & ~n22879;
  assign n25162 = n22879 & ~n23645;
  assign n25163 = ~n25161 & ~n25162;
  assign n25164 = n22860 & ~n25163;
  assign po2389 = n25160 | n25164;
  assign n25166 = ~pi2214 & ~n22860;
  assign n25167 = ~pi2214 & ~n22900;
  assign n25168 = n22900 & ~n23408;
  assign n25169 = ~n25167 & ~n25168;
  assign n25170 = n22860 & ~n25169;
  assign po2390 = n25166 | n25170;
  assign n25172 = ~pi2215 & ~n22860;
  assign n25173 = ~pi2215 & ~n22879;
  assign n25174 = n22879 & ~n23638;
  assign n25175 = ~n25173 & ~n25174;
  assign n25176 = n22860 & ~n25175;
  assign po2391 = n25172 | n25176;
  assign n25178 = ~pi2216 & ~n22860;
  assign n25179 = ~pi2216 & ~n22879;
  assign n25180 = n22879 & ~n23664;
  assign n25181 = ~n25179 & ~n25180;
  assign n25182 = n22860 & ~n25181;
  assign po2392 = n25178 | n25182;
  assign n25184 = ~pi2217 & ~n22860;
  assign n25185 = ~pi2217 & ~n22900;
  assign n25186 = pi2975 & n22900;
  assign n25187 = ~n25185 & ~n25186;
  assign n25188 = n22860 & ~n25187;
  assign po2393 = n25184 | n25188;
  assign n25190 = ~pi2218 & ~n22860;
  assign n25191 = ~pi2218 & ~n22879;
  assign n25192 = n22879 & ~n23557;
  assign n25193 = ~n25191 & ~n25192;
  assign n25194 = n22860 & ~n25193;
  assign po2394 = n25190 | n25194;
  assign n25196 = ~pi2219 & ~n22860;
  assign n25197 = ~pi2219 & ~n22900;
  assign n25198 = n22900 & ~n23557;
  assign n25199 = ~n25197 & ~n25198;
  assign n25200 = n22860 & ~n25199;
  assign po2395 = n25196 | n25200;
  assign n25202 = ~pi2220 & ~n22860;
  assign n25203 = ~pi2220 & ~n22900;
  assign n25204 = n22900 & ~n23570;
  assign n25205 = ~n25203 & ~n25204;
  assign n25206 = n22860 & ~n25205;
  assign po2396 = n25202 | n25206;
  assign n25208 = ~pi2221 & ~n22860;
  assign n25209 = ~pi2221 & ~n22879;
  assign n25210 = n22879 & ~n23518;
  assign n25211 = ~n25209 & ~n25210;
  assign n25212 = n22860 & ~n25211;
  assign po2397 = n25208 | n25212;
  assign n25214 = ~pi2222 & ~n22860;
  assign n25215 = ~pi2222 & ~n22900;
  assign n25216 = n22900 & ~n23537;
  assign n25217 = ~n25215 & ~n25216;
  assign n25218 = n22860 & ~n25217;
  assign po2398 = n25214 | n25218;
  assign n25220 = ~pi2223 & ~n22860;
  assign n25221 = ~pi2223 & ~n22900;
  assign n25222 = n22900 & ~n23550;
  assign n25223 = ~n25221 & ~n25222;
  assign n25224 = n22860 & ~n25223;
  assign po2399 = n25220 | n25224;
  assign n25226 = ~pi2224 & ~n22860;
  assign n25227 = ~pi2224 & ~n22900;
  assign n25228 = n22900 & ~n23448;
  assign n25229 = ~n25227 & ~n25228;
  assign n25230 = n22860 & ~n25229;
  assign po2400 = n25226 | n25230;
  assign n25232 = ~pi2225 & ~n22860;
  assign n25233 = ~pi2225 & ~n22879;
  assign n25234 = n22879 & ~n23428;
  assign n25235 = ~n25233 & ~n25234;
  assign n25236 = n22860 & ~n25235;
  assign po2401 = n25232 | n25236;
  assign n25238 = ~pi2226 & ~n22860;
  assign n25239 = ~pi2226 & ~n22900;
  assign n25240 = n22900 & ~n23862;
  assign n25241 = ~n25239 & ~n25240;
  assign n25242 = n22860 & ~n25241;
  assign po2402 = n25238 | n25242;
  assign n25244 = ~pi2227 & ~n22860;
  assign n25245 = ~pi2227 & ~n22900;
  assign n25246 = n22900 & ~n23415;
  assign n25247 = ~n25245 & ~n25246;
  assign n25248 = n22860 & ~n25247;
  assign po2403 = n25244 | n25248;
  assign n25250 = ~pi2228 & ~n22860;
  assign n25251 = ~pi2228 & ~n22879;
  assign n25252 = n22879 & ~n23348;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = n22860 & ~n25253;
  assign po2404 = n25250 | n25254;
  assign n25256 = ~pi2229 & ~n22860;
  assign n25257 = ~pi2229 & ~n22879;
  assign n25258 = n22879 & ~n23461;
  assign n25259 = ~n25257 & ~n25258;
  assign n25260 = n22860 & ~n25259;
  assign po2405 = n25256 | n25260;
  assign n25262 = ~pi2230 & ~n22860;
  assign n25263 = ~pi2230 & ~n22900;
  assign n25264 = n22900 & ~n23664;
  assign n25265 = ~n25263 & ~n25264;
  assign n25266 = n22860 & ~n25265;
  assign po2406 = n25262 | n25266;
  assign n25268 = ~pi2231 & ~n22860;
  assign n25269 = ~pi2231 & ~n22879;
  assign n25270 = n22879 & ~n23448;
  assign n25271 = ~n25269 & ~n25270;
  assign n25272 = n22860 & ~n25271;
  assign po2407 = n25268 | n25272;
  assign n25274 = ~pi2232 & ~n22860;
  assign n25275 = ~pi2232 & ~n22900;
  assign n25276 = n22900 & ~n23511;
  assign n25277 = ~n25275 & ~n25276;
  assign n25278 = n22860 & ~n25277;
  assign po2408 = n25274 | n25278;
  assign n25280 = ~pi2233 & ~n22860;
  assign n25281 = ~pi2233 & ~n22900;
  assign n25282 = n22900 & ~n23461;
  assign n25283 = ~n25281 & ~n25282;
  assign n25284 = n22860 & ~n25283;
  assign po2409 = n25280 | n25284;
  assign n25286 = ~pi2234 & ~n22860;
  assign n25287 = ~pi2234 & ~n22900;
  assign n25288 = n22900 & ~n23381;
  assign n25289 = ~n25287 & ~n25288;
  assign n25290 = n22860 & ~n25289;
  assign po2410 = n25286 | n25290;
  assign n25292 = ~pi2235 & ~n22860;
  assign n25293 = ~pi2235 & ~n22900;
  assign n25294 = n22900 & ~n23395;
  assign n25295 = ~n25293 & ~n25294;
  assign n25296 = n22860 & ~n25295;
  assign po2411 = n25292 | n25296;
  assign n25298 = ~pi2236 & ~n22860;
  assign n25299 = ~pi2236 & ~n22900;
  assign n25300 = n22900 & ~n23645;
  assign n25301 = ~n25299 & ~n25300;
  assign n25302 = n22860 & ~n25301;
  assign po2412 = n25298 | n25302;
  assign n25304 = ~pi2237 & ~n22860;
  assign n25305 = ~pi2237 & ~n22900;
  assign n25306 = n22900 & ~n23518;
  assign n25307 = ~n25305 & ~n25306;
  assign n25308 = n22860 & ~n25307;
  assign po2413 = n25304 | n25308;
  assign n25310 = ~pi2238 & ~n22860;
  assign n25311 = ~pi2238 & ~n22900;
  assign n25312 = n22900 & ~n23428;
  assign n25313 = ~n25311 & ~n25312;
  assign n25314 = n22860 & ~n25313;
  assign po2414 = n25310 | n25314;
  assign n25316 = ~pi2239 & ~n22860;
  assign n25317 = ~pi2239 & ~n22900;
  assign n25318 = n22900 & ~n23368;
  assign n25319 = ~n25317 & ~n25318;
  assign n25320 = n22860 & ~n25319;
  assign po2415 = n25316 | n25320;
  assign n25322 = ~pi2240 & ~n22860;
  assign n25323 = ~pi2240 & ~n22900;
  assign n25324 = n22900 & ~n23320;
  assign n25325 = ~n25323 & ~n25324;
  assign n25326 = n22860 & ~n25325;
  assign po2416 = n25322 | n25326;
  assign n25328 = ~pi2241 & ~n22860;
  assign n25329 = n22931 & ~n23327;
  assign n25330 = ~pi2241 & ~n22931;
  assign n25331 = ~n25329 & ~n25330;
  assign n25332 = n22860 & ~n25331;
  assign po2417 = n25328 | n25332;
  assign n25334 = ~pi2242 & ~n22860;
  assign n25335 = n22945 & ~n23388;
  assign n25336 = ~pi2242 & ~n22945;
  assign n25337 = ~n25335 & ~n25336;
  assign n25338 = n22860 & ~n25337;
  assign po2418 = n25334 | n25338;
  assign n25340 = ~pi2243 & ~n22860;
  assign n25341 = n22945 & ~n23341;
  assign n25342 = ~pi2243 & ~n22945;
  assign n25343 = ~n25341 & ~n25342;
  assign n25344 = n22860 & ~n25343;
  assign po2419 = n25340 | n25344;
  assign n25346 = ~pi2244 & ~n22860;
  assign n25347 = n22924 & ~n23518;
  assign n25348 = ~pi2244 & ~n22924;
  assign n25349 = ~n25347 & ~n25348;
  assign n25350 = n22860 & ~n25349;
  assign po2420 = n25346 | n25350;
  assign n25352 = ~pi2245 & ~n22860;
  assign n25353 = n22973 & ~n23953;
  assign n25354 = ~pi2245 & ~n22973;
  assign n25355 = ~n25353 & ~n25354;
  assign n25356 = n22860 & ~n25355;
  assign po2421 = n25352 | n25356;
  assign n25358 = ~pi2246 & ~n22860;
  assign n25359 = n22959 & ~n23341;
  assign n25360 = ~pi2246 & ~n22959;
  assign n25361 = ~n25359 & ~n25360;
  assign n25362 = n22860 & ~n25361;
  assign po2422 = n25358 | n25362;
  assign n25364 = ~pi2247 & ~n22860;
  assign n25365 = n22973 & ~n23638;
  assign n25366 = ~pi2247 & ~n22973;
  assign n25367 = ~n25365 & ~n25366;
  assign n25368 = n22860 & ~n25367;
  assign po2423 = n25364 | n25368;
  assign n25370 = ~pi2248 & ~n22860;
  assign n25371 = n22945 & ~n24002;
  assign n25372 = ~pi2248 & ~n22945;
  assign n25373 = ~n25371 & ~n25372;
  assign n25374 = n22860 & ~n25373;
  assign po2424 = n25370 | n25374;
  assign n25376 = ~pi2249 & ~n22860;
  assign n25377 = n22931 & ~n24002;
  assign n25378 = ~pi2249 & ~n22931;
  assign n25379 = ~n25377 & ~n25378;
  assign n25380 = n22860 & ~n25379;
  assign po2425 = n25376 | n25380;
  assign n25382 = ~pi2250 & ~n22860;
  assign n25383 = n22959 & ~n24002;
  assign n25384 = ~pi2250 & ~n22959;
  assign n25385 = ~n25383 & ~n25384;
  assign n25386 = n22860 & ~n25385;
  assign po2426 = n25382 | n25386;
  assign n25388 = ~pi2251 & ~n22860;
  assign n25389 = n22959 & ~n23334;
  assign n25390 = ~pi2251 & ~n22959;
  assign n25391 = ~n25389 & ~n25390;
  assign n25392 = n22860 & ~n25391;
  assign po2427 = n25388 | n25392;
  assign n25394 = pi1701 & n22080;
  assign n25395 = pi2252 & ~n23726;
  assign n25396 = ~pi2252 & n23740;
  assign n25397 = pi2252 & ~n23740;
  assign n25398 = ~n25396 & ~n25397;
  assign n25399 = n23726 & ~n25398;
  assign n25400 = ~n25395 & ~n25399;
  assign n25401 = ~n22080 & ~n25400;
  assign po2428 = n25394 | n25401;
  assign n25403 = ~pi2253 & ~n22860;
  assign n25404 = n22945 & ~n23306;
  assign n25405 = ~pi2253 & ~n22945;
  assign n25406 = ~n25404 & ~n25405;
  assign n25407 = n22860 & ~n25406;
  assign po2429 = n25403 | n25407;
  assign n25409 = ~pi2254 & ~n22860;
  assign n25410 = n22945 & ~n23334;
  assign n25411 = ~pi2254 & ~n22945;
  assign n25412 = ~n25410 & ~n25411;
  assign n25413 = n22860 & ~n25412;
  assign po2430 = n25409 | n25413;
  assign n25415 = ~pi2255 & ~n22860;
  assign n25416 = n22952 & ~n23537;
  assign n25417 = ~pi2255 & ~n22952;
  assign n25418 = ~n25416 & ~n25417;
  assign n25419 = n22860 & ~n25418;
  assign po2431 = n25415 | n25419;
  assign n25421 = ~pi2256 & ~n22860;
  assign n25422 = n22952 & ~n23355;
  assign n25423 = ~pi2256 & ~n22952;
  assign n25424 = ~n25422 & ~n25423;
  assign n25425 = n22860 & ~n25424;
  assign po2432 = n25421 | n25425;
  assign n25427 = ~pi2257 & ~n22860;
  assign n25428 = n22952 & ~n23388;
  assign n25429 = ~pi2257 & ~n22952;
  assign n25430 = ~n25428 & ~n25429;
  assign n25431 = n22860 & ~n25430;
  assign po2433 = n25427 | n25431;
  assign n25433 = ~pi2258 & ~n22860;
  assign n25434 = n22952 & ~n23313;
  assign n25435 = ~pi2258 & ~n22952;
  assign n25436 = ~n25434 & ~n25435;
  assign n25437 = n22860 & ~n25436;
  assign po2434 = n25433 | n25437;
  assign n25439 = ~pi2259 & ~n22860;
  assign n25440 = n22952 & ~n23408;
  assign n25441 = ~pi2259 & ~n22952;
  assign n25442 = ~n25440 & ~n25441;
  assign n25443 = n22860 & ~n25442;
  assign po2435 = n25439 | n25443;
  assign n25445 = ~pi2260 & ~n22860;
  assign n25446 = n22952 & ~n23625;
  assign n25447 = ~pi2260 & ~n22952;
  assign n25448 = ~n25446 & ~n25447;
  assign n25449 = n22860 & ~n25448;
  assign po2436 = n25445 | n25449;
  assign n25451 = ~pi2261 & ~n22860;
  assign n25452 = n22952 & ~n23953;
  assign n25453 = ~pi2261 & ~n22952;
  assign n25454 = ~n25452 & ~n25453;
  assign n25455 = n22860 & ~n25454;
  assign po2437 = n25451 | n25455;
  assign n25457 = ~pi2262 & ~n22860;
  assign n25458 = n22952 & ~n23557;
  assign n25459 = ~pi2262 & ~n22952;
  assign n25460 = ~n25458 & ~n25459;
  assign n25461 = n22860 & ~n25460;
  assign po2438 = n25457 | n25461;
  assign n25463 = ~pi2263 & ~n22860;
  assign n25464 = n22952 & ~n23511;
  assign n25465 = ~pi2263 & ~n22952;
  assign n25466 = ~n25464 & ~n25465;
  assign n25467 = n22860 & ~n25466;
  assign po2439 = n25463 | n25467;
  assign n25469 = ~pi2264 & ~n22860;
  assign n25470 = n22952 & ~n23415;
  assign n25471 = ~pi2264 & ~n22952;
  assign n25472 = ~n25470 & ~n25471;
  assign n25473 = n22860 & ~n25472;
  assign po2440 = n25469 | n25473;
  assign n25475 = ~pi2265 & ~n22860;
  assign n25476 = n22952 & ~n23664;
  assign n25477 = ~pi2265 & ~n22952;
  assign n25478 = ~n25476 & ~n25477;
  assign n25479 = n22860 & ~n25478;
  assign po2441 = n25475 | n25479;
  assign n25481 = ~pi2266 & ~n22860;
  assign n25482 = n22952 & ~n23638;
  assign n25483 = ~pi2266 & ~n22952;
  assign n25484 = ~n25482 & ~n25483;
  assign n25485 = n22860 & ~n25484;
  assign po2442 = n25481 | n25485;
  assign n25487 = ~pi2267 & ~n22860;
  assign n25488 = n22959 & ~n23625;
  assign n25489 = ~pi2267 & ~n22959;
  assign n25490 = ~n25488 & ~n25489;
  assign n25491 = n22860 & ~n25490;
  assign po2443 = n25487 | n25491;
  assign n25493 = ~pi2268 & ~n22860;
  assign n25494 = n22959 & ~n23327;
  assign n25495 = ~pi2268 & ~n22959;
  assign n25496 = ~n25494 & ~n25495;
  assign n25497 = n22860 & ~n25496;
  assign po2444 = n25493 | n25497;
  assign n25499 = ~pi2269 & ~n22860;
  assign n25500 = n22952 & ~n23381;
  assign n25501 = ~pi2269 & ~n22952;
  assign n25502 = ~n25500 & ~n25501;
  assign n25503 = n22860 & ~n25502;
  assign po2445 = n25499 | n25503;
  assign n25505 = ~pi2270 & ~n22860;
  assign n25506 = n22924 & ~n23448;
  assign n25507 = ~pi2270 & ~n22924;
  assign n25508 = ~n25506 & ~n25507;
  assign n25509 = n22860 & ~n25508;
  assign po2446 = n25505 | n25509;
  assign n25511 = ~pi2271 & ~n22860;
  assign n25512 = n22924 & ~n23461;
  assign n25513 = ~pi2271 & ~n22924;
  assign n25514 = ~n25512 & ~n25513;
  assign n25515 = n22860 & ~n25514;
  assign po2447 = n25511 | n25515;
  assign n25517 = ~pi2272 & ~n22860;
  assign n25518 = n22924 & ~n23428;
  assign n25519 = ~pi2272 & ~n22924;
  assign n25520 = ~n25518 & ~n25519;
  assign n25521 = n22860 & ~n25520;
  assign po2448 = n25517 | n25521;
  assign n25523 = ~pi2273 & ~n22860;
  assign n25524 = n22931 & ~n23395;
  assign n25525 = ~pi2273 & ~n22931;
  assign n25526 = ~n25524 & ~n25525;
  assign n25527 = n22860 & ~n25526;
  assign po2449 = n25523 | n25527;
  assign n25529 = ~pi2274 & ~n22860;
  assign n25530 = n22917 & ~n23862;
  assign n25531 = ~pi2274 & ~n22917;
  assign n25532 = ~n25530 & ~n25531;
  assign n25533 = n22860 & ~n25532;
  assign po2450 = n25529 | n25533;
  assign n25535 = ~pi2275 & ~n22860;
  assign n25536 = n22959 & ~n23368;
  assign n25537 = ~pi2275 & ~n22959;
  assign n25538 = ~n25536 & ~n25537;
  assign n25539 = n22860 & ~n25538;
  assign po2451 = n25535 | n25539;
  assign n25541 = ~pi2276 & ~n22860;
  assign n25542 = n22931 & ~n23625;
  assign n25543 = ~pi2276 & ~n22931;
  assign n25544 = ~n25542 & ~n25543;
  assign n25545 = n22860 & ~n25544;
  assign po2452 = n25541 | n25545;
  assign n25547 = ~pi2277 & ~n22860;
  assign n25548 = n22959 & ~n23474;
  assign n25549 = ~pi2277 & ~n22959;
  assign n25550 = ~n25548 & ~n25549;
  assign n25551 = n22860 & ~n25550;
  assign po2453 = n25547 | n25551;
  assign n25553 = ~pi2278 & ~n22860;
  assign n25554 = ~pi2278 & ~n22893;
  assign n25555 = n22893 & ~n24002;
  assign n25556 = ~n25554 & ~n25555;
  assign n25557 = n22860 & ~n25556;
  assign po2454 = n25553 | n25557;
  assign n25559 = ~pi2279 & ~n22860;
  assign n25560 = n22945 & ~n23327;
  assign n25561 = ~pi2279 & ~n22945;
  assign n25562 = ~n25560 & ~n25561;
  assign n25563 = n22860 & ~n25562;
  assign po2455 = n25559 | n25563;
  assign n25565 = ~pi2280 & ~n22860;
  assign n25566 = n22952 & ~n23645;
  assign n25567 = ~pi2280 & ~n22952;
  assign n25568 = ~n25566 & ~n25567;
  assign n25569 = n22860 & ~n25568;
  assign po2456 = n25565 | n25569;
  assign n25571 = ~pi2281 & ~n22860;
  assign n25572 = n22952 & ~n23368;
  assign n25573 = ~pi2281 & ~n22952;
  assign n25574 = ~n25572 & ~n25573;
  assign n25575 = n22860 & ~n25574;
  assign po2457 = n25571 | n25575;
  assign n25577 = ~pi2282 & ~n22860;
  assign n25578 = n22952 & ~n23395;
  assign n25579 = ~pi2282 & ~n22952;
  assign n25580 = ~n25578 & ~n25579;
  assign n25581 = n22860 & ~n25580;
  assign po2458 = n25577 | n25581;
  assign n25583 = ~pi2283 & ~n22860;
  assign n25584 = ~pi2283 & ~n22938;
  assign n25585 = n22938 & ~n23313;
  assign n25586 = ~n25584 & ~n25585;
  assign n25587 = n22860 & ~n25586;
  assign po2459 = n25583 | n25587;
  assign n25589 = pi2988 & n22561;
  assign n25590 = ~pi2284 & ~n22561;
  assign n25591 = ~n25589 & ~n25590;
  assign n25592 = n22306 & ~n25591;
  assign n25593 = ~pi2284 & ~n22306;
  assign po2460 = n25592 | n25593;
  assign n25595 = pi2285 & ~n20262;
  assign n25596 = n19955 & n20262;
  assign po2461 = n25595 | n25596;
  assign n25598 = ~pi2286 & ~n22860;
  assign n25599 = ~pi2286 & ~n22938;
  assign n25600 = n22938 & ~n24002;
  assign n25601 = ~n25599 & ~n25600;
  assign n25602 = n22860 & ~n25601;
  assign po2462 = n25598 | n25602;
  assign n25604 = ~pi2287 & ~n22860;
  assign n25605 = n22917 & ~n23511;
  assign n25606 = ~pi2287 & ~n22917;
  assign n25607 = ~n25605 & ~n25606;
  assign n25608 = n22860 & ~n25607;
  assign po2463 = n25604 | n25608;
  assign n25610 = ~pi2288 & ~n22860;
  assign n25611 = n22973 & ~n23348;
  assign n25612 = ~pi2288 & ~n22973;
  assign n25613 = ~n25611 & ~n25612;
  assign n25614 = n22860 & ~n25613;
  assign po2464 = n25610 | n25614;
  assign n25616 = pi2987 & n22302;
  assign n25617 = ~pi2289 & ~n22302;
  assign n25618 = ~n25616 & ~n25617;
  assign n25619 = n22306 & ~n25618;
  assign n25620 = ~pi2289 & ~n22306;
  assign po2465 = n25619 | n25620;
  assign n25622 = ~pi2290 & ~n22860;
  assign n25623 = n22959 & ~n23395;
  assign n25624 = ~pi2290 & ~n22959;
  assign n25625 = ~n25623 & ~n25624;
  assign n25626 = n22860 & ~n25625;
  assign po2466 = n25622 | n25626;
  assign n25628 = ~pi2291 & ~n22860;
  assign n25629 = n22917 & ~n23570;
  assign n25630 = ~pi2291 & ~n22917;
  assign n25631 = ~n25629 & ~n25630;
  assign n25632 = n22860 & ~n25631;
  assign po2467 = n25628 | n25632;
  assign n25634 = pi2987 & n22311;
  assign n25635 = ~pi2292 & ~n22311;
  assign n25636 = ~n25634 & ~n25635;
  assign n25637 = n22306 & ~n25636;
  assign n25638 = ~pi2292 & ~n22306;
  assign po2468 = n25637 | n25638;
  assign n25640 = pi2988 & n22554;
  assign n25641 = ~pi2293 & ~n22554;
  assign n25642 = ~n25640 & ~n25641;
  assign n25643 = n22306 & ~n25642;
  assign n25644 = ~pi2293 & ~n22306;
  assign po2469 = n25643 | n25644;
  assign n25646 = pi1699 & n22080;
  assign n25647 = pi2294 & ~n23726;
  assign n25648 = ~pi2294 & n23726;
  assign n25649 = ~n25647 & ~n25648;
  assign n25650 = ~n22080 & ~n25649;
  assign po2470 = n25646 | n25650;
  assign n25652 = pi2988 & n22302;
  assign n25653 = ~pi2295 & ~n22302;
  assign n25654 = ~n25652 & ~n25653;
  assign n25655 = n22306 & ~n25654;
  assign n25656 = ~pi2295 & ~n22306;
  assign po2471 = n25655 | n25656;
  assign n25658 = ~pi2296 & ~n22860;
  assign n25659 = ~pi2296 & ~n22938;
  assign n25660 = n22938 & ~n23341;
  assign n25661 = ~n25659 & ~n25660;
  assign n25662 = n22860 & ~n25661;
  assign po2472 = n25658 | n25662;
  assign n25664 = ~pi2297 & ~n22860;
  assign n25665 = pi2975 & n22945;
  assign n25666 = ~pi2297 & ~n22945;
  assign n25667 = ~n25665 & ~n25666;
  assign n25668 = n22860 & ~n25667;
  assign po2473 = n25664 | n25668;
  assign n25670 = ~pi2298 & ~n22860;
  assign n25671 = n22945 & ~n23570;
  assign n25672 = ~pi2298 & ~n22945;
  assign n25673 = ~n25671 & ~n25672;
  assign n25674 = n22860 & ~n25673;
  assign po2474 = n25670 | n25674;
  assign n25676 = ~pi2299 & ~n22860;
  assign n25677 = n22917 & ~n23415;
  assign n25678 = ~pi2299 & ~n22917;
  assign n25679 = ~n25677 & ~n25678;
  assign n25680 = n22860 & ~n25679;
  assign po2475 = n25676 | n25680;
  assign n25682 = ~pi2300 & ~n22860;
  assign n25683 = n22973 & ~n23461;
  assign n25684 = ~pi2300 & ~n22973;
  assign n25685 = ~n25683 & ~n25684;
  assign n25686 = n22860 & ~n25685;
  assign po2476 = n25682 | n25686;
  assign n25688 = ~pi2301 & ~n22860;
  assign n25689 = n22973 & ~n23395;
  assign n25690 = ~pi2301 & ~n22973;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = n22860 & ~n25691;
  assign po2477 = n25688 | n25692;
  assign n25694 = ~pi2302 & ~n22860;
  assign n25695 = n22945 & ~n23408;
  assign n25696 = ~pi2302 & ~n22945;
  assign n25697 = ~n25695 & ~n25696;
  assign n25698 = n22860 & ~n25697;
  assign po2478 = n25694 | n25698;
  assign n25700 = ~pi2303 & ~n22860;
  assign n25701 = ~pi2303 & ~n22938;
  assign n25702 = n22938 & ~n23334;
  assign n25703 = ~n25701 & ~n25702;
  assign n25704 = n22860 & ~n25703;
  assign po2479 = n25700 | n25704;
  assign n25706 = ~pi2304 & ~n22860;
  assign n25707 = n22917 & ~n24002;
  assign n25708 = ~pi2304 & ~n22917;
  assign n25709 = ~n25707 & ~n25708;
  assign n25710 = n22860 & ~n25709;
  assign po2480 = n25706 | n25710;
  assign n25712 = ~pi2305 & ~n22860;
  assign n25713 = n22945 & ~n23862;
  assign n25714 = ~pi2305 & ~n22945;
  assign n25715 = ~n25713 & ~n25714;
  assign n25716 = n22860 & ~n25715;
  assign po2481 = n25712 | n25716;
  assign n25718 = ~pi2306 & ~n22860;
  assign n25719 = n22931 & ~n23550;
  assign n25720 = ~pi2306 & ~n22931;
  assign n25721 = ~n25719 & ~n25720;
  assign n25722 = n22860 & ~n25721;
  assign po2482 = n25718 | n25722;
  assign n25724 = ~pi2307 & ~n22860;
  assign n25725 = n22973 & ~n23645;
  assign n25726 = ~pi2307 & ~n22973;
  assign n25727 = ~n25725 & ~n25726;
  assign n25728 = n22860 & ~n25727;
  assign po2483 = n25724 | n25728;
  assign n25730 = ~pi2308 & ~n22860;
  assign n25731 = n22945 & ~n23625;
  assign n25732 = ~pi2308 & ~n22945;
  assign n25733 = ~n25731 & ~n25732;
  assign n25734 = n22860 & ~n25733;
  assign po2484 = n25730 | n25734;
  assign n25736 = ~pi2309 & ~n22860;
  assign n25737 = n22931 & ~n23570;
  assign n25738 = ~pi2309 & ~n22931;
  assign n25739 = ~n25737 & ~n25738;
  assign n25740 = n22860 & ~n25739;
  assign po2485 = n25736 | n25740;
  assign n25742 = ~pi2310 & ~n22860;
  assign n25743 = n22959 & ~n23570;
  assign n25744 = ~pi2310 & ~n22959;
  assign n25745 = ~n25743 & ~n25744;
  assign n25746 = n22860 & ~n25745;
  assign po2486 = n25742 | n25746;
  assign n25748 = ~pi2311 & ~n22860;
  assign n25749 = n22917 & ~n23334;
  assign n25750 = ~pi2311 & ~n22917;
  assign n25751 = ~n25749 & ~n25750;
  assign n25752 = n22860 & ~n25751;
  assign po2487 = n25748 | n25752;
  assign n25754 = ~pi2312 & ~n22860;
  assign n25755 = n22973 & ~n23355;
  assign n25756 = ~pi2312 & ~n22973;
  assign n25757 = ~n25755 & ~n25756;
  assign n25758 = n22860 & ~n25757;
  assign po2488 = n25754 | n25758;
  assign n25760 = ~pi2313 & ~n22860;
  assign n25761 = n22931 & ~n23953;
  assign n25762 = ~pi2313 & ~n22931;
  assign n25763 = ~n25761 & ~n25762;
  assign n25764 = n22860 & ~n25763;
  assign po2489 = n25760 | n25764;
  assign n25766 = ~pi2314 & ~n22860;
  assign n25767 = n22973 & ~n23368;
  assign n25768 = ~pi2314 & ~n22973;
  assign n25769 = ~n25767 & ~n25768;
  assign n25770 = n22860 & ~n25769;
  assign po2490 = n25766 | n25770;
  assign n25772 = ~pi2315 & ~n22860;
  assign n25773 = n22945 & ~n23474;
  assign n25774 = ~pi2315 & ~n22945;
  assign n25775 = ~n25773 & ~n25774;
  assign n25776 = n22860 & ~n25775;
  assign po2491 = n25772 | n25776;
  assign n25778 = ~pi2316 & ~n22860;
  assign n25779 = n22959 & ~n23638;
  assign n25780 = ~pi2316 & ~n22959;
  assign n25781 = ~n25779 & ~n25780;
  assign n25782 = n22860 & ~n25781;
  assign po2492 = n25778 | n25782;
  assign n25784 = ~pi2317 & ~n22860;
  assign n25785 = n22917 & ~n23550;
  assign n25786 = ~pi2317 & ~n22917;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = n22860 & ~n25787;
  assign po2493 = n25784 | n25788;
  assign n25790 = ~pi2318 & ~n22860;
  assign n25791 = ~pi2318 & ~n22938;
  assign n25792 = n22938 & ~n23388;
  assign n25793 = ~n25791 & ~n25792;
  assign n25794 = n22860 & ~n25793;
  assign po2494 = n25790 | n25794;
  assign n25796 = ~pi2319 & ~n22860;
  assign n25797 = n22959 & ~n23355;
  assign n25798 = ~pi2319 & ~n22959;
  assign n25799 = ~n25797 & ~n25798;
  assign n25800 = n22860 & ~n25799;
  assign po2495 = n25796 | n25800;
  assign n25802 = ~pi2320 & ~n22860;
  assign n25803 = n22973 & ~n23381;
  assign n25804 = ~pi2320 & ~n22973;
  assign n25805 = ~n25803 & ~n25804;
  assign n25806 = n22860 & ~n25805;
  assign po2496 = n25802 | n25806;
  assign n25808 = ~pi2321 & ~n22860;
  assign n25809 = n22931 & ~n23862;
  assign n25810 = ~pi2321 & ~n22931;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = n22860 & ~n25811;
  assign po2497 = n25808 | n25812;
  assign n25814 = ~pi2322 & ~n22860;
  assign n25815 = n22945 & ~n23537;
  assign n25816 = ~pi2322 & ~n22945;
  assign n25817 = ~n25815 & ~n25816;
  assign n25818 = n22860 & ~n25817;
  assign po2498 = n25814 | n25818;
  assign n25820 = ~pi2323 & ~n22860;
  assign n25821 = n22917 & ~n23327;
  assign n25822 = ~pi2323 & ~n22917;
  assign n25823 = ~n25821 & ~n25822;
  assign n25824 = n22860 & ~n25823;
  assign po2499 = n25820 | n25824;
  assign n25826 = ~pi2324 & ~n22860;
  assign n25827 = n22917 & ~n23481;
  assign n25828 = ~pi2324 & ~n22917;
  assign n25829 = ~n25827 & ~n25828;
  assign n25830 = n22860 & ~n25829;
  assign po2500 = n25826 | n25830;
  assign n25832 = ~pi2325 & ~n22860;
  assign n25833 = n22973 & ~n23320;
  assign n25834 = ~pi2325 & ~n22973;
  assign n25835 = ~n25833 & ~n25834;
  assign n25836 = n22860 & ~n25835;
  assign po2501 = n25832 | n25836;
  assign n25838 = ~pi2326 & ~n22860;
  assign n25839 = n22973 & ~n23518;
  assign n25840 = ~pi2326 & ~n22973;
  assign n25841 = ~n25839 & ~n25840;
  assign n25842 = n22860 & ~n25841;
  assign po2502 = n25838 | n25842;
  assign n25844 = ~pi2327 & ~n22860;
  assign n25845 = n22917 & ~n23474;
  assign n25846 = ~pi2327 & ~n22917;
  assign n25847 = ~n25845 & ~n25846;
  assign n25848 = n22860 & ~n25847;
  assign po2503 = n25844 | n25848;
  assign n25850 = ~pi2328 & ~n22860;
  assign n25851 = n22945 & ~n23550;
  assign n25852 = ~pi2328 & ~n22945;
  assign n25853 = ~n25851 & ~n25852;
  assign n25854 = n22860 & ~n25853;
  assign po2504 = n25850 | n25854;
  assign n25856 = ~pi2329 & ~n22860;
  assign n25857 = n22959 & ~n23953;
  assign n25858 = ~pi2329 & ~n22959;
  assign n25859 = ~n25857 & ~n25858;
  assign n25860 = n22860 & ~n25859;
  assign po2505 = n25856 | n25860;
  assign n25862 = ~pi2330 & ~n22860;
  assign n25863 = n22886 & ~n23481;
  assign n25864 = ~pi2330 & ~n22886;
  assign n25865 = ~n25863 & ~n25864;
  assign n25866 = n22860 & ~n25865;
  assign po2506 = n25862 | n25866;
  assign n25868 = ~pi2331 & ~n22860;
  assign n25869 = n22966 & ~n23334;
  assign n25870 = ~pi2331 & ~n22966;
  assign n25871 = ~n25869 & ~n25870;
  assign n25872 = n22860 & ~n25871;
  assign po2507 = n25868 | n25872;
  assign n25874 = ~pi2332 & ~n22860;
  assign n25875 = n22973 & ~n23306;
  assign n25876 = ~pi2332 & ~n22973;
  assign n25877 = ~n25875 & ~n25876;
  assign n25878 = n22860 & ~n25877;
  assign po2508 = n25874 | n25878;
  assign n25880 = ~pi2333 & ~n22860;
  assign n25881 = n22952 & ~n23448;
  assign n25882 = ~pi2333 & ~n22952;
  assign n25883 = ~n25881 & ~n25882;
  assign n25884 = n22860 & ~n25883;
  assign po2509 = n25880 | n25884;
  assign n25886 = ~pi2334 & ~n22860;
  assign n25887 = n22917 & ~n23461;
  assign n25888 = ~pi2334 & ~n22917;
  assign n25889 = ~n25887 & ~n25888;
  assign n25890 = n22860 & ~n25889;
  assign po2510 = n25886 | n25890;
  assign n25892 = ~pi2335 & ~n22860;
  assign n25893 = n22917 & ~n23953;
  assign n25894 = ~pi2335 & ~n22917;
  assign n25895 = ~n25893 & ~n25894;
  assign n25896 = n22860 & ~n25895;
  assign po2511 = n25892 | n25896;
  assign n25898 = ~pi2336 & ~n22860;
  assign n25899 = n22966 & ~n23625;
  assign n25900 = ~pi2336 & ~n22966;
  assign n25901 = ~n25899 & ~n25900;
  assign n25902 = n22860 & ~n25901;
  assign po2512 = n25898 | n25902;
  assign n25904 = ~pi2337 & ~n22860;
  assign n25905 = n22924 & ~n23557;
  assign n25906 = ~pi2337 & ~n22924;
  assign n25907 = ~n25905 & ~n25906;
  assign n25908 = n22860 & ~n25907;
  assign po2513 = n25904 | n25908;
  assign n25910 = ~pi2338 & ~n22860;
  assign n25911 = n22945 & ~n23395;
  assign n25912 = ~pi2338 & ~n22945;
  assign n25913 = ~n25911 & ~n25912;
  assign n25914 = n22860 & ~n25913;
  assign po2514 = n25910 | n25914;
  assign n25916 = ~pi2339 & ~n22860;
  assign n25917 = n22924 & ~n23537;
  assign n25918 = ~pi2339 & ~n22924;
  assign n25919 = ~n25917 & ~n25918;
  assign n25920 = n22860 & ~n25919;
  assign po2515 = n25916 | n25920;
  assign n25922 = ~pi2340 & ~n22860;
  assign n25923 = ~pi2340 & ~n22938;
  assign n25924 = n22938 & ~n23570;
  assign n25925 = ~n25923 & ~n25924;
  assign n25926 = n22860 & ~n25925;
  assign po2516 = n25922 | n25926;
  assign n25928 = ~pi2341 & ~n22860;
  assign n25929 = n22973 & ~n23570;
  assign n25930 = ~pi2341 & ~n22973;
  assign n25931 = ~n25929 & ~n25930;
  assign n25932 = n22860 & ~n25931;
  assign po2517 = n25928 | n25932;
  assign n25934 = ~pi2342 & ~n22860;
  assign n25935 = n22931 & ~n23348;
  assign n25936 = ~pi2342 & ~n22931;
  assign n25937 = ~n25935 & ~n25936;
  assign n25938 = n22860 & ~n25937;
  assign po2518 = n25934 | n25938;
  assign n25940 = ~pi2343 & ~n22860;
  assign n25941 = n22931 & ~n23341;
  assign n25942 = ~pi2343 & ~n22931;
  assign n25943 = ~n25941 & ~n25942;
  assign n25944 = n22860 & ~n25943;
  assign po2519 = n25940 | n25944;
  assign n25946 = ~pi2344 & ~n22860;
  assign n25947 = n22973 & ~n23550;
  assign n25948 = ~pi2344 & ~n22973;
  assign n25949 = ~n25947 & ~n25948;
  assign n25950 = n22860 & ~n25949;
  assign po2520 = n25946 | n25950;
  assign n25952 = ~pi2345 & ~n22860;
  assign n25953 = n22924 & ~n23645;
  assign n25954 = ~pi2345 & ~n22924;
  assign n25955 = ~n25953 & ~n25954;
  assign n25956 = n22860 & ~n25955;
  assign po2521 = n25952 | n25956;
  assign n25958 = ~pi2346 & ~n22860;
  assign n25959 = n22966 & ~n23306;
  assign n25960 = ~pi2346 & ~n22966;
  assign n25961 = ~n25959 & ~n25960;
  assign n25962 = n22860 & ~n25961;
  assign po2522 = n25958 | n25962;
  assign n25964 = ~pi2347 & ~n22860;
  assign n25965 = n22945 & ~n23953;
  assign n25966 = ~pi2347 & ~n22945;
  assign n25967 = ~n25965 & ~n25966;
  assign n25968 = n22860 & ~n25967;
  assign po2523 = n25964 | n25968;
  assign n25970 = ~pi2348 & ~n22860;
  assign n25971 = n22917 & ~n23664;
  assign n25972 = ~pi2348 & ~n22917;
  assign n25973 = ~n25971 & ~n25972;
  assign n25974 = n22860 & ~n25973;
  assign po2524 = n25970 | n25974;
  assign n25976 = ~pi2349 & ~n22860;
  assign n25977 = n22959 & ~n23320;
  assign n25978 = ~pi2349 & ~n22959;
  assign n25979 = ~n25977 & ~n25978;
  assign n25980 = n22860 & ~n25979;
  assign po2525 = n25976 | n25980;
  assign n25982 = ~pi2350 & ~n22860;
  assign n25983 = n22917 & ~n23638;
  assign n25984 = ~pi2350 & ~n22917;
  assign n25985 = ~n25983 & ~n25984;
  assign n25986 = n22860 & ~n25985;
  assign po2526 = n25982 | n25986;
  assign n25988 = ~pi2351 & ~n22860;
  assign n25989 = n22966 & ~n24002;
  assign n25990 = ~pi2351 & ~n22966;
  assign n25991 = ~n25989 & ~n25990;
  assign n25992 = n22860 & ~n25991;
  assign po2527 = n25988 | n25992;
  assign n25994 = ~pi2352 & ~n22860;
  assign n25995 = n22931 & ~n23320;
  assign n25996 = ~pi2352 & ~n22931;
  assign n25997 = ~n25995 & ~n25996;
  assign n25998 = n22860 & ~n25997;
  assign po2528 = n25994 | n25998;
  assign n26000 = ~pi2353 & ~n22860;
  assign n26001 = n22966 & ~n23327;
  assign n26002 = ~pi2353 & ~n22966;
  assign n26003 = ~n26001 & ~n26002;
  assign n26004 = n22860 & ~n26003;
  assign po2529 = n26000 | n26004;
  assign n26006 = ~pi2354 & ~n22860;
  assign n26007 = n22931 & ~n23461;
  assign n26008 = ~pi2354 & ~n22931;
  assign n26009 = ~n26007 & ~n26008;
  assign n26010 = n22860 & ~n26009;
  assign po2530 = n26006 | n26010;
  assign n26012 = ~pi2355 & ~n22860;
  assign n26013 = n22924 & ~n23395;
  assign n26014 = ~pi2355 & ~n22924;
  assign n26015 = ~n26013 & ~n26014;
  assign n26016 = n22860 & ~n26015;
  assign po2531 = n26012 | n26016;
  assign n26018 = ~pi2356 & ~n22860;
  assign n26019 = n22959 & ~n23461;
  assign n26020 = ~pi2356 & ~n22959;
  assign n26021 = ~n26019 & ~n26020;
  assign n26022 = n22860 & ~n26021;
  assign po2532 = n26018 | n26022;
  assign n26024 = ~pi2357 & ~n22860;
  assign n26025 = n22966 & ~n23313;
  assign n26026 = ~pi2357 & ~n22966;
  assign n26027 = ~n26025 & ~n26026;
  assign n26028 = n22860 & ~n26027;
  assign po2533 = n26024 | n26028;
  assign n26030 = ~pi2358 & ~n22860;
  assign n26031 = ~pi1983 & pi1985;
  assign n26032 = pi1983 & ~pi1985;
  assign n26033 = ~n26031 & ~n26032;
  assign n26034 = n22860 & ~n26033;
  assign po2534 = n26030 | n26034;
  assign n26036 = ~pi2359 & ~n22860;
  assign n26037 = n22917 & ~n23645;
  assign n26038 = ~pi2359 & ~n22917;
  assign n26039 = ~n26037 & ~n26038;
  assign n26040 = n22860 & ~n26039;
  assign po2535 = n26036 | n26040;
  assign n26042 = ~pi2360 & ~n22860;
  assign n26043 = n22966 & ~n23408;
  assign n26044 = ~pi2360 & ~n22966;
  assign n26045 = ~n26043 & ~n26044;
  assign n26046 = n22860 & ~n26045;
  assign po2536 = n26042 | n26046;
  assign n26048 = ~pi2361 & ~n22860;
  assign n26049 = n22924 & ~n23306;
  assign n26050 = ~pi2361 & ~n22924;
  assign n26051 = ~n26049 & ~n26050;
  assign n26052 = n22860 & ~n26051;
  assign po2537 = n26048 | n26052;
  assign n26054 = ~pi2362 & ~n22860;
  assign n26055 = n22966 & ~n23557;
  assign n26056 = ~pi2362 & ~n22966;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = n22860 & ~n26057;
  assign po2538 = n26054 | n26058;
  assign n26060 = ~pi2363 & ~n22860;
  assign n26061 = n22973 & ~n23334;
  assign n26062 = ~pi2363 & ~n22973;
  assign n26063 = ~n26061 & ~n26062;
  assign n26064 = n22860 & ~n26063;
  assign po2539 = n26060 | n26064;
  assign n26066 = ~pi2364 & ~n22860;
  assign n26067 = ~pi2364 & ~n22938;
  assign n26068 = n22938 & ~n23408;
  assign n26069 = ~n26067 & ~n26068;
  assign n26070 = n22860 & ~n26069;
  assign po2540 = n26066 | n26070;
  assign n26072 = ~pi2365 & ~n22860;
  assign n26073 = n22945 & ~n23320;
  assign n26074 = ~pi2365 & ~n22945;
  assign n26075 = ~n26073 & ~n26074;
  assign n26076 = n22860 & ~n26075;
  assign po2541 = n26072 | n26076;
  assign n26078 = ~pi2366 & ~n22860;
  assign n26079 = n22917 & ~n23355;
  assign n26080 = ~pi2366 & ~n22917;
  assign n26081 = ~n26079 & ~n26080;
  assign n26082 = n22860 & ~n26081;
  assign po2542 = n26078 | n26082;
  assign n26084 = ~pi2367 & ~n22860;
  assign n26085 = n22924 & ~n23388;
  assign n26086 = ~pi2367 & ~n22924;
  assign n26087 = ~n26085 & ~n26086;
  assign n26088 = n22860 & ~n26087;
  assign po2543 = n26084 | n26088;
  assign n26090 = ~pi2368 & ~n22860;
  assign n26091 = n22945 & ~n23368;
  assign n26092 = ~pi2368 & ~n22945;
  assign n26093 = ~n26091 & ~n26092;
  assign n26094 = n22860 & ~n26093;
  assign po2544 = n26090 | n26094;
  assign n26096 = ~pi2369 & ~n22860;
  assign n26097 = n22924 & ~n23313;
  assign n26098 = ~pi2369 & ~n22924;
  assign n26099 = ~n26097 & ~n26098;
  assign n26100 = n22860 & ~n26099;
  assign po2545 = n26096 | n26100;
  assign n26102 = ~pi2370 & ~n22860;
  assign n26103 = n22973 & ~n23388;
  assign n26104 = ~pi2370 & ~n22973;
  assign n26105 = ~n26103 & ~n26104;
  assign n26106 = n22860 & ~n26105;
  assign po2546 = n26102 | n26106;
  assign n26108 = ~pi2371 & ~n22860;
  assign n26109 = n22917 & ~n23395;
  assign n26110 = ~pi2371 & ~n22917;
  assign n26111 = ~n26109 & ~n26110;
  assign n26112 = n22860 & ~n26111;
  assign po2547 = n26108 | n26112;
  assign n26114 = ~pi2372 & ~n22860;
  assign n26115 = n22924 & ~n23481;
  assign n26116 = ~pi2372 & ~n22924;
  assign n26117 = ~n26115 & ~n26116;
  assign n26118 = n22860 & ~n26117;
  assign po2548 = n26114 | n26118;
  assign n26120 = ~pi2373 & ~n22860;
  assign n26121 = n22966 & ~n23537;
  assign n26122 = ~pi2373 & ~n22966;
  assign n26123 = ~n26121 & ~n26122;
  assign n26124 = n22860 & ~n26123;
  assign po2549 = n26120 | n26124;
  assign n26126 = ~pi2374 & ~n22860;
  assign n26127 = ~pi2374 & ~n22938;
  assign n26128 = n22938 & ~n23625;
  assign n26129 = ~n26127 & ~n26128;
  assign n26130 = n22860 & ~n26129;
  assign po2550 = n26126 | n26130;
  assign n26132 = ~pi2375 & ~n22860;
  assign n26133 = n22945 & ~n23461;
  assign n26134 = ~pi2375 & ~n22945;
  assign n26135 = ~n26133 & ~n26134;
  assign n26136 = n22860 & ~n26135;
  assign po2551 = n26132 | n26136;
  assign n26138 = ~pi2376 & ~n22860;
  assign n26139 = n22973 & ~n23341;
  assign n26140 = ~pi2376 & ~n22973;
  assign n26141 = ~n26139 & ~n26140;
  assign n26142 = n22860 & ~n26141;
  assign po2552 = n26138 | n26142;
  assign n26144 = ~pi2377 & ~n22860;
  assign n26145 = n22924 & ~n23625;
  assign n26146 = ~pi2377 & ~n22924;
  assign n26147 = ~n26145 & ~n26146;
  assign n26148 = n22860 & ~n26147;
  assign po2553 = n26144 | n26148;
  assign n26150 = ~pi2378 & ~n22860;
  assign n26151 = n22966 & ~n23415;
  assign n26152 = ~pi2378 & ~n22966;
  assign n26153 = ~n26151 & ~n26152;
  assign n26154 = n22860 & ~n26153;
  assign po2554 = n26150 | n26154;
  assign n26156 = ~pi2379 & ~n22860;
  assign n26157 = n22917 & ~n23368;
  assign n26158 = ~pi2379 & ~n22917;
  assign n26159 = ~n26157 & ~n26158;
  assign n26160 = n22860 & ~n26159;
  assign po2555 = n26156 | n26160;
  assign n26162 = ~pi2380 & ~n22860;
  assign n26163 = n22966 & ~n23511;
  assign n26164 = ~pi2380 & ~n22966;
  assign n26165 = ~n26163 & ~n26164;
  assign n26166 = n22860 & ~n26165;
  assign po2556 = n26162 | n26166;
  assign n26168 = ~pi2381 & ~n22860;
  assign n26169 = n22945 & ~n23348;
  assign n26170 = ~pi2381 & ~n22945;
  assign n26171 = ~n26169 & ~n26170;
  assign n26172 = n22860 & ~n26171;
  assign po2557 = n26168 | n26172;
  assign n26174 = ~pi2382 & ~n22860;
  assign n26175 = n22973 & ~n23474;
  assign n26176 = ~pi2382 & ~n22973;
  assign n26177 = ~n26175 & ~n26176;
  assign n26178 = n22860 & ~n26177;
  assign po2558 = n26174 | n26178;
  assign n26180 = ~pi2383 & ~n22860;
  assign n26181 = ~pi2383 & ~n22893;
  assign n26182 = n22893 & ~n23625;
  assign n26183 = ~n26181 & ~n26182;
  assign n26184 = n22860 & ~n26183;
  assign po2559 = n26180 | n26184;
  assign n26186 = ~pi2384 & ~n22860;
  assign n26187 = ~n19071 & ~n22865;
  assign n26188 = n22860 & ~n26187;
  assign po2560 = n26186 | n26188;
  assign n26190 = ~pi2385 & ~n22860;
  assign n26191 = n22973 & ~n24002;
  assign n26192 = ~pi2385 & ~n22973;
  assign n26193 = ~n26191 & ~n26192;
  assign n26194 = n22860 & ~n26193;
  assign po2561 = n26190 | n26194;
  assign n26196 = ~pi2386 & ~n22860;
  assign n26197 = n22973 & ~n23327;
  assign n26198 = ~pi2386 & ~n22973;
  assign n26199 = ~n26197 & ~n26198;
  assign n26200 = n22860 & ~n26199;
  assign po2562 = n26196 | n26200;
  assign n26202 = ~pi2387 & ~n22860;
  assign n26203 = n22966 & ~n23381;
  assign n26204 = ~pi2387 & ~n22966;
  assign n26205 = ~n26203 & ~n26204;
  assign n26206 = n22860 & ~n26205;
  assign po2563 = n26202 | n26206;
  assign n26208 = ~pi2388 & ~n22860;
  assign n26209 = n22909 & ~n23388;
  assign n26210 = ~pi2388 & ~n22909;
  assign n26211 = ~n26209 & ~n26210;
  assign n26212 = n22860 & ~n26211;
  assign po2564 = n26208 | n26212;
  assign n26214 = ~pi2389 & ~n22860;
  assign n26215 = n22966 & ~n23448;
  assign n26216 = ~pi2389 & ~n22966;
  assign n26217 = ~n26215 & ~n26216;
  assign n26218 = n22860 & ~n26217;
  assign po2565 = n26214 | n26218;
  assign n26220 = ~pi2390 & ~n22860;
  assign n26221 = n22924 & ~n23415;
  assign n26222 = ~pi2390 & ~n22924;
  assign n26223 = ~n26221 & ~n26222;
  assign n26224 = n22860 & ~n26223;
  assign po2566 = n26220 | n26224;
  assign n26226 = ~pi2391 & ~n22860;
  assign n26227 = n22973 & ~n23481;
  assign n26228 = ~pi2391 & ~n22973;
  assign n26229 = ~n26227 & ~n26228;
  assign n26230 = n22860 & ~n26229;
  assign po2567 = n26226 | n26230;
  assign n26232 = ~pi2392 & ~n22860;
  assign n26233 = n22917 & ~n23348;
  assign n26234 = ~pi2392 & ~n22917;
  assign n26235 = ~n26233 & ~n26234;
  assign n26236 = n22860 & ~n26235;
  assign po2568 = n26232 | n26236;
  assign n26238 = ~pi2393 & ~n22860;
  assign n26239 = ~pi2393 & ~n22893;
  assign n26240 = pi2975 & n22893;
  assign n26241 = ~n26239 & ~n26240;
  assign n26242 = n22860 & ~n26241;
  assign po2569 = n26238 | n26242;
  assign n26244 = ~pi2394 & ~n22860;
  assign n26245 = ~pi2394 & ~n22938;
  assign n26246 = n22938 & ~n23537;
  assign n26247 = ~n26245 & ~n26246;
  assign n26248 = n22860 & ~n26247;
  assign po2570 = n26244 | n26248;
  assign n26250 = ~pi2395 & ~n22860;
  assign n26251 = n22973 & ~n23625;
  assign n26252 = ~pi2395 & ~n22973;
  assign n26253 = ~n26251 & ~n26252;
  assign n26254 = n22860 & ~n26253;
  assign po2571 = n26250 | n26254;
  assign n26256 = ~pi2396 & ~n22860;
  assign n26257 = n22909 & ~n23313;
  assign n26258 = ~pi2396 & ~n22909;
  assign n26259 = ~n26257 & ~n26258;
  assign n26260 = n22860 & ~n26259;
  assign po2572 = n26256 | n26260;
  assign n26262 = ~pi2397 & ~n22860;
  assign n26263 = ~pi2397 & ~n22980;
  assign n26264 = n22980 & ~n23953;
  assign n26265 = ~n26263 & ~n26264;
  assign n26266 = n22860 & ~n26265;
  assign po2573 = n26262 | n26266;
  assign n26268 = ~pi2398 & ~n22860;
  assign n26269 = ~pi2398 & ~n22938;
  assign n26270 = n22938 & ~n23550;
  assign n26271 = ~n26269 & ~n26270;
  assign n26272 = n22860 & ~n26271;
  assign po2574 = n26268 | n26272;
  assign n26274 = ~pi2399 & ~n22860;
  assign n26275 = ~pi2399 & ~n22893;
  assign n26276 = n22893 & ~n23415;
  assign n26277 = ~n26275 & ~n26276;
  assign n26278 = n22860 & ~n26277;
  assign po2575 = n26274 | n26278;
  assign n26280 = ~pi2400 & ~n22860;
  assign n26281 = n22924 & ~n23664;
  assign n26282 = ~pi2400 & ~n22924;
  assign n26283 = ~n26281 & ~n26282;
  assign n26284 = n22860 & ~n26283;
  assign po2576 = n26280 | n26284;
  assign n26286 = ~pi2401 & ~n22860;
  assign n26287 = ~pi2401 & ~n22893;
  assign n26288 = n22893 & ~n23327;
  assign n26289 = ~n26287 & ~n26288;
  assign n26290 = n22860 & ~n26289;
  assign po2577 = n26286 | n26290;
  assign n26292 = ~pi2402 & ~n22860;
  assign n26293 = n22909 & ~n23537;
  assign n26294 = ~pi2402 & ~n22909;
  assign n26295 = ~n26293 & ~n26294;
  assign n26296 = n22860 & ~n26295;
  assign po2578 = n26292 | n26296;
  assign n26298 = ~pi2403 & ~n22860;
  assign n26299 = n22966 & ~n23428;
  assign n26300 = ~pi2403 & ~n22966;
  assign n26301 = ~n26299 & ~n26300;
  assign n26302 = n22860 & ~n26301;
  assign po2579 = n26298 | n26302;
  assign n26304 = ~pi2406 & ~n22860;
  assign n26305 = ~pi2406 & ~n22938;
  assign n26306 = n22938 & ~n23474;
  assign n26307 = ~n26305 & ~n26306;
  assign n26308 = n22860 & ~n26307;
  assign po2580 = n26304 | n26308;
  assign n26310 = ~pi2407 & ~n22860;
  assign n26311 = n22909 & ~n23481;
  assign n26312 = ~pi2407 & ~n22909;
  assign n26313 = ~n26311 & ~n26312;
  assign n26314 = n22860 & ~n26313;
  assign po2581 = n26310 | n26314;
  assign n26316 = ~pi2408 & ~n22860;
  assign n26317 = n22909 & ~n23408;
  assign n26318 = ~pi2408 & ~n22909;
  assign n26319 = ~n26317 & ~n26318;
  assign n26320 = n22860 & ~n26319;
  assign po2582 = n26316 | n26320;
  assign n26322 = ~pi2409 & ~n22860;
  assign n26323 = n22886 & ~n23408;
  assign n26324 = ~pi2409 & ~n22886;
  assign n26325 = ~n26323 & ~n26324;
  assign n26326 = n22860 & ~n26325;
  assign po2583 = n26322 | n26326;
  assign n26328 = ~pi2410 & ~n22860;
  assign n26329 = ~pi2410 & ~n22893;
  assign n26330 = n22893 & ~n23408;
  assign n26331 = ~n26329 & ~n26330;
  assign n26332 = n22860 & ~n26331;
  assign po2584 = n26328 | n26332;
  assign n26334 = ~pi2411 & ~n22860;
  assign n26335 = n22886 & ~n23625;
  assign n26336 = ~pi2411 & ~n22886;
  assign n26337 = ~n26335 & ~n26336;
  assign n26338 = n22860 & ~n26337;
  assign po2585 = n26334 | n26338;
  assign n26340 = ~pi2412 & ~n22860;
  assign n26341 = n22909 & ~n23664;
  assign n26342 = ~pi2412 & ~n22909;
  assign n26343 = ~n26341 & ~n26342;
  assign n26344 = n22860 & ~n26343;
  assign po2586 = n26340 | n26344;
  assign n26346 = ~pi2413 & ~n22860;
  assign n26347 = ~pi2413 & ~n22980;
  assign n26348 = n22980 & ~n23474;
  assign n26349 = ~n26347 & ~n26348;
  assign n26350 = n22860 & ~n26349;
  assign po2587 = n26346 | n26350;
  assign n26352 = ~pi2414 & ~n22860;
  assign n26353 = ~pi2414 & ~n22938;
  assign n26354 = n22938 & ~n23953;
  assign n26355 = ~n26353 & ~n26354;
  assign n26356 = n22860 & ~n26355;
  assign po2588 = n26352 | n26356;
  assign n26358 = ~pi2415 & ~n22860;
  assign n26359 = ~pi2415 & ~n22938;
  assign n26360 = n22938 & ~n23415;
  assign n26361 = ~n26359 & ~n26360;
  assign n26362 = n22860 & ~n26361;
  assign po2589 = n26358 | n26362;
  assign n26364 = ~pi2416 & ~n22860;
  assign n26365 = n22909 & ~n23511;
  assign n26366 = ~pi2416 & ~n22909;
  assign n26367 = ~n26365 & ~n26366;
  assign n26368 = n22860 & ~n26367;
  assign po2590 = n26364 | n26368;
  assign n26370 = ~pi2417 & ~n22860;
  assign n26371 = ~pi2417 & ~n22938;
  assign n26372 = n22938 & ~n23428;
  assign n26373 = ~n26371 & ~n26372;
  assign n26374 = n22860 & ~n26373;
  assign po2591 = n26370 | n26374;
  assign n26376 = ~pi2418 & ~n22860;
  assign n26377 = ~pi2418 & ~n22938;
  assign n26378 = n22938 & ~n23862;
  assign n26379 = ~n26377 & ~n26378;
  assign n26380 = n22860 & ~n26379;
  assign po2592 = n26376 | n26380;
  assign n26382 = ~pi2419 & ~n22860;
  assign n26383 = n22909 & ~n23428;
  assign n26384 = ~pi2419 & ~n22909;
  assign n26385 = ~n26383 & ~n26384;
  assign n26386 = n22860 & ~n26385;
  assign po2593 = n26382 | n26386;
  assign n26388 = ~pi2420 & ~n22860;
  assign n26389 = n22909 & ~n23557;
  assign n26390 = ~pi2420 & ~n22909;
  assign n26391 = ~n26389 & ~n26390;
  assign n26392 = n22860 & ~n26391;
  assign po2594 = n26388 | n26392;
  assign n26394 = ~pi2421 & ~n22860;
  assign n26395 = ~pi2421 & ~n22938;
  assign n26396 = n22938 & ~n23664;
  assign n26397 = ~n26395 & ~n26396;
  assign n26398 = n22860 & ~n26397;
  assign po2595 = n26394 | n26398;
  assign n26400 = ~pi2422 & ~n22860;
  assign n26401 = ~pi2422 & ~n22938;
  assign n26402 = n22938 & ~n23638;
  assign n26403 = ~n26401 & ~n26402;
  assign n26404 = n22860 & ~n26403;
  assign po2596 = n26400 | n26404;
  assign n26406 = ~pi2423 & ~n22860;
  assign n26407 = n22909 & ~n23518;
  assign n26408 = ~pi2423 & ~n22909;
  assign n26409 = ~n26407 & ~n26408;
  assign n26410 = n22860 & ~n26409;
  assign po2597 = n26406 | n26410;
  assign n26412 = ~pi2424 & ~n22860;
  assign n26413 = n22909 & ~n23381;
  assign n26414 = ~pi2424 & ~n22909;
  assign n26415 = ~n26413 & ~n26414;
  assign n26416 = n22860 & ~n26415;
  assign po2598 = n26412 | n26416;
  assign n26418 = ~pi2425 & ~n22860;
  assign n26419 = ~pi2425 & ~n22879;
  assign n26420 = n22879 & ~n23570;
  assign n26421 = ~n26419 & ~n26420;
  assign n26422 = n22860 & ~n26421;
  assign po2599 = n26418 | n26422;
  assign n26424 = ~pi2426 & ~n22860;
  assign n26425 = n22909 & ~n23448;
  assign n26426 = ~pi2426 & ~n22909;
  assign n26427 = ~n26425 & ~n26426;
  assign n26428 = n22860 & ~n26427;
  assign po2600 = n26424 | n26428;
  assign n26430 = ~pi2427 & ~n22860;
  assign n26431 = ~pi2427 & ~n22938;
  assign n26432 = n22938 & ~n23320;
  assign n26433 = ~n26431 & ~n26432;
  assign n26434 = n22860 & ~n26433;
  assign po2601 = n26430 | n26434;
  assign n26436 = ~pi2428 & ~n22860;
  assign n26437 = ~pi2428 & ~n22938;
  assign n26438 = n22938 & ~n23355;
  assign n26439 = ~n26437 & ~n26438;
  assign n26440 = n22860 & ~n26439;
  assign po2602 = n26436 | n26440;
  assign n26442 = ~pi2429 & ~n22860;
  assign n26443 = n22886 & ~n23388;
  assign n26444 = ~pi2429 & ~n22886;
  assign n26445 = ~n26443 & ~n26444;
  assign n26446 = n22860 & ~n26445;
  assign po2603 = n26442 | n26446;
  assign n26448 = ~pi2430 & ~n22860;
  assign n26449 = ~pi2430 & ~n22938;
  assign n26450 = n22938 & ~n23395;
  assign n26451 = ~n26449 & ~n26450;
  assign n26452 = n22860 & ~n26451;
  assign po2604 = n26448 | n26452;
  assign n26454 = ~pi2431 & ~n22860;
  assign n26455 = n22886 & ~n23313;
  assign n26456 = ~pi2431 & ~n22886;
  assign n26457 = ~n26455 & ~n26456;
  assign n26458 = n22860 & ~n26457;
  assign po2605 = n26454 | n26458;
  assign n26460 = ~pi2432 & ~n22539;
  assign n26461 = pi2988 & n22539;
  assign n26462 = ~n26460 & ~n26461;
  assign n26463 = n22306 & ~n26462;
  assign n26464 = ~pi2432 & ~n22306;
  assign po2606 = n26463 | n26464;
  assign n26466 = ~pi2433 & ~n22860;
  assign n26467 = n22886 & ~n23306;
  assign n26468 = ~pi2433 & ~n22886;
  assign n26469 = ~n26467 & ~n26468;
  assign n26470 = n22860 & ~n26469;
  assign po2607 = n26466 | n26470;
  assign n26472 = ~pi2434 & ~n22326;
  assign n26473 = pi2988 & n22326;
  assign n26474 = ~n26472 & ~n26473;
  assign n26475 = n22306 & ~n26474;
  assign n26476 = ~pi2434 & ~n22306;
  assign po2608 = n26475 | n26476;
  assign n26478 = ~pi2435 & ~n22860;
  assign n26479 = ~pi2435 & ~n22938;
  assign n26480 = n22938 & ~n23368;
  assign n26481 = ~n26479 & ~n26480;
  assign n26482 = n22860 & ~n26481;
  assign po2609 = n26478 | n26482;
  assign n26484 = ~pi2436 & ~n22318;
  assign n26485 = pi2988 & n22318;
  assign n26486 = ~n26484 & ~n26485;
  assign n26487 = n22306 & ~n26486;
  assign n26488 = ~pi2436 & ~n22306;
  assign po2610 = n26487 | n26488;
  assign n26490 = ~pi2437 & ~n22860;
  assign n26491 = ~pi2437 & ~n22938;
  assign n26492 = n22938 & ~n23381;
  assign n26493 = ~n26491 & ~n26492;
  assign n26494 = n22860 & ~n26493;
  assign po2611 = n26490 | n26494;
  assign n26496 = ~pi2438 & ~n22860;
  assign n26497 = ~pi2438 & ~n22980;
  assign n26498 = n22980 & ~n23341;
  assign n26499 = ~n26497 & ~n26498;
  assign n26500 = n22860 & ~n26499;
  assign po2612 = n26496 | n26500;
  assign n26502 = ~pi2439 & ~n22860;
  assign n26503 = ~pi2439 & ~n22938;
  assign n26504 = n22938 & ~n23461;
  assign n26505 = ~n26503 & ~n26504;
  assign n26506 = n22860 & ~n26505;
  assign po2613 = n26502 | n26506;
  assign n26508 = ~pi2440 & ~n22860;
  assign n26509 = ~pi2440 & ~n22938;
  assign n26510 = n22938 & ~n23348;
  assign n26511 = ~n26509 & ~n26510;
  assign n26512 = n22860 & ~n26511;
  assign po2614 = n26508 | n26512;
  assign n26514 = ~pi2441 & ~n22860;
  assign n26515 = pi2975 & n22917;
  assign n26516 = ~pi2441 & ~n22917;
  assign n26517 = ~n26515 & ~n26516;
  assign n26518 = n22860 & ~n26517;
  assign po2615 = n26514 | n26518;
  assign n26520 = ~pi2442 & ~n22860;
  assign n26521 = ~pi2442 & ~n22980;
  assign n26522 = n22980 & ~n23625;
  assign n26523 = ~n26521 & ~n26522;
  assign n26524 = n22860 & ~n26523;
  assign po2616 = n26520 | n26524;
  assign n26526 = ~pi2443 & ~n22860;
  assign n26527 = ~pi2443 & ~n22980;
  assign n26528 = n22980 & ~n23306;
  assign n26529 = ~n26527 & ~n26528;
  assign n26530 = n22860 & ~n26529;
  assign po2617 = n26526 | n26530;
  assign n26532 = ~pi2444 & ~n22860;
  assign n26533 = ~pi2444 & ~n22980;
  assign n26534 = n22980 & ~n23334;
  assign n26535 = ~n26533 & ~n26534;
  assign n26536 = n22860 & ~n26535;
  assign po2618 = n26532 | n26536;
  assign n26538 = ~pi2445 & ~n22860;
  assign n26539 = ~pi2445 & ~n22893;
  assign n26540 = n22893 & ~n23550;
  assign n26541 = ~n26539 & ~n26540;
  assign n26542 = n22860 & ~n26541;
  assign po2619 = n26538 | n26542;
  assign n26544 = ~pi2446 & ~n22860;
  assign n26545 = ~pi2446 & ~n22893;
  assign n26546 = n22893 & ~n23570;
  assign n26547 = ~n26545 & ~n26546;
  assign n26548 = n22860 & ~n26547;
  assign po2620 = n26544 | n26548;
  assign n26550 = ~pi2447 & ~n22860;
  assign n26551 = ~pi2447 & ~n22980;
  assign n26552 = n22980 & ~n23388;
  assign n26553 = ~n26551 & ~n26552;
  assign n26554 = n22860 & ~n26553;
  assign po2621 = n26550 | n26554;
  assign n26556 = ~pi2448 & ~n22860;
  assign n26557 = ~pi2448 & ~n22980;
  assign n26558 = n22980 & ~n24002;
  assign n26559 = ~n26557 & ~n26558;
  assign n26560 = n22860 & ~n26559;
  assign po2622 = n26556 | n26560;
  assign n26562 = ~pi2449 & ~n22860;
  assign n26563 = ~pi2449 & ~n22980;
  assign n26564 = n22980 & ~n23327;
  assign n26565 = ~n26563 & ~n26564;
  assign n26566 = n22860 & ~n26565;
  assign po2623 = n26562 | n26566;
  assign n26568 = ~pi2450 & ~n22860;
  assign n26569 = ~pi2450 & ~n22893;
  assign n26570 = n22893 & ~n23474;
  assign n26571 = ~n26569 & ~n26570;
  assign n26572 = n22860 & ~n26571;
  assign po2624 = n26568 | n26572;
  assign n26574 = ~pi2451 & ~n22860;
  assign n26575 = ~pi2451 & ~n22980;
  assign n26576 = n22980 & ~n23313;
  assign n26577 = ~n26575 & ~n26576;
  assign n26578 = n22860 & ~n26577;
  assign po2625 = n26574 | n26578;
  assign n26580 = ~pi2452 & ~n22860;
  assign n26581 = ~pi2452 & ~n22980;
  assign n26582 = n22980 & ~n23550;
  assign n26583 = ~n26581 & ~n26582;
  assign n26584 = n22860 & ~n26583;
  assign po2626 = n26580 | n26584;
  assign n26586 = ~pi2453 & ~n22860;
  assign n26587 = ~pi2453 & ~n22893;
  assign n26588 = n22893 & ~n23638;
  assign n26589 = ~n26587 & ~n26588;
  assign n26590 = n22860 & ~n26589;
  assign po2627 = n26586 | n26590;
  assign n26592 = ~pi2454 & ~n22860;
  assign n26593 = ~pi2454 & ~n22980;
  assign n26594 = n22980 & ~n23570;
  assign n26595 = ~n26593 & ~n26594;
  assign n26596 = n22860 & ~n26595;
  assign po2628 = n26592 | n26596;
  assign n26598 = ~pi2455 & ~n22860;
  assign n26599 = ~pi2455 & ~n22893;
  assign n26600 = n22893 & ~n23461;
  assign n26601 = ~n26599 & ~n26600;
  assign n26602 = n22860 & ~n26601;
  assign po2629 = n26598 | n26602;
  assign n26604 = ~pi2456 & ~n22860;
  assign n26605 = ~pi2456 & ~n22893;
  assign n26606 = n22893 & ~n23862;
  assign n26607 = ~n26605 & ~n26606;
  assign n26608 = n22860 & ~n26607;
  assign po2630 = n26604 | n26608;
  assign n26610 = ~pi2457 & ~n22860;
  assign n26611 = ~pi2457 & ~n22980;
  assign n26612 = n22980 & ~n23664;
  assign n26613 = ~n26611 & ~n26612;
  assign n26614 = n22860 & ~n26613;
  assign po2631 = n26610 | n26614;
  assign n26616 = ~pi2458 & ~n22860;
  assign n26617 = ~pi2458 & ~n22893;
  assign n26618 = n22893 & ~n23664;
  assign n26619 = ~n26617 & ~n26618;
  assign n26620 = n22860 & ~n26619;
  assign po2632 = n26616 | n26620;
  assign n26622 = ~pi2459 & ~n22860;
  assign n26623 = n22952 & ~n23461;
  assign n26624 = ~pi2459 & ~n22952;
  assign n26625 = ~n26623 & ~n26624;
  assign n26626 = n22860 & ~n26625;
  assign po2633 = n26622 | n26626;
  assign n26628 = ~pi2460 & ~n22860;
  assign n26629 = n22952 & ~n23428;
  assign n26630 = ~pi2460 & ~n22952;
  assign n26631 = ~n26629 & ~n26630;
  assign n26632 = n22860 & ~n26631;
  assign po2634 = n26628 | n26632;
  assign n26634 = pi1703 & n22080;
  assign n26635 = pi2461 & ~n23726;
  assign n26636 = ~pi2252 & n23728;
  assign n26637 = ~pi2526 & n26636;
  assign n26638 = ~pi1972 & n26637;
  assign n26639 = pi2461 & n26638;
  assign n26640 = ~pi2461 & ~n26638;
  assign n26641 = ~n26639 & ~n26640;
  assign n26642 = n23726 & n26641;
  assign n26643 = ~n26635 & ~n26642;
  assign n26644 = ~n22080 & ~n26643;
  assign po2635 = n26634 | n26644;
  assign n26646 = ~pi2462 & ~n22860;
  assign n26647 = ~pi2462 & ~n22893;
  assign n26648 = n22893 & ~n23428;
  assign n26649 = ~n26647 & ~n26648;
  assign n26650 = n22860 & ~n26649;
  assign po2636 = n26646 | n26650;
  assign n26652 = pi1670 & n22080;
  assign n26653 = pi2463 & ~n23726;
  assign n26654 = pi2294 & pi2463;
  assign n26655 = ~n23728 & ~n26654;
  assign n26656 = n23726 & ~n26655;
  assign n26657 = ~n26653 & ~n26656;
  assign n26658 = ~n22080 & ~n26657;
  assign po2637 = n26652 | n26658;
  assign n26660 = ~pi2464 & ~n22860;
  assign n26661 = ~pi2464 & ~n22980;
  assign n26662 = n22980 & ~n23638;
  assign n26663 = ~n26661 & ~n26662;
  assign n26664 = n22860 & ~n26663;
  assign po2638 = n26660 | n26664;
  assign n26666 = pi2465 & ~n14916;
  assign n26667 = ~pi3514 & ~pi3516;
  assign n26668 = ~pi3380 & ~pi3381;
  assign n26669 = ~pi3382 & n26668;
  assign n26670 = pi3518 & ~n26669;
  assign n26671 = ~pi3517 & ~n26670;
  assign n26672 = pi3517 & ~pi3518;
  assign n26673 = n26668 & n26672;
  assign n26674 = pi3517 & pi3518;
  assign n26675 = ~pi3383 & n26669;
  assign n26676 = n26674 & n26675;
  assign n26677 = ~n26673 & ~n26676;
  assign n26678 = ~n26671 & n26677;
  assign n26679 = n14916 & ~n26678;
  assign n26680 = n26667 & n26679;
  assign n26681 = pi3515 & n26680;
  assign po2639 = n26666 | n26681;
  assign n26683 = ~pi2466 & ~n22860;
  assign n26684 = ~pi2466 & ~n22893;
  assign n26685 = n22893 & ~n23645;
  assign n26686 = ~n26684 & ~n26685;
  assign n26687 = n22860 & ~n26686;
  assign po2640 = n26683 | n26687;
  assign n26689 = pi2988 & n22311;
  assign n26690 = ~pi2467 & ~n22311;
  assign n26691 = ~n26689 & ~n26690;
  assign n26692 = n22306 & ~n26691;
  assign n26693 = ~pi2467 & ~n22306;
  assign po2641 = n26692 | n26693;
  assign n26695 = ~pi2468 & ~n22860;
  assign n26696 = pi2975 & n22886;
  assign n26697 = ~pi2468 & ~n22886;
  assign n26698 = ~n26696 & ~n26697;
  assign n26699 = n22860 & ~n26698;
  assign po2642 = n26695 | n26699;
  assign n26701 = ~pi2469 & ~n22860;
  assign n26702 = ~pi2469 & ~n22893;
  assign n26703 = n22893 & ~n23953;
  assign n26704 = ~n26702 & ~n26703;
  assign n26705 = n22860 & ~n26704;
  assign po2643 = n26701 | n26705;
  assign n26707 = ~pi2470 & ~n22860;
  assign n26708 = ~pi2470 & ~n22980;
  assign n26709 = n22980 & ~n23511;
  assign n26710 = ~n26708 & ~n26709;
  assign n26711 = n22860 & ~n26710;
  assign po2644 = n26707 | n26711;
  assign n26713 = ~pi2471 & ~n22860;
  assign n26714 = ~pi2471 & ~n22893;
  assign n26715 = n22893 & ~n23320;
  assign n26716 = ~n26714 & ~n26715;
  assign n26717 = n22860 & ~n26716;
  assign po2645 = n26713 | n26717;
  assign n26719 = ~pi2472 & ~n22860;
  assign n26720 = ~pi2472 & ~n22893;
  assign n26721 = n22893 & ~n23355;
  assign n26722 = ~n26720 & ~n26721;
  assign n26723 = n22860 & ~n26722;
  assign po2646 = n26719 | n26723;
  assign n26725 = ~pi2473 & ~n22860;
  assign n26726 = ~pi2473 & ~n22980;
  assign n26727 = n22980 & ~n23862;
  assign n26728 = ~n26726 & ~n26727;
  assign n26729 = n22860 & ~n26728;
  assign po2647 = n26725 | n26729;
  assign n26731 = ~pi2474 & ~n22860;
  assign n26732 = pi2975 & n22867;
  assign n26733 = ~pi2474 & ~n22867;
  assign n26734 = ~n26732 & ~n26733;
  assign n26735 = n22860 & ~n26734;
  assign po2648 = n26731 | n26735;
  assign n26737 = ~pi2475 & ~n22860;
  assign n26738 = pi2975 & n22973;
  assign n26739 = ~pi2475 & ~n22973;
  assign n26740 = ~n26738 & ~n26739;
  assign n26741 = n22860 & ~n26740;
  assign po2649 = n26737 | n26741;
  assign n26743 = ~pi2476 & ~n22860;
  assign n26744 = ~pi2476 & ~n22893;
  assign n26745 = n22893 & ~n23395;
  assign n26746 = ~n26744 & ~n26745;
  assign n26747 = n22860 & ~n26746;
  assign po2650 = n26743 | n26747;
  assign n26749 = ~pi2477 & ~n22860;
  assign n26750 = ~pi2477 & ~n22893;
  assign n26751 = n22893 & ~n23368;
  assign n26752 = ~n26750 & ~n26751;
  assign n26753 = n22860 & ~n26752;
  assign po2651 = n26749 | n26753;
  assign n26755 = ~pi2478 & ~n22860;
  assign n26756 = ~pi2478 & ~n22893;
  assign n26757 = n22893 & ~n23381;
  assign n26758 = ~n26756 & ~n26757;
  assign n26759 = n22860 & ~n26758;
  assign po2652 = n26755 | n26759;
  assign n26761 = pi0325 & n20262;
  assign n26762 = pi2479 & ~n20262;
  assign po2653 = n26761 | n26762;
  assign n26764 = pi0201 & n20262;
  assign n26765 = pi2480 & ~n20262;
  assign po2654 = n26764 | n26765;
  assign n26767 = ~pi2481 & ~n22318;
  assign n26768 = pi3049 & n22318;
  assign n26769 = ~n26767 & ~n26768;
  assign n26770 = n22306 & ~n26769;
  assign n26771 = ~pi2481 & ~n22306;
  assign po2655 = n26770 | n26771;
  assign n26773 = pi0139 & n20262;
  assign n26774 = pi2482 & ~n20262;
  assign po2656 = n26773 | n26774;
  assign n26776 = pi0251 & n20262;
  assign n26777 = pi2483 & ~n20262;
  assign po2657 = n26776 | n26777;
  assign n26779 = ~pi2484 & ~n22318;
  assign n26780 = pi3100 & n22318;
  assign n26781 = ~n26779 & ~n26780;
  assign n26782 = n22306 & ~n26781;
  assign n26783 = ~pi2484 & ~n22306;
  assign po2658 = n26782 | n26783;
  assign n26785 = pi0024 & ~n23715;
  assign n26786 = pi2485 & n23715;
  assign po2659 = n26785 | n26786;
  assign n26788 = pi2486 & ~n10977;
  assign n26789 = ~pi1265 & n19974;
  assign n26790 = ~n19975 & ~n26789;
  assign n26791 = n10977 & ~n26790;
  assign po2660 = n26788 | n26791;
  assign n26793 = ~pi2487 & ~n22547;
  assign n26794 = pi3095 & n22547;
  assign n26795 = ~n26793 & ~n26794;
  assign n26796 = n22306 & ~n26795;
  assign n26797 = ~pi2487 & ~n22306;
  assign po2661 = n26796 | n26797;
  assign n26799 = pi0135 & n20262;
  assign n26800 = pi2488 & ~n20262;
  assign po2662 = n26799 | n26800;
  assign n26802 = pi0299 & n20262;
  assign n26803 = pi2489 & ~n20262;
  assign po2663 = n26802 | n26803;
  assign n26805 = ~pi2490 & ~n22318;
  assign n26806 = pi3086 & n22318;
  assign n26807 = ~n26805 & ~n26806;
  assign n26808 = n22306 & ~n26807;
  assign n26809 = ~pi2490 & ~n22306;
  assign po2664 = n26808 | n26809;
  assign n26811 = pi3053 & n22554;
  assign n26812 = ~pi2491 & ~n22554;
  assign n26813 = ~n26811 & ~n26812;
  assign n26814 = n22306 & ~n26813;
  assign n26815 = ~pi2491 & ~n22306;
  assign po2665 = n26814 | n26815;
  assign n26817 = ~pi2492 & ~n22318;
  assign n26818 = pi3098 & n22318;
  assign n26819 = ~n26817 & ~n26818;
  assign n26820 = n22306 & ~n26819;
  assign n26821 = ~pi2492 & ~n22306;
  assign po2666 = n26820 | n26821;
  assign n26823 = pi3060 & n22302;
  assign n26824 = ~pi2493 & ~n22302;
  assign n26825 = ~n26823 & ~n26824;
  assign n26826 = n22306 & ~n26825;
  assign n26827 = ~pi2493 & ~n22306;
  assign po2667 = n26826 | n26827;
  assign n26829 = pi3053 & n22311;
  assign n26830 = ~pi2494 & ~n22311;
  assign n26831 = ~n26829 & ~n26830;
  assign n26832 = n22306 & ~n26831;
  assign n26833 = ~pi2494 & ~n22306;
  assign po2668 = n26832 | n26833;
  assign n26835 = pi3058 & n22311;
  assign n26836 = ~pi2495 & ~n22311;
  assign n26837 = ~n26835 & ~n26836;
  assign n26838 = n22306 & ~n26837;
  assign n26839 = ~pi2495 & ~n22306;
  assign po2669 = n26838 | n26839;
  assign n26841 = pi0151 & n20262;
  assign n26842 = pi2496 & ~n20262;
  assign po2670 = n26841 | n26842;
  assign n26844 = ~pi2497 & ~n22318;
  assign n26845 = pi3047 & n22318;
  assign n26846 = ~n26844 & ~n26845;
  assign n26847 = n22306 & ~n26846;
  assign n26848 = ~pi2497 & ~n22306;
  assign po2671 = n26847 | n26848;
  assign n26850 = ~pi2498 & ~n22318;
  assign n26851 = pi3097 & n22318;
  assign n26852 = ~n26850 & ~n26851;
  assign n26853 = n22306 & ~n26852;
  assign n26854 = ~pi2498 & ~n22306;
  assign po2672 = n26853 | n26854;
  assign n26856 = pi0153 & n20262;
  assign n26857 = pi2499 & ~n20262;
  assign po2673 = n26856 | n26857;
  assign n26859 = pi3050 & n22311;
  assign n26860 = ~pi2500 & ~n22311;
  assign n26861 = ~n26859 & ~n26860;
  assign n26862 = n22306 & ~n26861;
  assign n26863 = ~pi2500 & ~n22306;
  assign po2674 = n26862 | n26863;
  assign n26865 = pi0192 & n20262;
  assign n26866 = pi2501 & ~n20262;
  assign po2675 = n26865 | n26866;
  assign n26868 = pi0149 & n20262;
  assign n26869 = pi2502 & ~n20262;
  assign po2676 = n26868 | n26869;
  assign n26871 = pi0130 & n20262;
  assign n26872 = pi2503 & ~n20262;
  assign po2677 = n26871 | n26872;
  assign n26874 = ~pi2504 & ~n22539;
  assign n26875 = pi3099 & n22539;
  assign n26876 = ~n26874 & ~n26875;
  assign n26877 = n22306 & ~n26876;
  assign n26878 = ~pi2504 & ~n22306;
  assign po2678 = n26877 | n26878;
  assign n26880 = pi0145 & n20262;
  assign n26881 = pi2505 & ~n20262;
  assign po2679 = n26880 | n26881;
  assign n26883 = pi0144 & n20262;
  assign n26884 = pi2506 & ~n20262;
  assign po2680 = n26883 | n26884;
  assign n26886 = pi3056 & n22311;
  assign n26887 = ~pi2507 & ~n22311;
  assign n26888 = ~n26886 & ~n26887;
  assign n26889 = n22306 & ~n26888;
  assign n26890 = ~pi2507 & ~n22306;
  assign po2681 = n26889 | n26890;
  assign n26892 = pi0143 & n20262;
  assign n26893 = pi2508 & ~n20262;
  assign po2682 = n26892 | n26893;
  assign n26895 = ~pi2509 & ~n22318;
  assign n26896 = pi3088 & n22318;
  assign n26897 = ~n26895 & ~n26896;
  assign n26898 = n22306 & ~n26897;
  assign n26899 = ~pi2509 & ~n22306;
  assign po2683 = n26898 | n26899;
  assign n26901 = ~pi2510 & ~n22539;
  assign n26902 = pi3060 & n22539;
  assign n26903 = ~n26901 & ~n26902;
  assign n26904 = n22306 & ~n26903;
  assign n26905 = ~pi2510 & ~n22306;
  assign po2684 = n26904 | n26905;
  assign n26907 = pi3061 & n22311;
  assign n26908 = ~pi2511 & ~n22311;
  assign n26909 = ~n26907 & ~n26908;
  assign n26910 = n22306 & ~n26909;
  assign n26911 = ~pi2511 & ~n22306;
  assign po2685 = n26910 | n26911;
  assign n26913 = pi3047 & n22311;
  assign n26914 = ~pi2512 & ~n22311;
  assign n26915 = ~n26913 & ~n26914;
  assign n26916 = n22306 & ~n26915;
  assign n26917 = ~pi2512 & ~n22306;
  assign po2686 = n26916 | n26917;
  assign n26919 = ~pi2513 & ~n22539;
  assign n26920 = pi3047 & n22539;
  assign n26921 = ~n26919 & ~n26920;
  assign n26922 = n22306 & ~n26921;
  assign n26923 = ~pi2513 & ~n22306;
  assign po2687 = n26922 | n26923;
  assign n26925 = ~pi2514 & ~n22539;
  assign n26926 = pi3086 & n22539;
  assign n26927 = ~n26925 & ~n26926;
  assign n26928 = n22306 & ~n26927;
  assign n26929 = ~pi2514 & ~n22306;
  assign po2688 = n26928 | n26929;
  assign n26931 = pi3062 & n22302;
  assign n26932 = ~pi2515 & ~n22302;
  assign n26933 = ~n26931 & ~n26932;
  assign n26934 = n22306 & ~n26933;
  assign n26935 = ~pi2515 & ~n22306;
  assign po2689 = n26934 | n26935;
  assign n26937 = pi3048 & n22561;
  assign n26938 = ~pi2516 & ~n22561;
  assign n26939 = ~n26937 & ~n26938;
  assign n26940 = n22306 & ~n26939;
  assign n26941 = ~pi2516 & ~n22306;
  assign po2690 = n26940 | n26941;
  assign n26943 = pi3059 & n22311;
  assign n26944 = ~pi2517 & ~n22311;
  assign n26945 = ~n26943 & ~n26944;
  assign n26946 = n22306 & ~n26945;
  assign n26947 = ~pi2517 & ~n22306;
  assign po2691 = n26946 | n26947;
  assign n26949 = pi0177 & n20262;
  assign n26950 = pi2518 & ~n20262;
  assign po2692 = n26949 | n26950;
  assign n26952 = ~pi1816 & n22621;
  assign n26953 = pi1337 & n26952;
  assign n26954 = pi1761 & n26953;
  assign n26955 = n19459 & ~n22621;
  assign po2693 = n26954 | n26955;
  assign n26957 = pi2520 & n23715;
  assign n26958 = n23714 & ~n23715;
  assign po2694 = n26957 | n26958;
  assign n26960 = pi2521 & n23715;
  assign po2695 = n26958 | n26960;
  assign n26962 = pi2522 & n23715;
  assign n26963 = ~pi0005 & ~n23715;
  assign po2696 = n26962 | n26963;
  assign n26965 = pi2523 & n23715;
  assign n26966 = ~pi0003 & ~n23715;
  assign po2697 = n26965 | n26966;
  assign n26968 = pi2524 & n23715;
  assign n26969 = ~pi0004 & ~n23715;
  assign po2698 = n26968 | n26969;
  assign n26971 = pi2525 & n22622;
  assign n26972 = pi2525 & pi2874;
  assign n26973 = ~n22632 & ~n26972;
  assign n26974 = pi1337 & ~n26973;
  assign n26975 = ~n22628 & ~n26974;
  assign n26976 = ~n22622 & ~n26975;
  assign po2699 = n26971 | n26976;
  assign n26978 = pi1702 & n22080;
  assign n26979 = pi2526 & ~n23729;
  assign n26980 = ~pi2526 & n23729;
  assign n26981 = ~n26979 & ~n26980;
  assign n26982 = n23726 & ~n26981;
  assign n26983 = pi2526 & ~n23726;
  assign n26984 = ~n26982 & ~n26983;
  assign n26985 = ~n22080 & ~n26984;
  assign po2700 = n26978 | n26985;
  assign n26987 = pi0069 & ~n23715;
  assign n26988 = pi2527 & n23715;
  assign po2701 = n26987 | n26988;
  assign n26990 = pi0052 & ~n23715;
  assign n26991 = pi2528 & n23715;
  assign po2702 = n26990 | n26991;
  assign n26993 = pi0053 & ~n23715;
  assign n26994 = pi2529 & n23715;
  assign po2703 = n26993 | n26994;
  assign n26996 = pi0067 & ~n23715;
  assign n26997 = pi2530 & n23715;
  assign po2704 = n26996 | n26997;
  assign n26999 = pi0039 & ~n23715;
  assign n27000 = pi2531 & n23715;
  assign po2705 = n26999 | n27000;
  assign n27002 = pi0042 & ~n23715;
  assign n27003 = pi2532 & n23715;
  assign po2706 = n27002 | n27003;
  assign n27005 = pi0040 & ~n23715;
  assign n27006 = pi2533 & n23715;
  assign po2707 = n27005 | n27006;
  assign n27008 = pi0058 & ~n23715;
  assign n27009 = pi2534 & n23715;
  assign po2708 = n27008 | n27009;
  assign n27011 = pi0047 & ~n23715;
  assign n27012 = pi2535 & n23715;
  assign po2709 = n27011 | n27012;
  assign n27014 = pi0065 & ~n23715;
  assign n27015 = pi2536 & n23715;
  assign po2710 = n27014 | n27015;
  assign n27017 = pi0048 & ~n23715;
  assign n27018 = pi2537 & n23715;
  assign po2711 = n27017 | n27018;
  assign n27020 = pi0060 & ~n23715;
  assign n27021 = pi2538 & n23715;
  assign po2712 = n27020 | n27021;
  assign n27023 = pi0062 & ~n23715;
  assign n27024 = pi2539 & n23715;
  assign po2713 = n27023 | n27024;
  assign n27026 = pi0063 & ~n23715;
  assign n27027 = pi2540 & n23715;
  assign po2714 = n27026 | n27027;
  assign n27029 = pi0007 & ~n23715;
  assign n27030 = pi2541 & n23715;
  assign po2715 = n27029 | n27030;
  assign n27032 = pi0009 & ~n23715;
  assign n27033 = pi2542 & n23715;
  assign po2716 = n27032 | n27033;
  assign n27035 = pi0011 & ~n23715;
  assign n27036 = pi2543 & n23715;
  assign po2717 = n27035 | n27036;
  assign n27038 = pi0038 & ~n23715;
  assign n27039 = pi2544 & n23715;
  assign po2718 = n27038 | n27039;
  assign n27041 = pi0013 & ~n23715;
  assign n27042 = pi2545 & n23715;
  assign po2719 = n27041 | n27042;
  assign n27044 = pi0014 & ~n23715;
  assign n27045 = pi2546 & n23715;
  assign po2720 = n27044 | n27045;
  assign n27047 = pi0017 & ~n23715;
  assign n27048 = pi2547 & n23715;
  assign po2721 = n27047 | n27048;
  assign n27050 = pi0021 & ~n23715;
  assign n27051 = pi2548 & n23715;
  assign po2722 = n27050 | n27051;
  assign n27053 = pi0025 & ~n23715;
  assign n27054 = pi2549 & n23715;
  assign po2723 = n27053 | n27054;
  assign n27056 = pi0027 & ~n23715;
  assign n27057 = pi2550 & n23715;
  assign po2724 = n27056 | n27057;
  assign n27059 = pi0028 & ~n23715;
  assign n27060 = pi2551 & n23715;
  assign po2725 = n27059 | n27060;
  assign n27062 = pi0037 & ~n23715;
  assign n27063 = pi2552 & n23715;
  assign po2726 = n27062 | n27063;
  assign n27065 = pi2553 & ~n8009;
  assign n27066 = ~pi3018 & pi3102;
  assign n27067 = pi3018 & ~pi3102;
  assign n27068 = ~n27066 & ~n27067;
  assign n27069 = pi3007 & ~pi3057;
  assign n27070 = ~pi3007 & pi3057;
  assign n27071 = ~n27069 & ~n27070;
  assign n27072 = n27068 & n27071;
  assign n27073 = ~pi3020 & pi3112;
  assign n27074 = pi3020 & ~pi3112;
  assign n27075 = ~n27073 & ~n27074;
  assign n27076 = ~pi2972 & pi3111;
  assign n27077 = pi2972 & ~pi3111;
  assign n27078 = ~n27076 & ~n27077;
  assign n27079 = n27075 & n27078;
  assign n27080 = n27072 & n27079;
  assign n27081 = pi3006 & ~pi3162;
  assign n27082 = ~pi3006 & pi3162;
  assign n27083 = ~n27081 & ~n27082;
  assign n27084 = pi3031 & ~pi3154;
  assign n27085 = ~pi3031 & pi3154;
  assign n27086 = ~n27084 & ~n27085;
  assign n27087 = n27083 & n27086;
  assign n27088 = pi3005 & ~pi3165;
  assign n27089 = ~pi3005 & pi3165;
  assign n27090 = ~n27088 & ~n27089;
  assign n27091 = pi3033 & ~pi3155;
  assign n27092 = ~pi3033 & pi3155;
  assign n27093 = ~n27091 & ~n27092;
  assign n27094 = n27090 & n27093;
  assign n27095 = pi3072 & ~pi3171;
  assign n27096 = ~pi3072 & pi3171;
  assign n27097 = ~n27095 & ~n27096;
  assign n27098 = pi3116 & ~pi3132;
  assign n27099 = ~pi3116 & pi3132;
  assign n27100 = ~n27098 & ~n27099;
  assign n27101 = n27097 & n27100;
  assign n27102 = pi3114 & ~pi3164;
  assign n27103 = ~pi3114 & pi3164;
  assign n27104 = ~n27102 & ~n27103;
  assign n27105 = pi3013 & ~pi3134;
  assign n27106 = ~pi3013 & pi3134;
  assign n27107 = ~n27105 & ~n27106;
  assign n27108 = n27104 & n27107;
  assign n27109 = n27101 & n27108;
  assign n27110 = n27094 & n27109;
  assign n27111 = n27087 & n27110;
  assign n27112 = pi3051 & ~pi3158;
  assign n27113 = ~pi3051 & pi3158;
  assign n27114 = ~n27112 & ~n27113;
  assign n27115 = pi3032 & ~pi3135;
  assign n27116 = ~pi3032 & pi3135;
  assign n27117 = ~n27115 & ~n27116;
  assign n27118 = n27114 & n27117;
  assign n27119 = pi3074 & ~pi3133;
  assign n27120 = ~pi3074 & pi3133;
  assign n27121 = ~n27119 & ~n27120;
  assign n27122 = pi3113 & ~pi3150;
  assign n27123 = ~pi3113 & pi3150;
  assign n27124 = ~n27122 & ~n27123;
  assign n27125 = n27121 & n27124;
  assign n27126 = pi3044 & ~pi3172;
  assign n27127 = ~pi3044 & pi3172;
  assign n27128 = ~n27126 & ~n27127;
  assign n27129 = pi3028 & ~pi3157;
  assign n27130 = ~pi3028 & pi3157;
  assign n27131 = ~n27129 & ~n27130;
  assign n27132 = n27128 & n27131;
  assign n27133 = pi3029 & ~pi3151;
  assign n27134 = ~pi3029 & pi3151;
  assign n27135 = ~n27133 & ~n27134;
  assign n27136 = pi3030 & ~pi3138;
  assign n27137 = ~pi3030 & pi3138;
  assign n27138 = ~n27136 & ~n27137;
  assign n27139 = n27135 & n27138;
  assign n27140 = n27132 & n27139;
  assign n27141 = n27125 & n27140;
  assign n27142 = n27118 & n27141;
  assign n27143 = n27111 & n27142;
  assign n27144 = pi3066 & ~pi3163;
  assign n27145 = ~pi3066 & pi3163;
  assign n27146 = ~n27144 & ~n27145;
  assign n27147 = pi3115 & ~pi3136;
  assign n27148 = ~pi3115 & pi3136;
  assign n27149 = ~n27147 & ~n27148;
  assign n27150 = n27146 & n27149;
  assign n27151 = pi3026 & ~pi3166;
  assign n27152 = ~pi3026 & pi3166;
  assign n27153 = ~n27151 & ~n27152;
  assign n27154 = pi3076 & ~pi3142;
  assign n27155 = ~pi3076 & pi3142;
  assign n27156 = ~n27154 & ~n27155;
  assign n27157 = n27153 & n27156;
  assign n27158 = pi3067 & ~pi3147;
  assign n27159 = ~pi3067 & pi3147;
  assign n27160 = ~n27158 & ~n27159;
  assign n27161 = pi3073 & ~pi3153;
  assign n27162 = ~pi3073 & pi3153;
  assign n27163 = ~n27161 & ~n27162;
  assign n27164 = n27160 & n27163;
  assign n27165 = pi3080 & ~pi3141;
  assign n27166 = ~pi3080 & pi3141;
  assign n27167 = ~n27165 & ~n27166;
  assign n27168 = pi3078 & ~pi3143;
  assign n27169 = ~pi3078 & pi3143;
  assign n27170 = ~n27168 & ~n27169;
  assign n27171 = n27167 & n27170;
  assign n27172 = n27164 & n27171;
  assign n27173 = n27157 & n27172;
  assign n27174 = n27150 & n27173;
  assign n27175 = pi3037 & ~pi3131;
  assign n27176 = ~pi3037 & pi3131;
  assign n27177 = ~n27175 & ~n27176;
  assign n27178 = pi3068 & ~pi3159;
  assign n27179 = ~pi3068 & pi3159;
  assign n27180 = ~n27178 & ~n27179;
  assign n27181 = n27177 & n27180;
  assign n27182 = pi3105 & ~pi3169;
  assign n27183 = ~pi3105 & pi3169;
  assign n27184 = ~n27182 & ~n27183;
  assign n27185 = pi3035 & ~pi3145;
  assign n27186 = ~pi3035 & pi3145;
  assign n27187 = ~n27185 & ~n27186;
  assign n27188 = n27184 & n27187;
  assign n27189 = pi3069 & ~pi3168;
  assign n27190 = ~pi3069 & pi3168;
  assign n27191 = ~n27189 & ~n27190;
  assign n27192 = pi3075 & ~pi3170;
  assign n27193 = ~pi3075 & pi3170;
  assign n27194 = ~n27192 & ~n27193;
  assign n27195 = n27191 & n27194;
  assign n27196 = pi3081 & ~pi3139;
  assign n27197 = ~pi3081 & pi3139;
  assign n27198 = ~n27196 & ~n27197;
  assign n27199 = pi3046 & ~pi3146;
  assign n27200 = ~pi3046 & pi3146;
  assign n27201 = ~n27199 & ~n27200;
  assign n27202 = n27198 & n27201;
  assign n27203 = n27195 & n27202;
  assign n27204 = n27188 & n27203;
  assign n27205 = n27181 & n27204;
  assign n27206 = n27174 & n27205;
  assign n27207 = n27143 & n27206;
  assign n27208 = n8009 & n27207;
  assign n27209 = n27080 & n27208;
  assign po2727 = n27065 | n27209;
  assign n27211 = pi1683 & n20262;
  assign n27212 = pi2554 & ~n20262;
  assign po2728 = n27211 | n27212;
  assign n27214 = pi0136 & n20262;
  assign n27215 = pi2555 & ~n20262;
  assign po2729 = n27214 | n27215;
  assign n27217 = pi0187 & n20262;
  assign n27218 = pi2556 & ~n20262;
  assign po2730 = n27217 | n27218;
  assign n27220 = pi0189 & n20262;
  assign n27221 = pi2557 & ~n20262;
  assign po2731 = n27220 | n27221;
  assign n27223 = pi0190 & n20262;
  assign n27224 = pi2558 & ~n20262;
  assign po2732 = n27223 | n27224;
  assign n27226 = pi0172 & n20262;
  assign n27227 = pi2559 & ~n20262;
  assign po2733 = n27226 | n27227;
  assign n27229 = pi0141 & n20262;
  assign n27230 = pi2560 & ~n20262;
  assign po2734 = n27229 | n27230;
  assign n27232 = pi0173 & n20262;
  assign n27233 = pi2561 & ~n20262;
  assign po2735 = n27232 | n27233;
  assign n27235 = pi0175 & n20262;
  assign n27236 = pi2562 & ~n20262;
  assign po2736 = n27235 | n27236;
  assign n27238 = pi0176 & n20262;
  assign n27239 = pi2563 & ~n20262;
  assign po2737 = n27238 | n27239;
  assign n27241 = pi0191 & n20262;
  assign n27242 = pi2564 & ~n20262;
  assign po2738 = n27241 | n27242;
  assign n27244 = pi0195 & n20262;
  assign n27245 = pi2565 & ~n20262;
  assign po2739 = n27244 | n27245;
  assign n27247 = pi0178 & n20262;
  assign n27248 = pi2566 & ~n20262;
  assign po2740 = n27247 | n27248;
  assign n27250 = pi0142 & n20262;
  assign n27251 = pi2567 & ~n20262;
  assign po2741 = n27250 | n27251;
  assign n27253 = pi0203 & n20262;
  assign n27254 = pi2568 & ~n20262;
  assign po2742 = n27253 | n27254;
  assign n27256 = pi0198 & n20262;
  assign n27257 = pi2569 & ~n20262;
  assign po2743 = n27256 | n27257;
  assign n27259 = pi0146 & n20262;
  assign n27260 = pi2570 & ~n20262;
  assign po2744 = n27259 | n27260;
  assign n27262 = pi0147 & n20262;
  assign n27263 = pi2571 & ~n20262;
  assign po2745 = n27262 | n27263;
  assign n27265 = pi0148 & n20262;
  assign n27266 = pi2572 & ~n20262;
  assign po2746 = n27265 | n27266;
  assign n27268 = pi0150 & n20262;
  assign n27269 = pi2573 & ~n20262;
  assign po2747 = n27268 | n27269;
  assign n27271 = pi0179 & n20262;
  assign n27272 = pi2574 & ~n20262;
  assign po2748 = n27271 | n27272;
  assign n27274 = pi0152 & n20262;
  assign n27275 = pi2575 & ~n20262;
  assign po2749 = n27274 | n27275;
  assign n27277 = pi0303 & n20262;
  assign n27278 = pi2576 & ~n20262;
  assign po2750 = n27277 | n27278;
  assign n27280 = pi0304 & n20262;
  assign n27281 = pi2577 & ~n20262;
  assign po2751 = n27280 | n27281;
  assign n27283 = pi0298 & n20262;
  assign n27284 = pi2578 & ~n20262;
  assign po2752 = n27283 | n27284;
  assign n27286 = pi0249 & n20262;
  assign n27287 = pi2579 & ~n20262;
  assign po2753 = n27286 | n27287;
  assign n27289 = pi0250 & n20262;
  assign n27290 = pi2580 & ~n20262;
  assign po2754 = n27289 | n27290;
  assign n27292 = pi0272 & n20262;
  assign n27293 = pi2581 & ~n20262;
  assign po2755 = n27292 | n27293;
  assign n27295 = pi0252 & n20262;
  assign n27296 = pi2582 & ~n20262;
  assign po2756 = n27295 | n27296;
  assign n27298 = pi0253 & n20262;
  assign n27299 = pi2583 & ~n20262;
  assign po2757 = n27298 | n27299;
  assign n27301 = pi0255 & n20262;
  assign n27302 = pi2584 & ~n20262;
  assign po2758 = n27301 | n27302;
  assign n27304 = pi0247 & n20262;
  assign n27305 = pi2585 & ~n20262;
  assign po2759 = n27304 | n27305;
  assign n27307 = pi0257 & n20262;
  assign n27308 = pi2586 & ~n20262;
  assign po2760 = n27307 | n27308;
  assign n27310 = pi0268 & n20262;
  assign n27311 = pi2587 & ~n20262;
  assign po2761 = n27310 | n27311;
  assign n27313 = ~pi0259 & n20262;
  assign n27314 = pi2588 & ~n20262;
  assign po2762 = n27313 | n27314;
  assign n27316 = pi0260 & n20262;
  assign n27317 = pi2589 & ~n20262;
  assign po2763 = n27316 | n27317;
  assign n27319 = pi0261 & n20262;
  assign n27320 = pi2590 & ~n20262;
  assign po2764 = n27319 | n27320;
  assign n27322 = pi0262 & n20262;
  assign n27323 = pi2591 & ~n20262;
  assign po2765 = n27322 | n27323;
  assign n27325 = pi0302 & n20262;
  assign n27326 = pi2592 & ~n20262;
  assign po2766 = n27325 | n27326;
  assign n27328 = ~pi3082 & n22306;
  assign n27329 = pi2593 & pi2906;
  assign n27330 = ~pi2593 & ~pi2906;
  assign n27331 = ~n27329 & ~n27330;
  assign n27332 = n27328 & ~n27331;
  assign n27333 = ~pi2593 & ~n27328;
  assign po2767 = n27332 | n27333;
  assign n27335 = ~pi2594 & ~n27328;
  assign po2768 = n27332 | n27335;
  assign n27337 = pi3101 & n22311;
  assign n27338 = ~pi2595 & ~n22311;
  assign n27339 = ~n27337 & ~n27338;
  assign n27340 = n22306 & ~n27339;
  assign n27341 = ~pi2595 & ~n22306;
  assign po2769 = n27340 | n27341;
  assign n27343 = pi3062 & n22311;
  assign n27344 = ~pi2596 & ~n22311;
  assign n27345 = ~n27343 & ~n27344;
  assign n27346 = n22306 & ~n27345;
  assign n27347 = ~pi2596 & ~n22306;
  assign po2770 = n27346 | n27347;
  assign n27349 = pi3085 & n22311;
  assign n27350 = ~pi2597 & ~n22311;
  assign n27351 = ~n27349 & ~n27350;
  assign n27352 = n22306 & ~n27351;
  assign n27353 = ~pi2597 & ~n22306;
  assign po2771 = n27352 | n27353;
  assign n27355 = pi3049 & n22311;
  assign n27356 = ~pi2598 & ~n22311;
  assign n27357 = ~n27355 & ~n27356;
  assign n27358 = n22306 & ~n27357;
  assign n27359 = ~pi2598 & ~n22306;
  assign po2772 = n27358 | n27359;
  assign n27361 = pi3094 & n22561;
  assign n27362 = ~pi2599 & ~n22561;
  assign n27363 = ~n27361 & ~n27362;
  assign n27364 = n22306 & ~n27363;
  assign n27365 = ~pi2599 & ~n22306;
  assign po2773 = n27364 | n27365;
  assign n27367 = pi3097 & n22311;
  assign n27368 = ~pi2600 & ~n22311;
  assign n27369 = ~n27367 & ~n27368;
  assign n27370 = n22306 & ~n27369;
  assign n27371 = ~pi2600 & ~n22306;
  assign po2774 = n27370 | n27371;
  assign n27373 = pi3092 & n22311;
  assign n27374 = ~pi2601 & ~n22311;
  assign n27375 = ~n27373 & ~n27374;
  assign n27376 = n22306 & ~n27375;
  assign n27377 = ~pi2601 & ~n22306;
  assign po2775 = n27376 | n27377;
  assign n27379 = pi3091 & n22561;
  assign n27380 = ~pi2602 & ~n22561;
  assign n27381 = ~n27379 & ~n27380;
  assign n27382 = n22306 & ~n27381;
  assign n27383 = ~pi2602 & ~n22306;
  assign po2776 = n27382 | n27383;
  assign n27385 = pi3055 & n22561;
  assign n27386 = ~pi2603 & ~n22561;
  assign n27387 = ~n27385 & ~n27386;
  assign n27388 = n22306 & ~n27387;
  assign n27389 = ~pi2603 & ~n22306;
  assign po2777 = n27388 | n27389;
  assign n27391 = pi3099 & n22554;
  assign n27392 = ~pi2604 & ~n22554;
  assign n27393 = ~n27391 & ~n27392;
  assign n27394 = n22306 & ~n27393;
  assign n27395 = ~pi2604 & ~n22306;
  assign po2778 = n27394 | n27395;
  assign n27397 = pi3056 & n22561;
  assign n27398 = ~pi2605 & ~n22561;
  assign n27399 = ~n27397 & ~n27398;
  assign n27400 = n22306 & ~n27399;
  assign n27401 = ~pi2605 & ~n22306;
  assign po2779 = n27400 | n27401;
  assign n27403 = pi3085 & n22302;
  assign n27404 = ~pi2606 & ~n22302;
  assign n27405 = ~n27403 & ~n27404;
  assign n27406 = n22306 & ~n27405;
  assign n27407 = ~pi2606 & ~n22306;
  assign po2780 = n27406 | n27407;
  assign n27409 = pi3045 & n22302;
  assign n27410 = ~pi2607 & ~n22302;
  assign n27411 = ~n27409 & ~n27410;
  assign n27412 = n22306 & ~n27411;
  assign n27413 = ~pi2607 & ~n22306;
  assign po2781 = n27412 | n27413;
  assign n27415 = pi3099 & n22302;
  assign n27416 = ~pi2608 & ~n22302;
  assign n27417 = ~n27415 & ~n27416;
  assign n27418 = n22306 & ~n27417;
  assign n27419 = ~pi2608 & ~n22306;
  assign po2782 = n27418 | n27419;
  assign n27421 = pi3101 & n22302;
  assign n27422 = ~pi2609 & ~n22302;
  assign n27423 = ~n27421 & ~n27422;
  assign n27424 = n22306 & ~n27423;
  assign n27425 = ~pi2609 & ~n22306;
  assign po2783 = n27424 | n27425;
  assign n27427 = pi3049 & n22302;
  assign n27428 = ~pi2610 & ~n22302;
  assign n27429 = ~n27427 & ~n27428;
  assign n27430 = n22306 & ~n27429;
  assign n27431 = ~pi2610 & ~n22306;
  assign po2784 = n27430 | n27431;
  assign n27433 = pi3088 & n22302;
  assign n27434 = ~pi2611 & ~n22302;
  assign n27435 = ~n27433 & ~n27434;
  assign n27436 = n22306 & ~n27435;
  assign n27437 = ~pi2611 & ~n22306;
  assign po2785 = n27436 | n27437;
  assign n27439 = pi3100 & n22302;
  assign n27440 = ~pi2612 & ~n22302;
  assign n27441 = ~n27439 & ~n27440;
  assign n27442 = n22306 & ~n27441;
  assign n27443 = ~pi2612 & ~n22306;
  assign po2786 = n27442 | n27443;
  assign n27445 = pi3089 & n22302;
  assign n27446 = ~pi2613 & ~n22302;
  assign n27447 = ~n27445 & ~n27446;
  assign n27448 = n22306 & ~n27447;
  assign n27449 = ~pi2613 & ~n22306;
  assign po2787 = n27448 | n27449;
  assign n27451 = pi3061 & n22302;
  assign n27452 = ~pi2614 & ~n22302;
  assign n27453 = ~n27451 & ~n27452;
  assign n27454 = n22306 & ~n27453;
  assign n27455 = ~pi2614 & ~n22306;
  assign po2788 = n27454 | n27455;
  assign n27457 = pi3058 & n22302;
  assign n27458 = ~pi2615 & ~n22302;
  assign n27459 = ~n27457 & ~n27458;
  assign n27460 = n22306 & ~n27459;
  assign n27461 = ~pi2615 & ~n22306;
  assign po2789 = n27460 | n27461;
  assign n27463 = pi3091 & n22302;
  assign n27464 = ~pi2616 & ~n22302;
  assign n27465 = ~n27463 & ~n27464;
  assign n27466 = n22306 & ~n27465;
  assign n27467 = ~pi2616 & ~n22306;
  assign po2790 = n27466 | n27467;
  assign n27469 = pi3048 & n22302;
  assign n27470 = ~pi2617 & ~n22302;
  assign n27471 = ~n27469 & ~n27470;
  assign n27472 = n22306 & ~n27471;
  assign n27473 = ~pi2617 & ~n22306;
  assign po2791 = n27472 | n27473;
  assign n27475 = pi3093 & n22302;
  assign n27476 = ~pi2618 & ~n22302;
  assign n27477 = ~n27475 & ~n27476;
  assign n27478 = n22306 & ~n27477;
  assign n27479 = ~pi2618 & ~n22306;
  assign po2792 = n27478 | n27479;
  assign n27481 = pi3094 & n22302;
  assign n27482 = ~pi2619 & ~n22302;
  assign n27483 = ~n27481 & ~n27482;
  assign n27484 = n22306 & ~n27483;
  assign n27485 = ~pi2619 & ~n22306;
  assign po2793 = n27484 | n27485;
  assign n27487 = pi3084 & n22561;
  assign n27488 = ~pi2620 & ~n22561;
  assign n27489 = ~n27487 & ~n27488;
  assign n27490 = n22306 & ~n27489;
  assign n27491 = ~pi2620 & ~n22306;
  assign po2794 = n27490 | n27491;
  assign n27493 = pi3062 & n22561;
  assign n27494 = ~pi2621 & ~n22561;
  assign n27495 = ~n27493 & ~n27494;
  assign n27496 = n22306 & ~n27495;
  assign n27497 = ~pi2621 & ~n22306;
  assign po2795 = n27496 | n27497;
  assign n27499 = pi3101 & n22561;
  assign n27500 = ~pi2622 & ~n22561;
  assign n27501 = ~n27499 & ~n27500;
  assign n27502 = n22306 & ~n27501;
  assign n27503 = ~pi2622 & ~n22306;
  assign po2796 = n27502 | n27503;
  assign n27505 = pi3060 & n22561;
  assign n27506 = ~pi2623 & ~n22561;
  assign n27507 = ~n27505 & ~n27506;
  assign n27508 = n22306 & ~n27507;
  assign n27509 = ~pi2623 & ~n22306;
  assign po2797 = n27508 | n27509;
  assign n27511 = pi3097 & n22561;
  assign n27512 = ~pi2624 & ~n22561;
  assign n27513 = ~n27511 & ~n27512;
  assign n27514 = n22306 & ~n27513;
  assign n27515 = ~pi2624 & ~n22306;
  assign po2798 = n27514 | n27515;
  assign n27517 = pi3096 & n22561;
  assign n27518 = ~pi2625 & ~n22561;
  assign n27519 = ~n27517 & ~n27518;
  assign n27520 = n22306 & ~n27519;
  assign n27521 = ~pi2625 & ~n22306;
  assign po2799 = n27520 | n27521;
  assign n27523 = pi3052 & n22561;
  assign n27524 = ~pi2626 & ~n22561;
  assign n27525 = ~n27523 & ~n27524;
  assign n27526 = n22306 & ~n27525;
  assign n27527 = ~pi2626 & ~n22306;
  assign po2800 = n27526 | n27527;
  assign n27529 = pi3086 & n22311;
  assign n27530 = ~pi2627 & ~n22311;
  assign n27531 = ~n27529 & ~n27530;
  assign n27532 = n22306 & ~n27531;
  assign n27533 = ~pi2627 & ~n22306;
  assign po2801 = n27532 | n27533;
  assign n27535 = pi3087 & n22311;
  assign n27536 = ~pi2628 & ~n22311;
  assign n27537 = ~n27535 & ~n27536;
  assign n27538 = n22306 & ~n27537;
  assign n27539 = ~pi2628 & ~n22306;
  assign po2802 = n27538 | n27539;
  assign n27541 = pi3060 & n22311;
  assign n27542 = ~pi2629 & ~n22311;
  assign n27543 = ~n27541 & ~n27542;
  assign n27544 = n22306 & ~n27543;
  assign n27545 = ~pi2629 & ~n22306;
  assign po2803 = n27544 | n27545;
  assign n27547 = pi3059 & n22302;
  assign n27548 = ~pi2630 & ~n22302;
  assign n27549 = ~n27547 & ~n27548;
  assign n27550 = n22306 & ~n27549;
  assign n27551 = ~pi2630 & ~n22306;
  assign po2804 = n27550 | n27551;
  assign n27553 = pi3090 & n22311;
  assign n27554 = ~pi2631 & ~n22311;
  assign n27555 = ~n27553 & ~n27554;
  assign n27556 = n22306 & ~n27555;
  assign n27557 = ~pi2631 & ~n22306;
  assign po2805 = n27556 | n27557;
  assign n27559 = pi3091 & n22311;
  assign n27560 = ~pi2632 & ~n22311;
  assign n27561 = ~n27559 & ~n27560;
  assign n27562 = n22306 & ~n27561;
  assign n27563 = ~pi2632 & ~n22306;
  assign po2806 = n27562 | n27563;
  assign n27565 = pi3055 & n22311;
  assign n27566 = ~pi2633 & ~n22311;
  assign n27567 = ~n27565 & ~n27566;
  assign n27568 = n22306 & ~n27567;
  assign n27569 = ~pi2633 & ~n22306;
  assign po2807 = n27568 | n27569;
  assign n27571 = pi3093 & n22311;
  assign n27572 = ~pi2634 & ~n22311;
  assign n27573 = ~n27571 & ~n27572;
  assign n27574 = n22306 & ~n27573;
  assign n27575 = ~pi2634 & ~n22306;
  assign po2808 = n27574 | n27575;
  assign n27577 = pi3094 & n22311;
  assign n27578 = ~pi2635 & ~n22311;
  assign n27579 = ~n27577 & ~n27578;
  assign n27580 = n22306 & ~n27579;
  assign n27581 = ~pi2635 & ~n22306;
  assign po2809 = n27580 | n27581;
  assign n27583 = pi3095 & n22311;
  assign n27584 = ~pi2636 & ~n22311;
  assign n27585 = ~n27583 & ~n27584;
  assign n27586 = n22306 & ~n27585;
  assign n27587 = ~pi2636 & ~n22306;
  assign po2810 = n27586 | n27587;
  assign n27589 = pi3098 & n22554;
  assign n27590 = ~pi2637 & ~n22554;
  assign n27591 = ~n27589 & ~n27590;
  assign n27592 = n22306 & ~n27591;
  assign n27593 = ~pi2637 & ~n22306;
  assign po2811 = n27592 | n27593;
  assign n27595 = pi3084 & n22311;
  assign n27596 = ~pi2638 & ~n22311;
  assign n27597 = ~n27595 & ~n27596;
  assign n27598 = n22306 & ~n27597;
  assign n27599 = ~pi2638 & ~n22306;
  assign po2812 = n27598 | n27599;
  assign n27601 = pi3101 & n22554;
  assign n27602 = ~pi2639 & ~n22554;
  assign n27603 = ~n27601 & ~n27602;
  assign n27604 = n22306 & ~n27603;
  assign n27605 = ~pi2639 & ~n22306;
  assign po2813 = n27604 | n27605;
  assign n27607 = pi3049 & n22554;
  assign n27608 = ~pi2640 & ~n22554;
  assign n27609 = ~n27607 & ~n27608;
  assign n27610 = n22306 & ~n27609;
  assign n27611 = ~pi2640 & ~n22306;
  assign po2814 = n27610 | n27611;
  assign n27613 = pi3060 & n22554;
  assign n27614 = ~pi2641 & ~n22554;
  assign n27615 = ~n27613 & ~n27614;
  assign n27616 = n22306 & ~n27615;
  assign n27617 = ~pi2641 & ~n22306;
  assign po2815 = n27616 | n27617;
  assign n27619 = pi3097 & n22302;
  assign n27620 = ~pi2642 & ~n22302;
  assign n27621 = ~n27619 & ~n27620;
  assign n27622 = n22306 & ~n27621;
  assign n27623 = ~pi2642 & ~n22306;
  assign po2816 = n27622 | n27623;
  assign n27625 = pi3088 & n22554;
  assign n27626 = ~pi2643 & ~n22554;
  assign n27627 = ~n27625 & ~n27626;
  assign n27628 = n22306 & ~n27627;
  assign n27629 = ~pi2643 & ~n22306;
  assign po2817 = n27628 | n27629;
  assign n27631 = pi3047 & n22302;
  assign n27632 = ~pi2644 & ~n22302;
  assign n27633 = ~n27631 & ~n27632;
  assign n27634 = n22306 & ~n27633;
  assign n27635 = ~pi2644 & ~n22306;
  assign po2818 = n27634 | n27635;
  assign n27637 = pi3100 & n22554;
  assign n27638 = ~pi2645 & ~n22554;
  assign n27639 = ~n27637 & ~n27638;
  assign n27640 = n22306 & ~n27639;
  assign n27641 = ~pi2645 & ~n22306;
  assign po2819 = n27640 | n27641;
  assign n27643 = ~pi2646 & ~n22539;
  assign n27644 = pi3062 & n22539;
  assign n27645 = ~n27643 & ~n27644;
  assign n27646 = n22306 & ~n27645;
  assign n27647 = ~pi2646 & ~n22306;
  assign po2820 = n27646 | n27647;
  assign n27649 = pi3091 & n22554;
  assign n27650 = ~pi2647 & ~n22554;
  assign n27651 = ~n27649 & ~n27650;
  assign n27652 = n22306 & ~n27651;
  assign n27653 = ~pi2647 & ~n22306;
  assign po2821 = n27652 | n27653;
  assign n27655 = pi3093 & n22554;
  assign n27656 = ~pi2648 & ~n22554;
  assign n27657 = ~n27655 & ~n27656;
  assign n27658 = n22306 & ~n27657;
  assign n27659 = ~pi2648 & ~n22306;
  assign po2822 = n27658 | n27659;
  assign n27661 = pi3094 & n22554;
  assign n27662 = ~pi2649 & ~n22554;
  assign n27663 = ~n27661 & ~n27662;
  assign n27664 = n22306 & ~n27663;
  assign n27665 = ~pi2649 & ~n22306;
  assign po2823 = n27664 | n27665;
  assign n27667 = pi3086 & n22561;
  assign n27668 = ~pi2650 & ~n22561;
  assign n27669 = ~n27667 & ~n27668;
  assign n27670 = n22306 & ~n27669;
  assign n27671 = ~pi2650 & ~n22306;
  assign po2824 = n27670 | n27671;
  assign n27673 = pi3088 & n22561;
  assign n27674 = ~pi2651 & ~n22561;
  assign n27675 = ~n27673 & ~n27674;
  assign n27676 = n22306 & ~n27675;
  assign n27677 = ~pi2651 & ~n22306;
  assign po2825 = n27676 | n27677;
  assign n27679 = pi3047 & n22561;
  assign n27680 = ~pi2652 & ~n22561;
  assign n27681 = ~n27679 & ~n27680;
  assign n27682 = n22306 & ~n27681;
  assign n27683 = ~pi2652 & ~n22306;
  assign po2826 = n27682 | n27683;
  assign n27685 = pi3098 & n22311;
  assign n27686 = ~pi2653 & ~n22311;
  assign n27687 = ~n27685 & ~n27686;
  assign n27688 = n22306 & ~n27687;
  assign n27689 = ~pi2653 & ~n22306;
  assign po2827 = n27688 | n27689;
  assign n27691 = ~pi2654 & ~n22318;
  assign n27692 = pi3085 & n22318;
  assign n27693 = ~n27691 & ~n27692;
  assign n27694 = n22306 & ~n27693;
  assign n27695 = ~pi2654 & ~n22306;
  assign po2828 = n27694 | n27695;
  assign n27697 = ~pi2655 & ~n22318;
  assign n27698 = pi3045 & n22318;
  assign n27699 = ~n27697 & ~n27698;
  assign n27700 = n22306 & ~n27699;
  assign n27701 = ~pi2655 & ~n22306;
  assign po2829 = n27700 | n27701;
  assign n27703 = ~pi2656 & ~n22318;
  assign n27704 = pi3099 & n22318;
  assign n27705 = ~n27703 & ~n27704;
  assign n27706 = n22306 & ~n27705;
  assign n27707 = ~pi2656 & ~n22306;
  assign po2830 = n27706 | n27707;
  assign n27709 = ~pi2657 & ~n22318;
  assign n27710 = pi3101 & n22318;
  assign n27711 = ~n27709 & ~n27710;
  assign n27712 = n22306 & ~n27711;
  assign n27713 = ~pi2657 & ~n22306;
  assign po2831 = n27712 | n27713;
  assign n27715 = ~pi2658 & ~n22318;
  assign n27716 = pi3087 & n22318;
  assign n27717 = ~n27715 & ~n27716;
  assign n27718 = n22306 & ~n27717;
  assign n27719 = ~pi2658 & ~n22306;
  assign po2832 = n27718 | n27719;
  assign n27721 = ~pi2659 & ~n22318;
  assign n27722 = pi3050 & n22318;
  assign n27723 = ~n27721 & ~n27722;
  assign n27724 = n22306 & ~n27723;
  assign n27725 = ~pi2659 & ~n22306;
  assign po2833 = n27724 | n27725;
  assign n27727 = ~pi2660 & ~n22318;
  assign n27728 = pi3090 & n22318;
  assign n27729 = ~n27727 & ~n27728;
  assign n27730 = n22306 & ~n27729;
  assign n27731 = ~pi2660 & ~n22306;
  assign po2834 = n27730 | n27731;
  assign n27733 = ~pi2661 & ~n22318;
  assign n27734 = pi3092 & n22318;
  assign n27735 = ~n27733 & ~n27734;
  assign n27736 = n22306 & ~n27735;
  assign n27737 = ~pi2661 & ~n22306;
  assign po2835 = n27736 | n27737;
  assign n27739 = ~pi2662 & ~n22318;
  assign n27740 = pi3053 & n22318;
  assign n27741 = ~n27739 & ~n27740;
  assign n27742 = n22306 & ~n27741;
  assign n27743 = ~pi2662 & ~n22306;
  assign po2836 = n27742 | n27743;
  assign n27745 = ~pi2663 & ~n22318;
  assign n27746 = pi3054 & n22318;
  assign n27747 = ~n27745 & ~n27746;
  assign n27748 = n22306 & ~n27747;
  assign n27749 = ~pi2663 & ~n22306;
  assign po2837 = n27748 | n27749;
  assign n27751 = ~pi2664 & ~n22318;
  assign n27752 = pi3094 & n22318;
  assign n27753 = ~n27751 & ~n27752;
  assign n27754 = n22306 & ~n27753;
  assign n27755 = ~pi2664 & ~n22306;
  assign po2838 = n27754 | n27755;
  assign n27757 = ~pi2665 & ~n22547;
  assign n27758 = pi3086 & n22547;
  assign n27759 = ~n27757 & ~n27758;
  assign n27760 = n22306 & ~n27759;
  assign n27761 = ~pi2665 & ~n22306;
  assign po2839 = n27760 | n27761;
  assign n27763 = ~pi2666 & ~n22547;
  assign n27764 = pi3049 & n22547;
  assign n27765 = ~n27763 & ~n27764;
  assign n27766 = n22306 & ~n27765;
  assign n27767 = ~pi2666 & ~n22306;
  assign po2840 = n27766 | n27767;
  assign n27769 = ~pi2667 & ~n22547;
  assign n27770 = pi3060 & n22547;
  assign n27771 = ~n27769 & ~n27770;
  assign n27772 = n22306 & ~n27771;
  assign n27773 = ~pi2667 & ~n22306;
  assign po2841 = n27772 | n27773;
  assign n27775 = ~pi2668 & ~n22547;
  assign n27776 = pi3050 & n22547;
  assign n27777 = ~n27775 & ~n27776;
  assign n27778 = n22306 & ~n27777;
  assign n27779 = ~pi2668 & ~n22306;
  assign po2842 = n27778 | n27779;
  assign n27781 = ~pi2669 & ~n22547;
  assign n27782 = pi3056 & n22547;
  assign n27783 = ~n27781 & ~n27782;
  assign n27784 = n22306 & ~n27783;
  assign n27785 = ~pi2669 & ~n22306;
  assign po2843 = n27784 | n27785;
  assign n27787 = ~pi2670 & ~n22547;
  assign n27788 = pi3055 & n22547;
  assign n27789 = ~n27787 & ~n27788;
  assign n27790 = n22306 & ~n27789;
  assign n27791 = ~pi2670 & ~n22306;
  assign po2844 = n27790 | n27791;
  assign n27793 = ~pi2671 & ~n22547;
  assign n27794 = pi3054 & n22547;
  assign n27795 = ~n27793 & ~n27794;
  assign n27796 = n22306 & ~n27795;
  assign n27797 = ~pi2671 & ~n22306;
  assign po2845 = n27796 | n27797;
  assign n27799 = ~pi2672 & ~n22547;
  assign n27800 = pi3052 & n22547;
  assign n27801 = ~n27799 & ~n27800;
  assign n27802 = n22306 & ~n27801;
  assign n27803 = ~pi2672 & ~n22306;
  assign po2846 = n27802 | n27803;
  assign n27805 = ~pi2673 & ~n22539;
  assign n27806 = pi3084 & n22539;
  assign n27807 = ~n27805 & ~n27806;
  assign n27808 = n22306 & ~n27807;
  assign n27809 = ~pi2673 & ~n22306;
  assign po2847 = n27808 | n27809;
  assign n27811 = ~pi2674 & ~n22539;
  assign n27812 = pi3098 & n22539;
  assign n27813 = ~n27811 & ~n27812;
  assign n27814 = n22306 & ~n27813;
  assign n27815 = ~pi2674 & ~n22306;
  assign po2848 = n27814 | n27815;
  assign n27817 = ~pi2675 & ~n22539;
  assign n27818 = pi3095 & n22539;
  assign n27819 = ~n27817 & ~n27818;
  assign n27820 = n22306 & ~n27819;
  assign n27821 = ~pi2675 & ~n22306;
  assign po2849 = n27820 | n27821;
  assign n27823 = ~pi2676 & ~n22539;
  assign n27824 = pi3087 & n22539;
  assign n27825 = ~n27823 & ~n27824;
  assign n27826 = n22306 & ~n27825;
  assign n27827 = ~pi2676 & ~n22306;
  assign po2850 = n27826 | n27827;
  assign n27829 = ~pi2677 & ~n22539;
  assign n27830 = pi3088 & n22539;
  assign n27831 = ~n27829 & ~n27830;
  assign n27832 = n22306 & ~n27831;
  assign n27833 = ~pi2677 & ~n22306;
  assign po2851 = n27832 | n27833;
  assign n27835 = ~pi2678 & ~n22539;
  assign n27836 = pi3089 & n22539;
  assign n27837 = ~n27835 & ~n27836;
  assign n27838 = n22306 & ~n27837;
  assign n27839 = ~pi2678 & ~n22306;
  assign po2852 = n27838 | n27839;
  assign n27841 = ~pi2679 & ~n22539;
  assign n27842 = pi3052 & n22539;
  assign n27843 = ~n27841 & ~n27842;
  assign n27844 = n22306 & ~n27843;
  assign n27845 = ~pi2679 & ~n22306;
  assign po2853 = n27844 | n27845;
  assign n27847 = ~pi2680 & ~n22326;
  assign n27848 = pi3085 & n22326;
  assign n27849 = ~n27847 & ~n27848;
  assign n27850 = n22306 & ~n27849;
  assign n27851 = ~pi2680 & ~n22306;
  assign po2854 = n27850 | n27851;
  assign n27853 = ~pi2681 & ~n22326;
  assign n27854 = pi3047 & n22326;
  assign n27855 = ~n27853 & ~n27854;
  assign n27856 = n22306 & ~n27855;
  assign n27857 = ~pi2681 & ~n22306;
  assign po2855 = n27856 | n27857;
  assign n27859 = ~pi2682 & ~n22326;
  assign n27860 = pi3097 & n22326;
  assign n27861 = ~n27859 & ~n27860;
  assign n27862 = n22306 & ~n27861;
  assign n27863 = ~pi2682 & ~n22306;
  assign po2856 = n27862 | n27863;
  assign n27865 = ~pi2683 & ~n22326;
  assign n27866 = pi3050 & n22326;
  assign n27867 = ~n27865 & ~n27866;
  assign n27868 = n22306 & ~n27867;
  assign n27869 = ~pi2683 & ~n22306;
  assign po2857 = n27868 | n27869;
  assign n27871 = ~pi2684 & ~n22326;
  assign n27872 = pi3090 & n22326;
  assign n27873 = ~n27871 & ~n27872;
  assign n27874 = n22306 & ~n27873;
  assign n27875 = ~pi2684 & ~n22306;
  assign po2858 = n27874 | n27875;
  assign n27877 = ~pi2685 & ~n22318;
  assign n27878 = pi3061 & n22318;
  assign n27879 = ~n27877 & ~n27878;
  assign n27880 = n22306 & ~n27879;
  assign n27881 = ~pi2685 & ~n22306;
  assign po2859 = n27880 | n27881;
  assign n27883 = ~pi2686 & ~n22318;
  assign n27884 = pi3056 & n22318;
  assign n27885 = ~n27883 & ~n27884;
  assign n27886 = n22306 & ~n27885;
  assign n27887 = ~pi2686 & ~n22306;
  assign po2860 = n27886 | n27887;
  assign n27889 = ~pi2687 & ~n22326;
  assign n27890 = pi3048 & n22326;
  assign n27891 = ~n27889 & ~n27890;
  assign n27892 = n22306 & ~n27891;
  assign n27893 = ~pi2687 & ~n22306;
  assign po2861 = n27892 | n27893;
  assign n27895 = ~pi2688 & ~n22326;
  assign n27896 = pi3059 & n22326;
  assign n27897 = ~n27895 & ~n27896;
  assign n27898 = n22306 & ~n27897;
  assign n27899 = ~pi2688 & ~n22306;
  assign po2862 = n27898 | n27899;
  assign n27901 = pi3103 & n22561;
  assign n27902 = ~pi2689 & ~n22561;
  assign n27903 = ~n27901 & ~n27902;
  assign n27904 = n22306 & ~n27903;
  assign n27905 = ~pi2689 & ~n22306;
  assign po2863 = n27904 | n27905;
  assign n27907 = pi3103 & n22302;
  assign n27908 = ~pi2690 & ~n22302;
  assign n27909 = ~n27907 & ~n27908;
  assign n27910 = n22306 & ~n27909;
  assign n27911 = ~pi2690 & ~n22306;
  assign po2864 = n27910 | n27911;
  assign n27913 = ~pi2691 & ~n22318;
  assign n27914 = pi3103 & n22318;
  assign n27915 = ~n27913 & ~n27914;
  assign n27916 = n22306 & ~n27915;
  assign n27917 = ~pi2691 & ~n22306;
  assign po2865 = n27916 | n27917;
  assign n27919 = ~pi2692 & ~n22547;
  assign n27920 = pi3103 & n22547;
  assign n27921 = ~n27919 & ~n27920;
  assign n27922 = n22306 & ~n27921;
  assign n27923 = ~pi2692 & ~n22306;
  assign po2866 = n27922 | n27923;
  assign n27925 = ~pi2693 & ~n22539;
  assign n27926 = pi3045 & n22539;
  assign n27927 = ~n27925 & ~n27926;
  assign n27928 = n22306 & ~n27927;
  assign n27929 = ~pi2693 & ~n22306;
  assign po2867 = n27928 | n27929;
  assign n27931 = pi3061 & n22561;
  assign n27932 = ~pi2694 & ~n22561;
  assign n27933 = ~n27931 & ~n27932;
  assign n27934 = n22306 & ~n27933;
  assign n27935 = ~pi2694 & ~n22306;
  assign po2868 = n27934 | n27935;
  assign n27937 = pi3045 & n22311;
  assign n27938 = ~pi2695 & ~n22311;
  assign n27939 = ~n27937 & ~n27938;
  assign n27940 = n22306 & ~n27939;
  assign n27941 = ~pi2695 & ~n22306;
  assign po2869 = n27940 | n27941;
  assign n27943 = pi3100 & n22311;
  assign n27944 = ~pi2696 & ~n22311;
  assign n27945 = ~n27943 & ~n27944;
  assign n27946 = n22306 & ~n27945;
  assign n27947 = ~pi2696 & ~n22306;
  assign po2870 = n27946 | n27947;
  assign n27949 = pi3087 & n22561;
  assign n27950 = ~pi2697 & ~n22561;
  assign n27951 = ~n27949 & ~n27950;
  assign n27952 = n22306 & ~n27951;
  assign n27953 = ~pi2697 & ~n22306;
  assign po2871 = n27952 | n27953;
  assign n27955 = pi3099 & n22311;
  assign n27956 = ~pi2698 & ~n22311;
  assign n27957 = ~n27955 & ~n27956;
  assign n27958 = n22306 & ~n27957;
  assign n27959 = ~pi2698 & ~n22306;
  assign po2872 = n27958 | n27959;
  assign n27961 = pi3049 & n22561;
  assign n27962 = ~pi2699 & ~n22561;
  assign n27963 = ~n27961 & ~n27962;
  assign n27964 = n22306 & ~n27963;
  assign n27965 = ~pi2699 & ~n22306;
  assign po2873 = n27964 | n27965;
  assign n27967 = pi3089 & n22311;
  assign n27968 = ~pi2700 & ~n22311;
  assign n27969 = ~n27967 & ~n27968;
  assign n27970 = n22306 & ~n27969;
  assign n27971 = ~pi2700 & ~n22306;
  assign po2874 = n27970 | n27971;
  assign n27973 = pi3062 & n22554;
  assign n27974 = ~pi2701 & ~n22554;
  assign n27975 = ~n27973 & ~n27974;
  assign n27976 = n22306 & ~n27975;
  assign n27977 = ~pi2701 & ~n22306;
  assign po2875 = n27976 | n27977;
  assign n27979 = pi3098 & n22561;
  assign n27980 = ~pi2702 & ~n22561;
  assign n27981 = ~n27979 & ~n27980;
  assign n27982 = n22306 & ~n27981;
  assign n27983 = ~pi2702 & ~n22306;
  assign po2876 = n27982 | n27983;
  assign n27985 = pi3095 & n22554;
  assign n27986 = ~pi2703 & ~n22554;
  assign n27987 = ~n27985 & ~n27986;
  assign n27988 = n22306 & ~n27987;
  assign n27989 = ~pi2703 & ~n22306;
  assign po2877 = n27988 | n27989;
  assign n27991 = pi3061 & n22554;
  assign n27992 = ~pi2704 & ~n22554;
  assign n27993 = ~n27991 & ~n27992;
  assign n27994 = n22306 & ~n27993;
  assign n27995 = ~pi2704 & ~n22306;
  assign po2878 = n27994 | n27995;
  assign n27997 = pi1336 & n20262;
  assign n27998 = pi2705 & ~n20262;
  assign po2879 = n27997 | n27998;
  assign n28000 = pi3055 & n22302;
  assign n28001 = ~pi2706 & ~n22302;
  assign n28002 = ~n28000 & ~n28001;
  assign n28003 = n22306 & ~n28002;
  assign n28004 = ~pi2706 & ~n22306;
  assign po2880 = n28003 | n28004;
  assign n28006 = pi3050 & n22561;
  assign n28007 = ~pi2707 & ~n22561;
  assign n28008 = ~n28006 & ~n28007;
  assign n28009 = n22306 & ~n28008;
  assign n28010 = ~pi2707 & ~n22306;
  assign po2881 = n28009 | n28010;
  assign n28012 = pi3054 & n22554;
  assign n28013 = ~pi2708 & ~n22554;
  assign n28014 = ~n28012 & ~n28013;
  assign n28015 = n22306 & ~n28014;
  assign n28016 = ~pi2708 & ~n22306;
  assign po2882 = n28015 | n28016;
  assign n28018 = pi3048 & n22311;
  assign n28019 = ~pi2709 & ~n22311;
  assign n28020 = ~n28018 & ~n28019;
  assign n28021 = n22306 & ~n28020;
  assign n28022 = ~pi2709 & ~n22306;
  assign po2883 = n28021 | n28022;
  assign n28024 = pi3093 & n22561;
  assign n28025 = ~pi2710 & ~n22561;
  assign n28026 = ~n28024 & ~n28025;
  assign n28027 = n22306 & ~n28026;
  assign n28028 = ~pi2710 & ~n22306;
  assign po2884 = n28027 | n28028;
  assign n28030 = pi3054 & n22561;
  assign n28031 = ~pi2711 & ~n22561;
  assign n28032 = ~n28030 & ~n28031;
  assign n28033 = n22306 & ~n28032;
  assign n28034 = ~pi2711 & ~n22306;
  assign po2885 = n28033 | n28034;
  assign n28036 = pi3054 & n22302;
  assign n28037 = ~pi2712 & ~n22302;
  assign n28038 = ~n28036 & ~n28037;
  assign n28039 = n22306 & ~n28038;
  assign n28040 = ~pi2712 & ~n22306;
  assign po2886 = n28039 | n28040;
  assign n28042 = pi3092 & n22561;
  assign n28043 = ~pi2713 & ~n22561;
  assign n28044 = ~n28042 & ~n28043;
  assign n28045 = n22306 & ~n28044;
  assign n28046 = ~pi2713 & ~n22306;
  assign po2887 = n28045 | n28046;
  assign n28048 = pi3052 & n22554;
  assign n28049 = ~pi2714 & ~n22554;
  assign n28050 = ~n28048 & ~n28049;
  assign n28051 = n22306 & ~n28050;
  assign n28052 = ~pi2714 & ~n22306;
  assign po2888 = n28051 | n28052;
  assign n28054 = pi3088 & n22311;
  assign n28055 = ~pi2715 & ~n22311;
  assign n28056 = ~n28054 & ~n28055;
  assign n28057 = n22306 & ~n28056;
  assign n28058 = ~pi2715 & ~n22306;
  assign po2889 = n28057 | n28058;
  assign n28060 = ~pi2716 & ~n22318;
  assign n28061 = pi3060 & n22318;
  assign n28062 = ~n28060 & ~n28061;
  assign n28063 = n22306 & ~n28062;
  assign n28064 = ~pi2716 & ~n22306;
  assign po2890 = n28063 | n28064;
  assign n28066 = pi3053 & n22561;
  assign n28067 = ~pi2717 & ~n22561;
  assign n28068 = ~n28066 & ~n28067;
  assign n28069 = n22306 & ~n28068;
  assign n28070 = ~pi2717 & ~n22306;
  assign po2891 = n28069 | n28070;
  assign n28072 = pi3095 & n22302;
  assign n28073 = ~pi2718 & ~n22302;
  assign n28074 = ~n28072 & ~n28073;
  assign n28075 = n22306 & ~n28074;
  assign n28076 = ~pi2718 & ~n22306;
  assign po2892 = n28075 | n28076;
  assign n28078 = pi3054 & n22311;
  assign n28079 = ~pi2719 & ~n22311;
  assign n28080 = ~n28078 & ~n28079;
  assign n28081 = n22306 & ~n28080;
  assign n28082 = ~pi2719 & ~n22306;
  assign po2893 = n28081 | n28082;
  assign n28084 = pi3099 & n22561;
  assign n28085 = ~pi2720 & ~n22561;
  assign n28086 = ~n28084 & ~n28085;
  assign n28087 = n22306 & ~n28086;
  assign n28088 = ~pi2720 & ~n22306;
  assign po2894 = n28087 | n28088;
  assign n28090 = pi3058 & n22554;
  assign n28091 = ~pi2721 & ~n22554;
  assign n28092 = ~n28090 & ~n28091;
  assign n28093 = n22306 & ~n28092;
  assign n28094 = ~pi2721 & ~n22306;
  assign po2895 = n28093 | n28094;
  assign n28096 = pi3052 & n22311;
  assign n28097 = ~pi2722 & ~n22311;
  assign n28098 = ~n28096 & ~n28097;
  assign n28099 = n22306 & ~n28098;
  assign n28100 = ~pi2722 & ~n22306;
  assign po2896 = n28099 | n28100;
  assign n28102 = pi3085 & n22561;
  assign n28103 = ~pi2723 & ~n22561;
  assign n28104 = ~n28102 & ~n28103;
  assign n28105 = n22306 & ~n28104;
  assign n28106 = ~pi2723 & ~n22306;
  assign po2897 = n28105 | n28106;
  assign n28108 = pi3045 & n22561;
  assign n28109 = ~pi2724 & ~n22561;
  assign n28110 = ~n28108 & ~n28109;
  assign n28111 = n22306 & ~n28110;
  assign n28112 = ~pi2724 & ~n22306;
  assign po2898 = n28111 | n28112;
  assign n28114 = pi3095 & n22561;
  assign n28115 = ~pi2725 & ~n22561;
  assign n28116 = ~n28114 & ~n28115;
  assign n28117 = n22306 & ~n28116;
  assign n28118 = ~pi2725 & ~n22306;
  assign po2899 = n28117 | n28118;
  assign n28120 = pi3098 & n22302;
  assign n28121 = ~pi2726 & ~n22302;
  assign n28122 = ~n28120 & ~n28121;
  assign n28123 = n22306 & ~n28122;
  assign n28124 = ~pi2726 & ~n22306;
  assign po2900 = n28123 | n28124;
  assign n28126 = pi3087 & n22302;
  assign n28127 = ~pi2727 & ~n22302;
  assign n28128 = ~n28126 & ~n28127;
  assign n28129 = n22306 & ~n28128;
  assign n28130 = ~pi2727 & ~n22306;
  assign po2901 = n28129 | n28130;
  assign n28132 = pi3053 & n22302;
  assign n28133 = ~pi2728 & ~n22302;
  assign n28134 = ~n28132 & ~n28133;
  assign n28135 = n22306 & ~n28134;
  assign n28136 = ~pi2728 & ~n22306;
  assign po2902 = n28135 | n28136;
  assign n28138 = pi3092 & n22302;
  assign n28139 = ~pi2729 & ~n22302;
  assign n28140 = ~n28138 & ~n28139;
  assign n28141 = n22306 & ~n28140;
  assign n28142 = ~pi2729 & ~n22306;
  assign po2903 = n28141 | n28142;
  assign n28144 = pi3055 & n22554;
  assign n28145 = ~pi2730 & ~n22554;
  assign n28146 = ~n28144 & ~n28145;
  assign n28147 = n22306 & ~n28146;
  assign n28148 = ~pi2730 & ~n22306;
  assign po2904 = n28147 | n28148;
  assign n28150 = pi3090 & n22302;
  assign n28151 = ~pi2731 & ~n22302;
  assign n28152 = ~n28150 & ~n28151;
  assign n28153 = n22306 & ~n28152;
  assign n28154 = ~pi2731 & ~n22306;
  assign po2905 = n28153 | n28154;
  assign n28156 = pi3096 & n22302;
  assign n28157 = ~pi2732 & ~n22302;
  assign n28158 = ~n28156 & ~n28157;
  assign n28159 = n22306 & ~n28158;
  assign n28160 = ~pi2732 & ~n22306;
  assign po2906 = n28159 | n28160;
  assign n28162 = pi0171 & n20262;
  assign n28163 = pi2733 & ~n20262;
  assign po2907 = n28162 | n28163;
  assign n28165 = pi3050 & n22302;
  assign n28166 = ~pi2734 & ~n22302;
  assign n28167 = ~n28165 & ~n28166;
  assign n28168 = n22306 & ~n28167;
  assign n28169 = ~pi2734 & ~n22306;
  assign po2908 = n28168 | n28169;
  assign n28171 = pi3056 & n22302;
  assign n28172 = ~pi2735 & ~n22302;
  assign n28173 = ~n28171 & ~n28172;
  assign n28174 = n22306 & ~n28173;
  assign n28175 = ~pi2735 & ~n22306;
  assign po2909 = n28174 | n28175;
  assign n28177 = pi0307 & n20262;
  assign n28178 = pi2736 & ~n20262;
  assign po2910 = n28177 | n28178;
  assign n28180 = pi0306 & n20262;
  assign n28181 = pi2737 & ~n20262;
  assign po2911 = n28180 | n28181;
  assign n28183 = pi0305 & n20262;
  assign n28184 = pi2738 & ~n20262;
  assign po2912 = n28183 | n28184;
  assign n28186 = ~pi2739 & ~n22318;
  assign n28187 = pi3062 & n22318;
  assign n28188 = ~n28186 & ~n28187;
  assign n28189 = n22306 & ~n28188;
  assign n28190 = ~pi2739 & ~n22306;
  assign po2913 = n28189 | n28190;
  assign n28192 = ~pi2740 & ~n22547;
  assign n28193 = pi3092 & n22547;
  assign n28194 = ~n28192 & ~n28193;
  assign n28195 = n22306 & ~n28194;
  assign n28196 = ~pi2740 & ~n22306;
  assign po2914 = n28195 | n28196;
  assign n28198 = ~pi2741 & ~n22318;
  assign n28199 = pi3084 & n22318;
  assign n28200 = ~n28198 & ~n28199;
  assign n28201 = n22306 & ~n28200;
  assign n28202 = ~pi2741 & ~n22306;
  assign po2915 = n28201 | n28202;
  assign n28204 = ~pi2742 & ~n22547;
  assign n28205 = pi3094 & n22547;
  assign n28206 = ~n28204 & ~n28205;
  assign n28207 = n22306 & ~n28206;
  assign n28208 = ~pi2742 & ~n22306;
  assign po2916 = n28207 | n28208;
  assign n28210 = ~pi2743 & ~n22547;
  assign n28211 = pi3053 & n22547;
  assign n28212 = ~n28210 & ~n28211;
  assign n28213 = n22306 & ~n28212;
  assign n28214 = ~pi2743 & ~n22306;
  assign po2917 = n28213 | n28214;
  assign n28216 = ~pi2744 & ~n22326;
  assign n28217 = pi3056 & n22326;
  assign n28218 = ~n28216 & ~n28217;
  assign n28219 = n22306 & ~n28218;
  assign n28220 = ~pi2744 & ~n22306;
  assign po2918 = n28219 | n28220;
  assign n28222 = ~pi2745 & ~n22539;
  assign n28223 = pi3085 & n22539;
  assign n28224 = ~n28222 & ~n28223;
  assign n28225 = n22306 & ~n28224;
  assign n28226 = ~pi2745 & ~n22306;
  assign po2919 = n28225 | n28226;
  assign n28228 = ~pi2746 & ~n22547;
  assign n28229 = pi3089 & n22547;
  assign n28230 = ~n28228 & ~n28229;
  assign n28231 = n22306 & ~n28230;
  assign n28232 = ~pi2746 & ~n22306;
  assign po2920 = n28231 | n28232;
  assign n28234 = ~pi2747 & ~n22547;
  assign n28235 = pi3093 & n22547;
  assign n28236 = ~n28234 & ~n28235;
  assign n28237 = n22306 & ~n28236;
  assign n28238 = ~pi2747 & ~n22306;
  assign po2921 = n28237 | n28238;
  assign n28240 = pi3086 & n22302;
  assign n28241 = ~pi2748 & ~n22302;
  assign n28242 = ~n28240 & ~n28241;
  assign n28243 = n22306 & ~n28242;
  assign n28244 = ~pi2748 & ~n22306;
  assign po2922 = n28243 | n28244;
  assign n28246 = pi0174 & n20262;
  assign n28247 = pi2749 & ~n20262;
  assign po2923 = n28246 | n28247;
  assign n28249 = ~pi2750 & ~n22539;
  assign n28250 = pi3053 & n22539;
  assign n28251 = ~n28249 & ~n28250;
  assign n28252 = n22306 & ~n28251;
  assign n28253 = ~pi2750 & ~n22306;
  assign po2924 = n28252 | n28253;
  assign n28255 = ~pi2751 & ~n22547;
  assign n28256 = pi3096 & n22547;
  assign n28257 = ~n28255 & ~n28256;
  assign n28258 = n22306 & ~n28257;
  assign n28259 = ~pi2751 & ~n22306;
  assign po2925 = n28258 | n28259;
  assign n28261 = pi0026 & ~n23715;
  assign n28262 = pi2752 & n23715;
  assign po2926 = n28261 | n28262;
  assign n28264 = ~pi2753 & ~n22547;
  assign n28265 = pi3048 & n22547;
  assign n28266 = ~n28264 & ~n28265;
  assign n28267 = n22306 & ~n28266;
  assign n28268 = ~pi2753 & ~n22306;
  assign po2927 = n28267 | n28268;
  assign n28270 = ~pi2754 & ~n22539;
  assign n28271 = pi3096 & n22539;
  assign n28272 = ~n28270 & ~n28271;
  assign n28273 = n22306 & ~n28272;
  assign n28274 = ~pi2754 & ~n22306;
  assign po2928 = n28273 | n28274;
  assign n28276 = n10695 & ~n10704;
  assign n28277 = n20262 & n28276;
  assign n28278 = pi2755 & ~n20262;
  assign po2929 = n28277 | n28278;
  assign n28280 = ~pi2756 & ~n22326;
  assign n28281 = pi3060 & n22326;
  assign n28282 = ~n28280 & ~n28281;
  assign n28283 = n22306 & ~n28282;
  assign n28284 = ~pi2756 & ~n22306;
  assign po2930 = n28283 | n28284;
  assign n28286 = pi1705 & n22080;
  assign n28287 = n19465 & n25396;
  assign n28288 = pi2757 & ~n28287;
  assign n28289 = ~pi2757 & n28287;
  assign n28290 = ~n28288 & ~n28289;
  assign n28291 = n23726 & ~n28290;
  assign n28292 = pi2757 & ~n23726;
  assign n28293 = ~n28291 & ~n28292;
  assign n28294 = ~n22080 & ~n28293;
  assign po2931 = n28286 | n28294;
  assign n28296 = pi2758 & ~n8009;
  assign po2932 = n27209 | n28296;
  assign n28298 = ~pi2759 & ~n22547;
  assign n28299 = pi3091 & n22547;
  assign n28300 = ~n28298 & ~n28299;
  assign n28301 = n22306 & ~n28300;
  assign n28302 = ~pi2759 & ~n22306;
  assign po2933 = n28301 | n28302;
  assign n28304 = pi0032 & ~n23715;
  assign n28305 = pi2760 & n23715;
  assign po2934 = n28304 | n28305;
  assign n28307 = pi0034 & ~n23715;
  assign n28308 = pi2761 & n23715;
  assign po2935 = n28307 | n28308;
  assign n28310 = pi0033 & ~n23715;
  assign n28311 = pi2762 & n23715;
  assign po2936 = n28310 | n28311;
  assign n28313 = ~pi2763 & ~n22326;
  assign n28314 = pi3045 & n22326;
  assign n28315 = ~n28313 & ~n28314;
  assign n28316 = n22306 & ~n28315;
  assign n28317 = ~pi2763 & ~n22306;
  assign po2937 = n28316 | n28317;
  assign n28319 = ~pi2764 & ~n22539;
  assign n28320 = pi3049 & n22539;
  assign n28321 = ~n28319 & ~n28320;
  assign n28322 = n22306 & ~n28321;
  assign n28323 = ~pi2764 & ~n22306;
  assign po2938 = n28322 | n28323;
  assign n28325 = pi0030 & ~n23715;
  assign n28326 = pi2765 & n23715;
  assign po2939 = n28325 | n28326;
  assign n28328 = pi0031 & ~n23715;
  assign n28329 = pi2766 & n23715;
  assign po2940 = n28328 | n28329;
  assign n28331 = pi0029 & ~n23715;
  assign n28332 = pi2767 & n23715;
  assign po2941 = n28331 | n28332;
  assign n28334 = ~pi2768 & ~n22539;
  assign n28335 = pi3054 & n22539;
  assign n28336 = ~n28334 & ~n28335;
  assign n28337 = n22306 & ~n28336;
  assign n28338 = ~pi2768 & ~n22306;
  assign po2942 = n28337 | n28338;
  assign n28340 = ~pi2769 & ~n22547;
  assign n28341 = pi3090 & n22547;
  assign n28342 = ~n28340 & ~n28341;
  assign n28343 = n22306 & ~n28342;
  assign n28344 = ~pi2769 & ~n22306;
  assign po2943 = n28343 | n28344;
  assign n28346 = ~pi2770 & ~n22547;
  assign n28347 = pi3058 & n22547;
  assign n28348 = ~n28346 & ~n28347;
  assign n28349 = n22306 & ~n28348;
  assign n28350 = ~pi2770 & ~n22306;
  assign po2944 = n28349 | n28350;
  assign n28352 = ~pi2771 & ~n22326;
  assign n28353 = pi3088 & n22326;
  assign n28354 = ~n28352 & ~n28353;
  assign n28355 = n22306 & ~n28354;
  assign n28356 = ~pi2771 & ~n22306;
  assign po2945 = n28355 | n28356;
  assign n28358 = ~pi2772 & ~n22326;
  assign n28359 = pi3053 & n22326;
  assign n28360 = ~n28358 & ~n28359;
  assign n28361 = n22306 & ~n28360;
  assign n28362 = ~pi2772 & ~n22306;
  assign po2946 = n28361 | n28362;
  assign n28364 = ~pi2773 & ~n22547;
  assign n28365 = pi3059 & n22547;
  assign n28366 = ~n28364 & ~n28365;
  assign n28367 = n22306 & ~n28366;
  assign n28368 = ~pi2773 & ~n22306;
  assign po2947 = n28367 | n28368;
  assign n28370 = ~pi2774 & ~n22326;
  assign n28371 = pi3094 & n22326;
  assign n28372 = ~n28370 & ~n28371;
  assign n28373 = n22306 & ~n28372;
  assign n28374 = ~pi2774 & ~n22306;
  assign po2948 = n28373 | n28374;
  assign n28376 = ~pi2775 & ~n22539;
  assign n28377 = pi3097 & n22539;
  assign n28378 = ~n28376 & ~n28377;
  assign n28379 = n22306 & ~n28378;
  assign n28380 = ~pi2775 & ~n22306;
  assign po2949 = n28379 | n28380;
  assign n28382 = ~pi2776 & ~n22318;
  assign n28383 = pi3059 & n22318;
  assign n28384 = ~n28382 & ~n28383;
  assign n28385 = n22306 & ~n28384;
  assign n28386 = ~pi2776 & ~n22306;
  assign po2950 = n28385 | n28386;
  assign n28388 = ~pi2777 & ~n22318;
  assign n28389 = pi3096 & n22318;
  assign n28390 = ~n28388 & ~n28389;
  assign n28391 = n22306 & ~n28390;
  assign n28392 = ~pi2777 & ~n22306;
  assign po2951 = n28391 | n28392;
  assign n28394 = pi3056 & n22554;
  assign n28395 = ~pi2778 & ~n22554;
  assign n28396 = ~n28394 & ~n28395;
  assign n28397 = n22306 & ~n28396;
  assign n28398 = ~pi2778 & ~n22306;
  assign po2952 = n28397 | n28398;
  assign n28400 = pi0019 & ~n23715;
  assign n28401 = pi2779 & n23715;
  assign po2953 = n28400 | n28401;
  assign n28403 = pi3059 & n22561;
  assign n28404 = ~pi2780 & ~n22561;
  assign n28405 = ~n28403 & ~n28404;
  assign n28406 = n22306 & ~n28405;
  assign n28407 = ~pi2780 & ~n22306;
  assign po2954 = n28406 | n28407;
  assign n28409 = pi3100 & n22561;
  assign n28410 = ~pi2781 & ~n22561;
  assign n28411 = ~n28409 & ~n28410;
  assign n28412 = n22306 & ~n28411;
  assign n28413 = ~pi2781 & ~n22306;
  assign po2955 = n28412 | n28413;
  assign n28415 = ~pi2782 & ~n22547;
  assign n28416 = pi3088 & n22547;
  assign n28417 = ~n28415 & ~n28416;
  assign n28418 = n22306 & ~n28417;
  assign n28419 = ~pi2782 & ~n22306;
  assign po2956 = n28418 | n28419;
  assign n28421 = ~pi2783 & ~n22326;
  assign n28422 = pi3093 & n22326;
  assign n28423 = ~n28421 & ~n28422;
  assign n28424 = n22306 & ~n28423;
  assign n28425 = ~pi2783 & ~n22306;
  assign po2957 = n28424 | n28425;
  assign n28427 = pi3084 & n22302;
  assign n28428 = ~pi2784 & ~n22302;
  assign n28429 = ~n28427 & ~n28428;
  assign n28430 = n22306 & ~n28429;
  assign n28431 = ~pi2784 & ~n22306;
  assign po2958 = n28430 | n28431;
  assign n28433 = pi3096 & n22554;
  assign n28434 = ~pi2785 & ~n22554;
  assign n28435 = ~n28433 & ~n28434;
  assign n28436 = n22306 & ~n28435;
  assign n28437 = ~pi2785 & ~n22306;
  assign po2959 = n28436 | n28437;
  assign n28439 = pi3090 & n22554;
  assign n28440 = ~pi2786 & ~n22554;
  assign n28441 = ~n28439 & ~n28440;
  assign n28442 = n22306 & ~n28441;
  assign n28443 = ~pi2786 & ~n22306;
  assign po2960 = n28442 | n28443;
  assign n28445 = pi0300 & n20262;
  assign n28446 = pi2787 & ~n20262;
  assign po2961 = n28445 | n28446;
  assign n28448 = ~pi2788 & ~n22547;
  assign n28449 = pi3100 & n22547;
  assign n28450 = ~n28448 & ~n28449;
  assign n28451 = n22306 & ~n28450;
  assign n28452 = ~pi2788 & ~n22306;
  assign po2962 = n28451 | n28452;
  assign n28454 = ~pi2789 & ~n22326;
  assign n28455 = pi3095 & n22326;
  assign n28456 = ~n28454 & ~n28455;
  assign n28457 = n22306 & ~n28456;
  assign n28458 = ~pi2789 & ~n22306;
  assign po2963 = n28457 | n28458;
  assign n28460 = ~pi2790 & ~n22326;
  assign n28461 = pi3054 & n22326;
  assign n28462 = ~n28460 & ~n28461;
  assign n28463 = n22306 & ~n28462;
  assign n28464 = ~pi2790 & ~n22306;
  assign po2964 = n28463 | n28464;
  assign n28466 = ~pi2791 & ~n22547;
  assign n28467 = pi3097 & n22547;
  assign n28468 = ~n28466 & ~n28467;
  assign n28469 = n22306 & ~n28468;
  assign n28470 = ~pi2791 & ~n22306;
  assign po2965 = n28469 | n28470;
  assign n28472 = ~pi2792 & ~n22326;
  assign n28473 = pi3052 & n22326;
  assign n28474 = ~n28472 & ~n28473;
  assign n28475 = n22306 & ~n28474;
  assign n28476 = ~pi2792 & ~n22306;
  assign po2966 = n28475 | n28476;
  assign n28478 = ~pi2793 & ~n22547;
  assign n28479 = pi3101 & n22547;
  assign n28480 = ~n28478 & ~n28479;
  assign n28481 = n22306 & ~n28480;
  assign n28482 = ~pi2793 & ~n22306;
  assign po2967 = n28481 | n28482;
  assign n28484 = ~pi2794 & ~n22326;
  assign n28485 = pi3096 & n22326;
  assign n28486 = ~n28484 & ~n28485;
  assign n28487 = n22306 & ~n28486;
  assign n28488 = ~pi2794 & ~n22306;
  assign po2968 = n28487 | n28488;
  assign n28490 = pi0020 & ~n23715;
  assign n28491 = pi2795 & n23715;
  assign po2969 = n28490 | n28491;
  assign n28493 = ~pi2796 & ~n22318;
  assign n28494 = pi3055 & n22318;
  assign n28495 = ~n28493 & ~n28494;
  assign n28496 = n22306 & ~n28495;
  assign n28497 = ~pi2796 & ~n22306;
  assign po2970 = n28496 | n28497;
  assign n28499 = ~pi2797 & ~n22318;
  assign n28500 = pi3095 & n22318;
  assign n28501 = ~n28499 & ~n28500;
  assign n28502 = n22306 & ~n28501;
  assign n28503 = ~pi2797 & ~n22306;
  assign po2971 = n28502 | n28503;
  assign n28505 = ~pi2798 & ~n22547;
  assign n28506 = pi3061 & n22547;
  assign n28507 = ~n28505 & ~n28506;
  assign n28508 = n22306 & ~n28507;
  assign n28509 = ~pi2798 & ~n22306;
  assign po2972 = n28508 | n28509;
  assign n28511 = ~pi2799 & ~n22547;
  assign n28512 = pi3047 & n22547;
  assign n28513 = ~n28511 & ~n28512;
  assign n28514 = n22306 & ~n28513;
  assign n28515 = ~pi2799 & ~n22306;
  assign po2973 = n28514 | n28515;
  assign n28517 = ~pi2800 & ~n22547;
  assign n28518 = pi3087 & n22547;
  assign n28519 = ~n28517 & ~n28518;
  assign n28520 = n22306 & ~n28519;
  assign n28521 = ~pi2800 & ~n22306;
  assign po2974 = n28520 | n28521;
  assign n28523 = ~pi2801 & ~n22326;
  assign n28524 = pi3055 & n22326;
  assign n28525 = ~n28523 & ~n28524;
  assign n28526 = n22306 & ~n28525;
  assign n28527 = ~pi2801 & ~n22306;
  assign po2975 = n28526 | n28527;
  assign n28529 = ~pi2802 & ~n22547;
  assign n28530 = pi3084 & n22547;
  assign n28531 = ~n28529 & ~n28530;
  assign n28532 = n22306 & ~n28531;
  assign n28533 = ~pi2802 & ~n22306;
  assign po2976 = n28532 | n28533;
  assign n28535 = ~pi2803 & ~n22326;
  assign n28536 = pi3099 & n22326;
  assign n28537 = ~n28535 & ~n28536;
  assign n28538 = n22306 & ~n28537;
  assign n28539 = ~pi2803 & ~n22306;
  assign po2977 = n28538 | n28539;
  assign n28541 = ~pi2804 & ~n22326;
  assign n28542 = pi3092 & n22326;
  assign n28543 = ~n28541 & ~n28542;
  assign n28544 = n22306 & ~n28543;
  assign n28545 = ~pi2804 & ~n22306;
  assign po2978 = n28544 | n28545;
  assign n28547 = ~pi2805 & ~n22547;
  assign n28548 = pi3099 & n22547;
  assign n28549 = ~n28547 & ~n28548;
  assign n28550 = n22306 & ~n28549;
  assign n28551 = ~pi2805 & ~n22306;
  assign po2979 = n28550 | n28551;
  assign n28553 = ~pi2806 & ~n22547;
  assign n28554 = pi3098 & n22547;
  assign n28555 = ~n28553 & ~n28554;
  assign n28556 = n22306 & ~n28555;
  assign n28557 = ~pi2806 & ~n22306;
  assign po2980 = n28556 | n28557;
  assign n28559 = ~pi2807 & ~n22326;
  assign n28560 = pi3091 & n22326;
  assign n28561 = ~n28559 & ~n28560;
  assign n28562 = n22306 & ~n28561;
  assign n28563 = ~pi2807 & ~n22306;
  assign po2981 = n28562 | n28563;
  assign n28565 = ~pi2808 & ~n22547;
  assign n28566 = pi3085 & n22547;
  assign n28567 = ~n28565 & ~n28566;
  assign n28568 = n22306 & ~n28567;
  assign n28569 = ~pi2808 & ~n22306;
  assign po2982 = n28568 | n28569;
  assign n28571 = ~pi2809 & ~n22547;
  assign n28572 = pi3062 & n22547;
  assign n28573 = ~n28571 & ~n28572;
  assign n28574 = n22306 & ~n28573;
  assign n28575 = ~pi2809 & ~n22306;
  assign po2983 = n28574 | n28575;
  assign n28577 = ~pi2810 & ~n22539;
  assign n28578 = pi3091 & n22539;
  assign n28579 = ~n28577 & ~n28578;
  assign n28580 = n22306 & ~n28579;
  assign n28581 = ~pi2810 & ~n22306;
  assign po2984 = n28580 | n28581;
  assign n28583 = ~pi2811 & ~n22547;
  assign n28584 = pi3045 & n22547;
  assign n28585 = ~n28583 & ~n28584;
  assign n28586 = n22306 & ~n28585;
  assign n28587 = ~pi2811 & ~n22306;
  assign po2985 = n28586 | n28587;
  assign n28589 = ~pi2812 & ~n22318;
  assign n28590 = pi3052 & n22318;
  assign n28591 = ~n28589 & ~n28590;
  assign n28592 = n22306 & ~n28591;
  assign n28593 = ~pi2812 & ~n22306;
  assign po2986 = n28592 | n28593;
  assign n28595 = ~pi2813 & ~n22326;
  assign n28596 = pi3087 & n22326;
  assign n28597 = ~n28595 & ~n28596;
  assign n28598 = n22306 & ~n28597;
  assign n28599 = ~pi2813 & ~n22306;
  assign po2987 = n28598 | n28599;
  assign n28601 = ~pi2814 & ~n22326;
  assign n28602 = pi3100 & n22326;
  assign n28603 = ~n28601 & ~n28602;
  assign n28604 = n22306 & ~n28603;
  assign n28605 = ~pi2814 & ~n22306;
  assign po2988 = n28604 | n28605;
  assign n28607 = ~pi2815 & ~n22326;
  assign n28608 = pi3101 & n22326;
  assign n28609 = ~n28607 & ~n28608;
  assign n28610 = n22306 & ~n28609;
  assign n28611 = ~pi2815 & ~n22306;
  assign po2989 = n28610 | n28611;
  assign n28613 = ~pi2816 & ~n22326;
  assign n28614 = pi3058 & n22326;
  assign n28615 = ~n28613 & ~n28614;
  assign n28616 = n22306 & ~n28615;
  assign n28617 = ~pi2816 & ~n22306;
  assign po2990 = n28616 | n28617;
  assign n28619 = ~pi2817 & ~n22318;
  assign n28620 = pi3093 & n22318;
  assign n28621 = ~n28619 & ~n28620;
  assign n28622 = n22306 & ~n28621;
  assign n28623 = ~pi2817 & ~n22306;
  assign po2991 = n28622 | n28623;
  assign n28625 = pi0022 & ~n23715;
  assign n28626 = pi2818 & n23715;
  assign po2992 = n28625 | n28626;
  assign n28628 = pi0023 & ~n23715;
  assign n28629 = pi2819 & n23715;
  assign po2993 = n28628 | n28629;
  assign n28631 = ~pi2820 & ~n22318;
  assign n28632 = pi3091 & n22318;
  assign n28633 = ~n28631 & ~n28632;
  assign n28634 = n22306 & ~n28633;
  assign n28635 = ~pi2820 & ~n22306;
  assign po2994 = n28634 | n28635;
  assign n28637 = ~pi2821 & ~n22539;
  assign n28638 = pi3048 & n22539;
  assign n28639 = ~n28637 & ~n28638;
  assign n28640 = n22306 & ~n28639;
  assign n28641 = ~pi2821 & ~n22306;
  assign po2995 = n28640 | n28641;
  assign n28643 = ~pi2822 & ~n22326;
  assign n28644 = pi3089 & n22326;
  assign n28645 = ~n28643 & ~n28644;
  assign n28646 = n22306 & ~n28645;
  assign n28647 = ~pi2822 & ~n22306;
  assign po2996 = n28646 | n28647;
  assign n28649 = ~pi2823 & ~n22318;
  assign n28650 = pi3048 & n22318;
  assign n28651 = ~n28649 & ~n28650;
  assign n28652 = n22306 & ~n28651;
  assign n28653 = ~pi2823 & ~n22306;
  assign po2997 = n28652 | n28653;
  assign n28655 = ~pi2824 & ~n22539;
  assign n28656 = pi3103 & n22539;
  assign n28657 = ~n28655 & ~n28656;
  assign n28658 = n22306 & ~n28657;
  assign n28659 = ~pi2824 & ~n22306;
  assign po2998 = n28658 | n28659;
  assign n28661 = pi3089 & n22561;
  assign n28662 = ~pi2825 & ~n22561;
  assign n28663 = ~n28661 & ~n28662;
  assign n28664 = n22306 & ~n28663;
  assign n28665 = ~pi2825 & ~n22306;
  assign po2999 = n28664 | n28665;
  assign n28667 = ~pi2826 & ~n22326;
  assign n28668 = pi3086 & n22326;
  assign n28669 = ~n28667 & ~n28668;
  assign n28670 = n22306 & ~n28669;
  assign n28671 = ~pi2826 & ~n22306;
  assign po3000 = n28670 | n28671;
  assign n28673 = pi3059 & n22554;
  assign n28674 = ~pi2827 & ~n22554;
  assign n28675 = ~n28673 & ~n28674;
  assign n28676 = n22306 & ~n28675;
  assign n28677 = ~pi2827 & ~n22306;
  assign po3001 = n28676 | n28677;
  assign n28679 = pi3050 & n22554;
  assign n28680 = ~pi2828 & ~n22554;
  assign n28681 = ~n28679 & ~n28680;
  assign n28682 = n22306 & ~n28681;
  assign n28683 = ~pi2828 & ~n22306;
  assign po3002 = n28682 | n28683;
  assign n28685 = pi3084 & n22554;
  assign n28686 = ~pi2829 & ~n22554;
  assign n28687 = ~n28685 & ~n28686;
  assign n28688 = n22306 & ~n28687;
  assign n28689 = ~pi2829 & ~n22306;
  assign po3003 = n28688 | n28689;
  assign n28691 = ~pi2830 & ~n22539;
  assign n28692 = pi3094 & n22539;
  assign n28693 = ~n28691 & ~n28692;
  assign n28694 = n22306 & ~n28693;
  assign n28695 = ~pi2830 & ~n22306;
  assign po3004 = n28694 | n28695;
  assign n28697 = pi3052 & n22302;
  assign n28698 = ~pi2831 & ~n22302;
  assign n28699 = ~n28697 & ~n28698;
  assign n28700 = n22306 & ~n28699;
  assign n28701 = ~pi2831 & ~n22306;
  assign po3005 = n28700 | n28701;
  assign n28703 = ~pi2832 & ~n22326;
  assign n28704 = pi3061 & n22326;
  assign n28705 = ~n28703 & ~n28704;
  assign n28706 = n22306 & ~n28705;
  assign n28707 = ~pi2832 & ~n22306;
  assign po3006 = n28706 | n28707;
  assign n28709 = ~pi2833 & ~n22539;
  assign n28710 = pi3061 & n22539;
  assign n28711 = ~n28709 & ~n28710;
  assign n28712 = n22306 & ~n28711;
  assign n28713 = ~pi2833 & ~n22306;
  assign po3007 = n28712 | n28713;
  assign n28715 = pi0068 & ~n23715;
  assign n28716 = pi2834 & n23715;
  assign po3008 = n28715 | n28716;
  assign n28718 = ~pi2835 & ~n22326;
  assign n28719 = pi3049 & n22326;
  assign n28720 = ~n28718 & ~n28719;
  assign n28721 = n22306 & ~n28720;
  assign n28722 = ~pi2835 & ~n22306;
  assign po3009 = n28721 | n28722;
  assign n28724 = ~pi2836 & ~n22326;
  assign n28725 = pi3103 & n22326;
  assign n28726 = ~n28724 & ~n28725;
  assign n28727 = n22306 & ~n28726;
  assign n28728 = ~pi2836 & ~n22306;
  assign po3010 = n28727 | n28728;
  assign n28730 = ~pi2837 & ~n22326;
  assign n28731 = pi3098 & n22326;
  assign n28732 = ~n28730 & ~n28731;
  assign n28733 = n22306 & ~n28732;
  assign n28734 = ~pi2837 & ~n22306;
  assign po3011 = n28733 | n28734;
  assign n28736 = pi0064 & ~n23715;
  assign n28737 = pi2838 & n23715;
  assign po3012 = n28736 | n28737;
  assign n28739 = ~pi2839 & ~n22326;
  assign n28740 = pi3062 & n22326;
  assign n28741 = ~n28739 & ~n28740;
  assign n28742 = n22306 & ~n28741;
  assign n28743 = ~pi2839 & ~n22306;
  assign po3013 = n28742 | n28743;
  assign n28745 = pi0036 & ~n23715;
  assign n28746 = pi2840 & n23715;
  assign po3014 = n28745 | n28746;
  assign n28748 = pi0015 & ~n23715;
  assign n28749 = pi2841 & n23715;
  assign po3015 = n28748 | n28749;
  assign n28751 = pi0016 & ~n23715;
  assign n28752 = pi2842 & n23715;
  assign po3016 = n28751 | n28752;
  assign n28754 = pi0018 & ~n23715;
  assign n28755 = pi2843 & n23715;
  assign po3017 = n28754 | n28755;
  assign n28757 = ~pi2844 & ~n22326;
  assign n28758 = pi3084 & n22326;
  assign n28759 = ~n28757 & ~n28758;
  assign n28760 = n22306 & ~n28759;
  assign n28761 = ~pi2844 & ~n22306;
  assign po3018 = n28760 | n28761;
  assign n28763 = pi0035 & ~n23715;
  assign n28764 = pi2845 & n23715;
  assign po3019 = n28763 | n28764;
  assign n28766 = ~pi0072 & ~n23715;
  assign n28767 = pi2846 & n23715;
  assign po3020 = n28766 | n28767;
  assign n28769 = pi0012 & ~n23715;
  assign n28770 = pi2847 & n23715;
  assign po3021 = n28769 | n28770;
  assign n28772 = ~pi0073 & ~n23715;
  assign n28773 = pi2848 & n23715;
  assign po3022 = n28772 | n28773;
  assign n28775 = pi0008 & ~n23715;
  assign n28776 = pi2849 & n23715;
  assign po3023 = n28775 | n28776;
  assign n28778 = pi0010 & ~n23715;
  assign n28779 = pi2850 & n23715;
  assign po3024 = n28778 | n28779;
  assign n28781 = ~pi0074 & ~n23715;
  assign n28782 = pi2851 & n23715;
  assign po3025 = n28781 | n28782;
  assign n28784 = ~pi0075 & ~n23715;
  assign n28785 = pi2852 & n23715;
  assign po3026 = n28784 | n28785;
  assign n28787 = pi0059 & ~n23715;
  assign n28788 = pi2853 & n23715;
  assign po3027 = n28787 | n28788;
  assign n28790 = pi0051 & ~n23715;
  assign n28791 = pi2854 & n23715;
  assign po3028 = n28790 | n28791;
  assign n28793 = ~pi2855 & ~n22539;
  assign n28794 = pi3093 & n22539;
  assign n28795 = ~n28793 & ~n28794;
  assign n28796 = n22306 & ~n28795;
  assign n28797 = ~pi2855 & ~n22306;
  assign po3029 = n28796 | n28797;
  assign n28799 = pi0269 & n20262;
  assign n28800 = pi2856 & ~n20262;
  assign po3030 = n28799 | n28800;
  assign n28802 = pi3103 & n22554;
  assign n28803 = ~pi2857 & ~n22554;
  assign n28804 = ~n28802 & ~n28803;
  assign n28805 = n22306 & ~n28804;
  assign n28806 = ~pi2857 & ~n22306;
  assign po3031 = n28805 | n28806;
  assign n28808 = pi0061 & ~n23715;
  assign n28809 = pi2858 & n23715;
  assign po3032 = n28808 | n28809;
  assign n28811 = pi0045 & ~n23715;
  assign n28812 = pi2859 & n23715;
  assign po3033 = n28811 | n28812;
  assign n28814 = pi3085 & n22554;
  assign n28815 = ~pi2860 & ~n22554;
  assign n28816 = ~n28814 & ~n28815;
  assign n28817 = n22306 & ~n28816;
  assign n28818 = ~pi2860 & ~n22306;
  assign po3034 = n28817 | n28818;
  assign n28820 = pi0043 & ~n23715;
  assign n28821 = pi2861 & n23715;
  assign po3035 = n28820 | n28821;
  assign n28823 = pi0049 & ~n23715;
  assign n28824 = pi2862 & n23715;
  assign po3036 = n28823 | n28824;
  assign n28826 = pi0046 & ~n23715;
  assign n28827 = pi2863 & n23715;
  assign po3037 = n28826 | n28827;
  assign n28829 = pi0070 & ~n23715;
  assign n28830 = pi2864 & n23715;
  assign po3038 = n28829 | n28830;
  assign n28832 = pi0057 & ~n23715;
  assign n28833 = pi2865 & n23715;
  assign po3039 = n28832 | n28833;
  assign n28835 = pi0041 & ~n23715;
  assign n28836 = pi2866 & n23715;
  assign po3040 = n28835 | n28836;
  assign n28838 = pi0044 & ~n23715;
  assign n28839 = pi2867 & n23715;
  assign po3041 = n28838 | n28839;
  assign n28841 = pi0056 & ~n23715;
  assign n28842 = pi2868 & n23715;
  assign po3042 = n28841 | n28842;
  assign n28844 = pi0066 & ~n23715;
  assign n28845 = pi2869 & n23715;
  assign po3043 = n28844 | n28845;
  assign n28847 = pi0050 & ~n23715;
  assign n28848 = pi2870 & n23715;
  assign po3044 = n28847 | n28848;
  assign n28850 = pi0055 & ~n23715;
  assign n28851 = pi2871 & n23715;
  assign po3045 = n28850 | n28851;
  assign n28853 = pi0054 & ~n23715;
  assign n28854 = pi2872 & n23715;
  assign po3046 = n28853 | n28854;
  assign n28856 = pi2873 & n23715;
  assign n28857 = ~pi0006 & ~n23715;
  assign po3047 = n28856 | n28857;
  assign n28859 = pi2874 & n22622;
  assign n28860 = pi1337 & ~pi2874;
  assign n28861 = ~n22628 & ~n28860;
  assign n28862 = ~n22622 & ~n28861;
  assign po3048 = n28859 | n28862;
  assign n28864 = ~pi2875 & ~n22539;
  assign n28865 = pi3092 & n22539;
  assign n28866 = ~n28864 & ~n28865;
  assign n28867 = n22306 & ~n28866;
  assign n28868 = ~pi2875 & ~n22306;
  assign po3049 = n28867 | n28868;
  assign n28870 = ~pi2876 & ~n22539;
  assign n28871 = pi3100 & n22539;
  assign n28872 = ~n28870 & ~n28871;
  assign n28873 = n22306 & ~n28872;
  assign n28874 = ~pi2876 & ~n22306;
  assign po3050 = n28873 | n28874;
  assign n28876 = ~pi2877 & ~n22539;
  assign n28877 = pi3055 & n22539;
  assign n28878 = ~n28876 & ~n28877;
  assign n28879 = n22306 & ~n28878;
  assign n28880 = ~pi2877 & ~n22306;
  assign po3051 = n28879 | n28880;
  assign n28882 = pi3096 & n22311;
  assign n28883 = ~pi2878 & ~n22311;
  assign n28884 = ~n28882 & ~n28883;
  assign n28885 = n22306 & ~n28884;
  assign n28886 = ~pi2878 & ~n22306;
  assign po3052 = n28885 | n28886;
  assign n28888 = pi3090 & n22561;
  assign n28889 = ~pi2879 & ~n22561;
  assign n28890 = ~n28888 & ~n28889;
  assign n28891 = n22306 & ~n28890;
  assign n28892 = ~pi2879 & ~n22306;
  assign po3053 = n28891 | n28892;
  assign n28894 = pi3097 & n22554;
  assign n28895 = ~pi2880 & ~n22554;
  assign n28896 = ~n28894 & ~n28895;
  assign n28897 = n22306 & ~n28896;
  assign n28898 = ~pi2880 & ~n22306;
  assign po3054 = n28897 | n28898;
  assign n28900 = pi3045 & n22554;
  assign n28901 = ~pi2881 & ~n22554;
  assign n28902 = ~n28900 & ~n28901;
  assign n28903 = n22306 & ~n28902;
  assign n28904 = ~pi2881 & ~n22306;
  assign po3055 = n28903 | n28904;
  assign n28906 = pi3047 & n22554;
  assign n28907 = ~pi2882 & ~n22554;
  assign n28908 = ~n28906 & ~n28907;
  assign n28909 = n22306 & ~n28908;
  assign n28910 = ~pi2882 & ~n22306;
  assign po3056 = n28909 | n28910;
  assign n28912 = ~pi2883 & ~n22539;
  assign n28913 = pi3059 & n22539;
  assign n28914 = ~n28912 & ~n28913;
  assign n28915 = n22306 & ~n28914;
  assign n28916 = ~pi2883 & ~n22306;
  assign po3057 = n28915 | n28916;
  assign n28918 = pi0263 & n20262;
  assign n28919 = pi2884 & ~n20262;
  assign po3058 = n28918 | n28919;
  assign n28921 = pi0248 & n20262;
  assign n28922 = pi2885 & ~n20262;
  assign po3059 = n28921 | n28922;
  assign n28924 = pi3058 & n22561;
  assign n28925 = ~pi2886 & ~n22561;
  assign n28926 = ~n28924 & ~n28925;
  assign n28927 = n22306 & ~n28926;
  assign n28928 = ~pi2886 & ~n22306;
  assign po3060 = n28927 | n28928;
  assign n28930 = ~pi2887 & ~n22539;
  assign n28931 = pi3058 & n22539;
  assign n28932 = ~n28930 & ~n28931;
  assign n28933 = n22306 & ~n28932;
  assign n28934 = ~pi2887 & ~n22306;
  assign po3061 = n28933 | n28934;
  assign n28936 = pi0301 & n20262;
  assign n28937 = pi2888 & ~n20262;
  assign po3062 = n28936 | n28937;
  assign n28939 = pi0254 & n20262;
  assign n28940 = pi2889 & ~n20262;
  assign po3063 = n28939 | n28940;
  assign n28942 = ~pi2890 & ~n22539;
  assign n28943 = pi3050 & n22539;
  assign n28944 = ~n28942 & ~n28943;
  assign n28945 = n22306 & ~n28944;
  assign n28946 = ~pi2890 & ~n22306;
  assign po3064 = n28945 | n28946;
  assign n28948 = ~pi2891 & ~n22318;
  assign n28949 = pi3058 & n22318;
  assign n28950 = ~n28948 & ~n28949;
  assign n28951 = n22306 & ~n28950;
  assign n28952 = ~pi2891 & ~n22306;
  assign po3065 = n28951 | n28952;
  assign n28954 = pi3089 & n22554;
  assign n28955 = ~pi2892 & ~n22554;
  assign n28956 = ~n28954 & ~n28955;
  assign n28957 = n22306 & ~n28956;
  assign n28958 = ~pi2892 & ~n22306;
  assign po3066 = n28957 | n28958;
  assign n28960 = ~pi2893 & ~n22539;
  assign n28961 = pi3056 & n22539;
  assign n28962 = ~n28960 & ~n28961;
  assign n28963 = n22306 & ~n28962;
  assign n28964 = ~pi2893 & ~n22306;
  assign po3067 = n28963 | n28964;
  assign n28966 = pi0271 & n20262;
  assign n28967 = pi2894 & ~n20262;
  assign po3068 = n28966 | n28967;
  assign n28969 = pi0258 & n20262;
  assign n28970 = pi2895 & ~n20262;
  assign po3069 = n28969 | n28970;
  assign n28972 = pi3087 & n22554;
  assign n28973 = ~pi2896 & ~n22554;
  assign n28974 = ~n28972 & ~n28973;
  assign n28975 = n22306 & ~n28974;
  assign n28976 = ~pi2896 & ~n22306;
  assign po3070 = n28975 | n28976;
  assign n28978 = pi3048 & n22554;
  assign n28979 = ~pi2897 & ~n22554;
  assign n28980 = ~n28978 & ~n28979;
  assign n28981 = n22306 & ~n28980;
  assign n28982 = ~pi2897 & ~n22306;
  assign po3071 = n28981 | n28982;
  assign n28984 = pi3086 & n22554;
  assign n28985 = ~pi2898 & ~n22554;
  assign n28986 = ~n28984 & ~n28985;
  assign n28987 = n22306 & ~n28986;
  assign n28988 = ~pi2898 & ~n22306;
  assign po3072 = n28987 | n28988;
  assign n28990 = ~pi2899 & ~n22318;
  assign n28991 = pi3089 & n22318;
  assign n28992 = ~n28990 & ~n28991;
  assign n28993 = n22306 & ~n28992;
  assign n28994 = ~pi2899 & ~n22306;
  assign po3073 = n28993 | n28994;
  assign n28996 = ~pi2900 & ~n22539;
  assign n28997 = pi3101 & n22539;
  assign n28998 = ~n28996 & ~n28997;
  assign n28999 = n22306 & ~n28998;
  assign n29000 = ~pi2900 & ~n22306;
  assign po3074 = n28999 | n29000;
  assign n29002 = pi0270 & n20262;
  assign n29003 = pi2901 & ~n20262;
  assign po3075 = n29002 | n29003;
  assign n29005 = ~pi2902 & ~n22539;
  assign n29006 = pi3090 & n22539;
  assign n29007 = ~n29005 & ~n29006;
  assign n29008 = n22306 & ~n29007;
  assign n29009 = ~pi2902 & ~n22306;
  assign po3076 = n29008 | n29009;
  assign n29011 = pi3092 & n22554;
  assign n29012 = ~pi2903 & ~n22554;
  assign n29013 = ~n29011 & ~n29012;
  assign n29014 = n22306 & ~n29013;
  assign n29015 = ~pi2903 & ~n22306;
  assign po3077 = n29014 | n29015;
  assign n29017 = pi0256 & n20262;
  assign n29018 = pi2904 & ~n20262;
  assign po3078 = n29017 | n29018;
  assign n29020 = pi3103 & n22311;
  assign n29021 = ~pi2905 & ~n22311;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = n22306 & ~n29022;
  assign n29024 = ~pi2905 & ~n22306;
  assign po3079 = n29023 | n29024;
  assign n29026 = pi2906 & ~n27328;
  assign n29027 = ~pi2906 & n27328;
  assign po3080 = n29026 | n29027;
  assign n29029 = ~pi2907 & ~n27328;
  assign n29030 = ~pi2593 & n27328;
  assign po3081 = n29029 | n29030;
  assign n29032 = pi2908 & pi3175;
  assign n29033 = ~pi2908 & n22297;
  assign n29034 = pi1686 & n29033;
  assign po3082 = n29032 | n29034;
  assign n29036 = ~pi2919 & ~pi2925;
  assign n29037 = pi2909 & ~n29036;
  assign n29038 = ~pi2909 & ~pi2919;
  assign n29039 = ~pi2925 & n29038;
  assign n29040 = ~n29037 & ~n29039;
  assign n29041 = ~pi1220 & pi3373;
  assign n29042 = ~n20029 & ~n29041;
  assign n29043 = n9391 & n15368;
  assign n29044 = ~n29042 & n29043;
  assign po3083 = ~n29040 | ~n29044;
  assign n29046 = pi3210 & pi3351;
  assign n29047 = ~pi2910 & ~n29046;
  assign po3084 = n23716 | n29047;
  assign n29049 = ~pi1337 & n19974;
  assign n29050 = ~pi1858 & n29049;
  assign n29051 = ~pi1265 & n29050;
  assign n29052 = ~pi2911 & n29051;
  assign n29053 = pi2911 & ~n19958;
  assign po3085 = n29052 | n29053;
  assign n29055 = pi2961 & n19402;
  assign n29056 = n7250 & n29055;
  assign n29057 = ~n8057 & n29056;
  assign po3087 = ~pi3203 | n29057;
  assign n29059 = ~n22310 & ~n22546;
  assign n29060 = n22306 & ~n29059;
  assign n29061 = pi2914 & ~n22306;
  assign po3088 = n29060 | n29061;
  assign n29063 = pi2915 & ~n22306;
  assign n29064 = ~pi2915 & ~pi2917;
  assign n29065 = pi2915 & pi2917;
  assign n29066 = ~n29064 & ~n29065;
  assign n29067 = n22306 & n29066;
  assign po3089 = n29063 | n29067;
  assign n29069 = pi2916 & ~n22306;
  assign po3090 = n29067 | n29069;
  assign n29071 = pi2917 & ~n22306;
  assign n29072 = ~pi2917 & n22306;
  assign po3091 = n29071 | n29072;
  assign n29074 = pi1965 & ~n29056;
  assign n29075 = ~pi2918 & n29074;
  assign po3092 = ~pi3189 & ~n29075;
  assign n29077 = pi2919 & pi2925;
  assign n29078 = ~n29036 & ~n29077;
  assign po3093 = n29044 & ~n29078;
  assign n29080 = pi3166 & n8009;
  assign n29081 = pi2920 & ~n8009;
  assign po3094 = n29080 | n29081;
  assign n29083 = pi2921 & ~n22306;
  assign n29084 = ~pi2923 & pi2949;
  assign n29085 = pi2923 & ~pi2949;
  assign n29086 = ~n29084 & ~n29085;
  assign n29087 = n22306 & ~n29086;
  assign po3095 = n29083 | n29087;
  assign n29089 = pi2922 & ~n22306;
  assign n29090 = ~pi2922 & n22306;
  assign po3096 = n29089 | n29090;
  assign n29092 = pi2923 & ~n22306;
  assign po3097 = n29060 | n29092;
  assign n29094 = ~pi1232 & n19470;
  assign n29095 = ~pi2924 & ~n29094;
  assign po3098 = n9402 & ~n29095;
  assign po3099 = ~pi2925 & n29044;
  assign n29098 = ~pi2926 & ~n22326;
  assign n29099 = pi3128 & n22326;
  assign n29100 = ~n29098 & ~n29099;
  assign n29101 = n22306 & ~n29100;
  assign n29102 = ~pi2926 & ~n22306;
  assign po3100 = n29101 | n29102;
  assign n29104 = ~pi2927 & ~n22547;
  assign n29105 = pi3128 & n22547;
  assign n29106 = ~n29104 & ~n29105;
  assign n29107 = n22306 & ~n29106;
  assign n29108 = ~pi2927 & ~n22306;
  assign po3101 = n29107 | n29108;
  assign n29110 = pi3128 & n22554;
  assign n29111 = ~pi2928 & ~n22554;
  assign n29112 = ~n29110 & ~n29111;
  assign n29113 = n22306 & ~n29112;
  assign n29114 = ~pi2928 & ~n22306;
  assign po3102 = n29113 | n29114;
  assign n29116 = ~pi2929 & ~n22539;
  assign n29117 = pi3128 & n22539;
  assign n29118 = ~n29116 & ~n29117;
  assign n29119 = n22306 & ~n29118;
  assign n29120 = ~pi2929 & ~n22306;
  assign po3103 = n29119 | n29120;
  assign n29122 = ~pi2930 & ~n22318;
  assign n29123 = pi3128 & n22318;
  assign n29124 = ~n29122 & ~n29123;
  assign n29125 = n22306 & ~n29124;
  assign n29126 = ~pi2930 & ~n22306;
  assign po3104 = n29125 | n29126;
  assign n29128 = pi3128 & n22561;
  assign n29129 = ~pi2931 & ~n22561;
  assign n29130 = ~n29128 & ~n29129;
  assign n29131 = n22306 & ~n29130;
  assign n29132 = ~pi2931 & ~n22306;
  assign po3105 = n29131 | n29132;
  assign n29134 = pi3128 & n22311;
  assign n29135 = ~pi2932 & ~n22311;
  assign n29136 = ~n29134 & ~n29135;
  assign n29137 = n22306 & ~n29136;
  assign n29138 = ~pi2932 & ~n22306;
  assign po3106 = n29137 | n29138;
  assign n29140 = pi3128 & n22302;
  assign n29141 = ~pi2933 & ~n22302;
  assign n29142 = ~n29140 & ~n29141;
  assign n29143 = n22306 & ~n29142;
  assign n29144 = ~pi2933 & ~n22306;
  assign po3107 = n29143 | n29144;
  assign n29146 = pi2936 & n22306;
  assign n29147 = pi2934 & ~n22306;
  assign po3108 = n29146 | n29147;
  assign n29149 = pi2914 & n22306;
  assign n29150 = pi2935 & ~n22306;
  assign po3109 = n29149 | n29150;
  assign n29152 = pi2940 & n22306;
  assign n29153 = pi2936 & ~n22306;
  assign po3110 = n29152 | n29153;
  assign n29155 = pi2937 & ~n8009;
  assign po3111 = n19906 | n29155;
  assign n29157 = pi3378 & n14916;
  assign n29158 = pi2938 & ~n14916;
  assign po3112 = n29157 | n29158;
  assign n29160 = pi2977 & n23688;
  assign n29161 = pi2970 & n29160;
  assign n29162 = pi2979 & pi2986;
  assign n29163 = n23689 & n23691;
  assign n29164 = n29162 & n29163;
  assign n29165 = n29161 & n29164;
  assign n29166 = pi2957 & pi2962;
  assign n29167 = n29165 & n29166;
  assign n29168 = pi2947 & n29167;
  assign n29169 = pi2974 & n29168;
  assign n29170 = pi2939 & n29169;
  assign n29171 = ~pi2939 & ~n29169;
  assign n29172 = ~n29170 & ~n29171;
  assign po3113 = n23709 & n29172;
  assign n29174 = pi2949 & n22306;
  assign n29175 = pi2940 & ~n22306;
  assign po3114 = n29174 | n29175;
  assign n29177 = pi3379 & n14916;
  assign n29178 = pi2941 & ~n14916;
  assign po3115 = n29177 | n29178;
  assign n29180 = pi2953 & n22306;
  assign n29181 = pi2942 & ~n22306;
  assign po3116 = n29180 | n29181;
  assign n29183 = ~pi2918 & pi3231;
  assign n29184 = pi2918 & pi2943;
  assign n29185 = ~n29183 & ~n29184;
  assign po3117 = n29074 & ~n29185;
  assign n29187 = n9396 & n29042;
  assign n29188 = ~pi2944 & ~n29187;
  assign po3118 = n9391 & ~n29188;
  assign n29190 = pi2921 & n22306;
  assign n29191 = pi2945 & ~n22306;
  assign po3119 = n29190 | n29191;
  assign n29193 = pi0120 & pi3207;
  assign n29194 = pi3057 & ~n20042;
  assign n29195 = ~pi3057 & n20042;
  assign n29196 = ~n29194 & ~n29195;
  assign n29197 = pi2972 & ~n20045;
  assign n29198 = ~pi2972 & n20045;
  assign n29199 = ~n29197 & ~n29198;
  assign n29200 = pi3018 & ~n20051;
  assign n29201 = ~pi3018 & n20051;
  assign n29202 = ~n29200 & ~n29201;
  assign n29203 = pi3020 & ~n20054;
  assign n29204 = ~pi3020 & n20054;
  assign n29205 = ~n29203 & ~n29204;
  assign n29206 = ~n29202 & ~n29205;
  assign n29207 = ~n29199 & n29206;
  assign n29208 = ~n29196 & n29207;
  assign po3120 = n29193 & ~n29208;
  assign n29210 = pi2983 & n29160;
  assign n29211 = n23690 & n29162;
  assign n29212 = pi2998 & n29211;
  assign n29213 = pi2991 & n29212;
  assign n29214 = n29210 & n29213;
  assign n29215 = pi2970 & n29214;
  assign n29216 = n23699 & n29215;
  assign n29217 = pi2962 & n29216;
  assign n29218 = pi2947 & n29217;
  assign n29219 = ~pi2947 & ~n29217;
  assign n29220 = ~n29218 & ~n29219;
  assign po3121 = n23709 & n29220;
  assign po3122 = pi2948 & pi2985;
  assign n29223 = ~pi2922 & pi2949;
  assign n29224 = ~n29084 & ~n29223;
  assign n29225 = ~n22326 & n29224;
  assign n29226 = n22306 & ~n29225;
  assign n29227 = pi2949 & ~n22306;
  assign po3123 = n29226 | n29227;
  assign n29229 = n8031 & n11053;
  assign n29230 = pi3020 & n29229;
  assign po3124 = pi3018 & n29230;
  assign n29232 = ~pi2915 & pi2953;
  assign n29233 = pi2915 & ~pi2953;
  assign n29234 = ~n29232 & ~n29233;
  assign n29235 = n22306 & ~n29234;
  assign n29236 = pi2951 & ~n22306;
  assign po3125 = n29235 | n29236;
  assign n29238 = pi3508 & n14916;
  assign n29239 = pi2952 & ~n14916;
  assign po3126 = n29238 | n29239;
  assign n29241 = ~pi2917 & pi2953;
  assign n29242 = pi2917 & n29233;
  assign n29243 = ~n29241 & ~n29242;
  assign n29244 = ~n29232 & n29243;
  assign n29245 = n22306 & ~n29244;
  assign n29246 = pi2953 & ~n22306;
  assign po3127 = n29245 | n29246;
  assign n29248 = pi2945 & n22306;
  assign n29249 = pi2954 & ~n22306;
  assign po3128 = n29248 | n29249;
  assign n29251 = pi3506 & n14916;
  assign n29252 = pi2955 & ~n14916;
  assign po3129 = n29251 | n29252;
  assign n29254 = pi2935 & n22306;
  assign n29255 = pi2956 & ~n22306;
  assign po3130 = n29254 | n29255;
  assign n29257 = pi2957 & n23698;
  assign n29258 = ~pi2957 & ~n23698;
  assign n29259 = ~n29257 & ~n29258;
  assign po3131 = n23709 & n29259;
  assign n29261 = pi3507 & n14916;
  assign n29262 = pi2958 & ~n14916;
  assign po3132 = n29261 | n29262;
  assign n29264 = pi3509 & n14916;
  assign n29265 = pi2959 & ~n14916;
  assign po3133 = n29264 | n29265;
  assign n29267 = pi3363 & n14916;
  assign n29268 = pi2960 & ~n14916;
  assign po3134 = n29267 | n29268;
  assign n29270 = pi2961 & ~n19402;
  assign n29271 = pi0126 & ~pi0128;
  assign n29272 = ~n29270 & ~n29271;
  assign n29273 = ~pi0120 & n29272;
  assign po3135 = pi2758 & ~n29273;
  assign n29275 = pi2962 & n29165;
  assign n29276 = ~pi2962 & ~n29165;
  assign n29277 = ~n29275 & ~n29276;
  assign po3136 = n23709 & n29277;
  assign n29279 = pi2963 & ~n8009;
  assign po3137 = n19634 | n29279;
  assign n29281 = pi2964 & ~pi3160;
  assign n29282 = pi3126 & pi3160;
  assign po3138 = n29281 | n29282;
  assign n29284 = pi2965 & ~n8009;
  assign n29285 = pi2972 & n8009;
  assign po3139 = n29284 | n29285;
  assign n29287 = pi2966 & ~n8009;
  assign n29288 = pi3142 & n8009;
  assign po3140 = n29287 | n29288;
  assign po3141 = n22296 | n23713;
  assign po3168 = n7078 & n7101;
  assign po3142 = n7496 | po3168;
  assign n29293 = pi2969 & ~n8009;
  assign po3143 = n29285 | n29293;
  assign n29295 = ~pi2970 & ~n29214;
  assign n29296 = ~n29215 & ~n29295;
  assign po3144 = n23709 & n29296;
  assign n29298 = ~pi3120 & ~pi3123;
  assign n29299 = pi1344 & n29298;
  assign n29300 = ~po3339 & n29299;
  assign n29301 = ~pi3123 & n29300;
  assign n29302 = pi2972 & n29301;
  assign n29303 = ~pi2971 & ~n29301;
  assign po3145 = n29302 | n29303;
  assign n29305 = pi2972 & ~pi3160;
  assign n29306 = pi3160 & ~n20045;
  assign po3146 = n29305 | n29306;
  assign n29308 = pi2973 & n23695;
  assign n29309 = ~pi2973 & ~n23695;
  assign n29310 = ~n29308 & ~n29309;
  assign po3147 = n23709 & n29310;
  assign n29312 = pi2999 & n29162;
  assign n29313 = pi3002 & n29312;
  assign n29314 = pi2991 & n29313;
  assign n29315 = pi2977 & n23689;
  assign n29316 = pi2973 & n29315;
  assign n29317 = n29314 & n29316;
  assign n29318 = n29166 & n29317;
  assign n29319 = pi2978 & n29318;
  assign n29320 = pi2970 & n29319;
  assign n29321 = pi2974 & n29320;
  assign n29322 = ~pi2974 & ~n29320;
  assign n29323 = ~n29321 & ~n29322;
  assign po3148 = n23709 & n29323;
  assign n29325 = pi1805 & n9396;
  assign po3149 = n9402 & n29325;
  assign n29327 = pi2965 & ~pi3207;
  assign n29328 = pi2972 & pi3207;
  assign po3150 = n29327 | n29328;
  assign n29330 = pi2977 & n29164;
  assign n29331 = ~pi2977 & ~n29164;
  assign n29332 = ~n29330 & ~n29331;
  assign po3151 = n23709 & n29332;
  assign n29334 = pi2978 & n29317;
  assign n29335 = ~pi2978 & ~n29317;
  assign n29336 = ~n29334 & ~n29335;
  assign po3152 = n23709 & n29336;
  assign n29338 = ~pi2979 & ~n23692;
  assign n29339 = ~n23693 & ~n29338;
  assign po3153 = n23709 & n29339;
  assign n29341 = pi3163 & n8009;
  assign n29342 = pi2980 & ~n8009;
  assign po3154 = n29341 | n29342;
  assign n29344 = pi2981 & ~n8009;
  assign n29345 = pi3170 & n8009;
  assign po3155 = n29344 | n29345;
  assign n29347 = pi2982 & ~n8009;
  assign n29348 = pi3159 & n8009;
  assign po3156 = n29347 | n29348;
  assign n29350 = pi2983 & n29213;
  assign n29351 = ~pi2983 & ~n29213;
  assign n29352 = ~n29350 & ~n29351;
  assign po3157 = n23709 & n29352;
  assign n29354 = pi2984 & ~n8009;
  assign po3158 = n9001 | n29354;
  assign n29356 = ~pi2986 & ~n23691;
  assign n29357 = ~n23692 & ~n29356;
  assign po3160 = n23709 & n29357;
  assign n29359 = ~pi3207 & n8147;
  assign n29360 = ~pi3107 & n29359;
  assign n29361 = pi3136 & pi3207;
  assign po3161 = n29360 | n29361;
  assign n29363 = ~pi2990 & n29359;
  assign n29364 = pi3163 & pi3207;
  assign po3162 = n29363 | n29364;
  assign n29366 = pi3179 & po3351;
  assign po3163 = pi1337 | n29366;
  assign n29368 = ~pi2990 & ~n8009;
  assign po3164 = n29341 | n29368;
  assign n29370 = ~pi2991 & ~n23690;
  assign n29371 = ~n23691 & ~n29370;
  assign po3165 = n23709 & n29371;
  assign n29373 = ~pi2992 & ~n8009;
  assign po3166 = n29288 | n29373;
  assign n29375 = pi2993 & ~n8009;
  assign n29376 = pi3057 & n8009;
  assign po3167 = n29375 | n29376;
  assign n29378 = pi2995 & ~n8009;
  assign n29379 = pi3145 & n8009;
  assign po3169 = n29378 | n29379;
  assign n29381 = pi2996 & ~n8009;
  assign n29382 = pi3131 & n8009;
  assign po3170 = n29381 | n29382;
  assign n29384 = pi2997 & ~n8009;
  assign n29385 = pi3146 & n8009;
  assign po3171 = n29384 | n29385;
  assign n29387 = pi2998 & n29314;
  assign n29388 = ~pi2998 & ~n29314;
  assign n29389 = ~n29387 & ~n29388;
  assign po3172 = n23709 & n29389;
  assign n29391 = ~pi2999 & ~pi3002;
  assign n29392 = ~n23690 & ~n29391;
  assign po3173 = n23709 & n29392;
  assign n29394 = ~pi3000 & ~n8009;
  assign po3174 = n29348 | n29394;
  assign n29396 = pi3001 & ~n8009;
  assign n29397 = pi3169 & n8009;
  assign po3175 = n29396 | n29397;
  assign po3176 = ~pi3002 & n23709;
  assign n29400 = ~pi3003 & ~n8009;
  assign po3177 = n29080 | n29400;
  assign n29402 = pi3168 & n8009;
  assign n29403 = pi3004 & ~n8009;
  assign po3178 = n29402 | n29403;
  assign n29405 = pi3009 & n29301;
  assign n29406 = pi3005 & ~n29301;
  assign po3179 = n29405 | n29406;
  assign n29408 = pi3038 & n29301;
  assign n29409 = pi3006 & ~n29301;
  assign po3180 = n29408 | n29409;
  assign n29411 = pi2993 & n29301;
  assign n29412 = pi3007 & ~n29301;
  assign po3181 = n29411 | n29412;
  assign n29414 = pi3134 & n8009;
  assign n29415 = pi3008 & ~n8009;
  assign po3182 = n29414 | n29415;
  assign n29417 = pi3165 & n8009;
  assign n29418 = pi3009 & ~n8009;
  assign po3183 = n29417 | n29418;
  assign n29420 = pi3154 & n8009;
  assign n29421 = pi3010 & ~n8009;
  assign po3184 = n29420 | n29421;
  assign n29423 = pi3138 & n8009;
  assign n29424 = pi3011 & ~n8009;
  assign po3185 = n29423 | n29424;
  assign n29426 = pi3151 & n8009;
  assign n29427 = pi3012 & ~n8009;
  assign po3186 = n29426 | n29427;
  assign n29429 = pi3008 & n29301;
  assign n29430 = pi3013 & ~n29301;
  assign po3187 = n29429 | n29430;
  assign n29432 = pi3132 & n8009;
  assign n29433 = pi3014 & ~n8009;
  assign po3188 = n29432 | n29433;
  assign n29435 = pi3139 & n8009;
  assign n29436 = pi3015 & ~n8009;
  assign po3189 = n29435 | n29436;
  assign n29438 = pi3057 & n29301;
  assign n29439 = ~pi3016 & ~n29301;
  assign po3190 = n29438 | n29439;
  assign n29441 = pi3133 & n8009;
  assign n29442 = pi3017 & ~n8009;
  assign po3191 = n29441 | n29442;
  assign n29444 = pi3018 & ~pi3160;
  assign n29445 = pi3160 & ~n20051;
  assign po3192 = n29444 | n29445;
  assign n29447 = pi3147 & n8009;
  assign n29448 = pi3019 & ~n8009;
  assign po3193 = n29447 | n29448;
  assign n29450 = pi3020 & ~pi3160;
  assign n29451 = pi3160 & ~n20054;
  assign po3194 = n29450 | n29451;
  assign n29453 = pi3135 & n8009;
  assign n29454 = pi3021 & ~n8009;
  assign po3195 = n29453 | n29454;
  assign n29456 = pi3172 & n8009;
  assign n29457 = pi3022 & ~n8009;
  assign po3196 = n29456 | n29457;
  assign n29459 = pi3143 & n8009;
  assign n29460 = pi3023 & ~n8009;
  assign po3197 = n29459 | n29460;
  assign n29462 = pi3024 & ~n8009;
  assign n29463 = pi3018 & n8009;
  assign po3198 = n29462 | n29463;
  assign n29465 = pi3025 & ~n8009;
  assign n29466 = pi3020 & n8009;
  assign po3199 = n29465 | n29466;
  assign n29468 = ~pi3003 & n29301;
  assign n29469 = pi3026 & ~n29301;
  assign po3200 = n29468 | n29469;
  assign n29471 = n15368 & n29038;
  assign po3201 = ~n29042 & n29471;
  assign n29473 = pi3041 & n29301;
  assign n29474 = pi3028 & ~n29301;
  assign po3202 = n29473 | n29474;
  assign n29476 = pi3012 & n29301;
  assign n29477 = pi3029 & ~n29301;
  assign po3203 = n29476 | n29477;
  assign n29479 = pi3011 & n29301;
  assign n29480 = pi3030 & ~n29301;
  assign po3204 = n29479 | n29480;
  assign n29482 = pi3010 & n29301;
  assign n29483 = pi3031 & ~n29301;
  assign po3205 = n29482 | n29483;
  assign n29485 = pi3021 & n29301;
  assign n29486 = pi3032 & ~n29301;
  assign po3206 = n29485 | n29486;
  assign n29488 = pi3065 & n29301;
  assign n29489 = pi3033 & ~n29301;
  assign po3207 = n29488 | n29489;
  assign n29491 = n8153 & n29301;
  assign n29492 = pi3034 & ~n29301;
  assign po3208 = n29491 | n29492;
  assign n29494 = ~pi3106 & n29301;
  assign n29495 = pi3035 & ~n29301;
  assign po3209 = n29494 | n29495;
  assign n29497 = ~pi3036 & ~n8009;
  assign po3210 = n29397 | n29497;
  assign n29499 = ~pi3110 & n29301;
  assign n29500 = pi3037 & ~n29301;
  assign po3211 = n29499 | n29500;
  assign n29502 = pi3162 & n8009;
  assign n29503 = pi3038 & ~n8009;
  assign po3212 = n29502 | n29503;
  assign n29505 = pi3141 & n8009;
  assign n29506 = pi3039 & ~n8009;
  assign po3213 = n29505 | n29506;
  assign n29508 = pi3158 & n8009;
  assign n29509 = pi3040 & ~n8009;
  assign po3214 = n29508 | n29509;
  assign n29511 = pi3157 & n8009;
  assign n29512 = pi3041 & ~n8009;
  assign po3215 = n29511 | n29512;
  assign n29514 = pi3042 & ~pi3160;
  assign n29515 = pi3160 & ~n9396;
  assign po3216 = n29514 | n29515;
  assign n29517 = pi3153 & n8009;
  assign n29518 = pi3043 & ~n8009;
  assign po3217 = n29517 | n29518;
  assign n29520 = pi3022 & n29301;
  assign n29521 = pi3044 & ~n29301;
  assign po3218 = n29520 | n29521;
  assign n29523 = pi3023 & ~pi3207;
  assign n29524 = pi3143 & pi3207;
  assign po3219 = n29523 | n29524;
  assign n29526 = ~pi3104 & n29301;
  assign n29527 = pi3046 & ~n29301;
  assign po3220 = n29526 | n29527;
  assign n29529 = pi3038 & ~pi3207;
  assign n29530 = pi3162 & pi3207;
  assign po3221 = n29529 | n29530;
  assign n29532 = pi3024 & ~pi3207;
  assign n29533 = pi3018 & pi3207;
  assign po3222 = n29532 | n29533;
  assign n29535 = pi3065 & ~pi3207;
  assign n29536 = pi3155 & pi3207;
  assign po3223 = n29535 | n29536;
  assign n29538 = pi3022 & ~pi3207;
  assign n29539 = pi3172 & pi3207;
  assign po3224 = n29538 | n29539;
  assign n29541 = pi3040 & n29301;
  assign n29542 = pi3051 & ~n29301;
  assign po3225 = n29541 | n29542;
  assign n29544 = ~pi3108 & ~pi3207;
  assign n29545 = pi3170 & pi3207;
  assign po3226 = n29544 | n29545;
  assign n29547 = ~pi3106 & ~pi3207;
  assign n29548 = pi3145 & pi3207;
  assign po3227 = n29547 | n29548;
  assign n29550 = ~pi3000 & ~pi3207;
  assign n29551 = pi3159 & pi3207;
  assign po3228 = n29550 | n29551;
  assign n29553 = pi2993 & ~pi3207;
  assign n29554 = pi3057 & pi3207;
  assign po3229 = n29553 | n29554;
  assign n29556 = pi3063 & ~pi3207;
  assign n29557 = pi3150 & pi3207;
  assign po3230 = n29556 | n29557;
  assign n29559 = pi3057 & ~pi3160;
  assign n29560 = pi3160 & ~n20042;
  assign po3231 = n29559 | n29560;
  assign n29562 = pi3017 & ~pi3207;
  assign n29563 = pi3133 & pi3207;
  assign po3232 = n29562 | n29563;
  assign n29565 = pi3041 & ~pi3207;
  assign n29566 = pi3157 & pi3207;
  assign po3233 = n29565 | n29566;
  assign n29568 = pi3009 & ~pi3207;
  assign n29569 = pi3165 & pi3207;
  assign po3234 = n29568 | n29569;
  assign n29571 = pi3079 & ~pi3207;
  assign n29572 = pi3164 & pi3207;
  assign po3235 = n29571 | n29572;
  assign n29574 = pi3039 & ~pi3207;
  assign n29575 = pi3141 & pi3207;
  assign po3236 = n29574 | n29575;
  assign n29577 = pi3150 & n8009;
  assign n29578 = pi3063 & ~n8009;
  assign po3237 = n29577 | n29578;
  assign n29580 = pi3020 & n29301;
  assign n29581 = ~pi3064 & ~n29301;
  assign po3238 = n29580 | n29581;
  assign n29583 = pi3155 & n8009;
  assign n29584 = pi3065 & ~n8009;
  assign po3239 = n29583 | n29584;
  assign n29586 = ~pi2990 & n29301;
  assign n29587 = pi3066 & ~n29301;
  assign po3240 = n29586 | n29587;
  assign n29589 = pi3019 & n29301;
  assign n29590 = pi3067 & ~n29301;
  assign po3241 = n29589 | n29590;
  assign n29592 = ~pi3000 & n29301;
  assign n29593 = pi3068 & ~n29301;
  assign po3242 = n29592 | n29593;
  assign n29595 = pi3004 & n29301;
  assign n29596 = pi3069 & ~n29301;
  assign po3243 = n29595 | n29596;
  assign n29598 = pi3018 & n29301;
  assign n29599 = ~pi3070 & ~n29301;
  assign po3244 = n29598 | n29599;
  assign n29601 = pi3077 & n29301;
  assign n29602 = pi3072 & ~n29301;
  assign po3246 = n29601 | n29602;
  assign n29604 = pi3043 & n29301;
  assign n29605 = pi3073 & ~n29301;
  assign po3247 = n29604 | n29605;
  assign n29607 = pi3017 & n29301;
  assign n29608 = pi3074 & ~n29301;
  assign po3248 = n29607 | n29608;
  assign n29610 = ~pi3108 & n29301;
  assign n29611 = pi3075 & ~n29301;
  assign po3249 = n29610 | n29611;
  assign n29613 = ~pi2992 & n29301;
  assign n29614 = pi3076 & ~n29301;
  assign po3250 = n29613 | n29614;
  assign n29616 = pi3171 & n8009;
  assign n29617 = pi3077 & ~n8009;
  assign po3251 = n29616 | n29617;
  assign n29619 = pi3023 & n29301;
  assign n29620 = pi3078 & ~n29301;
  assign po3252 = n29619 | n29620;
  assign n29622 = pi3164 & n8009;
  assign n29623 = pi3079 & ~n8009;
  assign po3253 = n29622 | n29623;
  assign n29625 = pi3039 & n29301;
  assign n29626 = pi3080 & ~n29301;
  assign po3254 = n29625 | n29626;
  assign n29628 = pi3015 & n29301;
  assign n29629 = pi3081 & ~n29301;
  assign po3255 = n29628 | n29629;
  assign n29631 = ~pi3117 & ~n20028;
  assign po3256 = pi3207 & ~n29631;
  assign n29633 = pi3015 & ~pi3207;
  assign n29634 = pi3139 & pi3207;
  assign po3258 = n29633 | n29634;
  assign n29636 = pi3004 & ~pi3207;
  assign n29637 = pi3168 & pi3207;
  assign po3259 = n29636 | n29637;
  assign n29639 = pi3008 & ~pi3207;
  assign n29640 = pi3134 & pi3207;
  assign po3260 = n29639 | n29640;
  assign n29642 = pi3077 & ~pi3207;
  assign n29643 = pi3171 & pi3207;
  assign po3261 = n29642 | n29643;
  assign n29645 = pi3010 & ~pi3207;
  assign n29646 = pi3154 & pi3207;
  assign po3262 = n29645 | n29646;
  assign n29648 = pi3021 & ~pi3207;
  assign n29649 = pi3135 & pi3207;
  assign po3263 = n29648 | n29649;
  assign n29651 = ~pi3003 & ~pi3207;
  assign n29652 = pi3166 & pi3207;
  assign po3264 = n29651 | n29652;
  assign n29654 = pi3025 & ~pi3207;
  assign n29655 = pi3020 & pi3207;
  assign po3265 = n29654 | n29655;
  assign n29657 = ~pi2992 & ~pi3207;
  assign n29658 = pi3142 & pi3207;
  assign po3266 = n29657 | n29658;
  assign n29660 = ~pi3036 & ~pi3207;
  assign n29661 = pi3169 & pi3207;
  assign po3267 = n29660 | n29661;
  assign n29663 = ~pi3110 & ~pi3207;
  assign n29664 = pi3131 & pi3207;
  assign po3268 = n29663 | n29664;
  assign n29666 = ~pi3104 & ~pi3207;
  assign n29667 = pi3146 & pi3207;
  assign po3269 = n29666 | n29667;
  assign n29669 = pi3040 & ~pi3207;
  assign n29670 = pi3158 & pi3207;
  assign po3270 = n29669 | n29670;
  assign n29672 = pi3011 & ~pi3207;
  assign n29673 = pi3138 & pi3207;
  assign po3271 = n29672 | n29673;
  assign n29675 = pi3019 & ~pi3207;
  assign n29676 = pi3147 & pi3207;
  assign po3272 = n29675 | n29676;
  assign n29678 = pi3043 & ~pi3207;
  assign n29679 = pi3153 & pi3207;
  assign po3273 = n29678 | n29679;
  assign n29681 = pi3012 & ~pi3207;
  assign n29682 = pi3151 & pi3207;
  assign po3274 = n29681 | n29682;
  assign n29684 = pi3014 & ~pi3207;
  assign n29685 = pi3132 & pi3207;
  assign po3275 = n29684 | n29685;
  assign n29687 = pi3024 & n29301;
  assign n29688 = pi3102 & ~n29301;
  assign po3276 = n29687 | n29688;
  assign po3277 = ~pi3117 & pi3207;
  assign n29691 = ~pi3104 & ~n8009;
  assign po3278 = n29385 | n29691;
  assign n29693 = ~pi3036 & n29301;
  assign n29694 = pi3105 & ~n29301;
  assign po3279 = n29693 | n29694;
  assign n29696 = ~pi3106 & ~n8009;
  assign po3280 = n29379 | n29696;
  assign n29698 = pi3136 & n8009;
  assign n29699 = ~pi3107 & ~n8009;
  assign po3281 = n29698 | n29699;
  assign n29701 = ~pi3108 & ~n8009;
  assign po3282 = n29345 | n29701;
  assign n29703 = pi3109 & ~n8009;
  assign po3283 = n29698 | n29703;
  assign n29705 = ~pi3110 & ~n8009;
  assign po3284 = n29382 | n29705;
  assign n29707 = pi2965 & n29301;
  assign n29708 = pi3111 & ~n29301;
  assign po3285 = n29707 | n29708;
  assign n29710 = pi3025 & n29301;
  assign n29711 = pi3112 & ~n29301;
  assign po3286 = n29710 | n29711;
  assign n29713 = pi3063 & n29301;
  assign n29714 = pi3113 & ~n29301;
  assign po3287 = n29713 | n29714;
  assign n29716 = pi3079 & n29301;
  assign n29717 = pi3114 & ~n29301;
  assign po3288 = n29716 | n29717;
  assign n29719 = ~pi3107 & n29301;
  assign n29720 = pi3115 & ~n29301;
  assign po3289 = n29719 | n29720;
  assign n29722 = pi3014 & n29301;
  assign n29723 = pi3116 & ~n29301;
  assign po3290 = n29722 | n29723;
  assign n29725 = pi3117 & ~pi3160;
  assign n29726 = pi3160 & ~n8078;
  assign po3291 = n29725 | n29726;
  assign n29728 = pi3118 & ~pi3160;
  assign n29729 = pi3160 & ~n29042;
  assign po3292 = n29728 | n29729;
  assign n29731 = pi1232 & ~n15368;
  assign po3293 = ~n15354 | n29731;
  assign n29733 = pi3120 & ~pi3160;
  assign n29734 = pi3160 & ~n8170;
  assign po3294 = n29733 | n29734;
  assign po3295 = ~pi3156 & pi3249;
  assign n29737 = pi3184 & pi3239;
  assign n29738 = ~pi2943 & ~n29737;
  assign n29739 = ~pi3123 & ~n29299;
  assign po3296 = n29738 & ~n29739;
  assign n29741 = pi3124 & ~pi3160;
  assign n29742 = pi3160 & ~n15367;
  assign po3297 = n29741 | n29742;
  assign n29744 = pi3131 & ~pi3160;
  assign n29745 = pi3160 & pi3481;
  assign po3304 = n29744 | n29745;
  assign n29747 = pi3132 & ~pi3160;
  assign n29748 = pi3160 & pi3491;
  assign po3305 = n29747 | n29748;
  assign n29750 = pi3133 & ~pi3160;
  assign n29751 = pi3160 & pi3504;
  assign po3306 = n29750 | n29751;
  assign n29753 = pi3134 & ~pi3160;
  assign n29754 = pi3160 & pi3490;
  assign po3307 = n29753 | n29754;
  assign n29756 = pi3135 & ~pi3160;
  assign n29757 = pi3160 & pi3502;
  assign po3308 = n29756 | n29757;
  assign n29759 = pi3136 & ~pi3160;
  assign n29760 = pi3160 & pi3474;
  assign po3309 = n29759 | n29760;
  assign po3393 = pi1405 & ~pi1966;
  assign n29763 = ~pi1373 & ~po3393;
  assign po3384 = pi1395 & pi3360;
  assign po3310 = ~n29763 | po3384;
  assign n29766 = pi3138 & ~pi3160;
  assign n29767 = pi3160 & pi3498;
  assign po3311 = n29766 | n29767;
  assign n29769 = pi3139 & ~pi3160;
  assign n29770 = pi3160 & pi3484;
  assign po3312 = n29769 | n29770;
  assign n29772 = ~pi1706 & ~pi1708;
  assign n29773 = ~pi1400 & ~pi1709;
  assign n29774 = n22626 & n29773;
  assign po3313 = n29772 & ~n29774;
  assign n29776 = pi3141 & ~pi3160;
  assign n29777 = pi3160 & pi3486;
  assign po3314 = n29776 | n29777;
  assign n29779 = pi3142 & ~pi3160;
  assign n29780 = pi3160 & pi3477;
  assign po3315 = n29779 | n29780;
  assign n29782 = pi3143 & ~pi3160;
  assign n29783 = pi3160 & pi3487;
  assign po3316 = n29782 | n29783;
  assign n29785 = pi3145 & ~pi3160;
  assign n29786 = pi3160 & pi3478;
  assign po3318 = n29785 | n29786;
  assign n29788 = pi3146 & ~pi3160;
  assign n29789 = pi3160 & pi3483;
  assign po3319 = n29788 | n29789;
  assign n29791 = pi3147 & ~pi3160;
  assign n29792 = pi3160 & pi3488;
  assign po3320 = n29791 | n29792;
  assign n29794 = pi3150 & ~pi3160;
  assign n29795 = pi3160 & pi3503;
  assign po3323 = n29794 | n29795;
  assign n29797 = pi3151 & ~pi3160;
  assign n29798 = pi3160 & pi3499;
  assign po3324 = n29797 | n29798;
  assign n29800 = pi3153 & ~pi3160;
  assign n29801 = pi3160 & pi3489;
  assign po3325 = n29800 | n29801;
  assign n29803 = pi3154 & ~pi3160;
  assign n29804 = pi3160 & pi3497;
  assign po3326 = n29803 | n29804;
  assign n29806 = pi3155 & ~pi3160;
  assign n29807 = pi3160 & pi3494;
  assign po3327 = n29806 | n29807;
  assign n29809 = pi3157 & ~pi3160;
  assign n29810 = pi3160 & pi3500;
  assign po3329 = n29809 | n29810;
  assign n29812 = pi3158 & ~pi3160;
  assign n29813 = pi3160 & pi3505;
  assign po3330 = n29812 | n29813;
  assign n29815 = pi3159 & ~pi3160;
  assign n29816 = pi3160 & pi3480;
  assign po3331 = n29815 | n29816;
  assign po3332 = pi3160 | pi3241;
  assign n29819 = ~pi3160 & pi3161;
  assign n29820 = pi3160 & pi3372;
  assign po3333 = n29819 | n29820;
  assign n29822 = ~pi3160 & pi3162;
  assign n29823 = pi3160 & pi3495;
  assign po3334 = n29822 | n29823;
  assign n29825 = ~pi3160 & pi3163;
  assign n29826 = pi3160 & pi3475;
  assign po3335 = n29825 | n29826;
  assign n29828 = ~pi3160 & pi3164;
  assign n29829 = pi3160 & pi3492;
  assign po3336 = n29828 | n29829;
  assign n29831 = ~pi3160 & pi3165;
  assign n29832 = pi3160 & pi3496;
  assign po3337 = n29831 | n29832;
  assign n29834 = ~pi3160 & pi3166;
  assign n29835 = pi3160 & pi3476;
  assign po3338 = n29834 | n29835;
  assign n29837 = ~pi3160 & pi3168;
  assign n29838 = pi3160 & pi3485;
  assign po3340 = n29837 | n29838;
  assign n29840 = ~pi3160 & pi3169;
  assign n29841 = pi3160 & pi3479;
  assign po3341 = n29840 | n29841;
  assign n29843 = ~pi3160 & pi3170;
  assign n29844 = pi3160 & pi3482;
  assign po3342 = n29843 | n29844;
  assign n29846 = ~pi3160 & pi3171;
  assign n29847 = pi3160 & pi3493;
  assign po3343 = n29846 | n29847;
  assign n29849 = ~pi3160 & pi3172;
  assign n29850 = pi3160 & pi3501;
  assign po3344 = n29849 | n29850;
  assign po3368 = pi3184 & ~pi3239;
  assign po3383 = pi1973 & pi3227;
  assign po3387 = pi1406 & ~pi2910;
  assign po0007 = 1'b1;
  assign po0203 = 1'b1;
  assign po0004 = ~pi0339;
  assign po0332 = ~po0335;
  assign po0423 = ~po0431;
  assign po0580 = ~pi0411;
  assign po0611 = ~po0645;
  assign po1400 = ~po1405;
  assign po2055 = ~po2158;
  assign po2150 = ~po2036;
  assign po3301 = ~pi3207;
  assign po3321 = ~pi3191;
  assign po3355 = ~pi3160;
  assign po3367 = ~pi1973;
  assign po3369 = ~pi1877;
  assign po3374 = ~pi0078;
  assign po3375 = ~pi1965;
  assign po3378 = ~pi1318;
  assign po3379 = ~pi0120;
  assign po3402 = ~pi1374;
  assign po3408 = ~pi1405;
  assign po3424 = ~pi0319;
  assign po3425 = ~pi1208;
  assign po3427 = ~pi1196;
  assign po3428 = ~pi1409;
  assign po3429 = ~pi1248;
  assign po3430 = ~pi0320;
  assign po3431 = ~pi1383;
  assign po3432 = ~pi1986;
  assign po3433 = ~pi1253;
  assign po3434 = ~pi2384;
  assign po3435 = ~pi2907;
  assign po3436 = ~pi0318;
  assign po3437 = ~pi1408;
  assign po3438 = ~pi2594;
  assign po3439 = ~pi1249;
  assign po3440 = ~pi2358;
  assign po3441 = ~pi1406;
  assign po3442 = ~pi1247;
  assign po3443 = ~pi1194;
  assign po0001 = pi0988;
  assign po0002 = pi1312;
  assign po0003 = pi1210;
  assign po0005 = pi0340;
  assign po0006 = pi0336;
  assign po0008 = pi2964;
  assign po0009 = pi3127;
  assign po0010 = pi3183;
  assign po0011 = pi1259;
  assign po0012 = pi1859;
  assign po0013 = pi3195;
  assign po0014 = pi1227;
  assign po0015 = pi1225;
  assign po0016 = pi1226;
  assign po0017 = pi3119;
  assign po0018 = pi0127;
  assign po0019 = pi0121;
  assign po0020 = pi0125;
  assign po0021 = pi1347;
  assign po0022 = pi0445;
  assign po0023 = pi0219;
  assign po0024 = pi0132;
  assign po0025 = pi0221;
  assign po0026 = pi0220;
  assign po0027 = pi0231;
  assign po0028 = pi0213;
  assign po0029 = pi0229;
  assign po0030 = pi0242;
  assign po0031 = pi0243;
  assign po0032 = pi0217;
  assign po0033 = pi0218;
  assign po0034 = pi0244;
  assign po0035 = pi0245;
  assign po0036 = pi0246;
  assign po0037 = pi0208;
  assign po0038 = pi0209;
  assign po0039 = pi0232;
  assign po0040 = pi0233;
  assign po0041 = pi0234;
  assign po0042 = pi0225;
  assign po0043 = pi0210;
  assign po0044 = pi0235;
  assign po0045 = pi0211;
  assign po0046 = pi0212;
  assign po0047 = pi0236;
  assign po0048 = pi0214;
  assign po0049 = pi0215;
  assign po0050 = pi0237;
  assign po0051 = pi0226;
  assign po0052 = pi0227;
  assign po0053 = pi0238;
  assign po0054 = pi0228;
  assign po0055 = pi0239;
  assign po0056 = pi0240;
  assign po0057 = pi0216;
  assign po0058 = pi0241;
  assign po0059 = pi0069;
  assign po0060 = pi0070;
  assign po0061 = pi0065;
  assign po0062 = pi0059;
  assign po0063 = pi0060;
  assign po0064 = pi0061;
  assign po0065 = pi0062;
  assign po0066 = pi0068;
  assign po0067 = pi0063;
  assign po0068 = pi0064;
  assign po0069 = pi0051;
  assign po0070 = pi0052;
  assign po0071 = pi0053;
  assign po0072 = pi0056;
  assign po0073 = pi0055;
  assign po0074 = pi0067;
  assign po0075 = pi0054;
  assign po0076 = pi0050;
  assign po0077 = pi0066;
  assign po0078 = pi0039;
  assign po0079 = pi0042;
  assign po0080 = pi0044;
  assign po0081 = pi0040;
  assign po0082 = pi0057;
  assign po0083 = pi0041;
  assign po0084 = pi0046;
  assign po0085 = pi0058;
  assign po0086 = pi0043;
  assign po0087 = pi0047;
  assign po0088 = pi0049;
  assign po0089 = pi0045;
  assign po0090 = pi0048;
  assign po0091 = pi0007;
  assign po0092 = pi0015;
  assign po0093 = pi0026;
  assign po0094 = pi0028;
  assign po0095 = pi0029;
  assign po0096 = pi0030;
  assign po0097 = pi0031;
  assign po0098 = pi0037;
  assign po0099 = pi0032;
  assign po0100 = pi0033;
  assign po0101 = pi0008;
  assign po0102 = pi0009;
  assign po0103 = pi0010;
  assign po0104 = pi0011;
  assign po0105 = pi0035;
  assign po0106 = pi0038;
  assign po0107 = pi0012;
  assign po0108 = pi0013;
  assign po0109 = pi0036;
  assign po0110 = pi0014;
  assign po0111 = pi0016;
  assign po0112 = pi0017;
  assign po0113 = pi0018;
  assign po0114 = pi0019;
  assign po0115 = pi0020;
  assign po0116 = pi0021;
  assign po0117 = pi0022;
  assign po0118 = pi0023;
  assign po0119 = pi0024;
  assign po0120 = pi0025;
  assign po0121 = pi0034;
  assign po0122 = pi0027;
  assign po0123 = pi0930;
  assign po0124 = pi0536;
  assign po0125 = pi0537;
  assign po0126 = pi0534;
  assign po0127 = pi0535;
  assign po0128 = pi0533;
  assign po0129 = pi0931;
  assign po0130 = pi0531;
  assign po0131 = pi0530;
  assign po0132 = pi0532;
  assign po0133 = pi0934;
  assign po0134 = pi0528;
  assign po0135 = pi0933;
  assign po0136 = pi0527;
  assign po0137 = pi0526;
  assign po0138 = pi0525;
  assign po0139 = pi0935;
  assign po0140 = pi0523;
  assign po0141 = pi0524;
  assign po0142 = pi0522;
  assign po0143 = pi0938;
  assign po0144 = pi0521;
  assign po0145 = pi0520;
  assign po0146 = pi0519;
  assign po0147 = pi0939;
  assign po0148 = pi0529;
  assign po0149 = pi0538;
  assign po0150 = pi0542;
  assign po0151 = pi0541;
  assign po0152 = pi0540;
  assign po0153 = pi0928;
  assign po0154 = pi0539;
  assign po0155 = pi0200;
  assign po0156 = pi0193;
  assign po0157 = pi0163;
  assign po0158 = pi0170;
  assign po0159 = pi0164;
  assign po0160 = pi0165;
  assign po0161 = pi0166;
  assign po0162 = pi0167;
  assign po0163 = pi0169;
  assign po0164 = pi0188;
  assign po0165 = pi0180;
  assign po0166 = pi0154;
  assign po0167 = pi0155;
  assign po0168 = pi0156;
  assign po0169 = pi0157;
  assign po0170 = pi0158;
  assign po0171 = pi0181;
  assign po0172 = pi0182;
  assign po0173 = pi0183;
  assign po0174 = pi0184;
  assign po0175 = pi0186;
  assign po0176 = pi0196;
  assign po0177 = pi0185;
  assign po0178 = pi0168;
  assign po0179 = pi0159;
  assign po0180 = pi0204;
  assign po0181 = pi0199;
  assign po0182 = pi0160;
  assign po0183 = pi0162;
  assign po0184 = pi0161;
  assign po0185 = pi0194;
  assign po0186 = pi0131;
  assign po0187 = pi0003;
  assign po0188 = pi0004;
  assign po0189 = pi0005;
  assign po0190 = pi0006;
  assign po0191 = pi2405;
  assign po0192 = pi2404;
  assign po0193 = pi1982;
  assign po0194 = pi1981;
  assign po0195 = pi0137;
  assign po0196 = pi1343;
  assign po0197 = pi0138;
  assign po0198 = pi0140;
  assign po0199 = pi0000;
  assign po0200 = pi0080;
  assign po0201 = pi0001;
  assign po0202 = pi3368;
  assign po0204 = pi3359;
  assign po0207 = pi3367;
  assign po0720 = po0719;
  assign po0721 = po0719;
  assign po0722 = po0719;
  assign po0723 = po0719;
  assign po0724 = po0719;
  assign po0725 = po0719;
  assign po0726 = po0719;
  assign po0727 = po0719;
  assign po0728 = po0719;
  assign po0729 = po0719;
  assign po0730 = po0719;
  assign po3159 = pi3122;
  assign po3298 = pi3140;
  assign po3299 = pi3137;
  assign po3303 = pi3117;
  assign po3317 = pi3173;
  assign po3322 = pi3181;
  assign po3328 = pi3249;
  assign po3345 = pi3211;
  assign po3346 = pi3202;
  assign po3347 = pi3196;
  assign po3348 = pi3215;
  assign po3349 = pi3221;
  assign po3350 = pi3212;
  assign po3352 = pi3197;
  assign po3353 = pi3160;
  assign po3354 = pi3236;
  assign po3356 = pi3234;
  assign po3357 = pi3250;
  assign po3358 = pi3248;
  assign po3359 = pi3230;
  assign po3360 = pi3251;
  assign po3361 = pi3231;
  assign po3362 = pi3123;
  assign po3363 = pi3238;
  assign po3364 = pi3267;
  assign po3365 = pi3265;
  assign po3366 = pi3270;
  assign po3370 = pi3257;
  assign po3371 = pi3252;
  assign po3372 = pi1353;
  assign po3373 = pi3027;
  assign po3376 = pi3256;
  assign po3377 = pi3264;
  assign po3380 = pi3258;
  assign po3381 = pi3261;
  assign po3382 = pi3269;
  assign po3385 = pi3253;
  assign po3386 = pi3255;
  assign po3388 = pi3260;
  assign po3389 = pi3266;
  assign po3390 = pi3263;
  assign po3391 = pi3268;
  assign po3392 = pi3259;
  assign po3394 = pi3262;
  assign po3395 = pi3271;
  assign po3396 = pi3284;
  assign po3397 = pi3331;
  assign po3398 = pi3339;
  assign po3399 = pi1973;
  assign po3400 = pi3302;
  assign po3401 = pi3323;
  assign po3403 = pi1685;
  assign po3404 = pi3342;
  assign po3405 = pi3324;
  assign po3406 = pi2908;
  assign po3407 = pi3285;
  assign po3409 = pi3309;
  assign po3410 = pi2918;
  assign po3411 = pi3184;
  assign po3412 = pi3289;
  assign po3413 = pi3317;
  assign po3414 = pi3296;
  assign po3415 = pi3322;
  assign po3416 = pi3319;
  assign po3417 = pi3352;
  assign po3418 = pi3338;
  assign po3419 = pi3308;
  assign po3420 = pi3297;
  assign po3421 = pi3325;
  assign po3422 = pi3345;
  assign po3423 = pi1400;
  assign po3426 = pi0076;
  assign po3444 = pi3272;
  assign po3445 = pi3273;
  assign po3446 = pi3274;
  assign po3447 = pi3275;
  assign po3448 = pi3276;
  assign po3449 = pi3277;
  assign po3450 = pi3278;
  assign po3451 = pi3279;
  assign po3452 = pi3280;
  assign po3453 = pi3281;
  assign po3454 = pi3282;
  assign po3455 = pi3283;
  assign po3456 = pi1214;
  assign po3457 = pi2936;
  assign po3458 = pi3455;
  assign po3459 = pi3453;
  assign po3460 = pi3452;
  assign po3461 = pi1222;
  assign po3462 = pi3457;
  assign po3463 = pi3291;
  assign po3464 = pi3292;
  assign po3465 = pi3448;
  assign po3466 = pi3294;
  assign po3467 = pi3467;
  assign po3468 = pi1709;
  assign po3469 = pi3182;
  assign po3470 = pi3461;
  assign po3471 = pi3472;
  assign po3472 = pi3300;
  assign po3473 = pi3301;
  assign po3474 = pi1175;
  assign po3475 = pi3303;
  assign po3476 = pi3304;
  assign po3477 = pi3305;
  assign po3478 = pi3306;
  assign po3479 = pi3307;
  assign po3480 = pi1712;
  assign po3481 = pi1172;
  assign po3482 = pi3310;
  assign po3483 = pi3446;
  assign po3484 = pi3312;
  assign po3485 = pi3450;
  assign po3486 = pi3458;
  assign po3487 = pi3459;
  assign po3488 = pi3443;
  assign po3489 = pi3468;
  assign po3490 = pi1589;
  assign po3491 = pi3464;
  assign po3492 = pi1404;
  assign po3493 = pi2945;
  assign po3494 = pi1215;
  assign po3495 = pi2948;
  assign po3496 = pi3465;
  assign po3497 = pi3327;
  assign po3498 = pi3454;
  assign po3499 = pi3329;
  assign po3500 = pi3463;
  assign po3501 = pi2935;
  assign po3502 = pi3332;
  assign po3503 = pi3462;
  assign po3504 = pi3334;
  assign po3505 = pi3451;
  assign po3506 = pi3466;
  assign po3507 = pi3449;
  assign po3508 = pi1362;
  assign po3509 = pi1153;
  assign po3510 = pi3456;
  assign po3511 = pi3473;
  assign po3512 = pi1166;
  assign po3513 = pi3442;
  assign po3514 = pi3344;
  assign po3515 = pi3210;
  assign po3516 = pi3445;
  assign po3517 = pi3460;
  assign po3518 = pi3174;
  assign po3519 = pi3469;
  assign po3520 = pi3470;
  assign po3521 = pi1403;
  assign po3522 = pi3447;
  assign po3523 = pi3471;
  assign po3524 = pi3444;
  assign po3525 = pi3356;
  assign po3526 = pi3357;
  assign po3527 = pi3358;
endmodule


