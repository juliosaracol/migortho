module top (
            pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518, pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526, pi3527, pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535, pi3536, pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544, pi3545, pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553, pi3554, pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562, pi3563, pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571, pi3572, pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580, pi3581, pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589, pi3590, pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598, pi3599, pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607, pi3608, pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616, pi3617, pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625, pi3626, pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634, pi3635, pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643, pi3644, pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652, pi3653, pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661, pi3662, pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670, pi3671, pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679, pi3680, pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688, pi3689, pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697, pi3698, pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706, pi3707, pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715, pi3716, pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724, pi3725, pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733, pi3734, pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742, pi3743, pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751, pi3752, pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760, pi3761, pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769, pi3770, pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778, pi3779, pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787, pi3788, pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796, pi3797, pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805, pi3806, pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814, pi3815, pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823, pi3824, pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832, pi3833, pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841, pi3842, pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850, pi3851, pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859, pi3860, pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868, pi3869, pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877, pi3878, pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886, pi3887, pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895, pi3896, pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904, pi3905, pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913, pi3914, pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922, pi3923, pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931, pi3932, pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940, pi3941, pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949, pi3950, pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958, pi3959, pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967, pi3968, pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976, pi3977, pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985, pi3986, pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994, pi3995, pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003, pi4004, pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012, pi4013, pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021, pi4022, pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030, pi4031, pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039, pi4040, pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048, pi4049, pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057, pi4058, pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066, pi4067, pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075, pi4076, pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084, pi4085, pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093, pi4094, pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102, pi4103, pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111, pi4112, pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120, pi4121, pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129, pi4130, pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138, pi4139, pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147, pi4148, pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156, pi4157, pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165, pi4166, pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174, pi4175, pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183, pi4184, pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192, pi4193, pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201, pi4202, pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210, pi4211, pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219, pi4220, pi4221, pi4222, pi4223, pi4224, pi4225, pi4226, pi4227, pi4228, pi4229, pi4230, pi4231, pi4232, pi4233, pi4234, pi4235, pi4236, pi4237, pi4238, pi4239, pi4240, pi4241, pi4242, pi4243, pi4244, pi4245, pi4246, pi4247, pi4248, pi4249, pi4250, pi4251, pi4252, pi4253, pi4254, pi4255, pi4256, pi4257, pi4258, pi4259, pi4260, pi4261, pi4262, pi4263, pi4264, pi4265, pi4266, pi4267, pi4268, pi4269, pi4270, pi4271, pi4272, pi4273, pi4274, pi4275, pi4276, pi4277, pi4278, pi4279, pi4280, pi4281, pi4282, pi4283, pi4284, pi4285, pi4286, pi4287, pi4288, pi4289, pi4290, pi4291, pi4292, pi4293, pi4294, pi4295, pi4296, pi4297, pi4298, pi4299, pi4300, pi4301, pi4302, pi4303, pi4304, pi4305, pi4306, pi4307, pi4308, pi4309, pi4310, pi4311, pi4312, pi4313, pi4314, pi4315, pi4316, pi4317, pi4318, pi4319, pi4320, pi4321, pi4322, pi4323, pi4324, pi4325, pi4326, pi4327, pi4328, pi4329, pi4330, pi4331, pi4332, pi4333, pi4334, pi4335, pi4336, pi4337, pi4338, pi4339, pi4340, pi4341, pi4342, pi4343, pi4344, pi4345, pi4346, pi4347, pi4348, pi4349, pi4350, pi4351, pi4352, pi4353, pi4354, pi4355, pi4356, pi4357, pi4358, pi4359, pi4360, pi4361, pi4362, pi4363, pi4364, pi4365, pi4366, pi4367, pi4368, pi4369, pi4370, pi4371, pi4372, pi4373, pi4374, pi4375, pi4376, pi4377, pi4378, pi4379, pi4380, pi4381, pi4382, pi4383, pi4384, pi4385, pi4386, pi4387, pi4388, pi4389, pi4390, pi4391, pi4392, pi4393, pi4394, pi4395, pi4396, pi4397, pi4398, pi4399, pi4400, pi4401, pi4402, pi4403, pi4404, pi4405, pi4406, pi4407, pi4408, pi4409, pi4410, pi4411, pi4412, pi4413, pi4414, pi4415, pi4416, pi4417, pi4418, pi4419, pi4420, pi4421, pi4422, pi4423, pi4424, pi4425, pi4426, pi4427, pi4428, pi4429, pi4430, pi4431, pi4432, pi4433, pi4434, pi4435, pi4436, pi4437, pi4438, pi4439, pi4440, pi4441, pi4442, pi4443, pi4444, pi4445, pi4446, pi4447, pi4448, pi4449, pi4450, pi4451, pi4452, pi4453, pi4454, pi4455, pi4456, pi4457, pi4458, pi4459, pi4460, pi4461, pi4462, pi4463, pi4464, pi4465, pi4466, pi4467, pi4468, pi4469, pi4470, pi4471, pi4472, pi4473, pi4474, pi4475, pi4476, pi4477, pi4478, pi4479, pi4480, pi4481, pi4482, pi4483, pi4484, pi4485, pi4486, pi4487, pi4488, pi4489, pi4490, pi4491, pi4492, pi4493, pi4494, pi4495, pi4496, pi4497, pi4498, pi4499, pi4500, pi4501, pi4502, pi4503, pi4504, pi4505, pi4506, pi4507, pi4508, pi4509, pi4510, pi4511, pi4512, pi4513, pi4514, pi4515, pi4516, pi4517, pi4518, pi4519, pi4520, pi4521, pi4522, pi4523, pi4524, pi4525, pi4526, pi4527, pi4528, pi4529, pi4530, pi4531, pi4532, pi4533, pi4534, pi4535, pi4536, pi4537, pi4538, pi4539, pi4540, pi4541, pi4542, pi4543, pi4544, pi4545, pi4546, pi4547, pi4548, pi4549, pi4550, pi4551, pi4552, pi4553, pi4554, pi4555, pi4556, pi4557, pi4558, pi4559, pi4560, pi4561, pi4562, pi4563, pi4564, pi4565, pi4566, pi4567, pi4568, pi4569, pi4570, pi4571, pi4572, pi4573, pi4574, pi4575, pi4576, pi4577, pi4578, pi4579, pi4580, pi4581, pi4582, pi4583, pi4584, pi4585, pi4586, pi4587, pi4588, pi4589, pi4590, pi4591, pi4592, pi4593, pi4594, pi4595, pi4596, pi4597, pi4598, pi4599, pi4600, pi4601, pi4602, pi4603, pi4604, pi4605, pi4606, pi4607, pi4608, pi4609, pi4610, pi4611, pi4612, pi4613, pi4614, pi4615, pi4616, pi4617, pi4618, pi4619, pi4620, pi4621, pi4622, pi4623, pi4624, pi4625, pi4626, pi4627, pi4628, pi4629, pi4630, pi4631, pi4632, pi4633, pi4634, pi4635, pi4636, pi4637, pi4638, pi4639, pi4640, pi4641, pi4642, pi4643, pi4644, pi4645, pi4646, pi4647, pi4648, pi4649, pi4650, pi4651, pi4652, pi4653, pi4654, pi4655, pi4656, pi4657, pi4658, pi4659, pi4660, pi4661, pi4662, pi4663, pi4664, pi4665, pi4666, pi4667, pi4668, pi4669, pi4670, pi4671, pi4672, pi4673, pi4674, pi4675, pi4676, pi4677, pi4678, pi4679, pi4680, pi4681, pi4682, pi4683, pi4684, pi4685, pi4686, pi4687, pi4688, pi4689, pi4690, pi4691, pi4692, pi4693, pi4694, pi4695, pi4696, pi4697, pi4698, pi4699, pi4700, pi4701, pi4702, pi4703, pi4704, pi4705, pi4706, pi4707, pi4708, pi4709, pi4710, pi4711, pi4712, pi4713, pi4714, pi4715, pi4716, pi4717, pi4718, pi4719, pi4720, pi4721, pi4722, pi4723, pi4724, pi4725, pi4726, pi4727, pi4728, pi4729, pi4730, pi4731, pi4732, pi4733, pi4734, pi4735, pi4736, pi4737, pi4738, pi4739, pi4740, pi4741, pi4742, pi4743, pi4744, pi4745, pi4746, pi4747, pi4748, pi4749, pi4750, pi4751, pi4752, pi4753, pi4754, pi4755, pi4756, pi4757, pi4758, pi4759, pi4760, pi4761, pi4762, pi4763, pi4764, pi4765, pi4766, pi4767, pi4768, pi4769, pi4770, pi4771, pi4772, pi4773, pi4774, pi4775, pi4776, pi4777, pi4778, pi4779, pi4780, pi4781, pi4782, pi4783, pi4784, pi4785, pi4786, pi4787, pi4788, pi4789, pi4790, pi4791, pi4792, pi4793, pi4794, pi4795, pi4796, pi4797, pi4798, pi4799, pi4800, pi4801, pi4802, pi4803, pi4804, pi4805, pi4806, pi4807, pi4808, pi4809, pi4810, pi4811, pi4812, pi4813, pi4814, pi4815, pi4816, pi4817, pi4818, pi4819, pi4820, pi4821, pi4822, pi4823, pi4824, pi4825, pi4826, pi4827, pi4828, pi4829, pi4830, pi4831, pi4832, pi4833, pi4834, pi4835, pi4836, pi4837, pi4838, pi4839, pi4840, pi4841, pi4842, pi4843, pi4844, pi4845, pi4846, pi4847, pi4848, pi4849, pi4850, pi4851, pi4852, pi4853, pi4854, pi4855, pi4856, pi4857, pi4858, pi4859, pi4860, pi4861, pi4862, pi4863, pi4864, pi4865, pi4866, pi4867, pi4868, pi4869, pi4870, pi4871, pi4872, pi4873, pi4874, pi4875, pi4876, pi4877, pi4878, pi4879, pi4880, pi4881, pi4882, pi4883, pi4884, pi4885, pi4886, pi4887, pi4888, pi4889, pi4890, pi4891, pi4892, pi4893, pi4894, pi4895, pi4896, pi4897, pi4898, pi4899, pi4900, pi4901, pi4902, pi4903, pi4904, pi4905, pi4906, pi4907, pi4908, pi4909, pi4910, pi4911, pi4912, pi4913, pi4914, pi4915, pi4916, pi4917, pi4918, pi4919, pi4920, pi4921, pi4922, pi4923, pi4924, pi4925, pi4926, pi4927, pi4928, pi4929, pi4930, pi4931, pi4932, pi4933, pi4934, pi4935, pi4936, pi4937, pi4938, pi4939, pi4940, pi4941, pi4942, pi4943, pi4944, pi4945, pi4946, pi4947, pi4948, pi4949, pi4950, pi4951, pi4952, pi4953, pi4954, pi4955, pi4956, pi4957, pi4958, pi4959, pi4960, pi4961, pi4962, pi4963, pi4964, pi4965, pi4966, pi4967, pi4968, pi4969, pi4970, pi4971, pi4972, pi4973, pi4974, pi4975, pi4976, pi4977, pi4978, pi4979, pi4980, pi4981, pi4982, pi4983, pi4984, pi4985, pi4986, pi4987, pi4988, pi4989, pi4990, pi4991, pi4992, pi4993, pi4994, pi4995, pi4996, pi4997, pi4998, pi4999, pi5000, pi5001, pi5002, pi5003, pi5004, pi5005, pi5006, pi5007, pi5008, pi5009, pi5010, pi5011, pi5012, pi5013, pi5014, pi5015, pi5016, pi5017, pi5018, pi5019, pi5020, pi5021, pi5022, pi5023, pi5024, pi5025, pi5026, pi5027, pi5028, pi5029, pi5030, pi5031, pi5032, pi5033, pi5034, pi5035, pi5036, pi5037, pi5038, pi5039, pi5040, pi5041, pi5042, pi5043, pi5044, pi5045, pi5046, pi5047, pi5048, pi5049, pi5050, pi5051, pi5052, pi5053, pi5054, pi5055, pi5056, pi5057, pi5058, pi5059, pi5060, pi5061, pi5062, pi5063, pi5064, pi5065, pi5066, pi5067, pi5068, pi5069, pi5070, pi5071, pi5072, pi5073, pi5074, pi5075, pi5076, pi5077, pi5078, pi5079, pi5080, pi5081, pi5082, pi5083, pi5084, pi5085, pi5086, pi5087, pi5088, pi5089, pi5090, pi5091, pi5092, pi5093, pi5094, pi5095, pi5096, pi5097, pi5098, pi5099, pi5100, pi5101, pi5102, pi5103, pi5104, pi5105, pi5106, pi5107, pi5108, pi5109, pi5110, pi5111, pi5112, pi5113, pi5114, pi5115, pi5116, pi5117, pi5118, pi5119, pi5120, pi5121, pi5122, pi5123, pi5124, pi5125, pi5126, pi5127, pi5128, pi5129, pi5130, pi5131, pi5132, pi5133, pi5134, pi5135, pi5136, pi5137, pi5138, pi5139, pi5140, pi5141, pi5142, pi5143, pi5144, pi5145, pi5146, pi5147, pi5148, pi5149, pi5150, pi5151, pi5152, pi5153, pi5154, pi5155, pi5156, pi5157, pi5158, pi5159, pi5160, pi5161, pi5162, pi5163, pi5164, pi5165, pi5166, pi5167, pi5168, pi5169, pi5170, pi5171, pi5172, pi5173, pi5174, pi5175, pi5176, pi5177, pi5178, pi5179, pi5180, pi5181, pi5182, pi5183, pi5184, pi5185, pi5186, pi5187, pi5188, pi5189, pi5190, pi5191, pi5192, pi5193, pi5194, pi5195, pi5196, pi5197, pi5198, pi5199, pi5200, pi5201, pi5202, pi5203, pi5204, pi5205, pi5206, pi5207, pi5208, pi5209, pi5210, pi5211, pi5212, pi5213, pi5214, pi5215, pi5216, pi5217, pi5218, pi5219, pi5220, pi5221, pi5222, pi5223, pi5224, pi5225, pi5226, pi5227, pi5228, pi5229, pi5230, pi5231, pi5232, pi5233, pi5234, pi5235, pi5236, pi5237, pi5238, pi5239, pi5240, pi5241, pi5242, pi5243, pi5244, pi5245, pi5246, pi5247, pi5248, pi5249, pi5250, pi5251, pi5252, pi5253, pi5254, pi5255, pi5256, pi5257, pi5258, pi5259, pi5260, pi5261, pi5262, pi5263, pi5264, pi5265, pi5266, pi5267, pi5268, pi5269, pi5270, pi5271, pi5272, pi5273, pi5274, pi5275, pi5276, pi5277, pi5278, pi5279, pi5280, pi5281, pi5282, pi5283, pi5284, pi5285, pi5286, pi5287, pi5288, pi5289, pi5290, pi5291, pi5292, pi5293, pi5294, pi5295, pi5296, pi5297, pi5298, pi5299, pi5300, pi5301, pi5302, pi5303, pi5304, pi5305, pi5306, pi5307, pi5308, pi5309, pi5310, pi5311, pi5312, pi5313, pi5314, pi5315, pi5316, pi5317, pi5318, pi5319, pi5320, pi5321, pi5322, pi5323, pi5324, pi5325, pi5326, pi5327, pi5328, pi5329, pi5330, pi5331, pi5332, pi5333, pi5334, pi5335, pi5336, pi5337, pi5338, pi5339, pi5340, pi5341, pi5342, pi5343, pi5344, pi5345, pi5346, pi5347, pi5348, pi5349, pi5350, pi5351, pi5352, pi5353, pi5354, pi5355, pi5356, pi5357, pi5358, pi5359, pi5360, pi5361, pi5362, pi5363, pi5364, pi5365, pi5366, pi5367, pi5368, pi5369, pi5370, pi5371, pi5372, pi5373, pi5374, pi5375, pi5376, pi5377, pi5378, pi5379, pi5380, pi5381, pi5382, pi5383, pi5384, pi5385, pi5386, pi5387, pi5388, pi5389, pi5390, pi5391, pi5392, pi5393, pi5394, pi5395, pi5396, pi5397, pi5398, pi5399, pi5400, pi5401, pi5402, pi5403, pi5404, pi5405, pi5406, pi5407, pi5408, pi5409, pi5410, pi5411, pi5412, pi5413, pi5414, pi5415, pi5416, pi5417, pi5418, pi5419, pi5420, pi5421, pi5422, pi5423, pi5424, pi5425, pi5426, pi5427, pi5428, pi5429, pi5430, pi5431, pi5432, pi5433, pi5434, pi5435, pi5436, pi5437, pi5438, pi5439, pi5440, pi5441, pi5442, pi5443, pi5444, pi5445, pi5446, pi5447, pi5448, pi5449, pi5450, pi5451, pi5452, pi5453, pi5454, pi5455, pi5456, pi5457, pi5458, pi5459, pi5460, pi5461, pi5462, pi5463, pi5464, pi5465, pi5466, pi5467, pi5468, pi5469, pi5470, pi5471, pi5472, pi5473, pi5474, pi5475, pi5476, pi5477, pi5478, pi5479, pi5480, pi5481, pi5482, pi5483, pi5484, pi5485, pi5486, pi5487, pi5488, pi5489, pi5490, pi5491, pi5492, pi5493, pi5494, pi5495, pi5496, pi5497, pi5498, pi5499, pi5500, pi5501, pi5502, pi5503, pi5504, pi5505, pi5506, pi5507, pi5508, pi5509, pi5510, pi5511, pi5512, pi5513, pi5514, pi5515, pi5516, pi5517, pi5518, pi5519, pi5520, pi5521, pi5522, pi5523, pi5524, pi5525, pi5526, pi5527, pi5528, pi5529, pi5530, pi5531, pi5532, pi5533, pi5534, pi5535, pi5536, pi5537, pi5538, pi5539, pi5540, pi5541, pi5542, pi5543, pi5544, pi5545, pi5546, pi5547, pi5548, pi5549, pi5550, pi5551, pi5552, pi5553, pi5554, pi5555, pi5556, pi5557, pi5558, pi5559, pi5560, pi5561, pi5562, pi5563, pi5564, pi5565, pi5566, pi5567, pi5568, pi5569, pi5570, pi5571, pi5572, pi5573, pi5574, pi5575, pi5576, pi5577, pi5578, pi5579, pi5580, pi5581, pi5582, pi5583, pi5584, pi5585, pi5586, pi5587, pi5588, pi5589, pi5590, pi5591, pi5592, pi5593, pi5594, pi5595, pi5596, pi5597, pi5598, pi5599, pi5600, pi5601, pi5602, pi5603, pi5604, pi5605, pi5606, pi5607, pi5608, pi5609, pi5610, pi5611, pi5612, pi5613, pi5614, pi5615, pi5616, pi5617, pi5618, pi5619, pi5620, pi5621, pi5622, pi5623, pi5624, pi5625, pi5626, pi5627, pi5628, pi5629, pi5630, pi5631, pi5632, pi5633, pi5634, pi5635, pi5636, pi5637, pi5638, pi5639, pi5640, pi5641, pi5642, pi5643, pi5644, pi5645, pi5646, pi5647, pi5648, pi5649, pi5650, pi5651, pi5652, pi5653, pi5654, pi5655, pi5656, pi5657, pi5658, pi5659, pi5660, pi5661, pi5662, pi5663, pi5664, pi5665, pi5666, pi5667, pi5668, pi5669, pi5670, pi5671, pi5672, pi5673, pi5674, pi5675, pi5676, pi5677, pi5678, pi5679, pi5680, pi5681, pi5682, pi5683, pi5684, pi5685, pi5686, pi5687, pi5688, pi5689, pi5690, pi5691, pi5692, pi5693, pi5694, pi5695, pi5696, pi5697, pi5698, pi5699, pi5700, pi5701, pi5702, pi5703, pi5704, pi5705, pi5706, pi5707, pi5708, pi5709, pi5710, pi5711, pi5712, pi5713, pi5714, pi5715, pi5716, pi5717, pi5718, pi5719, pi5720, pi5721, pi5722, pi5723, pi5724, pi5725, pi5726, pi5727, pi5728, pi5729, pi5730, pi5731, pi5732, pi5733, pi5734, pi5735, pi5736, pi5737, pi5738, pi5739, pi5740, pi5741, pi5742, pi5743, pi5744, pi5745, pi5746, pi5747, pi5748, pi5749, pi5750, pi5751, pi5752, pi5753, pi5754, pi5755, pi5756, pi5757, pi5758, pi5759, pi5760, pi5761, pi5762, pi5763, pi5764, pi5765, pi5766, pi5767, pi5768, pi5769, pi5770, pi5771, pi5772, pi5773, pi5774, pi5775, pi5776, pi5777, pi5778, pi5779, pi5780, pi5781, pi5782, pi5783, pi5784, pi5785, pi5786, pi5787, pi5788, pi5789, pi5790, pi5791, pi5792, pi5793, pi5794, pi5795, pi5796, pi5797, pi5798, pi5799, pi5800, pi5801, pi5802, pi5803, pi5804, pi5805, pi5806, pi5807, pi5808, pi5809, pi5810, pi5811, pi5812, pi5813, pi5814, pi5815, pi5816, pi5817, pi5818, pi5819, pi5820, pi5821, pi5822, pi5823, pi5824, pi5825, pi5826, pi5827, pi5828, pi5829, pi5830, pi5831, pi5832, pi5833, pi5834, pi5835, pi5836, pi5837, pi5838, pi5839, pi5840, pi5841, pi5842, pi5843, pi5844, pi5845, pi5846, pi5847, pi5848, pi5849, pi5850, pi5851, pi5852, pi5853, pi5854, pi5855, pi5856, pi5857, pi5858, pi5859, pi5860, pi5861, pi5862, pi5863, pi5864, pi5865, pi5866, pi5867, pi5868, pi5869, pi5870, pi5871, pi5872, pi5873, pi5874, pi5875, pi5876, pi5877, pi5878, pi5879, pi5880, pi5881, pi5882, pi5883, pi5884, pi5885, pi5886, pi5887, pi5888, pi5889, pi5890, pi5891, pi5892, pi5893, pi5894, pi5895, pi5896, pi5897, pi5898, pi5899, pi5900, pi5901, pi5902, pi5903, pi5904, pi5905, pi5906, pi5907, pi5908, pi5909, pi5910, pi5911, pi5912, pi5913, pi5914, pi5915, pi5916, pi5917, pi5918, pi5919, pi5920, pi5921, pi5922, pi5923, pi5924, pi5925, pi5926, pi5927, pi5928, pi5929, pi5930, pi5931, pi5932, pi5933, pi5934, pi5935, pi5936, pi5937, pi5938, pi5939, pi5940, pi5941, pi5942, pi5943, pi5944, pi5945, pi5946, pi5947, pi5948, pi5949, pi5950, pi5951, pi5952, pi5953, pi5954, pi5955, pi5956, pi5957, pi5958, pi5959, pi5960, pi5961, pi5962, pi5963, pi5964, pi5965, pi5966, pi5967, pi5968, pi5969, pi5970, pi5971, pi5972, pi5973, pi5974, pi5975, pi5976, pi5977, pi5978, pi5979, pi5980, pi5981, pi5982, pi5983, pi5984, pi5985, pi5986, pi5987, pi5988, pi5989, pi5990, pi5991, pi5992, pi5993, pi5994, pi5995, pi5996, pi5997, pi5998, pi5999, pi6000, pi6001, pi6002, pi6003, pi6004, pi6005, pi6006, pi6007, pi6008, pi6009, pi6010, pi6011, pi6012, pi6013, pi6014, pi6015, pi6016, pi6017, pi6018, pi6019, pi6020, pi6021, pi6022, pi6023, pi6024, pi6025, pi6026, pi6027, pi6028, pi6029, pi6030, pi6031, pi6032, pi6033, pi6034, pi6035, pi6036, pi6037, pi6038, pi6039, pi6040, pi6041, pi6042, pi6043, pi6044, pi6045, pi6046, pi6047, pi6048, pi6049, pi6050, pi6051, pi6052, pi6053, pi6054, pi6055, pi6056, pi6057, pi6058, pi6059, pi6060, pi6061, pi6062, pi6063, pi6064, pi6065, pi6066, pi6067, pi6068, pi6069, pi6070, pi6071, pi6072, pi6073, pi6074, pi6075, pi6076, pi6077, pi6078, pi6079, pi6080, pi6081, pi6082, pi6083, pi6084, pi6085, pi6086, pi6087, pi6088, pi6089, pi6090, pi6091, pi6092, pi6093, pi6094, pi6095, pi6096, pi6097, pi6098, pi6099, pi6100, pi6101, pi6102, pi6103, pi6104, pi6105, pi6106, pi6107, pi6108, pi6109, pi6110, pi6111, pi6112, pi6113, pi6114, pi6115, pi6116, pi6117, pi6118, pi6119, pi6120, pi6121, pi6122, pi6123, pi6124, pi6125, pi6126, pi6127, pi6128, pi6129, pi6130, pi6131, pi6132, pi6133, pi6134, pi6135, pi6136, pi6137, pi6138, pi6139, pi6140, pi6141, pi6142, pi6143, pi6144, pi6145, pi6146, pi6147, pi6148, pi6149, pi6150, pi6151, pi6152, pi6153, pi6154, pi6155, pi6156, pi6157, pi6158, pi6159, pi6160, pi6161, pi6162, pi6163, pi6164, pi6165, pi6166, pi6167, pi6168, pi6169, pi6170, pi6171, pi6172, pi6173, pi6174, pi6175, pi6176, pi6177, pi6178, pi6179, pi6180, pi6181, pi6182, pi6183, pi6184, pi6185, pi6186, pi6187, pi6188, pi6189, pi6190, pi6191, pi6192, pi6193, pi6194, pi6195, pi6196, pi6197, pi6198, pi6199, pi6200, pi6201, pi6202, pi6203, pi6204, pi6205, pi6206, pi6207, pi6208, pi6209, pi6210, pi6211, pi6212, pi6213, pi6214, pi6215, pi6216, pi6217, pi6218, pi6219, pi6220, pi6221, pi6222, pi6223, pi6224, pi6225, pi6226, pi6227, pi6228, pi6229, pi6230, pi6231, pi6232, pi6233, pi6234, pi6235, pi6236, pi6237, pi6238, pi6239, pi6240, pi6241, pi6242, pi6243, pi6244, pi6245, pi6246, pi6247, pi6248, pi6249, pi6250, pi6251, pi6252, pi6253, pi6254, pi6255, pi6256, pi6257, pi6258, pi6259, pi6260, pi6261, pi6262, pi6263, pi6264, pi6265, pi6266, pi6267, pi6268, pi6269, pi6270, pi6271, pi6272, pi6273, pi6274, pi6275, pi6276, pi6277, pi6278, pi6279, pi6280, pi6281, pi6282, pi6283, pi6284, pi6285, pi6286, pi6287, pi6288, pi6289, pi6290, pi6291, pi6292, pi6293, pi6294, pi6295, pi6296, pi6297, pi6298, pi6299, pi6300, pi6301, pi6302, pi6303, pi6304, pi6305, pi6306, pi6307, pi6308, pi6309, pi6310, pi6311, pi6312, pi6313, pi6314, pi6315, pi6316, pi6317, pi6318, pi6319, pi6320, pi6321, pi6322, pi6323, pi6324, pi6325, pi6326, pi6327, pi6328, pi6329, pi6330, pi6331, pi6332, pi6333, pi6334, pi6335, pi6336, pi6337, pi6338, pi6339, pi6340, pi6341, pi6342, pi6343, pi6344, pi6345, pi6346, pi6347, pi6348, pi6349, pi6350, pi6351, pi6352, pi6353, pi6354, pi6355, pi6356, pi6357, pi6358, pi6359, pi6360, pi6361, pi6362, pi6363, pi6364, pi6365, pi6366, pi6367, pi6368, pi6369, pi6370, pi6371, pi6372, pi6373, pi6374, pi6375, pi6376, pi6377, pi6378, pi6379, pi6380, pi6381, pi6382, pi6383, pi6384, pi6385, pi6386, pi6387, pi6388, pi6389, pi6390, pi6391, pi6392, pi6393, pi6394, pi6395, pi6396, pi6397, pi6398, pi6399, pi6400, pi6401, pi6402, pi6403, pi6404, pi6405, pi6406, pi6407, pi6408, pi6409, pi6410, pi6411, pi6412, pi6413, pi6414, pi6415, pi6416, pi6417, pi6418, pi6419, pi6420, pi6421, pi6422, pi6423, pi6424, pi6425, pi6426, pi6427, pi6428, pi6429, pi6430, pi6431, pi6432, pi6433, pi6434, pi6435, pi6436, pi6437, pi6438, pi6439, pi6440, pi6441, pi6442, pi6443, pi6444, pi6445, pi6446, pi6447, pi6448, pi6449, pi6450, pi6451, pi6452, pi6453, pi6454, pi6455, pi6456, pi6457, pi6458, pi6459, pi6460, pi6461, pi6462, pi6463, pi6464, pi6465, pi6466, pi6467, pi6468, pi6469, pi6470, pi6471, pi6472, pi6473, pi6474, pi6475, pi6476, pi6477, pi6478, pi6479, pi6480, pi6481, pi6482, pi6483, pi6484, pi6485, pi6486, pi6487, pi6488, pi6489, pi6490, pi6491, pi6492, pi6493, pi6494, pi6495, pi6496, pi6497, pi6498, pi6499, pi6500, pi6501, pi6502, pi6503, pi6504, pi6505, pi6506, pi6507, pi6508, pi6509, pi6510, pi6511, pi6512, pi6513, pi6514, pi6515, pi6516, pi6517, pi6518, pi6519, pi6520, pi6521, pi6522, pi6523, pi6524, pi6525, pi6526, pi6527, pi6528, pi6529, pi6530, pi6531, pi6532, pi6533, pi6534, pi6535, pi6536, pi6537, pi6538, pi6539, pi6540, pi6541, pi6542, pi6543, pi6544, pi6545, pi6546, pi6547, pi6548, pi6549, pi6550, pi6551, pi6552, pi6553, pi6554, pi6555, pi6556, pi6557, pi6558, pi6559, pi6560, pi6561, pi6562, pi6563, pi6564, pi6565, pi6566, pi6567, pi6568, pi6569, pi6570, pi6571, pi6572, pi6573, pi6574, pi6575, pi6576, pi6577, pi6578, pi6579, pi6580, pi6581, pi6582, pi6583, pi6584, pi6585, pi6586, pi6587, pi6588, pi6589, pi6590, pi6591, pi6592, pi6593, pi6594, pi6595, pi6596, pi6597, pi6598, pi6599, pi6600, pi6601, pi6602, pi6603, pi6604, pi6605, pi6606, pi6607, pi6608, pi6609, pi6610, pi6611, pi6612, pi6613, pi6614, pi6615, pi6616, pi6617, pi6618, pi6619, pi6620, pi6621, pi6622, pi6623, pi6624, pi6625, pi6626, pi6627, pi6628, pi6629, pi6630, pi6631, pi6632, pi6633, pi6634, pi6635, pi6636, pi6637, pi6638, pi6639, pi6640, pi6641, pi6642, pi6643, pi6644, pi6645, pi6646, pi6647, pi6648, pi6649, pi6650, pi6651, pi6652, pi6653, pi6654, pi6655, pi6656, pi6657, pi6658, pi6659, pi6660, pi6661, pi6662, pi6663, pi6664, pi6665, pi6666, pi6667, pi6668, pi6669, pi6670, pi6671, pi6672, pi6673, pi6674, pi6675, pi6676, pi6677, pi6678, pi6679, pi6680, pi6681, pi6682, pi6683, pi6684, pi6685, pi6686, pi6687, pi6688, pi6689, pi6690, pi6691, pi6692, pi6693, pi6694, pi6695, pi6696, pi6697, pi6698, pi6699, pi6700, pi6701, pi6702, pi6703, pi6704, pi6705, pi6706, pi6707, pi6708, pi6709, pi6710, pi6711, pi6712, pi6713, pi6714, pi6715, pi6716, pi6717, pi6718, pi6719, pi6720, pi6721, pi6722, pi6723, pi6724, pi6725, pi6726, pi6727, pi6728, pi6729, pi6730, pi6731, pi6732, pi6733, pi6734, pi6735, pi6736, pi6737, pi6738, pi6739, pi6740, pi6741, pi6742, pi6743, pi6744, pi6745, pi6746, pi6747, pi6748, pi6749, pi6750, pi6751, pi6752, pi6753, pi6754, pi6755, pi6756, pi6757, pi6758, pi6759, pi6760, pi6761, pi6762, pi6763, pi6764, pi6765, pi6766, pi6767, pi6768, pi6769, pi6770, pi6771, pi6772, pi6773, pi6774, pi6775, pi6776, pi6777, pi6778, pi6779, pi6780, pi6781, pi6782, pi6783, pi6784, pi6785, pi6786, pi6787, pi6788, pi6789, pi6790, pi6791, pi6792, pi6793, pi6794, pi6795, pi6796, pi6797, pi6798, pi6799, pi6800, pi6801, pi6802, pi6803, pi6804, pi6805, pi6806, pi6807, pi6808, pi6809, pi6810, pi6811, pi6812, pi6813, pi6814, pi6815, pi6816, pi6817, pi6818, pi6819, pi6820, pi6821, pi6822, pi6823, pi6824, pi6825, pi6826, pi6827, pi6828, pi6829, pi6830, pi6831, pi6832, pi6833, pi6834, pi6835, pi6836, pi6837, pi6838, pi6839, pi6840, pi6841, pi6842, pi6843, pi6844, pi6845, pi6846, pi6847, pi6848, pi6849, pi6850, pi6851, pi6852, pi6853, pi6854, pi6855, pi6856, pi6857, pi6858, pi6859, pi6860, pi6861, pi6862, pi6863, pi6864, pi6865, pi6866, pi6867, pi6868, pi6869, pi6870, pi6871, pi6872, pi6873, pi6874, pi6875, pi6876, pi6877, pi6878, pi6879, pi6880, pi6881, pi6882, pi6883, pi6884, pi6885, pi6886, pi6887, pi6888, pi6889, pi6890, pi6891, pi6892, pi6893, pi6894, pi6895, pi6896, pi6897, pi6898, pi6899, pi6900, pi6901, pi6902, pi6903, pi6904, pi6905, pi6906, pi6907, pi6908, pi6909, pi6910, pi6911, pi6912, pi6913, pi6914, pi6915, pi6916, pi6917, pi6918, pi6919, pi6920, pi6921, pi6922, pi6923, pi6924, pi6925, pi6926, pi6927, pi6928, pi6929, pi6930, pi6931, pi6932, pi6933, pi6934, pi6935, pi6936, pi6937, pi6938, pi6939, pi6940, pi6941, pi6942, pi6943, pi6944, pi6945, pi6946, pi6947, pi6948, pi6949, pi6950, pi6951, pi6952, pi6953, pi6954, pi6955, pi6956, pi6957, pi6958, pi6959, pi6960, pi6961, pi6962, pi6963, pi6964, pi6965, pi6966, pi6967, pi6968, pi6969, pi6970, pi6971, pi6972, pi6973, pi6974, pi6975, pi6976, pi6977, pi6978, pi6979, pi6980, pi6981, pi6982, pi6983, pi6984, pi6985, pi6986, pi6987, pi6988, pi6989, pi6990, pi6991, pi6992, pi6993, pi6994, pi6995, pi6996, pi6997, pi6998, pi6999, pi7000, pi7001, pi7002, pi7003, pi7004, pi7005, pi7006, pi7007, pi7008, pi7009, pi7010, pi7011, pi7012, pi7013, pi7014, pi7015, pi7016, pi7017, pi7018, pi7019, pi7020, pi7021, pi7022, pi7023, pi7024, pi7025, pi7026, pi7027, pi7028, pi7029, pi7030, pi7031, pi7032, pi7033, pi7034, pi7035, pi7036, pi7037, pi7038, pi7039, pi7040, pi7041, pi7042, pi7043, pi7044, pi7045, pi7046, pi7047, pi7048, pi7049, pi7050, pi7051, pi7052, pi7053, pi7054, pi7055, pi7056, pi7057, pi7058, pi7059, pi7060, pi7061, pi7062, pi7063, pi7064, pi7065, pi7066, pi7067, pi7068, pi7069, pi7070, pi7071, pi7072, pi7073, pi7074, pi7075, pi7076, pi7077, pi7078, pi7079, pi7080, pi7081, pi7082, pi7083, pi7084, pi7085, pi7086, pi7087, pi7088, pi7089, pi7090, pi7091, pi7092, pi7093, pi7094, pi7095, pi7096, pi7097, pi7098, pi7099, pi7100, pi7101, pi7102, pi7103, pi7104, pi7105, pi7106, pi7107, pi7108, pi7109, pi7110, pi7111, pi7112, pi7113, pi7114, pi7115, pi7116, pi7117, pi7118, pi7119, pi7120, pi7121, pi7122, pi7123, pi7124, pi7125, pi7126, pi7127, pi7128, pi7129, pi7130, pi7131, pi7132, pi7133, pi7134, pi7135, pi7136, pi7137, pi7138, pi7139, pi7140, pi7141, pi7142, pi7143, pi7144, pi7145, pi7146, pi7147, pi7148, pi7149, pi7150, pi7151, pi7152, pi7153, pi7154, pi7155, pi7156, pi7157, pi7158, pi7159, pi7160, pi7161, pi7162, pi7163, pi7164, pi7165, pi7166, pi7167, pi7168, pi7169, pi7170, pi7171, pi7172, pi7173, pi7174, pi7175, pi7176, pi7177, pi7178, pi7179, pi7180, pi7181, pi7182, pi7183, pi7184, pi7185, pi7186, pi7187, pi7188, pi7189, pi7190, pi7191, pi7192, pi7193, pi7194, pi7195, pi7196, pi7197, pi7198, pi7199, pi7200, pi7201, pi7202, pi7203, pi7204, pi7205, pi7206, pi7207, pi7208, pi7209, pi7210, pi7211, pi7212, pi7213, pi7214, pi7215, pi7216, pi7217, pi7218, pi7219, pi7220, pi7221, pi7222, pi7223, pi7224, pi7225, pi7226, pi7227, pi7228, pi7229, pi7230, pi7231, pi7232, pi7233, pi7234, pi7235, pi7236, pi7237, pi7238, pi7239, pi7240, pi7241, pi7242, pi7243, pi7244, pi7245, pi7246, pi7247, pi7248, pi7249, pi7250, pi7251, pi7252, pi7253, pi7254, pi7255, pi7256, pi7257, pi7258, pi7259, pi7260, pi7261, pi7262, pi7263, pi7264, pi7265, pi7266, pi7267, pi7268, pi7269, pi7270, pi7271, pi7272, pi7273, pi7274, pi7275, pi7276, pi7277, pi7278, pi7279, pi7280, pi7281, pi7282, pi7283, pi7284, pi7285, pi7286, pi7287, pi7288, pi7289, pi7290, pi7291, pi7292, pi7293, pi7294, pi7295, pi7296, pi7297, pi7298, pi7299, pi7300, pi7301, pi7302, pi7303, pi7304, pi7305, pi7306, pi7307, pi7308, pi7309, pi7310, pi7311, pi7312, pi7313, pi7314, pi7315, pi7316, pi7317, pi7318, pi7319, pi7320, pi7321, pi7322, pi7323, pi7324, pi7325, pi7326, pi7327, pi7328, pi7329, pi7330, pi7331, pi7332, pi7333, pi7334, pi7335, pi7336, pi7337, pi7338, pi7339, pi7340, pi7341, pi7342, pi7343, pi7344, pi7345, pi7346, pi7347, pi7348, pi7349, pi7350, pi7351, pi7352, pi7353, pi7354, pi7355, pi7356, pi7357, pi7358, pi7359, pi7360, pi7361, pi7362, pi7363, pi7364, pi7365, pi7366, pi7367, pi7368, pi7369, pi7370, pi7371, pi7372, pi7373, pi7374, pi7375, pi7376, pi7377, pi7378, pi7379, pi7380, pi7381, pi7382, pi7383, pi7384, pi7385, pi7386, pi7387, pi7388, pi7389, pi7390, pi7391, pi7392, pi7393, pi7394, pi7395, pi7396, pi7397, pi7398, pi7399, pi7400, pi7401, pi7402, pi7403, pi7404, pi7405, pi7406, pi7407, pi7408, pi7409, pi7410, pi7411, pi7412, pi7413, pi7414, pi7415, pi7416, pi7417, pi7418, pi7419, pi7420, pi7421, pi7422, pi7423, pi7424, pi7425, pi7426, pi7427, pi7428, pi7429, pi7430, pi7431, pi7432, pi7433, pi7434, pi7435, pi7436, pi7437, pi7438, pi7439, pi7440, pi7441, pi7442, pi7443, pi7444, pi7445, pi7446, pi7447, pi7448, pi7449, pi7450, pi7451, pi7452, pi7453, pi7454, pi7455, pi7456, pi7457, pi7458, pi7459, pi7460, pi7461, pi7462, pi7463, pi7464, pi7465, pi7466, pi7467, pi7468, pi7469, pi7470, pi7471, pi7472, pi7473, pi7474, pi7475, pi7476, pi7477, pi7478, pi7479, pi7480, pi7481, pi7482, pi7483, pi7484, pi7485, pi7486, pi7487, pi7488, pi7489, pi7490, pi7491, pi7492, pi7493, pi7494, pi7495, pi7496, pi7497, pi7498, pi7499, pi7500, pi7501, pi7502, pi7503, pi7504, pi7505, pi7506, pi7507, pi7508, pi7509, pi7510, pi7511, pi7512, pi7513, pi7514, pi7515, pi7516, pi7517, pi7518, pi7519, pi7520, pi7521, pi7522, pi7523, pi7524, pi7525, pi7526, pi7527, pi7528, pi7529, pi7530, pi7531, pi7532, pi7533, pi7534, pi7535, pi7536, pi7537, pi7538, pi7539, pi7540, pi7541, pi7542, pi7543, pi7544, pi7545, pi7546, pi7547, pi7548, pi7549, pi7550, pi7551, pi7552, pi7553, pi7554, pi7555, pi7556, pi7557, pi7558, pi7559, pi7560, pi7561, pi7562, pi7563, pi7564, pi7565, pi7566, pi7567, pi7568, pi7569, pi7570, pi7571, pi7572, pi7573, pi7574, pi7575, pi7576, pi7577, pi7578, pi7579, pi7580, pi7581, pi7582, pi7583, pi7584, pi7585, pi7586, pi7587, pi7588, pi7589, pi7590, pi7591, pi7592, pi7593, pi7594, pi7595, pi7596, pi7597, pi7598, pi7599, pi7600, pi7601, pi7602, pi7603, pi7604, pi7605, pi7606, pi7607, pi7608, pi7609, pi7610, pi7611, pi7612, pi7613, pi7614, pi7615, pi7616, pi7617, pi7618, pi7619, pi7620, pi7621, pi7622, pi7623, pi7624, pi7625, pi7626, pi7627, pi7628, pi7629, pi7630, pi7631, pi7632, pi7633, pi7634, pi7635, pi7636, pi7637, pi7638, pi7639, pi7640, pi7641, pi7642, pi7643, pi7644, pi7645, pi7646, pi7647, pi7648, pi7649, pi7650, pi7651, pi7652, pi7653, pi7654, pi7655, pi7656, pi7657, pi7658, pi7659, pi7660, pi7661, pi7662, pi7663, pi7664, pi7665, pi7666, pi7667, pi7668, pi7669, pi7670, pi7671, pi7672, pi7673, pi7674, pi7675, pi7676, pi7677, pi7678, pi7679, pi7680, pi7681, pi7682, pi7683, pi7684, pi7685, pi7686, pi7687, pi7688, pi7689, pi7690, pi7691, pi7692, pi7693, pi7694, pi7695, pi7696, pi7697, pi7698, pi7699, pi7700, pi7701, pi7702, pi7703, pi7704, pi7705, pi7706, pi7707, pi7708, pi7709, pi7710, pi7711, pi7712, pi7713, pi7714, pi7715, pi7716, pi7717, pi7718, pi7719, pi7720, pi7721, pi7722, pi7723, pi7724, pi7725, pi7726, pi7727, pi7728, pi7729, pi7730, pi7731, pi7732, pi7733, pi7734, pi7735, pi7736, pi7737, pi7738, pi7739, pi7740, pi7741, pi7742, pi7743, pi7744, pi7745, pi7746, pi7747, pi7748, pi7749, pi7750, pi7751, pi7752, pi7753, pi7754, pi7755, pi7756, pi7757, pi7758, pi7759, pi7760, pi7761, pi7762, pi7763, pi7764, pi7765, pi7766, pi7767, pi7768, pi7769, pi7770, pi7771, pi7772, pi7773, pi7774, pi7775, pi7776, pi7777, pi7778, pi7779, pi7780, pi7781, pi7782, pi7783, pi7784, pi7785, pi7786, pi7787, pi7788, pi7789, pi7790, pi7791, pi7792, pi7793, pi7794, pi7795, pi7796, pi7797, pi7798, pi7799, pi7800, pi7801, pi7802, pi7803, pi7804, pi7805, pi7806, pi7807, pi7808, pi7809, pi7810, pi7811, pi7812, pi7813, pi7814, pi7815, pi7816, pi7817, pi7818, pi7819, pi7820, pi7821, pi7822, pi7823, pi7824, pi7825, pi7826, pi7827, pi7828, pi7829, pi7830, pi7831, pi7832, pi7833, pi7834, pi7835, pi7836, pi7837, pi7838, pi7839, pi7840, pi7841, pi7842, pi7843, pi7844, pi7845, pi7846, pi7847, pi7848, pi7849, pi7850, pi7851, pi7852, pi7853, pi7854, pi7855, pi7856, pi7857, pi7858, pi7859, pi7860, pi7861, pi7862, pi7863, pi7864, pi7865, pi7866, pi7867, pi7868, pi7869, pi7870, pi7871, pi7872, pi7873, pi7874, pi7875, pi7876, pi7877, pi7878, pi7879, pi7880, pi7881, pi7882, pi7883, pi7884, pi7885, pi7886, pi7887, pi7888, pi7889, pi7890, pi7891, pi7892, pi7893, pi7894, pi7895, pi7896, pi7897, pi7898, pi7899, pi7900, pi7901, pi7902, pi7903, pi7904, pi7905, pi7906, pi7907, pi7908, pi7909, pi7910, pi7911, pi7912, pi7913, pi7914, pi7915, pi7916, pi7917, pi7918, pi7919, pi7920, pi7921, pi7922, pi7923, pi7924, pi7925, pi7926, pi7927, pi7928, pi7929, pi7930, pi7931, pi7932, pi7933, pi7934, pi7935, pi7936, pi7937, pi7938, pi7939, pi7940, pi7941, pi7942, pi7943, pi7944, pi7945, pi7946, pi7947, pi7948, pi7949, pi7950, pi7951, pi7952, pi7953, pi7954, pi7955, pi7956, pi7957, pi7958, pi7959, pi7960, pi7961, pi7962, pi7963, pi7964, pi7965, pi7966, pi7967, pi7968, pi7969, pi7970, pi7971, pi7972, pi7973, pi7974, pi7975, pi7976, pi7977, pi7978, pi7979, pi7980, pi7981, pi7982, pi7983, pi7984, pi7985, pi7986, pi7987, pi7988, pi7989, pi7990, pi7991, pi7992, pi7993, pi7994, pi7995, pi7996, pi7997, pi7998, pi7999, pi8000, pi8001, pi8002, pi8003, pi8004, pi8005, pi8006, pi8007, pi8008, pi8009, pi8010, pi8011, pi8012, pi8013, pi8014, pi8015, pi8016, pi8017, pi8018, pi8019, pi8020, pi8021, pi8022, pi8023, pi8024, pi8025, pi8026, pi8027, pi8028, pi8029, pi8030, pi8031, pi8032, pi8033, pi8034, pi8035, pi8036, pi8037, pi8038, pi8039, pi8040, pi8041, pi8042, pi8043, pi8044, pi8045, pi8046, pi8047, pi8048, pi8049, pi8050, pi8051, pi8052, pi8053, pi8054, pi8055, pi8056, pi8057, pi8058, pi8059, pi8060, pi8061, pi8062, pi8063, pi8064, pi8065, pi8066, pi8067, pi8068, pi8069, pi8070, pi8071, pi8072, pi8073, pi8074, pi8075, pi8076, pi8077, pi8078, pi8079, pi8080, pi8081, pi8082, pi8083, pi8084, pi8085, pi8086, pi8087, pi8088, pi8089, pi8090, pi8091, pi8092, pi8093, pi8094, pi8095, pi8096, pi8097, pi8098, pi8099, pi8100, pi8101, pi8102, pi8103, pi8104, pi8105, pi8106, pi8107, pi8108, pi8109, pi8110, pi8111, pi8112, pi8113, pi8114, pi8115, pi8116, pi8117, pi8118, pi8119, pi8120, pi8121, pi8122, pi8123, pi8124, pi8125, pi8126, pi8127, pi8128, pi8129, pi8130, pi8131, pi8132, pi8133, pi8134, pi8135, pi8136, pi8137, pi8138, pi8139, pi8140, pi8141, pi8142, pi8143, pi8144, pi8145, pi8146, pi8147, pi8148, pi8149, pi8150, pi8151, pi8152, pi8153, pi8154, pi8155, pi8156, pi8157, pi8158, pi8159, pi8160, pi8161, pi8162, pi8163, pi8164, pi8165, pi8166, pi8167, pi8168, pi8169, pi8170, pi8171, pi8172, pi8173, pi8174, pi8175, pi8176, pi8177, pi8178, pi8179, pi8180, pi8181, pi8182, pi8183, pi8184, pi8185, pi8186, pi8187, pi8188, pi8189, pi8190, pi8191, pi8192, pi8193, pi8194, pi8195, pi8196, pi8197, pi8198, pi8199, pi8200, pi8201, pi8202, pi8203, pi8204, pi8205, pi8206, pi8207, pi8208, pi8209, pi8210, pi8211, pi8212, pi8213, pi8214, pi8215, pi8216, pi8217, pi8218, pi8219, pi8220, pi8221, pi8222, pi8223, pi8224, pi8225, pi8226, pi8227, pi8228, pi8229, pi8230, pi8231, pi8232, pi8233, pi8234, pi8235, pi8236, pi8237, pi8238, pi8239, pi8240, pi8241, pi8242, pi8243, pi8244, pi8245, pi8246, pi8247, pi8248, pi8249, pi8250, pi8251, pi8252, pi8253, pi8254, pi8255, pi8256, pi8257, pi8258, pi8259, pi8260, pi8261, pi8262, pi8263, pi8264, pi8265, pi8266, pi8267, pi8268, pi8269, pi8270, pi8271, pi8272, pi8273, pi8274, pi8275, pi8276, pi8277, pi8278, pi8279, pi8280, pi8281, pi8282, pi8283, pi8284, pi8285, pi8286, pi8287, pi8288, pi8289, pi8290, pi8291, pi8292, pi8293, pi8294, pi8295, pi8296, pi8297, pi8298, pi8299, pi8300, pi8301, pi8302, pi8303, pi8304, pi8305, pi8306, pi8307, pi8308, pi8309, pi8310, pi8311, pi8312, pi8313, pi8314, pi8315, pi8316, pi8317, pi8318, pi8319, pi8320, pi8321, pi8322, pi8323, pi8324, pi8325, pi8326, pi8327, pi8328, pi8329, pi8330, pi8331, pi8332, pi8333, pi8334, pi8335, pi8336, pi8337, pi8338, pi8339, pi8340, pi8341, pi8342, pi8343, pi8344, pi8345, pi8346, pi8347, pi8348, pi8349, pi8350, pi8351, pi8352, pi8353, pi8354, pi8355, pi8356, pi8357, pi8358, pi8359, pi8360, pi8361, pi8362, pi8363, pi8364, pi8365, pi8366, pi8367, pi8368, pi8369, pi8370, pi8371, pi8372, pi8373, pi8374, pi8375, pi8376, pi8377, pi8378, pi8379, pi8380, pi8381, pi8382, pi8383, pi8384, pi8385, pi8386, pi8387, pi8388, pi8389, pi8390, pi8391, pi8392, pi8393, pi8394, pi8395, pi8396, pi8397, pi8398, pi8399, pi8400, pi8401, pi8402, pi8403, pi8404, pi8405, pi8406, pi8407, pi8408, pi8409, pi8410, pi8411, pi8412, pi8413, pi8414, pi8415, pi8416, pi8417, pi8418, pi8419, pi8420, pi8421, pi8422, pi8423, pi8424, pi8425, pi8426, pi8427, pi8428, pi8429, pi8430, pi8431, pi8432, pi8433, pi8434, pi8435, pi8436, pi8437, pi8438, pi8439, pi8440, pi8441, pi8442, pi8443, pi8444, pi8445, pi8446, pi8447, pi8448, pi8449, pi8450, pi8451, pi8452, pi8453, pi8454, pi8455, pi8456, pi8457, pi8458, pi8459, pi8460, pi8461, pi8462, pi8463, pi8464, pi8465, pi8466, pi8467, pi8468, pi8469, pi8470, pi8471, pi8472, pi8473, pi8474, pi8475, pi8476, pi8477, pi8478, pi8479, pi8480, pi8481, pi8482, pi8483, pi8484, pi8485, pi8486, pi8487, pi8488, pi8489, pi8490, pi8491, pi8492, pi8493, pi8494, pi8495, pi8496, pi8497, pi8498, pi8499, pi8500, pi8501, pi8502, pi8503, pi8504, pi8505, pi8506, pi8507, pi8508, pi8509, pi8510, pi8511, pi8512, pi8513, pi8514, pi8515, pi8516, pi8517, pi8518, pi8519, pi8520, pi8521, pi8522, pi8523, pi8524, pi8525, pi8526, pi8527, pi8528, pi8529, pi8530, pi8531, pi8532, pi8533, pi8534, pi8535, pi8536, pi8537, pi8538, pi8539, pi8540, pi8541, pi8542, pi8543, pi8544, pi8545, pi8546, pi8547, pi8548, pi8549, pi8550, pi8551, pi8552, pi8553, pi8554, pi8555, pi8556, pi8557, pi8558, pi8559, pi8560, pi8561, pi8562, pi8563, pi8564, pi8565, pi8566, pi8567, pi8568, pi8569, pi8570, pi8571, pi8572, pi8573, pi8574, pi8575, pi8576, pi8577, pi8578, pi8579, pi8580, pi8581, pi8582, pi8583, pi8584, pi8585, pi8586, pi8587, pi8588, pi8589, pi8590, pi8591, pi8592, pi8593, pi8594, pi8595, pi8596, pi8597, pi8598, pi8599, pi8600, pi8601, pi8602, pi8603, pi8604, pi8605, pi8606, pi8607, pi8608, pi8609, pi8610, pi8611, pi8612, pi8613, pi8614, pi8615, pi8616, pi8617, pi8618, pi8619, pi8620, pi8621, pi8622, pi8623, pi8624, pi8625, pi8626, pi8627, pi8628, pi8629, pi8630, pi8631, pi8632, pi8633, pi8634, pi8635, pi8636, pi8637, pi8638, pi8639, pi8640, pi8641, pi8642, pi8643, pi8644, pi8645, pi8646, pi8647, pi8648, pi8649, pi8650, pi8651, pi8652, pi8653, pi8654, pi8655, pi8656, pi8657, pi8658, pi8659, pi8660, pi8661, pi8662, pi8663, pi8664, pi8665, pi8666, pi8667, pi8668, pi8669, pi8670, pi8671, pi8672, pi8673, pi8674, pi8675, pi8676, pi8677, pi8678, pi8679, pi8680, pi8681, pi8682, pi8683, pi8684, pi8685, pi8686, pi8687, pi8688, pi8689, pi8690, pi8691, pi8692, pi8693, pi8694, pi8695, pi8696, pi8697, pi8698, pi8699, pi8700, pi8701, pi8702, pi8703, pi8704, pi8705, pi8706, pi8707, pi8708, pi8709, pi8710, pi8711, pi8712, pi8713, pi8714, pi8715, pi8716, pi8717, pi8718, pi8719, pi8720, pi8721, pi8722, pi8723, pi8724, pi8725, pi8726, pi8727, pi8728, pi8729, pi8730, pi8731, pi8732, pi8733, pi8734, pi8735, pi8736, pi8737, pi8738, pi8739, pi8740, pi8741, pi8742, pi8743, pi8744, pi8745, pi8746, pi8747, pi8748, pi8749, pi8750, pi8751, pi8752, pi8753, pi8754, pi8755, pi8756, pi8757, pi8758, pi8759, pi8760, pi8761, pi8762, pi8763, pi8764, pi8765, pi8766, pi8767, pi8768, pi8769, pi8770, pi8771, pi8772, pi8773, pi8774, pi8775, pi8776, pi8777, pi8778, pi8779, pi8780, pi8781, pi8782, pi8783, pi8784, pi8785, pi8786, pi8787, pi8788, pi8789, pi8790, pi8791, pi8792, pi8793, pi8794, pi8795, pi8796, pi8797, pi8798, pi8799, pi8800, pi8801, pi8802, pi8803, pi8804, pi8805, pi8806, pi8807, pi8808, pi8809, pi8810, pi8811, pi8812, pi8813, pi8814, pi8815, pi8816, pi8817, pi8818, pi8819, pi8820, pi8821, pi8822, pi8823, pi8824, pi8825, pi8826, pi8827, pi8828, pi8829, pi8830, pi8831, pi8832, pi8833, pi8834, pi8835, pi8836, pi8837, pi8838, pi8839, pi8840, pi8841, pi8842, pi8843, pi8844, pi8845, pi8846, pi8847, pi8848, pi8849, pi8850, pi8851, pi8852, pi8853, pi8854, pi8855, pi8856, pi8857, pi8858, pi8859, pi8860, pi8861, pi8862, pi8863, pi8864, pi8865, pi8866, pi8867, pi8868, pi8869, pi8870, pi8871, pi8872, pi8873, pi8874, pi8875, pi8876, pi8877, pi8878, pi8879, pi8880, pi8881, pi8882, pi8883, pi8884, pi8885, pi8886, pi8887, pi8888, pi8889, pi8890, pi8891, pi8892, pi8893, pi8894, pi8895, pi8896, pi8897, pi8898, pi8899, pi8900, pi8901, pi8902, pi8903, pi8904, pi8905, pi8906, pi8907, pi8908, pi8909, pi8910, pi8911, pi8912, pi8913, pi8914, pi8915, pi8916, pi8917, pi8918, pi8919, pi8920, pi8921, pi8922, pi8923, pi8924, pi8925, pi8926, pi8927, pi8928, pi8929, pi8930, pi8931, pi8932, pi8933, pi8934, pi8935, pi8936, pi8937, pi8938, pi8939, pi8940, pi8941, pi8942, pi8943, pi8944, pi8945, pi8946, pi8947, pi8948, pi8949, pi8950, pi8951, pi8952, pi8953, pi8954, pi8955, pi8956, pi8957, pi8958, pi8959, pi8960, pi8961, pi8962, pi8963, pi8964, pi8965, pi8966, pi8967, pi8968, pi8969, pi8970, pi8971, pi8972, pi8973, pi8974, pi8975, pi8976, pi8977, pi8978, pi8979, pi8980, pi8981, pi8982, pi8983, pi8984, pi8985, pi8986, pi8987, pi8988, pi8989, pi8990, pi8991, pi8992, pi8993, pi8994, pi8995, pi8996, pi8997, pi8998, pi8999, pi9000, pi9001, pi9002, pi9003, pi9004, pi9005, pi9006, pi9007, pi9008, pi9009, pi9010, pi9011, pi9012, pi9013, pi9014, pi9015, pi9016, pi9017, pi9018, pi9019, pi9020, pi9021, pi9022, pi9023, pi9024, pi9025, pi9026, pi9027, pi9028, pi9029, pi9030, pi9031, pi9032, pi9033, pi9034, pi9035, pi9036, pi9037, pi9038, pi9039, pi9040, pi9041, 
            po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535, po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544, po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553, po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562, po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571, po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580, po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589, po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598, po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607, po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616, po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625, po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634, po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643, po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652, po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661, po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670, po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679, po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688, po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697, po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706, po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715, po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724, po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733, po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742, po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751, po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760, po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769, po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778, po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787, po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796, po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805, po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814, po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823, po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832, po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841, po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850, po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859, po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868, po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877, po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886, po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895, po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904, po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913, po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922, po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931, po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940, po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949, po3950, po3951, po3952, po3953, po3954, po3955, po3956, po3957, po3958, po3959, po3960, po3961, po3962, po3963, po3964, po3965, po3966, po3967, po3968, po3969, po3970, po3971, po3972, po3973, po3974, po3975, po3976, po3977, po3978, po3979, po3980, po3981, po3982, po3983, po3984, po3985, po3986, po3987, po3988, po3989, po3990, po3991, po3992, po3993, po3994, po3995, po3996, po3997, po3998, po3999, po4000, po4001, po4002, po4003, po4004, po4005, po4006, po4007, po4008, po4009, po4010, po4011, po4012, po4013, po4014, po4015, po4016, po4017, po4018, po4019, po4020, po4021, po4022, po4023, po4024, po4025, po4026, po4027, po4028, po4029, po4030, po4031, po4032, po4033, po4034, po4035, po4036, po4037, po4038, po4039, po4040, po4041, po4042, po4043, po4044, po4045, po4046, po4047, po4048, po4049, po4050, po4051, po4052, po4053, po4054, po4055, po4056, po4057, po4058, po4059, po4060, po4061, po4062, po4063, po4064, po4065, po4066, po4067, po4068, po4069, po4070, po4071, po4072, po4073, po4074, po4075, po4076, po4077, po4078, po4079, po4080, po4081, po4082, po4083, po4084, po4085, po4086, po4087, po4088, po4089, po4090, po4091, po4092, po4093, po4094, po4095, po4096, po4097, po4098, po4099, po4100, po4101, po4102, po4103, po4104, po4105, po4106, po4107, po4108, po4109, po4110, po4111, po4112, po4113, po4114, po4115, po4116, po4117, po4118, po4119, po4120, po4121, po4122, po4123, po4124, po4125, po4126, po4127, po4128, po4129, po4130, po4131, po4132, po4133, po4134, po4135, po4136, po4137, po4138, po4139, po4140, po4141, po4142, po4143, po4144, po4145, po4146, po4147, po4148, po4149, po4150, po4151, po4152, po4153, po4154, po4155, po4156, po4157, po4158, po4159, po4160, po4161, po4162, po4163, po4164, po4165, po4166, po4167, po4168, po4169, po4170, po4171, po4172, po4173, po4174, po4175, po4176, po4177, po4178, po4179, po4180, po4181, po4182, po4183, po4184, po4185, po4186, po4187, po4188, po4189, po4190, po4191, po4192, po4193, po4194, po4195, po4196, po4197, po4198, po4199, po4200, po4201, po4202, po4203, po4204, po4205, po4206, po4207, po4208, po4209, po4210, po4211, po4212, po4213, po4214, po4215, po4216, po4217, po4218, po4219, po4220, po4221, po4222, po4223, po4224, po4225, po4226, po4227, po4228, po4229, po4230, po4231, po4232, po4233, po4234, po4235, po4236, po4237, po4238, po4239, po4240, po4241, po4242, po4243, po4244, po4245, po4246, po4247, po4248, po4249, po4250, po4251, po4252, po4253, po4254, po4255, po4256, po4257, po4258, po4259, po4260, po4261, po4262, po4263, po4264, po4265, po4266, po4267, po4268, po4269, po4270, po4271, po4272, po4273, po4274, po4275, po4276, po4277, po4278, po4279, po4280, po4281, po4282, po4283, po4284, po4285, po4286, po4287, po4288, po4289, po4290, po4291, po4292, po4293, po4294, po4295, po4296, po4297, po4298, po4299, po4300, po4301, po4302, po4303, po4304, po4305, po4306, po4307, po4308, po4309, po4310, po4311, po4312, po4313, po4314, po4315, po4316, po4317, po4318, po4319, po4320, po4321, po4322, po4323, po4324, po4325, po4326, po4327, po4328, po4329, po4330, po4331, po4332, po4333, po4334, po4335, po4336, po4337, po4338, po4339, po4340, po4341, po4342, po4343, po4344, po4345, po4346, po4347, po4348, po4349, po4350, po4351, po4352, po4353, po4354, po4355, po4356, po4357, po4358, po4359, po4360, po4361, po4362, po4363, po4364, po4365, po4366, po4367, po4368, po4369, po4370, po4371, po4372, po4373, po4374, po4375, po4376, po4377, po4378, po4379, po4380, po4381, po4382, po4383, po4384, po4385, po4386, po4387, po4388, po4389, po4390, po4391, po4392, po4393, po4394, po4395, po4396, po4397, po4398, po4399, po4400, po4401, po4402, po4403, po4404, po4405, po4406, po4407, po4408, po4409, po4410, po4411, po4412, po4413, po4414, po4415, po4416, po4417, po4418, po4419, po4420, po4421, po4422, po4423, po4424, po4425, po4426, po4427, po4428, po4429, po4430, po4431, po4432, po4433, po4434, po4435, po4436, po4437, po4438, po4439, po4440, po4441, po4442, po4443, po4444, po4445, po4446, po4447, po4448, po4449, po4450, po4451, po4452, po4453, po4454, po4455, po4456, po4457, po4458, po4459, po4460, po4461, po4462, po4463, po4464, po4465, po4466, po4467, po4468, po4469, po4470, po4471, po4472, po4473, po4474, po4475, po4476, po4477, po4478, po4479, po4480, po4481, po4482, po4483, po4484, po4485, po4486, po4487, po4488, po4489, po4490, po4491, po4492, po4493, po4494, po4495, po4496, po4497, po4498, po4499, po4500, po4501, po4502, po4503, po4504, po4505, po4506, po4507, po4508, po4509, po4510, po4511, po4512, po4513, po4514, po4515, po4516, po4517, po4518, po4519, po4520, po4521, po4522, po4523, po4524, po4525, po4526, po4527, po4528, po4529, po4530, po4531, po4532, po4533, po4534, po4535, po4536, po4537, po4538, po4539, po4540, po4541, po4542, po4543, po4544, po4545, po4546, po4547, po4548, po4549, po4550, po4551, po4552, po4553, po4554, po4555, po4556, po4557, po4558, po4559, po4560, po4561, po4562, po4563, po4564, po4565, po4566, po4567, po4568, po4569, po4570, po4571, po4572, po4573, po4574, po4575, po4576, po4577, po4578, po4579, po4580, po4581, po4582, po4583, po4584, po4585, po4586, po4587, po4588, po4589, po4590, po4591, po4592, po4593, po4594, po4595, po4596, po4597, po4598, po4599, po4600, po4601, po4602, po4603, po4604, po4605, po4606, po4607, po4608, po4609, po4610, po4611, po4612, po4613, po4614, po4615, po4616, po4617, po4618, po4619, po4620, po4621, po4622, po4623, po4624, po4625, po4626, po4627, po4628, po4629, po4630, po4631, po4632, po4633, po4634, po4635, po4636, po4637, po4638, po4639, po4640, po4641, po4642, po4643, po4644, po4645, po4646, po4647, po4648, po4649, po4650, po4651, po4652, po4653, po4654, po4655, po4656, po4657, po4658, po4659, po4660, po4661, po4662, po4663, po4664, po4665, po4666, po4667, po4668, po4669, po4670, po4671, po4672, po4673, po4674, po4675, po4676, po4677, po4678, po4679, po4680, po4681, po4682, po4683, po4684, po4685, po4686, po4687, po4688, po4689, po4690, po4691, po4692, po4693, po4694, po4695, po4696, po4697, po4698, po4699, po4700, po4701, po4702, po4703, po4704, po4705, po4706, po4707, po4708, po4709, po4710, po4711, po4712, po4713, po4714, po4715, po4716, po4717, po4718, po4719, po4720, po4721, po4722, po4723, po4724, po4725, po4726, po4727, po4728, po4729, po4730, po4731, po4732, po4733, po4734, po4735, po4736, po4737, po4738, po4739, po4740, po4741, po4742, po4743, po4744, po4745, po4746, po4747, po4748, po4749, po4750, po4751, po4752, po4753, po4754, po4755, po4756, po4757, po4758, po4759, po4760, po4761, po4762, po4763, po4764, po4765, po4766, po4767, po4768, po4769, po4770, po4771, po4772, po4773, po4774, po4775, po4776, po4777, po4778, po4779, po4780, po4781, po4782, po4783, po4784, po4785, po4786, po4787, po4788, po4789, po4790, po4791, po4792, po4793, po4794, po4795, po4796, po4797, po4798, po4799, po4800, po4801, po4802, po4803, po4804, po4805, po4806, po4807, po4808, po4809, po4810, po4811, po4812, po4813, po4814, po4815, po4816, po4817, po4818, po4819, po4820, po4821, po4822, po4823, po4824, po4825, po4826, po4827, po4828, po4829, po4830, po4831, po4832, po4833, po4834, po4835, po4836, po4837, po4838, po4839, po4840, po4841, po4842, po4843, po4844, po4845, po4846, po4847, po4848, po4849, po4850, po4851, po4852, po4853, po4854, po4855, po4856, po4857, po4858, po4859, po4860, po4861, po4862, po4863, po4864, po4865, po4866, po4867, po4868, po4869, po4870, po4871, po4872, po4873, po4874, po4875, po4876, po4877, po4878, po4879, po4880, po4881, po4882, po4883, po4884, po4885, po4886, po4887, po4888, po4889, po4890, po4891, po4892, po4893, po4894, po4895, po4896, po4897, po4898, po4899, po4900, po4901, po4902, po4903, po4904, po4905, po4906, po4907, po4908, po4909, po4910, po4911, po4912, po4913, po4914, po4915, po4916, po4917, po4918, po4919, po4920, po4921, po4922, po4923, po4924, po4925, po4926, po4927, po4928, po4929, po4930, po4931, po4932, po4933, po4934, po4935, po4936, po4937, po4938, po4939, po4940, po4941, po4942, po4943, po4944, po4945, po4946, po4947, po4948, po4949, po4950, po4951, po4952, po4953, po4954, po4955, po4956, po4957, po4958, po4959, po4960, po4961, po4962, po4963, po4964, po4965, po4966, po4967, po4968, po4969, po4970, po4971, po4972, po4973, po4974, po4975, po4976, po4977, po4978, po4979, po4980, po4981, po4982, po4983, po4984, po4985, po4986, po4987, po4988, po4989, po4990, po4991, po4992, po4993, po4994, po4995, po4996, po4997, po4998, po4999, po5000, po5001, po5002, po5003, po5004, po5005, po5006, po5007, po5008, po5009, po5010, po5011, po5012, po5013, po5014, po5015, po5016, po5017, po5018, po5019, po5020, po5021, po5022, po5023, po5024, po5025, po5026, po5027, po5028, po5029, po5030, po5031, po5032, po5033, po5034, po5035, po5036, po5037, po5038, po5039, po5040, po5041, po5042, po5043, po5044, po5045, po5046, po5047, po5048, po5049, po5050, po5051, po5052, po5053, po5054, po5055, po5056, po5057, po5058, po5059, po5060, po5061, po5062, po5063, po5064, po5065, po5066, po5067, po5068, po5069, po5070, po5071, po5072, po5073, po5074, po5075, po5076, po5077, po5078, po5079, po5080, po5081, po5082, po5083, po5084, po5085, po5086, po5087, po5088, po5089, po5090, po5091, po5092, po5093, po5094, po5095, po5096, po5097, po5098, po5099, po5100, po5101, po5102, po5103, po5104, po5105, po5106, po5107, po5108, po5109, po5110, po5111, po5112, po5113, po5114, po5115, po5116, po5117, po5118, po5119, po5120, po5121, po5122, po5123, po5124, po5125, po5126, po5127, po5128, po5129, po5130, po5131, po5132, po5133, po5134, po5135, po5136, po5137, po5138, po5139, po5140, po5141, po5142, po5143, po5144, po5145, po5146, po5147, po5148, po5149, po5150, po5151, po5152, po5153, po5154, po5155, po5156, po5157, po5158, po5159, po5160, po5161, po5162, po5163, po5164, po5165, po5166, po5167, po5168, po5169, po5170, po5171, po5172, po5173, po5174, po5175, po5176, po5177, po5178, po5179, po5180, po5181, po5182, po5183, po5184, po5185, po5186, po5187, po5188, po5189, po5190, po5191, po5192, po5193, po5194, po5195, po5196, po5197, po5198, po5199, po5200, po5201, po5202, po5203, po5204, po5205, po5206, po5207, po5208, po5209, po5210, po5211, po5212, po5213, po5214, po5215, po5216, po5217, po5218, po5219, po5220, po5221, po5222, po5223, po5224, po5225, po5226, po5227, po5228, po5229, po5230, po5231, po5232, po5233, po5234, po5235, po5236, po5237, po5238, po5239, po5240, po5241, po5242, po5243, po5244, po5245, po5246, po5247, po5248, po5249, po5250, po5251, po5252, po5253, po5254, po5255, po5256, po5257, po5258, po5259, po5260, po5261, po5262, po5263, po5264, po5265, po5266, po5267, po5268, po5269, po5270, po5271, po5272, po5273, po5274, po5275, po5276, po5277, po5278, po5279, po5280, po5281, po5282, po5283, po5284, po5285, po5286, po5287, po5288, po5289, po5290, po5291, po5292, po5293, po5294, po5295, po5296, po5297, po5298, po5299, po5300, po5301, po5302, po5303, po5304, po5305, po5306, po5307, po5308, po5309, po5310, po5311, po5312, po5313, po5314, po5315, po5316, po5317, po5318, po5319, po5320, po5321, po5322, po5323, po5324, po5325, po5326, po5327, po5328, po5329, po5330, po5331, po5332, po5333, po5334, po5335, po5336, po5337, po5338, po5339, po5340, po5341, po5342, po5343, po5344, po5345, po5346, po5347, po5348, po5349, po5350, po5351, po5352, po5353, po5354, po5355, po5356, po5357, po5358, po5359, po5360, po5361, po5362, po5363, po5364, po5365, po5366, po5367, po5368, po5369, po5370, po5371, po5372, po5373, po5374, po5375, po5376, po5377, po5378, po5379, po5380, po5381, po5382, po5383, po5384, po5385, po5386, po5387, po5388, po5389, po5390, po5391, po5392, po5393, po5394, po5395, po5396, po5397, po5398, po5399, po5400, po5401, po5402, po5403, po5404, po5405, po5406, po5407, po5408, po5409, po5410, po5411, po5412, po5413, po5414, po5415, po5416, po5417, po5418, po5419, po5420, po5421, po5422, po5423, po5424, po5425, po5426, po5427, po5428, po5429, po5430, po5431, po5432, po5433, po5434, po5435, po5436, po5437, po5438, po5439, po5440, po5441, po5442, po5443, po5444, po5445, po5446, po5447, po5448, po5449, po5450, po5451, po5452, po5453, po5454, po5455, po5456, po5457, po5458, po5459, po5460, po5461, po5462, po5463, po5464, po5465, po5466, po5467, po5468, po5469, po5470, po5471, po5472, po5473, po5474, po5475, po5476, po5477, po5478, po5479, po5480, po5481, po5482, po5483, po5484, po5485, po5486, po5487, po5488, po5489, po5490, po5491, po5492, po5493, po5494, po5495, po5496, po5497, po5498, po5499, po5500, po5501, po5502, po5503, po5504, po5505, po5506, po5507, po5508, po5509, po5510, po5511, po5512, po5513, po5514, po5515, po5516, po5517, po5518, po5519, po5520, po5521, po5522, po5523, po5524, po5525, po5526, po5527, po5528, po5529, po5530, po5531, po5532, po5533, po5534, po5535, po5536, po5537, po5538, po5539, po5540, po5541, po5542, po5543, po5544, po5545, po5546, po5547, po5548, po5549, po5550, po5551, po5552, po5553, po5554, po5555, po5556, po5557, po5558, po5559, po5560, po5561, po5562, po5563, po5564, po5565, po5566, po5567, po5568, po5569, po5570, po5571, po5572, po5573, po5574, po5575, po5576, po5577, po5578, po5579, po5580, po5581, po5582, po5583, po5584, po5585, po5586, po5587, po5588, po5589, po5590, po5591, po5592, po5593, po5594, po5595, po5596, po5597, po5598, po5599, po5600, po5601, po5602, po5603, po5604, po5605, po5606, po5607, po5608, po5609, po5610, po5611, po5612, po5613, po5614, po5615, po5616, po5617, po5618, po5619, po5620, po5621, po5622, po5623, po5624, po5625, po5626, po5627, po5628, po5629, po5630, po5631, po5632, po5633, po5634, po5635, po5636, po5637, po5638, po5639, po5640, po5641, po5642, po5643, po5644, po5645, po5646, po5647, po5648, po5649, po5650, po5651, po5652, po5653, po5654, po5655, po5656, po5657, po5658, po5659, po5660, po5661, po5662, po5663, po5664, po5665, po5666, po5667, po5668, po5669, po5670, po5671, po5672, po5673, po5674, po5675, po5676, po5677, po5678, po5679, po5680, po5681, po5682, po5683, po5684, po5685, po5686, po5687, po5688, po5689, po5690, po5691, po5692, po5693, po5694, po5695, po5696, po5697, po5698, po5699, po5700, po5701, po5702, po5703, po5704, po5705, po5706, po5707, po5708, po5709, po5710, po5711, po5712, po5713, po5714, po5715, po5716, po5717, po5718, po5719, po5720, po5721, po5722, po5723, po5724, po5725, po5726, po5727, po5728, po5729, po5730, po5731, po5732, po5733, po5734, po5735, po5736, po5737, po5738, po5739, po5740, po5741, po5742, po5743, po5744, po5745, po5746, po5747, po5748, po5749, po5750, po5751, po5752, po5753, po5754, po5755, po5756, po5757, po5758, po5759, po5760, po5761, po5762, po5763, po5764, po5765, po5766, po5767, po5768, po5769, po5770, po5771, po5772, po5773, po5774, po5775, po5776, po5777, po5778, po5779, po5780, po5781, po5782, po5783, po5784, po5785, po5786, po5787, po5788, po5789, po5790, po5791, po5792, po5793, po5794, po5795, po5796, po5797, po5798, po5799, po5800, po5801, po5802, po5803, po5804, po5805, po5806, po5807, po5808, po5809, po5810, po5811, po5812, po5813, po5814, po5815, po5816, po5817, po5818, po5819, po5820, po5821, po5822, po5823, po5824, po5825, po5826, po5827, po5828, po5829, po5830, po5831, po5832, po5833, po5834, po5835, po5836, po5837, po5838, po5839, po5840, po5841, po5842, po5843, po5844, po5845, po5846, po5847, po5848, po5849, po5850, po5851, po5852, po5853, po5854, po5855, po5856, po5857, po5858, po5859, po5860, po5861, po5862, po5863, po5864, po5865, po5866, po5867, po5868, po5869, po5870, po5871, po5872, po5873, po5874, po5875, po5876, po5877, po5878, po5879, po5880, po5881, po5882, po5883, po5884, po5885, po5886, po5887, po5888, po5889, po5890, po5891, po5892, po5893, po5894, po5895, po5896, po5897, po5898, po5899, po5900, po5901, po5902, po5903, po5904, po5905, po5906, po5907, po5908, po5909, po5910, po5911, po5912, po5913, po5914, po5915, po5916, po5917, po5918, po5919, po5920, po5921, po5922, po5923, po5924, po5925, po5926, po5927, po5928, po5929, po5930, po5931, po5932, po5933, po5934, po5935, po5936, po5937, po5938, po5939, po5940, po5941, po5942, po5943, po5944, po5945, po5946, po5947, po5948, po5949, po5950, po5951, po5952, po5953, po5954, po5955, po5956, po5957, po5958, po5959, po5960, po5961, po5962, po5963, po5964, po5965, po5966, po5967, po5968, po5969, po5970, po5971, po5972, po5973, po5974, po5975, po5976, po5977, po5978, po5979, po5980, po5981, po5982, po5983, po5984, po5985, po5986, po5987, po5988, po5989, po5990, po5991, po5992, po5993, po5994, po5995, po5996, po5997, po5998, po5999, po6000, po6001, po6002, po6003, po6004, po6005, po6006, po6007, po6008, po6009, po6010, po6011, po6012, po6013, po6014, po6015, po6016, po6017, po6018, po6019, po6020, po6021, po6022, po6023, po6024, po6025, po6026, po6027, po6028, po6029, po6030, po6031, po6032, po6033, po6034, po6035, po6036, po6037, po6038, po6039, po6040, po6041, po6042, po6043, po6044, po6045, po6046, po6047, po6048, po6049, po6050, po6051, po6052, po6053, po6054, po6055, po6056, po6057, po6058, po6059, po6060, po6061, po6062, po6063, po6064, po6065, po6066, po6067, po6068, po6069, po6070, po6071, po6072, po6073, po6074, po6075, po6076, po6077, po6078, po6079, po6080, po6081, po6082, po6083, po6084, po6085, po6086, po6087, po6088, po6089, po6090, po6091, po6092, po6093, po6094, po6095, po6096, po6097, po6098, po6099, po6100, po6101, po6102, po6103, po6104, po6105, po6106, po6107, po6108, po6109, po6110, po6111, po6112, po6113, po6114, po6115, po6116, po6117, po6118, po6119, po6120, po6121, po6122, po6123, po6124, po6125, po6126, po6127, po6128, po6129, po6130, po6131, po6132, po6133, po6134, po6135, po6136, po6137, po6138, po6139, po6140, po6141, po6142, po6143, po6144, po6145, po6146, po6147, po6148, po6149, po6150, po6151, po6152, po6153, po6154, po6155, po6156, po6157, po6158, po6159, po6160, po6161, po6162, po6163, po6164, po6165, po6166, po6167, po6168, po6169, po6170, po6171, po6172, po6173, po6174, po6175, po6176, po6177, po6178, po6179, po6180, po6181, po6182, po6183, po6184, po6185, po6186, po6187, po6188, po6189, po6190, po6191, po6192, po6193, po6194, po6195, po6196, po6197, po6198, po6199, po6200, po6201, po6202, po6203, po6204, po6205, po6206, po6207, po6208, po6209, po6210, po6211, po6212, po6213, po6214, po6215, po6216, po6217, po6218, po6219, po6220, po6221, po6222, po6223, po6224, po6225, po6226, po6227, po6228, po6229, po6230, po6231, po6232, po6233, po6234, po6235, po6236, po6237, po6238, po6239, po6240, po6241, po6242, po6243, po6244, po6245, po6246, po6247, po6248, po6249, po6250, po6251, po6252, po6253, po6254, po6255, po6256, po6257, po6258, po6259, po6260, po6261, po6262, po6263, po6264, po6265, po6266, po6267, po6268, po6269, po6270, po6271, po6272, po6273, po6274, po6275, po6276, po6277, po6278, po6279, po6280, po6281, po6282, po6283, po6284, po6285, po6286, po6287, po6288, po6289, po6290, po6291, po6292, po6293, po6294, po6295, po6296, po6297, po6298, po6299, po6300, po6301, po6302, po6303, po6304, po6305, po6306, po6307, po6308, po6309, po6310, po6311, po6312, po6313, po6314, po6315, po6316, po6317, po6318, po6319, po6320, po6321, po6322, po6323, po6324, po6325, po6326, po6327, po6328, po6329, po6330, po6331, po6332, po6333, po6334, po6335, po6336, po6337, po6338, po6339, po6340, po6341, po6342, po6343, po6344, po6345, po6346, po6347, po6348, po6349, po6350, po6351, po6352, po6353, po6354, po6355, po6356, po6357, po6358, po6359, po6360, po6361, po6362, po6363, po6364, po6365, po6366, po6367, po6368, po6369, po6370, po6371, po6372, po6373, po6374, po6375, po6376, po6377, po6378, po6379, po6380, po6381, po6382, po6383, po6384, po6385, po6386, po6387, po6388, po6389, po6390, po6391, po6392, po6393, po6394, po6395, po6396, po6397, po6398, po6399, po6400, po6401, po6402, po6403, po6404, po6405, po6406, po6407, po6408, po6409, po6410, po6411, po6412, po6413, po6414, po6415, po6416, po6417, po6418, po6419, po6420, po6421, po6422, po6423, po6424, po6425, po6426, po6427, po6428, po6429, po6430, po6431, po6432, po6433, po6434, po6435, po6436, po6437, po6438, po6439, po6440, po6441, po6442, po6443, po6444, po6445, po6446, po6447, po6448, po6449, po6450, po6451, po6452, po6453, po6454, po6455, po6456, po6457, po6458, po6459, po6460, po6461, po6462, po6463, po6464, po6465, po6466, po6467, po6468, po6469, po6470, po6471, po6472, po6473, po6474, po6475, po6476, po6477, po6478, po6479, po6480, po6481, po6482, po6483, po6484, po6485, po6486, po6487, po6488, po6489, po6490, po6491, po6492, po6493, po6494, po6495, po6496, po6497, po6498, po6499, po6500, po6501, po6502, po6503, po6504, po6505, po6506, po6507, po6508, po6509, po6510, po6511, po6512, po6513, po6514, po6515, po6516, po6517, po6518, po6519, po6520, po6521, po6522, po6523, po6524, po6525, po6526, po6527, po6528, po6529, po6530, po6531, po6532, po6533, po6534, po6535, po6536, po6537, po6538, po6539, po6540, po6541, po6542, po6543, po6544, po6545, po6546, po6547, po6548, po6549, po6550, po6551, po6552, po6553, po6554, po6555, po6556, po6557, po6558, po6559, po6560, po6561, po6562, po6563, po6564, po6565, po6566, po6567, po6568, po6569, po6570, po6571, po6572, po6573, po6574, po6575, po6576, po6577, po6578, po6579, po6580, po6581, po6582, po6583, po6584, po6585, po6586, po6587, po6588, po6589, po6590, po6591, po6592, po6593, po6594, po6595, po6596, po6597, po6598, po6599, po6600, po6601, po6602, po6603, po6604, po6605, po6606, po6607, po6608, po6609, po6610, po6611, po6612, po6613, po6614, po6615, po6616, po6617, po6618, po6619, po6620, po6621, po6622, po6623, po6624, po6625, po6626, po6627, po6628, po6629, po6630, po6631, po6632, po6633, po6634, po6635, po6636, po6637, po6638, po6639, po6640, po6641, po6642, po6643, po6644, po6645, po6646, po6647, po6648, po6649, po6650, po6651, po6652, po6653, po6654, po6655, po6656, po6657, po6658, po6659, po6660, po6661, po6662, po6663, po6664, po6665, po6666, po6667, po6668, po6669, po6670, po6671, po6672, po6673, po6674, po6675, po6676, po6677, po6678, po6679, po6680, po6681, po6682, po6683, po6684, po6685, po6686, po6687, po6688, po6689, po6690, po6691, po6692, po6693, po6694, po6695, po6696, po6697, po6698, po6699, po6700, po6701, po6702, po6703, po6704, po6705, po6706, po6707, po6708, po6709, po6710, po6711, po6712, po6713, po6714, po6715, po6716, po6717, po6718, po6719, po6720, po6721, po6722, po6723, po6724, po6725, po6726, po6727, po6728, po6729, po6730, po6731, po6732, po6733, po6734, po6735, po6736, po6737, po6738, po6739, po6740, po6741, po6742, po6743, po6744, po6745, po6746, po6747, po6748, po6749, po6750, po6751, po6752, po6753, po6754, po6755, po6756, po6757, po6758, po6759, po6760, po6761, po6762, po6763, po6764, po6765, po6766, po6767, po6768, po6769, po6770, po6771, po6772, po6773, po6774, po6775, po6776, po6777, po6778, po6779, po6780, po6781, po6782, po6783, po6784, po6785, po6786, po6787, po6788, po6789, po6790, po6791, po6792, po6793, po6794, po6795, po6796, po6797, po6798, po6799, po6800, po6801, po6802, po6803, po6804, po6805, po6806, po6807, po6808, po6809, po6810, po6811, po6812, po6813, po6814, po6815, po6816, po6817, po6818, po6819, po6820, po6821, po6822, po6823, po6824, po6825, po6826, po6827, po6828, po6829, po6830, po6831, po6832, po6833, po6834, po6835, po6836, po6837, po6838, po6839, po6840, po6841, po6842, po6843, po6844, po6845, po6846, po6847, po6848, po6849, po6850, po6851, po6852, po6853, po6854, po6855, po6856, po6857, po6858, po6859, po6860, po6861, po6862, po6863, po6864, po6865, po6866, po6867, po6868, po6869, po6870, po6871, po6872, po6873, po6874, po6875, po6876, po6877, po6878, po6879, po6880, po6881, po6882, po6883, po6884, po6885, po6886, po6887, po6888, po6889, po6890, po6891, po6892, po6893, po6894, po6895, po6896, po6897, po6898, po6899, po6900, po6901, po6902, po6903, po6904, po6905, po6906, po6907, po6908, po6909, po6910, po6911, po6912, po6913, po6914, po6915, po6916, po6917, po6918, po6919, po6920, po6921, po6922, po6923, po6924, po6925, po6926, po6927, po6928, po6929, po6930, po6931, po6932, po6933, po6934, po6935, po6936, po6937, po6938, po6939, po6940, po6941, po6942, po6943, po6944, po6945, po6946, po6947, po6948, po6949, po6950, po6951, po6952, po6953, po6954, po6955, po6956, po6957, po6958, po6959, po6960, po6961, po6962, po6963, po6964, po6965, po6966, po6967, po6968, po6969, po6970, po6971, po6972, po6973, po6974, po6975, po6976, po6977, po6978, po6979, po6980, po6981, po6982, po6983, po6984, po6985, po6986, po6987, po6988, po6989, po6990, po6991, po6992, po6993, po6994, po6995, po6996, po6997, po6998, po6999, po7000, po7001, po7002, po7003, po7004, po7005, po7006, po7007, po7008, po7009, po7010, po7011, po7012, po7013, po7014, po7015, po7016, po7017, po7018, po7019, po7020, po7021, po7022, po7023, po7024, po7025, po7026, po7027, po7028, po7029, po7030, po7031, po7032, po7033, po7034, po7035, po7036, po7037, po7038, po7039, po7040, po7041, po7042, po7043, po7044, po7045, po7046, po7047, po7048, po7049, po7050, po7051, po7052, po7053, po7054, po7055, po7056, po7057, po7058, po7059, po7060, po7061, po7062, po7063, po7064, po7065, po7066, po7067, po7068, po7069, po7070, po7071, po7072, po7073, po7074, po7075, po7076, po7077, po7078, po7079, po7080, po7081, po7082, po7083, po7084, po7085, po7086, po7087, po7088, po7089, po7090, po7091, po7092, po7093, po7094, po7095, po7096, po7097, po7098, po7099, po7100, po7101, po7102, po7103, po7104, po7105, po7106, po7107, po7108, po7109, po7110, po7111, po7112, po7113, po7114, po7115, po7116, po7117, po7118, po7119, po7120, po7121, po7122, po7123, po7124, po7125, po7126, po7127, po7128, po7129, po7130, po7131, po7132, po7133, po7134, po7135, po7136, po7137, po7138, po7139, po7140, po7141, po7142, po7143, po7144, po7145, po7146, po7147, po7148, po7149, po7150, po7151, po7152, po7153, po7154, po7155, po7156, po7157, po7158, po7159, po7160, po7161, po7162, po7163, po7164, po7165, po7166, po7167, po7168, po7169, po7170, po7171, po7172, po7173, po7174, po7175, po7176, po7177, po7178, po7179, po7180, po7181, po7182, po7183, po7184, po7185, po7186, po7187, po7188, po7189, po7190, po7191, po7192, po7193, po7194, po7195, po7196, po7197, po7198, po7199, po7200, po7201, po7202, po7203, po7204, po7205, po7206, po7207, po7208, po7209, po7210, po7211, po7212, po7213, po7214, po7215, po7216, po7217, po7218, po7219, po7220, po7221, po7222, po7223, po7224, po7225, po7226, po7227, po7228, po7229, po7230, po7231, po7232, po7233, po7234, po7235, po7236, po7237, po7238, po7239, po7240, po7241, po7242, po7243, po7244, po7245, po7246, po7247, po7248, po7249, po7250, po7251, po7252, po7253, po7254, po7255, po7256, po7257, po7258, po7259, po7260, po7261, po7262, po7263, po7264, po7265, po7266, po7267, po7268, po7269, po7270, po7271, po7272, po7273, po7274, po7275, po7276, po7277, po7278, po7279, po7280, po7281, po7282, po7283, po7284, po7285, po7286, po7287, po7288, po7289, po7290, po7291, po7292, po7293, po7294, po7295, po7296, po7297, po7298, po7299, po7300, po7301, po7302, po7303, po7304, po7305, po7306, po7307, po7308, po7309, po7310, po7311, po7312, po7313, po7314, po7315, po7316, po7317, po7318, po7319, po7320, po7321, po7322, po7323, po7324, po7325, po7326, po7327, po7328, po7329, po7330, po7331, po7332, po7333, po7334, po7335, po7336, po7337, po7338, po7339, po7340, po7341, po7342, po7343, po7344, po7345, po7346, po7347, po7348, po7349, po7350, po7351, po7352, po7353, po7354, po7355, po7356, po7357, po7358, po7359, po7360, po7361, po7362, po7363, po7364, po7365, po7366, po7367, po7368, po7369, po7370, po7371, po7372, po7373, po7374, po7375, po7376, po7377, po7378, po7379, po7380, po7381, po7382, po7383, po7384, po7385, po7386, po7387, po7388, po7389, po7390, po7391, po7392, po7393, po7394, po7395, po7396, po7397, po7398, po7399, po7400, po7401, po7402, po7403, po7404, po7405, po7406, po7407, po7408, po7409, po7410, po7411, po7412, po7413, po7414, po7415, po7416, po7417, po7418, po7419, po7420, po7421, po7422, po7423, po7424, po7425, po7426, po7427, po7428, po7429, po7430, po7431, po7432, po7433, po7434, po7435, po7436, po7437, po7438, po7439, po7440, po7441, po7442, po7443, po7444, po7445, po7446, po7447, po7448, po7449, po7450, po7451, po7452, po7453, po7454, po7455, po7456, po7457, po7458, po7459, po7460, po7461, po7462, po7463, po7464, po7465, po7466, po7467, po7468, po7469, po7470, po7471, po7472, po7473, po7474, po7475, po7476, po7477, po7478, po7479, po7480, po7481, po7482, po7483, po7484, po7485, po7486, po7487, po7488, po7489, po7490, po7491, po7492, po7493, po7494, po7495, po7496, po7497, po7498, po7499, po7500, po7501, po7502, po7503, po7504, po7505, po7506, po7507, po7508, po7509, po7510, po7511, po7512, po7513, po7514, po7515, po7516, po7517, po7518, po7519, po7520, po7521, po7522, po7523, po7524, po7525, po7526, po7527, po7528, po7529, po7530, po7531, po7532, po7533, po7534, po7535, po7536, po7537, po7538, po7539, po7540, po7541, po7542, po7543, po7544, po7545, po7546, po7547, po7548, po7549, po7550, po7551, po7552, po7553, po7554, po7555, po7556, po7557, po7558, po7559, po7560, po7561, po7562, po7563, po7564, po7565, po7566, po7567, po7568, po7569, po7570, po7571, po7572, po7573, po7574, po7575, po7576, po7577, po7578, po7579, po7580, po7581, po7582, po7583, po7584, po7585, po7586, po7587, po7588, po7589, po7590, po7591, po7592, po7593, po7594, po7595, po7596, po7597, po7598, po7599, po7600, po7601, po7602, po7603, po7604, po7605, po7606, po7607, po7608, po7609, po7610, po7611, po7612, po7613, po7614, po7615, po7616, po7617, po7618, po7619, po7620, po7621, po7622, po7623, po7624, po7625, po7626, po7627, po7628, po7629, po7630, po7631, po7632, po7633, po7634, po7635, po7636, po7637, po7638, po7639, po7640, po7641, po7642, po7643, po7644, po7645, po7646, po7647, po7648, po7649, po7650, po7651, po7652, po7653, po7654, po7655, po7656, po7657, po7658, po7659, po7660, po7661, po7662, po7663, po7664, po7665, po7666, po7667, po7668, po7669, po7670, po7671, po7672, po7673, po7674, po7675, po7676, po7677, po7678, po7679, po7680, po7681, po7682, po7683, po7684, po7685, po7686, po7687, po7688, po7689, po7690, po7691, po7692, po7693, po7694, po7695, po7696, po7697, po7698, po7699, po7700, po7701, po7702, po7703, po7704, po7705, po7706, po7707, po7708, po7709, po7710, po7711, po7712, po7713, po7714, po7715, po7716, po7717, po7718, po7719, po7720, po7721, po7722, po7723, po7724, po7725, po7726, po7727, po7728, po7729, po7730, po7731, po7732, po7733, po7734, po7735, po7736, po7737, po7738, po7739, po7740, po7741, po7742, po7743, po7744, po7745, po7746, po7747, po7748, po7749, po7750, po7751, po7752, po7753, po7754, po7755, po7756, po7757, po7758, po7759, po7760, po7761, po7762, po7763, po7764, po7765, po7766, po7767, po7768, po7769, po7770, po7771, po7772, po7773, po7774, po7775, po7776, po7777, po7778, po7779, po7780, po7781, po7782, po7783, po7784, po7785, po7786, po7787, po7788, po7789, po7790, po7791, po7792, po7793, po7794, po7795, po7796, po7797, po7798, po7799, po7800, po7801, po7802, po7803, po7804, po7805, po7806, po7807, po7808, po7809, po7810, po7811, po7812, po7813, po7814, po7815, po7816, po7817, po7818, po7819, po7820, po7821, po7822, po7823, po7824, po7825, po7826, po7827, po7828, po7829, po7830, po7831, po7832, po7833, po7834, po7835, po7836, po7837, po7838, po7839, po7840, po7841, po7842, po7843, po7844, po7845, po7846, po7847, po7848, po7849, po7850, po7851, po7852, po7853, po7854, po7855, po7856, po7857, po7858, po7859, po7860, po7861, po7862, po7863, po7864, po7865, po7866, po7867, po7868, po7869, po7870, po7871, po7872, po7873, po7874, po7875, po7876, po7877, po7878, po7879, po7880, po7881, po7882, po7883, po7884, po7885, po7886, po7887, po7888, po7889, po7890, po7891, po7892, po7893, po7894, po7895, po7896, po7897, po7898, po7899, po7900, po7901, po7902, po7903, po7904, po7905, po7906, po7907, po7908, po7909, po7910, po7911, po7912, po7913, po7914, po7915, po7916, po7917, po7918, po7919, po7920, po7921, po7922, po7923, po7924, po7925, po7926, po7927, po7928, po7929, po7930, po7931, po7932, po7933, po7934, po7935, po7936, po7937, po7938, po7939, po7940, po7941, po7942, po7943, po7944, po7945, po7946, po7947, po7948, po7949, po7950, po7951, po7952, po7953, po7954, po7955, po7956, po7957, po7958, po7959, po7960, po7961, po7962, po7963, po7964, po7965, po7966, po7967, po7968, po7969, po7970, po7971, po7972, po7973, po7974, po7975, po7976, po7977, po7978, po7979, po7980, po7981, po7982, po7983, po7984, po7985, po7986, po7987, po7988, po7989, po7990, po7991, po7992, po7993, po7994, po7995, po7996, po7997, po7998, po7999, po8000, po8001, po8002, po8003, po8004, po8005, po8006, po8007, po8008, po8009, po8010, po8011, po8012, po8013, po8014, po8015, po8016, po8017, po8018, po8019, po8020, po8021, po8022, po8023, po8024, po8025, po8026, po8027, po8028, po8029, po8030, po8031, po8032, po8033, po8034, po8035, po8036, po8037, po8038, po8039, po8040, po8041, po8042, po8043, po8044, po8045, po8046, po8047, po8048, po8049, po8050, po8051, po8052, po8053, po8054, po8055, po8056, po8057, po8058, po8059, po8060, po8061, po8062, po8063, po8064, po8065, po8066, po8067, po8068, po8069, po8070, po8071, po8072, po8073, po8074, po8075, po8076, po8077, po8078, po8079, po8080, po8081, po8082, po8083, po8084, po8085, po8086, po8087, po8088, po8089, po8090, po8091, po8092, po8093, po8094, po8095, po8096, po8097, po8098, po8099, po8100, po8101, po8102, po8103, po8104, po8105, po8106, po8107, po8108, po8109, po8110, po8111, po8112, po8113, po8114, po8115, po8116, po8117, po8118, po8119, po8120, po8121, po8122, po8123, po8124, po8125, po8126, po8127, po8128, po8129, po8130, po8131, po8132, po8133, po8134, po8135, po8136, po8137, po8138, po8139, po8140, po8141, po8142, po8143, po8144, po8145, po8146, po8147, po8148, po8149, po8150, po8151, po8152, po8153, po8154, po8155, po8156, po8157, po8158, po8159, po8160, po8161, po8162, po8163, po8164, po8165, po8166, po8167, po8168, po8169, po8170, po8171, po8172, po8173, po8174, po8175, po8176, po8177, po8178, po8179, po8180, po8181, po8182, po8183, po8184, po8185, po8186, po8187, po8188, po8189, po8190, po8191, po8192, po8193, po8194, po8195, po8196, po8197, po8198, po8199, po8200, po8201, po8202, po8203, po8204, po8205, po8206, po8207, po8208, po8209, po8210, po8211, po8212, po8213, po8214, po8215, po8216, po8217, po8218, po8219, po8220, po8221, po8222, po8223, po8224, po8225, po8226, po8227, po8228, po8229, po8230, po8231, po8232, po8233, po8234, po8235, po8236, po8237, po8238, po8239, po8240, po8241, po8242, po8243, po8244, po8245, po8246, po8247, po8248, po8249, po8250, po8251, po8252, po8253, po8254, po8255, po8256, po8257, po8258, po8259, po8260, po8261, po8262, po8263, po8264, po8265, po8266, po8267, po8268, po8269, po8270, po8271, po8272, po8273, po8274, po8275, po8276, po8277, po8278, po8279, po8280, po8281, po8282, po8283, po8284, po8285, po8286, po8287, po8288, po8289, po8290, po8291, po8292, po8293, po8294, po8295, po8296, po8297, po8298, po8299, po8300, po8301, po8302, po8303, po8304, po8305, po8306, po8307, po8308, po8309, po8310, po8311, po8312, po8313, po8314, po8315, po8316, po8317, po8318, po8319, po8320, po8321, po8322, po8323, po8324, po8325, po8326, po8327, po8328, po8329, po8330, po8331, po8332, po8333, po8334, po8335, po8336, po8337, po8338, po8339, po8340, po8341, po8342, po8343, po8344, po8345, po8346, po8347, po8348, po8349, po8350, po8351, po8352, po8353, po8354, po8355, po8356, po8357, po8358, po8359, po8360, po8361, po8362, po8363, po8364, po8365, po8366, po8367, po8368, po8369, po8370, po8371, po8372, po8373, po8374, po8375, po8376, po8377, po8378, po8379, po8380, po8381, po8382, po8383, po8384, po8385, po8386, po8387, po8388, po8389, po8390, po8391, po8392, po8393, po8394, po8395, po8396, po8397, po8398, po8399, po8400, po8401, po8402, po8403, po8404, po8405, po8406, po8407, po8408, po8409, po8410, po8411, po8412, po8413, po8414, po8415, po8416, po8417, po8418, po8419, po8420, po8421, po8422, po8423, po8424, po8425, po8426, po8427, po8428, po8429, po8430, po8431, po8432, po8433, po8434, po8435, po8436, po8437, po8438, po8439, po8440, po8441, po8442, po8443, po8444, po8445, po8446, po8447, po8448, po8449, po8450, po8451, po8452, po8453, po8454, po8455, po8456, po8457, po8458, po8459, po8460, po8461, po8462, po8463, po8464, po8465, po8466, po8467, po8468, po8469, po8470, po8471, po8472, po8473, po8474, po8475, po8476, po8477, po8478, po8479, po8480, po8481, po8482, po8483, po8484, po8485, po8486, po8487, po8488, po8489, po8490, po8491, po8492, po8493, po8494, po8495, po8496, po8497, po8498, po8499, po8500, po8501, po8502, po8503, po8504, po8505, po8506, po8507, po8508, po8509, po8510, po8511, po8512, po8513, po8514, po8515, po8516, po8517, po8518, po8519, po8520, po8521, po8522, po8523, po8524, po8525, po8526, po8527, po8528, po8529, po8530, po8531, po8532, po8533, po8534, po8535, po8536, po8537, po8538, po8539, po8540, po8541, po8542, po8543, po8544, po8545, po8546, po8547, po8548, po8549, po8550, po8551, po8552, po8553, po8554, po8555, po8556, po8557, po8558, po8559, po8560, po8561, po8562, po8563, po8564, po8565, po8566, po8567, po8568, po8569, po8570, po8571, po8572, po8573, po8574, po8575, po8576, po8577, po8578, po8579, po8580, po8581, po8582, po8583, po8584, po8585, po8586, po8587, po8588, po8589, po8590, po8591, po8592, po8593, po8594, po8595, po8596, po8597, po8598, po8599, po8600, po8601, po8602, po8603, po8604, po8605, po8606, po8607, po8608, po8609, po8610, po8611, po8612, po8613, po8614, po8615, po8616, po8617, po8618, po8619, po8620, po8621, po8622, po8623, po8624, po8625, po8626, po8627, po8628, po8629, po8630, po8631, po8632, po8633, po8634, po8635, po8636, po8637, po8638, po8639, po8640, po8641, po8642, po8643, po8644, po8645, po8646, po8647, po8648, po8649, po8650, po8651, po8652, po8653, po8654, po8655, po8656, po8657, po8658, po8659, po8660, po8661, po8662, po8663, po8664, po8665, po8666, po8667, po8668, po8669, po8670, po8671, po8672, po8673, po8674, po8675, po8676, po8677, po8678, po8679, po8680, po8681, po8682, po8683, po8684, po8685, po8686, po8687, po8688, po8689, po8690, po8691, po8692, po8693, po8694, po8695, po8696, po8697, po8698, po8699, po8700, po8701, po8702, po8703, po8704, po8705, po8706, po8707, po8708, po8709, po8710, po8711, po8712, po8713, po8714, po8715, po8716, po8717, po8718, po8719, po8720, po8721, po8722, po8723, po8724, po8725, po8726, po8727, po8728, po8729, po8730, po8731, po8732, po8733, po8734, po8735, po8736, po8737, po8738, po8739, po8740, po8741, po8742, po8743, po8744, po8745, po8746, po8747, po8748, po8749, po8750, po8751, po8752, po8753, po8754, po8755, po8756, po8757, po8758, po8759, po8760, po8761, po8762, po8763, po8764, po8765, po8766, po8767, po8768, po8769, po8770, po8771, po8772, po8773, po8774, po8775, po8776, po8777, po8778, po8779, po8780, po8781, po8782, po8783, po8784, po8785, po8786, po8787, po8788, po8789, po8790, po8791, po8792, po8793, po8794, po8795, po8796, po8797, po8798, po8799, po8800, po8801, po8802, po8803, po8804, po8805, po8806, po8807, po8808, po8809, po8810, po8811, po8812, po8813, po8814, po8815, po8816, po8817, po8818, po8819, po8820, po8821, po8822, po8823, po8824, po8825, po8826, po8827, po8828, po8829, po8830, po8831, po8832, po8833, po8834, po8835, po8836, po8837, po8838, po8839, po8840, po8841, po8842, po8843, po8844, po8845, po8846, po8847, po8848, po8849, po8850, po8851, po8852, po8853, po8854, po8855, po8856, po8857, po8858, po8859, po8860, po8861, po8862, po8863, po8864, po8865, po8866, po8867, po8868, po8869, po8870, po8871, po8872, po8873, po8874, po8875, po8876, po8877, po8878, po8879, po8880, po8881, po8882, po8883, po8884, po8885, po8886, po8887, po8888, po8889, po8890, po8891, po8892, po8893, po8894, po8895, po8896, po8897, po8898, po8899, po8900, po8901, po8902, po8903, po8904, po8905, po8906, po8907, po8908, po8909, po8910, po8911, po8912, po8913, po8914, po8915, po8916, po8917, po8918, po8919, po8920, po8921, po8922, po8923, po8924, po8925, po8926, po8927, po8928, po8929, po8930, po8931, po8932, po8933, po8934, po8935, po8936, po8937, po8938, po8939, po8940, po8941, po8942, po8943, po8944, po8945, po8946, po8947, po8948, po8949, po8950, po8951, po8952, po8953, po8954, po8955, po8956, po8957, po8958, po8959, po8960, po8961, po8962, po8963, po8964, po8965, po8966, po8967, po8968, po8969, po8970, po8971, po8972, po8973, po8974, po8975, po8976, po8977, po8978, po8979, po8980, po8981, po8982, po8983, po8984, po8985, po8986, po8987, po8988, po8989, po8990, po8991, po8992, po8993, po8994, po8995, po8996, po8997, po8998, po8999, po9000, po9001, po9002, po9003, po9004, po9005, po9006, po9007, po9008, po9009, po9010, po9011, po9012, po9013, po9014, po9015, po9016, po9017, po9018, po9019, po9020, po9021, po9022, po9023, po9024, po9025, po9026, po9027, po9028, po9029, po9030, po9031, po9032, po9033, po9034, po9035, po9036, po9037);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518, pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526, pi3527, pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535, pi3536, pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544, pi3545, pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553, pi3554, pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562, pi3563, pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571, pi3572, pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580, pi3581, pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589, pi3590, pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598, pi3599, pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607, pi3608, pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616, pi3617, pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625, pi3626, pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634, pi3635, pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643, pi3644, pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652, pi3653, pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661, pi3662, pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670, pi3671, pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679, pi3680, pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688, pi3689, pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697, pi3698, pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706, pi3707, pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715, pi3716, pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724, pi3725, pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733, pi3734, pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742, pi3743, pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751, pi3752, pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760, pi3761, pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769, pi3770, pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778, pi3779, pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787, pi3788, pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796, pi3797, pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805, pi3806, pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814, pi3815, pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823, pi3824, pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832, pi3833, pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841, pi3842, pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850, pi3851, pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859, pi3860, pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868, pi3869, pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877, pi3878, pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886, pi3887, pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895, pi3896, pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904, pi3905, pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913, pi3914, pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922, pi3923, pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931, pi3932, pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940, pi3941, pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949, pi3950, pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958, pi3959, pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967, pi3968, pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976, pi3977, pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985, pi3986, pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994, pi3995, pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003, pi4004, pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012, pi4013, pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021, pi4022, pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030, pi4031, pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039, pi4040, pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048, pi4049, pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057, pi4058, pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066, pi4067, pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075, pi4076, pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084, pi4085, pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093, pi4094, pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102, pi4103, pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111, pi4112, pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120, pi4121, pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129, pi4130, pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138, pi4139, pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147, pi4148, pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156, pi4157, pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165, pi4166, pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174, pi4175, pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183, pi4184, pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192, pi4193, pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201, pi4202, pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210, pi4211, pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219, pi4220, pi4221, pi4222, pi4223, pi4224, pi4225, pi4226, pi4227, pi4228, pi4229, pi4230, pi4231, pi4232, pi4233, pi4234, pi4235, pi4236, pi4237, pi4238, pi4239, pi4240, pi4241, pi4242, pi4243, pi4244, pi4245, pi4246, pi4247, pi4248, pi4249, pi4250, pi4251, pi4252, pi4253, pi4254, pi4255, pi4256, pi4257, pi4258, pi4259, pi4260, pi4261, pi4262, pi4263, pi4264, pi4265, pi4266, pi4267, pi4268, pi4269, pi4270, pi4271, pi4272, pi4273, pi4274, pi4275, pi4276, pi4277, pi4278, pi4279, pi4280, pi4281, pi4282, pi4283, pi4284, pi4285, pi4286, pi4287, pi4288, pi4289, pi4290, pi4291, pi4292, pi4293, pi4294, pi4295, pi4296, pi4297, pi4298, pi4299, pi4300, pi4301, pi4302, pi4303, pi4304, pi4305, pi4306, pi4307, pi4308, pi4309, pi4310, pi4311, pi4312, pi4313, pi4314, pi4315, pi4316, pi4317, pi4318, pi4319, pi4320, pi4321, pi4322, pi4323, pi4324, pi4325, pi4326, pi4327, pi4328, pi4329, pi4330, pi4331, pi4332, pi4333, pi4334, pi4335, pi4336, pi4337, pi4338, pi4339, pi4340, pi4341, pi4342, pi4343, pi4344, pi4345, pi4346, pi4347, pi4348, pi4349, pi4350, pi4351, pi4352, pi4353, pi4354, pi4355, pi4356, pi4357, pi4358, pi4359, pi4360, pi4361, pi4362, pi4363, pi4364, pi4365, pi4366, pi4367, pi4368, pi4369, pi4370, pi4371, pi4372, pi4373, pi4374, pi4375, pi4376, pi4377, pi4378, pi4379, pi4380, pi4381, pi4382, pi4383, pi4384, pi4385, pi4386, pi4387, pi4388, pi4389, pi4390, pi4391, pi4392, pi4393, pi4394, pi4395, pi4396, pi4397, pi4398, pi4399, pi4400, pi4401, pi4402, pi4403, pi4404, pi4405, pi4406, pi4407, pi4408, pi4409, pi4410, pi4411, pi4412, pi4413, pi4414, pi4415, pi4416, pi4417, pi4418, pi4419, pi4420, pi4421, pi4422, pi4423, pi4424, pi4425, pi4426, pi4427, pi4428, pi4429, pi4430, pi4431, pi4432, pi4433, pi4434, pi4435, pi4436, pi4437, pi4438, pi4439, pi4440, pi4441, pi4442, pi4443, pi4444, pi4445, pi4446, pi4447, pi4448, pi4449, pi4450, pi4451, pi4452, pi4453, pi4454, pi4455, pi4456, pi4457, pi4458, pi4459, pi4460, pi4461, pi4462, pi4463, pi4464, pi4465, pi4466, pi4467, pi4468, pi4469, pi4470, pi4471, pi4472, pi4473, pi4474, pi4475, pi4476, pi4477, pi4478, pi4479, pi4480, pi4481, pi4482, pi4483, pi4484, pi4485, pi4486, pi4487, pi4488, pi4489, pi4490, pi4491, pi4492, pi4493, pi4494, pi4495, pi4496, pi4497, pi4498, pi4499, pi4500, pi4501, pi4502, pi4503, pi4504, pi4505, pi4506, pi4507, pi4508, pi4509, pi4510, pi4511, pi4512, pi4513, pi4514, pi4515, pi4516, pi4517, pi4518, pi4519, pi4520, pi4521, pi4522, pi4523, pi4524, pi4525, pi4526, pi4527, pi4528, pi4529, pi4530, pi4531, pi4532, pi4533, pi4534, pi4535, pi4536, pi4537, pi4538, pi4539, pi4540, pi4541, pi4542, pi4543, pi4544, pi4545, pi4546, pi4547, pi4548, pi4549, pi4550, pi4551, pi4552, pi4553, pi4554, pi4555, pi4556, pi4557, pi4558, pi4559, pi4560, pi4561, pi4562, pi4563, pi4564, pi4565, pi4566, pi4567, pi4568, pi4569, pi4570, pi4571, pi4572, pi4573, pi4574, pi4575, pi4576, pi4577, pi4578, pi4579, pi4580, pi4581, pi4582, pi4583, pi4584, pi4585, pi4586, pi4587, pi4588, pi4589, pi4590, pi4591, pi4592, pi4593, pi4594, pi4595, pi4596, pi4597, pi4598, pi4599, pi4600, pi4601, pi4602, pi4603, pi4604, pi4605, pi4606, pi4607, pi4608, pi4609, pi4610, pi4611, pi4612, pi4613, pi4614, pi4615, pi4616, pi4617, pi4618, pi4619, pi4620, pi4621, pi4622, pi4623, pi4624, pi4625, pi4626, pi4627, pi4628, pi4629, pi4630, pi4631, pi4632, pi4633, pi4634, pi4635, pi4636, pi4637, pi4638, pi4639, pi4640, pi4641, pi4642, pi4643, pi4644, pi4645, pi4646, pi4647, pi4648, pi4649, pi4650, pi4651, pi4652, pi4653, pi4654, pi4655, pi4656, pi4657, pi4658, pi4659, pi4660, pi4661, pi4662, pi4663, pi4664, pi4665, pi4666, pi4667, pi4668, pi4669, pi4670, pi4671, pi4672, pi4673, pi4674, pi4675, pi4676, pi4677, pi4678, pi4679, pi4680, pi4681, pi4682, pi4683, pi4684, pi4685, pi4686, pi4687, pi4688, pi4689, pi4690, pi4691, pi4692, pi4693, pi4694, pi4695, pi4696, pi4697, pi4698, pi4699, pi4700, pi4701, pi4702, pi4703, pi4704, pi4705, pi4706, pi4707, pi4708, pi4709, pi4710, pi4711, pi4712, pi4713, pi4714, pi4715, pi4716, pi4717, pi4718, pi4719, pi4720, pi4721, pi4722, pi4723, pi4724, pi4725, pi4726, pi4727, pi4728, pi4729, pi4730, pi4731, pi4732, pi4733, pi4734, pi4735, pi4736, pi4737, pi4738, pi4739, pi4740, pi4741, pi4742, pi4743, pi4744, pi4745, pi4746, pi4747, pi4748, pi4749, pi4750, pi4751, pi4752, pi4753, pi4754, pi4755, pi4756, pi4757, pi4758, pi4759, pi4760, pi4761, pi4762, pi4763, pi4764, pi4765, pi4766, pi4767, pi4768, pi4769, pi4770, pi4771, pi4772, pi4773, pi4774, pi4775, pi4776, pi4777, pi4778, pi4779, pi4780, pi4781, pi4782, pi4783, pi4784, pi4785, pi4786, pi4787, pi4788, pi4789, pi4790, pi4791, pi4792, pi4793, pi4794, pi4795, pi4796, pi4797, pi4798, pi4799, pi4800, pi4801, pi4802, pi4803, pi4804, pi4805, pi4806, pi4807, pi4808, pi4809, pi4810, pi4811, pi4812, pi4813, pi4814, pi4815, pi4816, pi4817, pi4818, pi4819, pi4820, pi4821, pi4822, pi4823, pi4824, pi4825, pi4826, pi4827, pi4828, pi4829, pi4830, pi4831, pi4832, pi4833, pi4834, pi4835, pi4836, pi4837, pi4838, pi4839, pi4840, pi4841, pi4842, pi4843, pi4844, pi4845, pi4846, pi4847, pi4848, pi4849, pi4850, pi4851, pi4852, pi4853, pi4854, pi4855, pi4856, pi4857, pi4858, pi4859, pi4860, pi4861, pi4862, pi4863, pi4864, pi4865, pi4866, pi4867, pi4868, pi4869, pi4870, pi4871, pi4872, pi4873, pi4874, pi4875, pi4876, pi4877, pi4878, pi4879, pi4880, pi4881, pi4882, pi4883, pi4884, pi4885, pi4886, pi4887, pi4888, pi4889, pi4890, pi4891, pi4892, pi4893, pi4894, pi4895, pi4896, pi4897, pi4898, pi4899, pi4900, pi4901, pi4902, pi4903, pi4904, pi4905, pi4906, pi4907, pi4908, pi4909, pi4910, pi4911, pi4912, pi4913, pi4914, pi4915, pi4916, pi4917, pi4918, pi4919, pi4920, pi4921, pi4922, pi4923, pi4924, pi4925, pi4926, pi4927, pi4928, pi4929, pi4930, pi4931, pi4932, pi4933, pi4934, pi4935, pi4936, pi4937, pi4938, pi4939, pi4940, pi4941, pi4942, pi4943, pi4944, pi4945, pi4946, pi4947, pi4948, pi4949, pi4950, pi4951, pi4952, pi4953, pi4954, pi4955, pi4956, pi4957, pi4958, pi4959, pi4960, pi4961, pi4962, pi4963, pi4964, pi4965, pi4966, pi4967, pi4968, pi4969, pi4970, pi4971, pi4972, pi4973, pi4974, pi4975, pi4976, pi4977, pi4978, pi4979, pi4980, pi4981, pi4982, pi4983, pi4984, pi4985, pi4986, pi4987, pi4988, pi4989, pi4990, pi4991, pi4992, pi4993, pi4994, pi4995, pi4996, pi4997, pi4998, pi4999, pi5000, pi5001, pi5002, pi5003, pi5004, pi5005, pi5006, pi5007, pi5008, pi5009, pi5010, pi5011, pi5012, pi5013, pi5014, pi5015, pi5016, pi5017, pi5018, pi5019, pi5020, pi5021, pi5022, pi5023, pi5024, pi5025, pi5026, pi5027, pi5028, pi5029, pi5030, pi5031, pi5032, pi5033, pi5034, pi5035, pi5036, pi5037, pi5038, pi5039, pi5040, pi5041, pi5042, pi5043, pi5044, pi5045, pi5046, pi5047, pi5048, pi5049, pi5050, pi5051, pi5052, pi5053, pi5054, pi5055, pi5056, pi5057, pi5058, pi5059, pi5060, pi5061, pi5062, pi5063, pi5064, pi5065, pi5066, pi5067, pi5068, pi5069, pi5070, pi5071, pi5072, pi5073, pi5074, pi5075, pi5076, pi5077, pi5078, pi5079, pi5080, pi5081, pi5082, pi5083, pi5084, pi5085, pi5086, pi5087, pi5088, pi5089, pi5090, pi5091, pi5092, pi5093, pi5094, pi5095, pi5096, pi5097, pi5098, pi5099, pi5100, pi5101, pi5102, pi5103, pi5104, pi5105, pi5106, pi5107, pi5108, pi5109, pi5110, pi5111, pi5112, pi5113, pi5114, pi5115, pi5116, pi5117, pi5118, pi5119, pi5120, pi5121, pi5122, pi5123, pi5124, pi5125, pi5126, pi5127, pi5128, pi5129, pi5130, pi5131, pi5132, pi5133, pi5134, pi5135, pi5136, pi5137, pi5138, pi5139, pi5140, pi5141, pi5142, pi5143, pi5144, pi5145, pi5146, pi5147, pi5148, pi5149, pi5150, pi5151, pi5152, pi5153, pi5154, pi5155, pi5156, pi5157, pi5158, pi5159, pi5160, pi5161, pi5162, pi5163, pi5164, pi5165, pi5166, pi5167, pi5168, pi5169, pi5170, pi5171, pi5172, pi5173, pi5174, pi5175, pi5176, pi5177, pi5178, pi5179, pi5180, pi5181, pi5182, pi5183, pi5184, pi5185, pi5186, pi5187, pi5188, pi5189, pi5190, pi5191, pi5192, pi5193, pi5194, pi5195, pi5196, pi5197, pi5198, pi5199, pi5200, pi5201, pi5202, pi5203, pi5204, pi5205, pi5206, pi5207, pi5208, pi5209, pi5210, pi5211, pi5212, pi5213, pi5214, pi5215, pi5216, pi5217, pi5218, pi5219, pi5220, pi5221, pi5222, pi5223, pi5224, pi5225, pi5226, pi5227, pi5228, pi5229, pi5230, pi5231, pi5232, pi5233, pi5234, pi5235, pi5236, pi5237, pi5238, pi5239, pi5240, pi5241, pi5242, pi5243, pi5244, pi5245, pi5246, pi5247, pi5248, pi5249, pi5250, pi5251, pi5252, pi5253, pi5254, pi5255, pi5256, pi5257, pi5258, pi5259, pi5260, pi5261, pi5262, pi5263, pi5264, pi5265, pi5266, pi5267, pi5268, pi5269, pi5270, pi5271, pi5272, pi5273, pi5274, pi5275, pi5276, pi5277, pi5278, pi5279, pi5280, pi5281, pi5282, pi5283, pi5284, pi5285, pi5286, pi5287, pi5288, pi5289, pi5290, pi5291, pi5292, pi5293, pi5294, pi5295, pi5296, pi5297, pi5298, pi5299, pi5300, pi5301, pi5302, pi5303, pi5304, pi5305, pi5306, pi5307, pi5308, pi5309, pi5310, pi5311, pi5312, pi5313, pi5314, pi5315, pi5316, pi5317, pi5318, pi5319, pi5320, pi5321, pi5322, pi5323, pi5324, pi5325, pi5326, pi5327, pi5328, pi5329, pi5330, pi5331, pi5332, pi5333, pi5334, pi5335, pi5336, pi5337, pi5338, pi5339, pi5340, pi5341, pi5342, pi5343, pi5344, pi5345, pi5346, pi5347, pi5348, pi5349, pi5350, pi5351, pi5352, pi5353, pi5354, pi5355, pi5356, pi5357, pi5358, pi5359, pi5360, pi5361, pi5362, pi5363, pi5364, pi5365, pi5366, pi5367, pi5368, pi5369, pi5370, pi5371, pi5372, pi5373, pi5374, pi5375, pi5376, pi5377, pi5378, pi5379, pi5380, pi5381, pi5382, pi5383, pi5384, pi5385, pi5386, pi5387, pi5388, pi5389, pi5390, pi5391, pi5392, pi5393, pi5394, pi5395, pi5396, pi5397, pi5398, pi5399, pi5400, pi5401, pi5402, pi5403, pi5404, pi5405, pi5406, pi5407, pi5408, pi5409, pi5410, pi5411, pi5412, pi5413, pi5414, pi5415, pi5416, pi5417, pi5418, pi5419, pi5420, pi5421, pi5422, pi5423, pi5424, pi5425, pi5426, pi5427, pi5428, pi5429, pi5430, pi5431, pi5432, pi5433, pi5434, pi5435, pi5436, pi5437, pi5438, pi5439, pi5440, pi5441, pi5442, pi5443, pi5444, pi5445, pi5446, pi5447, pi5448, pi5449, pi5450, pi5451, pi5452, pi5453, pi5454, pi5455, pi5456, pi5457, pi5458, pi5459, pi5460, pi5461, pi5462, pi5463, pi5464, pi5465, pi5466, pi5467, pi5468, pi5469, pi5470, pi5471, pi5472, pi5473, pi5474, pi5475, pi5476, pi5477, pi5478, pi5479, pi5480, pi5481, pi5482, pi5483, pi5484, pi5485, pi5486, pi5487, pi5488, pi5489, pi5490, pi5491, pi5492, pi5493, pi5494, pi5495, pi5496, pi5497, pi5498, pi5499, pi5500, pi5501, pi5502, pi5503, pi5504, pi5505, pi5506, pi5507, pi5508, pi5509, pi5510, pi5511, pi5512, pi5513, pi5514, pi5515, pi5516, pi5517, pi5518, pi5519, pi5520, pi5521, pi5522, pi5523, pi5524, pi5525, pi5526, pi5527, pi5528, pi5529, pi5530, pi5531, pi5532, pi5533, pi5534, pi5535, pi5536, pi5537, pi5538, pi5539, pi5540, pi5541, pi5542, pi5543, pi5544, pi5545, pi5546, pi5547, pi5548, pi5549, pi5550, pi5551, pi5552, pi5553, pi5554, pi5555, pi5556, pi5557, pi5558, pi5559, pi5560, pi5561, pi5562, pi5563, pi5564, pi5565, pi5566, pi5567, pi5568, pi5569, pi5570, pi5571, pi5572, pi5573, pi5574, pi5575, pi5576, pi5577, pi5578, pi5579, pi5580, pi5581, pi5582, pi5583, pi5584, pi5585, pi5586, pi5587, pi5588, pi5589, pi5590, pi5591, pi5592, pi5593, pi5594, pi5595, pi5596, pi5597, pi5598, pi5599, pi5600, pi5601, pi5602, pi5603, pi5604, pi5605, pi5606, pi5607, pi5608, pi5609, pi5610, pi5611, pi5612, pi5613, pi5614, pi5615, pi5616, pi5617, pi5618, pi5619, pi5620, pi5621, pi5622, pi5623, pi5624, pi5625, pi5626, pi5627, pi5628, pi5629, pi5630, pi5631, pi5632, pi5633, pi5634, pi5635, pi5636, pi5637, pi5638, pi5639, pi5640, pi5641, pi5642, pi5643, pi5644, pi5645, pi5646, pi5647, pi5648, pi5649, pi5650, pi5651, pi5652, pi5653, pi5654, pi5655, pi5656, pi5657, pi5658, pi5659, pi5660, pi5661, pi5662, pi5663, pi5664, pi5665, pi5666, pi5667, pi5668, pi5669, pi5670, pi5671, pi5672, pi5673, pi5674, pi5675, pi5676, pi5677, pi5678, pi5679, pi5680, pi5681, pi5682, pi5683, pi5684, pi5685, pi5686, pi5687, pi5688, pi5689, pi5690, pi5691, pi5692, pi5693, pi5694, pi5695, pi5696, pi5697, pi5698, pi5699, pi5700, pi5701, pi5702, pi5703, pi5704, pi5705, pi5706, pi5707, pi5708, pi5709, pi5710, pi5711, pi5712, pi5713, pi5714, pi5715, pi5716, pi5717, pi5718, pi5719, pi5720, pi5721, pi5722, pi5723, pi5724, pi5725, pi5726, pi5727, pi5728, pi5729, pi5730, pi5731, pi5732, pi5733, pi5734, pi5735, pi5736, pi5737, pi5738, pi5739, pi5740, pi5741, pi5742, pi5743, pi5744, pi5745, pi5746, pi5747, pi5748, pi5749, pi5750, pi5751, pi5752, pi5753, pi5754, pi5755, pi5756, pi5757, pi5758, pi5759, pi5760, pi5761, pi5762, pi5763, pi5764, pi5765, pi5766, pi5767, pi5768, pi5769, pi5770, pi5771, pi5772, pi5773, pi5774, pi5775, pi5776, pi5777, pi5778, pi5779, pi5780, pi5781, pi5782, pi5783, pi5784, pi5785, pi5786, pi5787, pi5788, pi5789, pi5790, pi5791, pi5792, pi5793, pi5794, pi5795, pi5796, pi5797, pi5798, pi5799, pi5800, pi5801, pi5802, pi5803, pi5804, pi5805, pi5806, pi5807, pi5808, pi5809, pi5810, pi5811, pi5812, pi5813, pi5814, pi5815, pi5816, pi5817, pi5818, pi5819, pi5820, pi5821, pi5822, pi5823, pi5824, pi5825, pi5826, pi5827, pi5828, pi5829, pi5830, pi5831, pi5832, pi5833, pi5834, pi5835, pi5836, pi5837, pi5838, pi5839, pi5840, pi5841, pi5842, pi5843, pi5844, pi5845, pi5846, pi5847, pi5848, pi5849, pi5850, pi5851, pi5852, pi5853, pi5854, pi5855, pi5856, pi5857, pi5858, pi5859, pi5860, pi5861, pi5862, pi5863, pi5864, pi5865, pi5866, pi5867, pi5868, pi5869, pi5870, pi5871, pi5872, pi5873, pi5874, pi5875, pi5876, pi5877, pi5878, pi5879, pi5880, pi5881, pi5882, pi5883, pi5884, pi5885, pi5886, pi5887, pi5888, pi5889, pi5890, pi5891, pi5892, pi5893, pi5894, pi5895, pi5896, pi5897, pi5898, pi5899, pi5900, pi5901, pi5902, pi5903, pi5904, pi5905, pi5906, pi5907, pi5908, pi5909, pi5910, pi5911, pi5912, pi5913, pi5914, pi5915, pi5916, pi5917, pi5918, pi5919, pi5920, pi5921, pi5922, pi5923, pi5924, pi5925, pi5926, pi5927, pi5928, pi5929, pi5930, pi5931, pi5932, pi5933, pi5934, pi5935, pi5936, pi5937, pi5938, pi5939, pi5940, pi5941, pi5942, pi5943, pi5944, pi5945, pi5946, pi5947, pi5948, pi5949, pi5950, pi5951, pi5952, pi5953, pi5954, pi5955, pi5956, pi5957, pi5958, pi5959, pi5960, pi5961, pi5962, pi5963, pi5964, pi5965, pi5966, pi5967, pi5968, pi5969, pi5970, pi5971, pi5972, pi5973, pi5974, pi5975, pi5976, pi5977, pi5978, pi5979, pi5980, pi5981, pi5982, pi5983, pi5984, pi5985, pi5986, pi5987, pi5988, pi5989, pi5990, pi5991, pi5992, pi5993, pi5994, pi5995, pi5996, pi5997, pi5998, pi5999, pi6000, pi6001, pi6002, pi6003, pi6004, pi6005, pi6006, pi6007, pi6008, pi6009, pi6010, pi6011, pi6012, pi6013, pi6014, pi6015, pi6016, pi6017, pi6018, pi6019, pi6020, pi6021, pi6022, pi6023, pi6024, pi6025, pi6026, pi6027, pi6028, pi6029, pi6030, pi6031, pi6032, pi6033, pi6034, pi6035, pi6036, pi6037, pi6038, pi6039, pi6040, pi6041, pi6042, pi6043, pi6044, pi6045, pi6046, pi6047, pi6048, pi6049, pi6050, pi6051, pi6052, pi6053, pi6054, pi6055, pi6056, pi6057, pi6058, pi6059, pi6060, pi6061, pi6062, pi6063, pi6064, pi6065, pi6066, pi6067, pi6068, pi6069, pi6070, pi6071, pi6072, pi6073, pi6074, pi6075, pi6076, pi6077, pi6078, pi6079, pi6080, pi6081, pi6082, pi6083, pi6084, pi6085, pi6086, pi6087, pi6088, pi6089, pi6090, pi6091, pi6092, pi6093, pi6094, pi6095, pi6096, pi6097, pi6098, pi6099, pi6100, pi6101, pi6102, pi6103, pi6104, pi6105, pi6106, pi6107, pi6108, pi6109, pi6110, pi6111, pi6112, pi6113, pi6114, pi6115, pi6116, pi6117, pi6118, pi6119, pi6120, pi6121, pi6122, pi6123, pi6124, pi6125, pi6126, pi6127, pi6128, pi6129, pi6130, pi6131, pi6132, pi6133, pi6134, pi6135, pi6136, pi6137, pi6138, pi6139, pi6140, pi6141, pi6142, pi6143, pi6144, pi6145, pi6146, pi6147, pi6148, pi6149, pi6150, pi6151, pi6152, pi6153, pi6154, pi6155, pi6156, pi6157, pi6158, pi6159, pi6160, pi6161, pi6162, pi6163, pi6164, pi6165, pi6166, pi6167, pi6168, pi6169, pi6170, pi6171, pi6172, pi6173, pi6174, pi6175, pi6176, pi6177, pi6178, pi6179, pi6180, pi6181, pi6182, pi6183, pi6184, pi6185, pi6186, pi6187, pi6188, pi6189, pi6190, pi6191, pi6192, pi6193, pi6194, pi6195, pi6196, pi6197, pi6198, pi6199, pi6200, pi6201, pi6202, pi6203, pi6204, pi6205, pi6206, pi6207, pi6208, pi6209, pi6210, pi6211, pi6212, pi6213, pi6214, pi6215, pi6216, pi6217, pi6218, pi6219, pi6220, pi6221, pi6222, pi6223, pi6224, pi6225, pi6226, pi6227, pi6228, pi6229, pi6230, pi6231, pi6232, pi6233, pi6234, pi6235, pi6236, pi6237, pi6238, pi6239, pi6240, pi6241, pi6242, pi6243, pi6244, pi6245, pi6246, pi6247, pi6248, pi6249, pi6250, pi6251, pi6252, pi6253, pi6254, pi6255, pi6256, pi6257, pi6258, pi6259, pi6260, pi6261, pi6262, pi6263, pi6264, pi6265, pi6266, pi6267, pi6268, pi6269, pi6270, pi6271, pi6272, pi6273, pi6274, pi6275, pi6276, pi6277, pi6278, pi6279, pi6280, pi6281, pi6282, pi6283, pi6284, pi6285, pi6286, pi6287, pi6288, pi6289, pi6290, pi6291, pi6292, pi6293, pi6294, pi6295, pi6296, pi6297, pi6298, pi6299, pi6300, pi6301, pi6302, pi6303, pi6304, pi6305, pi6306, pi6307, pi6308, pi6309, pi6310, pi6311, pi6312, pi6313, pi6314, pi6315, pi6316, pi6317, pi6318, pi6319, pi6320, pi6321, pi6322, pi6323, pi6324, pi6325, pi6326, pi6327, pi6328, pi6329, pi6330, pi6331, pi6332, pi6333, pi6334, pi6335, pi6336, pi6337, pi6338, pi6339, pi6340, pi6341, pi6342, pi6343, pi6344, pi6345, pi6346, pi6347, pi6348, pi6349, pi6350, pi6351, pi6352, pi6353, pi6354, pi6355, pi6356, pi6357, pi6358, pi6359, pi6360, pi6361, pi6362, pi6363, pi6364, pi6365, pi6366, pi6367, pi6368, pi6369, pi6370, pi6371, pi6372, pi6373, pi6374, pi6375, pi6376, pi6377, pi6378, pi6379, pi6380, pi6381, pi6382, pi6383, pi6384, pi6385, pi6386, pi6387, pi6388, pi6389, pi6390, pi6391, pi6392, pi6393, pi6394, pi6395, pi6396, pi6397, pi6398, pi6399, pi6400, pi6401, pi6402, pi6403, pi6404, pi6405, pi6406, pi6407, pi6408, pi6409, pi6410, pi6411, pi6412, pi6413, pi6414, pi6415, pi6416, pi6417, pi6418, pi6419, pi6420, pi6421, pi6422, pi6423, pi6424, pi6425, pi6426, pi6427, pi6428, pi6429, pi6430, pi6431, pi6432, pi6433, pi6434, pi6435, pi6436, pi6437, pi6438, pi6439, pi6440, pi6441, pi6442, pi6443, pi6444, pi6445, pi6446, pi6447, pi6448, pi6449, pi6450, pi6451, pi6452, pi6453, pi6454, pi6455, pi6456, pi6457, pi6458, pi6459, pi6460, pi6461, pi6462, pi6463, pi6464, pi6465, pi6466, pi6467, pi6468, pi6469, pi6470, pi6471, pi6472, pi6473, pi6474, pi6475, pi6476, pi6477, pi6478, pi6479, pi6480, pi6481, pi6482, pi6483, pi6484, pi6485, pi6486, pi6487, pi6488, pi6489, pi6490, pi6491, pi6492, pi6493, pi6494, pi6495, pi6496, pi6497, pi6498, pi6499, pi6500, pi6501, pi6502, pi6503, pi6504, pi6505, pi6506, pi6507, pi6508, pi6509, pi6510, pi6511, pi6512, pi6513, pi6514, pi6515, pi6516, pi6517, pi6518, pi6519, pi6520, pi6521, pi6522, pi6523, pi6524, pi6525, pi6526, pi6527, pi6528, pi6529, pi6530, pi6531, pi6532, pi6533, pi6534, pi6535, pi6536, pi6537, pi6538, pi6539, pi6540, pi6541, pi6542, pi6543, pi6544, pi6545, pi6546, pi6547, pi6548, pi6549, pi6550, pi6551, pi6552, pi6553, pi6554, pi6555, pi6556, pi6557, pi6558, pi6559, pi6560, pi6561, pi6562, pi6563, pi6564, pi6565, pi6566, pi6567, pi6568, pi6569, pi6570, pi6571, pi6572, pi6573, pi6574, pi6575, pi6576, pi6577, pi6578, pi6579, pi6580, pi6581, pi6582, pi6583, pi6584, pi6585, pi6586, pi6587, pi6588, pi6589, pi6590, pi6591, pi6592, pi6593, pi6594, pi6595, pi6596, pi6597, pi6598, pi6599, pi6600, pi6601, pi6602, pi6603, pi6604, pi6605, pi6606, pi6607, pi6608, pi6609, pi6610, pi6611, pi6612, pi6613, pi6614, pi6615, pi6616, pi6617, pi6618, pi6619, pi6620, pi6621, pi6622, pi6623, pi6624, pi6625, pi6626, pi6627, pi6628, pi6629, pi6630, pi6631, pi6632, pi6633, pi6634, pi6635, pi6636, pi6637, pi6638, pi6639, pi6640, pi6641, pi6642, pi6643, pi6644, pi6645, pi6646, pi6647, pi6648, pi6649, pi6650, pi6651, pi6652, pi6653, pi6654, pi6655, pi6656, pi6657, pi6658, pi6659, pi6660, pi6661, pi6662, pi6663, pi6664, pi6665, pi6666, pi6667, pi6668, pi6669, pi6670, pi6671, pi6672, pi6673, pi6674, pi6675, pi6676, pi6677, pi6678, pi6679, pi6680, pi6681, pi6682, pi6683, pi6684, pi6685, pi6686, pi6687, pi6688, pi6689, pi6690, pi6691, pi6692, pi6693, pi6694, pi6695, pi6696, pi6697, pi6698, pi6699, pi6700, pi6701, pi6702, pi6703, pi6704, pi6705, pi6706, pi6707, pi6708, pi6709, pi6710, pi6711, pi6712, pi6713, pi6714, pi6715, pi6716, pi6717, pi6718, pi6719, pi6720, pi6721, pi6722, pi6723, pi6724, pi6725, pi6726, pi6727, pi6728, pi6729, pi6730, pi6731, pi6732, pi6733, pi6734, pi6735, pi6736, pi6737, pi6738, pi6739, pi6740, pi6741, pi6742, pi6743, pi6744, pi6745, pi6746, pi6747, pi6748, pi6749, pi6750, pi6751, pi6752, pi6753, pi6754, pi6755, pi6756, pi6757, pi6758, pi6759, pi6760, pi6761, pi6762, pi6763, pi6764, pi6765, pi6766, pi6767, pi6768, pi6769, pi6770, pi6771, pi6772, pi6773, pi6774, pi6775, pi6776, pi6777, pi6778, pi6779, pi6780, pi6781, pi6782, pi6783, pi6784, pi6785, pi6786, pi6787, pi6788, pi6789, pi6790, pi6791, pi6792, pi6793, pi6794, pi6795, pi6796, pi6797, pi6798, pi6799, pi6800, pi6801, pi6802, pi6803, pi6804, pi6805, pi6806, pi6807, pi6808, pi6809, pi6810, pi6811, pi6812, pi6813, pi6814, pi6815, pi6816, pi6817, pi6818, pi6819, pi6820, pi6821, pi6822, pi6823, pi6824, pi6825, pi6826, pi6827, pi6828, pi6829, pi6830, pi6831, pi6832, pi6833, pi6834, pi6835, pi6836, pi6837, pi6838, pi6839, pi6840, pi6841, pi6842, pi6843, pi6844, pi6845, pi6846, pi6847, pi6848, pi6849, pi6850, pi6851, pi6852, pi6853, pi6854, pi6855, pi6856, pi6857, pi6858, pi6859, pi6860, pi6861, pi6862, pi6863, pi6864, pi6865, pi6866, pi6867, pi6868, pi6869, pi6870, pi6871, pi6872, pi6873, pi6874, pi6875, pi6876, pi6877, pi6878, pi6879, pi6880, pi6881, pi6882, pi6883, pi6884, pi6885, pi6886, pi6887, pi6888, pi6889, pi6890, pi6891, pi6892, pi6893, pi6894, pi6895, pi6896, pi6897, pi6898, pi6899, pi6900, pi6901, pi6902, pi6903, pi6904, pi6905, pi6906, pi6907, pi6908, pi6909, pi6910, pi6911, pi6912, pi6913, pi6914, pi6915, pi6916, pi6917, pi6918, pi6919, pi6920, pi6921, pi6922, pi6923, pi6924, pi6925, pi6926, pi6927, pi6928, pi6929, pi6930, pi6931, pi6932, pi6933, pi6934, pi6935, pi6936, pi6937, pi6938, pi6939, pi6940, pi6941, pi6942, pi6943, pi6944, pi6945, pi6946, pi6947, pi6948, pi6949, pi6950, pi6951, pi6952, pi6953, pi6954, pi6955, pi6956, pi6957, pi6958, pi6959, pi6960, pi6961, pi6962, pi6963, pi6964, pi6965, pi6966, pi6967, pi6968, pi6969, pi6970, pi6971, pi6972, pi6973, pi6974, pi6975, pi6976, pi6977, pi6978, pi6979, pi6980, pi6981, pi6982, pi6983, pi6984, pi6985, pi6986, pi6987, pi6988, pi6989, pi6990, pi6991, pi6992, pi6993, pi6994, pi6995, pi6996, pi6997, pi6998, pi6999, pi7000, pi7001, pi7002, pi7003, pi7004, pi7005, pi7006, pi7007, pi7008, pi7009, pi7010, pi7011, pi7012, pi7013, pi7014, pi7015, pi7016, pi7017, pi7018, pi7019, pi7020, pi7021, pi7022, pi7023, pi7024, pi7025, pi7026, pi7027, pi7028, pi7029, pi7030, pi7031, pi7032, pi7033, pi7034, pi7035, pi7036, pi7037, pi7038, pi7039, pi7040, pi7041, pi7042, pi7043, pi7044, pi7045, pi7046, pi7047, pi7048, pi7049, pi7050, pi7051, pi7052, pi7053, pi7054, pi7055, pi7056, pi7057, pi7058, pi7059, pi7060, pi7061, pi7062, pi7063, pi7064, pi7065, pi7066, pi7067, pi7068, pi7069, pi7070, pi7071, pi7072, pi7073, pi7074, pi7075, pi7076, pi7077, pi7078, pi7079, pi7080, pi7081, pi7082, pi7083, pi7084, pi7085, pi7086, pi7087, pi7088, pi7089, pi7090, pi7091, pi7092, pi7093, pi7094, pi7095, pi7096, pi7097, pi7098, pi7099, pi7100, pi7101, pi7102, pi7103, pi7104, pi7105, pi7106, pi7107, pi7108, pi7109, pi7110, pi7111, pi7112, pi7113, pi7114, pi7115, pi7116, pi7117, pi7118, pi7119, pi7120, pi7121, pi7122, pi7123, pi7124, pi7125, pi7126, pi7127, pi7128, pi7129, pi7130, pi7131, pi7132, pi7133, pi7134, pi7135, pi7136, pi7137, pi7138, pi7139, pi7140, pi7141, pi7142, pi7143, pi7144, pi7145, pi7146, pi7147, pi7148, pi7149, pi7150, pi7151, pi7152, pi7153, pi7154, pi7155, pi7156, pi7157, pi7158, pi7159, pi7160, pi7161, pi7162, pi7163, pi7164, pi7165, pi7166, pi7167, pi7168, pi7169, pi7170, pi7171, pi7172, pi7173, pi7174, pi7175, pi7176, pi7177, pi7178, pi7179, pi7180, pi7181, pi7182, pi7183, pi7184, pi7185, pi7186, pi7187, pi7188, pi7189, pi7190, pi7191, pi7192, pi7193, pi7194, pi7195, pi7196, pi7197, pi7198, pi7199, pi7200, pi7201, pi7202, pi7203, pi7204, pi7205, pi7206, pi7207, pi7208, pi7209, pi7210, pi7211, pi7212, pi7213, pi7214, pi7215, pi7216, pi7217, pi7218, pi7219, pi7220, pi7221, pi7222, pi7223, pi7224, pi7225, pi7226, pi7227, pi7228, pi7229, pi7230, pi7231, pi7232, pi7233, pi7234, pi7235, pi7236, pi7237, pi7238, pi7239, pi7240, pi7241, pi7242, pi7243, pi7244, pi7245, pi7246, pi7247, pi7248, pi7249, pi7250, pi7251, pi7252, pi7253, pi7254, pi7255, pi7256, pi7257, pi7258, pi7259, pi7260, pi7261, pi7262, pi7263, pi7264, pi7265, pi7266, pi7267, pi7268, pi7269, pi7270, pi7271, pi7272, pi7273, pi7274, pi7275, pi7276, pi7277, pi7278, pi7279, pi7280, pi7281, pi7282, pi7283, pi7284, pi7285, pi7286, pi7287, pi7288, pi7289, pi7290, pi7291, pi7292, pi7293, pi7294, pi7295, pi7296, pi7297, pi7298, pi7299, pi7300, pi7301, pi7302, pi7303, pi7304, pi7305, pi7306, pi7307, pi7308, pi7309, pi7310, pi7311, pi7312, pi7313, pi7314, pi7315, pi7316, pi7317, pi7318, pi7319, pi7320, pi7321, pi7322, pi7323, pi7324, pi7325, pi7326, pi7327, pi7328, pi7329, pi7330, pi7331, pi7332, pi7333, pi7334, pi7335, pi7336, pi7337, pi7338, pi7339, pi7340, pi7341, pi7342, pi7343, pi7344, pi7345, pi7346, pi7347, pi7348, pi7349, pi7350, pi7351, pi7352, pi7353, pi7354, pi7355, pi7356, pi7357, pi7358, pi7359, pi7360, pi7361, pi7362, pi7363, pi7364, pi7365, pi7366, pi7367, pi7368, pi7369, pi7370, pi7371, pi7372, pi7373, pi7374, pi7375, pi7376, pi7377, pi7378, pi7379, pi7380, pi7381, pi7382, pi7383, pi7384, pi7385, pi7386, pi7387, pi7388, pi7389, pi7390, pi7391, pi7392, pi7393, pi7394, pi7395, pi7396, pi7397, pi7398, pi7399, pi7400, pi7401, pi7402, pi7403, pi7404, pi7405, pi7406, pi7407, pi7408, pi7409, pi7410, pi7411, pi7412, pi7413, pi7414, pi7415, pi7416, pi7417, pi7418, pi7419, pi7420, pi7421, pi7422, pi7423, pi7424, pi7425, pi7426, pi7427, pi7428, pi7429, pi7430, pi7431, pi7432, pi7433, pi7434, pi7435, pi7436, pi7437, pi7438, pi7439, pi7440, pi7441, pi7442, pi7443, pi7444, pi7445, pi7446, pi7447, pi7448, pi7449, pi7450, pi7451, pi7452, pi7453, pi7454, pi7455, pi7456, pi7457, pi7458, pi7459, pi7460, pi7461, pi7462, pi7463, pi7464, pi7465, pi7466, pi7467, pi7468, pi7469, pi7470, pi7471, pi7472, pi7473, pi7474, pi7475, pi7476, pi7477, pi7478, pi7479, pi7480, pi7481, pi7482, pi7483, pi7484, pi7485, pi7486, pi7487, pi7488, pi7489, pi7490, pi7491, pi7492, pi7493, pi7494, pi7495, pi7496, pi7497, pi7498, pi7499, pi7500, pi7501, pi7502, pi7503, pi7504, pi7505, pi7506, pi7507, pi7508, pi7509, pi7510, pi7511, pi7512, pi7513, pi7514, pi7515, pi7516, pi7517, pi7518, pi7519, pi7520, pi7521, pi7522, pi7523, pi7524, pi7525, pi7526, pi7527, pi7528, pi7529, pi7530, pi7531, pi7532, pi7533, pi7534, pi7535, pi7536, pi7537, pi7538, pi7539, pi7540, pi7541, pi7542, pi7543, pi7544, pi7545, pi7546, pi7547, pi7548, pi7549, pi7550, pi7551, pi7552, pi7553, pi7554, pi7555, pi7556, pi7557, pi7558, pi7559, pi7560, pi7561, pi7562, pi7563, pi7564, pi7565, pi7566, pi7567, pi7568, pi7569, pi7570, pi7571, pi7572, pi7573, pi7574, pi7575, pi7576, pi7577, pi7578, pi7579, pi7580, pi7581, pi7582, pi7583, pi7584, pi7585, pi7586, pi7587, pi7588, pi7589, pi7590, pi7591, pi7592, pi7593, pi7594, pi7595, pi7596, pi7597, pi7598, pi7599, pi7600, pi7601, pi7602, pi7603, pi7604, pi7605, pi7606, pi7607, pi7608, pi7609, pi7610, pi7611, pi7612, pi7613, pi7614, pi7615, pi7616, pi7617, pi7618, pi7619, pi7620, pi7621, pi7622, pi7623, pi7624, pi7625, pi7626, pi7627, pi7628, pi7629, pi7630, pi7631, pi7632, pi7633, pi7634, pi7635, pi7636, pi7637, pi7638, pi7639, pi7640, pi7641, pi7642, pi7643, pi7644, pi7645, pi7646, pi7647, pi7648, pi7649, pi7650, pi7651, pi7652, pi7653, pi7654, pi7655, pi7656, pi7657, pi7658, pi7659, pi7660, pi7661, pi7662, pi7663, pi7664, pi7665, pi7666, pi7667, pi7668, pi7669, pi7670, pi7671, pi7672, pi7673, pi7674, pi7675, pi7676, pi7677, pi7678, pi7679, pi7680, pi7681, pi7682, pi7683, pi7684, pi7685, pi7686, pi7687, pi7688, pi7689, pi7690, pi7691, pi7692, pi7693, pi7694, pi7695, pi7696, pi7697, pi7698, pi7699, pi7700, pi7701, pi7702, pi7703, pi7704, pi7705, pi7706, pi7707, pi7708, pi7709, pi7710, pi7711, pi7712, pi7713, pi7714, pi7715, pi7716, pi7717, pi7718, pi7719, pi7720, pi7721, pi7722, pi7723, pi7724, pi7725, pi7726, pi7727, pi7728, pi7729, pi7730, pi7731, pi7732, pi7733, pi7734, pi7735, pi7736, pi7737, pi7738, pi7739, pi7740, pi7741, pi7742, pi7743, pi7744, pi7745, pi7746, pi7747, pi7748, pi7749, pi7750, pi7751, pi7752, pi7753, pi7754, pi7755, pi7756, pi7757, pi7758, pi7759, pi7760, pi7761, pi7762, pi7763, pi7764, pi7765, pi7766, pi7767, pi7768, pi7769, pi7770, pi7771, pi7772, pi7773, pi7774, pi7775, pi7776, pi7777, pi7778, pi7779, pi7780, pi7781, pi7782, pi7783, pi7784, pi7785, pi7786, pi7787, pi7788, pi7789, pi7790, pi7791, pi7792, pi7793, pi7794, pi7795, pi7796, pi7797, pi7798, pi7799, pi7800, pi7801, pi7802, pi7803, pi7804, pi7805, pi7806, pi7807, pi7808, pi7809, pi7810, pi7811, pi7812, pi7813, pi7814, pi7815, pi7816, pi7817, pi7818, pi7819, pi7820, pi7821, pi7822, pi7823, pi7824, pi7825, pi7826, pi7827, pi7828, pi7829, pi7830, pi7831, pi7832, pi7833, pi7834, pi7835, pi7836, pi7837, pi7838, pi7839, pi7840, pi7841, pi7842, pi7843, pi7844, pi7845, pi7846, pi7847, pi7848, pi7849, pi7850, pi7851, pi7852, pi7853, pi7854, pi7855, pi7856, pi7857, pi7858, pi7859, pi7860, pi7861, pi7862, pi7863, pi7864, pi7865, pi7866, pi7867, pi7868, pi7869, pi7870, pi7871, pi7872, pi7873, pi7874, pi7875, pi7876, pi7877, pi7878, pi7879, pi7880, pi7881, pi7882, pi7883, pi7884, pi7885, pi7886, pi7887, pi7888, pi7889, pi7890, pi7891, pi7892, pi7893, pi7894, pi7895, pi7896, pi7897, pi7898, pi7899, pi7900, pi7901, pi7902, pi7903, pi7904, pi7905, pi7906, pi7907, pi7908, pi7909, pi7910, pi7911, pi7912, pi7913, pi7914, pi7915, pi7916, pi7917, pi7918, pi7919, pi7920, pi7921, pi7922, pi7923, pi7924, pi7925, pi7926, pi7927, pi7928, pi7929, pi7930, pi7931, pi7932, pi7933, pi7934, pi7935, pi7936, pi7937, pi7938, pi7939, pi7940, pi7941, pi7942, pi7943, pi7944, pi7945, pi7946, pi7947, pi7948, pi7949, pi7950, pi7951, pi7952, pi7953, pi7954, pi7955, pi7956, pi7957, pi7958, pi7959, pi7960, pi7961, pi7962, pi7963, pi7964, pi7965, pi7966, pi7967, pi7968, pi7969, pi7970, pi7971, pi7972, pi7973, pi7974, pi7975, pi7976, pi7977, pi7978, pi7979, pi7980, pi7981, pi7982, pi7983, pi7984, pi7985, pi7986, pi7987, pi7988, pi7989, pi7990, pi7991, pi7992, pi7993, pi7994, pi7995, pi7996, pi7997, pi7998, pi7999, pi8000, pi8001, pi8002, pi8003, pi8004, pi8005, pi8006, pi8007, pi8008, pi8009, pi8010, pi8011, pi8012, pi8013, pi8014, pi8015, pi8016, pi8017, pi8018, pi8019, pi8020, pi8021, pi8022, pi8023, pi8024, pi8025, pi8026, pi8027, pi8028, pi8029, pi8030, pi8031, pi8032, pi8033, pi8034, pi8035, pi8036, pi8037, pi8038, pi8039, pi8040, pi8041, pi8042, pi8043, pi8044, pi8045, pi8046, pi8047, pi8048, pi8049, pi8050, pi8051, pi8052, pi8053, pi8054, pi8055, pi8056, pi8057, pi8058, pi8059, pi8060, pi8061, pi8062, pi8063, pi8064, pi8065, pi8066, pi8067, pi8068, pi8069, pi8070, pi8071, pi8072, pi8073, pi8074, pi8075, pi8076, pi8077, pi8078, pi8079, pi8080, pi8081, pi8082, pi8083, pi8084, pi8085, pi8086, pi8087, pi8088, pi8089, pi8090, pi8091, pi8092, pi8093, pi8094, pi8095, pi8096, pi8097, pi8098, pi8099, pi8100, pi8101, pi8102, pi8103, pi8104, pi8105, pi8106, pi8107, pi8108, pi8109, pi8110, pi8111, pi8112, pi8113, pi8114, pi8115, pi8116, pi8117, pi8118, pi8119, pi8120, pi8121, pi8122, pi8123, pi8124, pi8125, pi8126, pi8127, pi8128, pi8129, pi8130, pi8131, pi8132, pi8133, pi8134, pi8135, pi8136, pi8137, pi8138, pi8139, pi8140, pi8141, pi8142, pi8143, pi8144, pi8145, pi8146, pi8147, pi8148, pi8149, pi8150, pi8151, pi8152, pi8153, pi8154, pi8155, pi8156, pi8157, pi8158, pi8159, pi8160, pi8161, pi8162, pi8163, pi8164, pi8165, pi8166, pi8167, pi8168, pi8169, pi8170, pi8171, pi8172, pi8173, pi8174, pi8175, pi8176, pi8177, pi8178, pi8179, pi8180, pi8181, pi8182, pi8183, pi8184, pi8185, pi8186, pi8187, pi8188, pi8189, pi8190, pi8191, pi8192, pi8193, pi8194, pi8195, pi8196, pi8197, pi8198, pi8199, pi8200, pi8201, pi8202, pi8203, pi8204, pi8205, pi8206, pi8207, pi8208, pi8209, pi8210, pi8211, pi8212, pi8213, pi8214, pi8215, pi8216, pi8217, pi8218, pi8219, pi8220, pi8221, pi8222, pi8223, pi8224, pi8225, pi8226, pi8227, pi8228, pi8229, pi8230, pi8231, pi8232, pi8233, pi8234, pi8235, pi8236, pi8237, pi8238, pi8239, pi8240, pi8241, pi8242, pi8243, pi8244, pi8245, pi8246, pi8247, pi8248, pi8249, pi8250, pi8251, pi8252, pi8253, pi8254, pi8255, pi8256, pi8257, pi8258, pi8259, pi8260, pi8261, pi8262, pi8263, pi8264, pi8265, pi8266, pi8267, pi8268, pi8269, pi8270, pi8271, pi8272, pi8273, pi8274, pi8275, pi8276, pi8277, pi8278, pi8279, pi8280, pi8281, pi8282, pi8283, pi8284, pi8285, pi8286, pi8287, pi8288, pi8289, pi8290, pi8291, pi8292, pi8293, pi8294, pi8295, pi8296, pi8297, pi8298, pi8299, pi8300, pi8301, pi8302, pi8303, pi8304, pi8305, pi8306, pi8307, pi8308, pi8309, pi8310, pi8311, pi8312, pi8313, pi8314, pi8315, pi8316, pi8317, pi8318, pi8319, pi8320, pi8321, pi8322, pi8323, pi8324, pi8325, pi8326, pi8327, pi8328, pi8329, pi8330, pi8331, pi8332, pi8333, pi8334, pi8335, pi8336, pi8337, pi8338, pi8339, pi8340, pi8341, pi8342, pi8343, pi8344, pi8345, pi8346, pi8347, pi8348, pi8349, pi8350, pi8351, pi8352, pi8353, pi8354, pi8355, pi8356, pi8357, pi8358, pi8359, pi8360, pi8361, pi8362, pi8363, pi8364, pi8365, pi8366, pi8367, pi8368, pi8369, pi8370, pi8371, pi8372, pi8373, pi8374, pi8375, pi8376, pi8377, pi8378, pi8379, pi8380, pi8381, pi8382, pi8383, pi8384, pi8385, pi8386, pi8387, pi8388, pi8389, pi8390, pi8391, pi8392, pi8393, pi8394, pi8395, pi8396, pi8397, pi8398, pi8399, pi8400, pi8401, pi8402, pi8403, pi8404, pi8405, pi8406, pi8407, pi8408, pi8409, pi8410, pi8411, pi8412, pi8413, pi8414, pi8415, pi8416, pi8417, pi8418, pi8419, pi8420, pi8421, pi8422, pi8423, pi8424, pi8425, pi8426, pi8427, pi8428, pi8429, pi8430, pi8431, pi8432, pi8433, pi8434, pi8435, pi8436, pi8437, pi8438, pi8439, pi8440, pi8441, pi8442, pi8443, pi8444, pi8445, pi8446, pi8447, pi8448, pi8449, pi8450, pi8451, pi8452, pi8453, pi8454, pi8455, pi8456, pi8457, pi8458, pi8459, pi8460, pi8461, pi8462, pi8463, pi8464, pi8465, pi8466, pi8467, pi8468, pi8469, pi8470, pi8471, pi8472, pi8473, pi8474, pi8475, pi8476, pi8477, pi8478, pi8479, pi8480, pi8481, pi8482, pi8483, pi8484, pi8485, pi8486, pi8487, pi8488, pi8489, pi8490, pi8491, pi8492, pi8493, pi8494, pi8495, pi8496, pi8497, pi8498, pi8499, pi8500, pi8501, pi8502, pi8503, pi8504, pi8505, pi8506, pi8507, pi8508, pi8509, pi8510, pi8511, pi8512, pi8513, pi8514, pi8515, pi8516, pi8517, pi8518, pi8519, pi8520, pi8521, pi8522, pi8523, pi8524, pi8525, pi8526, pi8527, pi8528, pi8529, pi8530, pi8531, pi8532, pi8533, pi8534, pi8535, pi8536, pi8537, pi8538, pi8539, pi8540, pi8541, pi8542, pi8543, pi8544, pi8545, pi8546, pi8547, pi8548, pi8549, pi8550, pi8551, pi8552, pi8553, pi8554, pi8555, pi8556, pi8557, pi8558, pi8559, pi8560, pi8561, pi8562, pi8563, pi8564, pi8565, pi8566, pi8567, pi8568, pi8569, pi8570, pi8571, pi8572, pi8573, pi8574, pi8575, pi8576, pi8577, pi8578, pi8579, pi8580, pi8581, pi8582, pi8583, pi8584, pi8585, pi8586, pi8587, pi8588, pi8589, pi8590, pi8591, pi8592, pi8593, pi8594, pi8595, pi8596, pi8597, pi8598, pi8599, pi8600, pi8601, pi8602, pi8603, pi8604, pi8605, pi8606, pi8607, pi8608, pi8609, pi8610, pi8611, pi8612, pi8613, pi8614, pi8615, pi8616, pi8617, pi8618, pi8619, pi8620, pi8621, pi8622, pi8623, pi8624, pi8625, pi8626, pi8627, pi8628, pi8629, pi8630, pi8631, pi8632, pi8633, pi8634, pi8635, pi8636, pi8637, pi8638, pi8639, pi8640, pi8641, pi8642, pi8643, pi8644, pi8645, pi8646, pi8647, pi8648, pi8649, pi8650, pi8651, pi8652, pi8653, pi8654, pi8655, pi8656, pi8657, pi8658, pi8659, pi8660, pi8661, pi8662, pi8663, pi8664, pi8665, pi8666, pi8667, pi8668, pi8669, pi8670, pi8671, pi8672, pi8673, pi8674, pi8675, pi8676, pi8677, pi8678, pi8679, pi8680, pi8681, pi8682, pi8683, pi8684, pi8685, pi8686, pi8687, pi8688, pi8689, pi8690, pi8691, pi8692, pi8693, pi8694, pi8695, pi8696, pi8697, pi8698, pi8699, pi8700, pi8701, pi8702, pi8703, pi8704, pi8705, pi8706, pi8707, pi8708, pi8709, pi8710, pi8711, pi8712, pi8713, pi8714, pi8715, pi8716, pi8717, pi8718, pi8719, pi8720, pi8721, pi8722, pi8723, pi8724, pi8725, pi8726, pi8727, pi8728, pi8729, pi8730, pi8731, pi8732, pi8733, pi8734, pi8735, pi8736, pi8737, pi8738, pi8739, pi8740, pi8741, pi8742, pi8743, pi8744, pi8745, pi8746, pi8747, pi8748, pi8749, pi8750, pi8751, pi8752, pi8753, pi8754, pi8755, pi8756, pi8757, pi8758, pi8759, pi8760, pi8761, pi8762, pi8763, pi8764, pi8765, pi8766, pi8767, pi8768, pi8769, pi8770, pi8771, pi8772, pi8773, pi8774, pi8775, pi8776, pi8777, pi8778, pi8779, pi8780, pi8781, pi8782, pi8783, pi8784, pi8785, pi8786, pi8787, pi8788, pi8789, pi8790, pi8791, pi8792, pi8793, pi8794, pi8795, pi8796, pi8797, pi8798, pi8799, pi8800, pi8801, pi8802, pi8803, pi8804, pi8805, pi8806, pi8807, pi8808, pi8809, pi8810, pi8811, pi8812, pi8813, pi8814, pi8815, pi8816, pi8817, pi8818, pi8819, pi8820, pi8821, pi8822, pi8823, pi8824, pi8825, pi8826, pi8827, pi8828, pi8829, pi8830, pi8831, pi8832, pi8833, pi8834, pi8835, pi8836, pi8837, pi8838, pi8839, pi8840, pi8841, pi8842, pi8843, pi8844, pi8845, pi8846, pi8847, pi8848, pi8849, pi8850, pi8851, pi8852, pi8853, pi8854, pi8855, pi8856, pi8857, pi8858, pi8859, pi8860, pi8861, pi8862, pi8863, pi8864, pi8865, pi8866, pi8867, pi8868, pi8869, pi8870, pi8871, pi8872, pi8873, pi8874, pi8875, pi8876, pi8877, pi8878, pi8879, pi8880, pi8881, pi8882, pi8883, pi8884, pi8885, pi8886, pi8887, pi8888, pi8889, pi8890, pi8891, pi8892, pi8893, pi8894, pi8895, pi8896, pi8897, pi8898, pi8899, pi8900, pi8901, pi8902, pi8903, pi8904, pi8905, pi8906, pi8907, pi8908, pi8909, pi8910, pi8911, pi8912, pi8913, pi8914, pi8915, pi8916, pi8917, pi8918, pi8919, pi8920, pi8921, pi8922, pi8923, pi8924, pi8925, pi8926, pi8927, pi8928, pi8929, pi8930, pi8931, pi8932, pi8933, pi8934, pi8935, pi8936, pi8937, pi8938, pi8939, pi8940, pi8941, pi8942, pi8943, pi8944, pi8945, pi8946, pi8947, pi8948, pi8949, pi8950, pi8951, pi8952, pi8953, pi8954, pi8955, pi8956, pi8957, pi8958, pi8959, pi8960, pi8961, pi8962, pi8963, pi8964, pi8965, pi8966, pi8967, pi8968, pi8969, pi8970, pi8971, pi8972, pi8973, pi8974, pi8975, pi8976, pi8977, pi8978, pi8979, pi8980, pi8981, pi8982, pi8983, pi8984, pi8985, pi8986, pi8987, pi8988, pi8989, pi8990, pi8991, pi8992, pi8993, pi8994, pi8995, pi8996, pi8997, pi8998, pi8999, pi9000, pi9001, pi9002, pi9003, pi9004, pi9005, pi9006, pi9007, pi9008, pi9009, pi9010, pi9011, pi9012, pi9013, pi9014, pi9015, pi9016, pi9017, pi9018, pi9019, pi9020, pi9021, pi9022, pi9023, pi9024, pi9025, pi9026, pi9027, pi9028, pi9029, pi9030, pi9031, pi9032, pi9033, pi9034, pi9035, pi9036, pi9037, pi9038, pi9039, pi9040, pi9041;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535, po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544, po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553, po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562, po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571, po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580, po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589, po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598, po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607, po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616, po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625, po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634, po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643, po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652, po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661, po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670, po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679, po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688, po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697, po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706, po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715, po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724, po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733, po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742, po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751, po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760, po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769, po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778, po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787, po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796, po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805, po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814, po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823, po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832, po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841, po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850, po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859, po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868, po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877, po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886, po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895, po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904, po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913, po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922, po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931, po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940, po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949, po3950, po3951, po3952, po3953, po3954, po3955, po3956, po3957, po3958, po3959, po3960, po3961, po3962, po3963, po3964, po3965, po3966, po3967, po3968, po3969, po3970, po3971, po3972, po3973, po3974, po3975, po3976, po3977, po3978, po3979, po3980, po3981, po3982, po3983, po3984, po3985, po3986, po3987, po3988, po3989, po3990, po3991, po3992, po3993, po3994, po3995, po3996, po3997, po3998, po3999, po4000, po4001, po4002, po4003, po4004, po4005, po4006, po4007, po4008, po4009, po4010, po4011, po4012, po4013, po4014, po4015, po4016, po4017, po4018, po4019, po4020, po4021, po4022, po4023, po4024, po4025, po4026, po4027, po4028, po4029, po4030, po4031, po4032, po4033, po4034, po4035, po4036, po4037, po4038, po4039, po4040, po4041, po4042, po4043, po4044, po4045, po4046, po4047, po4048, po4049, po4050, po4051, po4052, po4053, po4054, po4055, po4056, po4057, po4058, po4059, po4060, po4061, po4062, po4063, po4064, po4065, po4066, po4067, po4068, po4069, po4070, po4071, po4072, po4073, po4074, po4075, po4076, po4077, po4078, po4079, po4080, po4081, po4082, po4083, po4084, po4085, po4086, po4087, po4088, po4089, po4090, po4091, po4092, po4093, po4094, po4095, po4096, po4097, po4098, po4099, po4100, po4101, po4102, po4103, po4104, po4105, po4106, po4107, po4108, po4109, po4110, po4111, po4112, po4113, po4114, po4115, po4116, po4117, po4118, po4119, po4120, po4121, po4122, po4123, po4124, po4125, po4126, po4127, po4128, po4129, po4130, po4131, po4132, po4133, po4134, po4135, po4136, po4137, po4138, po4139, po4140, po4141, po4142, po4143, po4144, po4145, po4146, po4147, po4148, po4149, po4150, po4151, po4152, po4153, po4154, po4155, po4156, po4157, po4158, po4159, po4160, po4161, po4162, po4163, po4164, po4165, po4166, po4167, po4168, po4169, po4170, po4171, po4172, po4173, po4174, po4175, po4176, po4177, po4178, po4179, po4180, po4181, po4182, po4183, po4184, po4185, po4186, po4187, po4188, po4189, po4190, po4191, po4192, po4193, po4194, po4195, po4196, po4197, po4198, po4199, po4200, po4201, po4202, po4203, po4204, po4205, po4206, po4207, po4208, po4209, po4210, po4211, po4212, po4213, po4214, po4215, po4216, po4217, po4218, po4219, po4220, po4221, po4222, po4223, po4224, po4225, po4226, po4227, po4228, po4229, po4230, po4231, po4232, po4233, po4234, po4235, po4236, po4237, po4238, po4239, po4240, po4241, po4242, po4243, po4244, po4245, po4246, po4247, po4248, po4249, po4250, po4251, po4252, po4253, po4254, po4255, po4256, po4257, po4258, po4259, po4260, po4261, po4262, po4263, po4264, po4265, po4266, po4267, po4268, po4269, po4270, po4271, po4272, po4273, po4274, po4275, po4276, po4277, po4278, po4279, po4280, po4281, po4282, po4283, po4284, po4285, po4286, po4287, po4288, po4289, po4290, po4291, po4292, po4293, po4294, po4295, po4296, po4297, po4298, po4299, po4300, po4301, po4302, po4303, po4304, po4305, po4306, po4307, po4308, po4309, po4310, po4311, po4312, po4313, po4314, po4315, po4316, po4317, po4318, po4319, po4320, po4321, po4322, po4323, po4324, po4325, po4326, po4327, po4328, po4329, po4330, po4331, po4332, po4333, po4334, po4335, po4336, po4337, po4338, po4339, po4340, po4341, po4342, po4343, po4344, po4345, po4346, po4347, po4348, po4349, po4350, po4351, po4352, po4353, po4354, po4355, po4356, po4357, po4358, po4359, po4360, po4361, po4362, po4363, po4364, po4365, po4366, po4367, po4368, po4369, po4370, po4371, po4372, po4373, po4374, po4375, po4376, po4377, po4378, po4379, po4380, po4381, po4382, po4383, po4384, po4385, po4386, po4387, po4388, po4389, po4390, po4391, po4392, po4393, po4394, po4395, po4396, po4397, po4398, po4399, po4400, po4401, po4402, po4403, po4404, po4405, po4406, po4407, po4408, po4409, po4410, po4411, po4412, po4413, po4414, po4415, po4416, po4417, po4418, po4419, po4420, po4421, po4422, po4423, po4424, po4425, po4426, po4427, po4428, po4429, po4430, po4431, po4432, po4433, po4434, po4435, po4436, po4437, po4438, po4439, po4440, po4441, po4442, po4443, po4444, po4445, po4446, po4447, po4448, po4449, po4450, po4451, po4452, po4453, po4454, po4455, po4456, po4457, po4458, po4459, po4460, po4461, po4462, po4463, po4464, po4465, po4466, po4467, po4468, po4469, po4470, po4471, po4472, po4473, po4474, po4475, po4476, po4477, po4478, po4479, po4480, po4481, po4482, po4483, po4484, po4485, po4486, po4487, po4488, po4489, po4490, po4491, po4492, po4493, po4494, po4495, po4496, po4497, po4498, po4499, po4500, po4501, po4502, po4503, po4504, po4505, po4506, po4507, po4508, po4509, po4510, po4511, po4512, po4513, po4514, po4515, po4516, po4517, po4518, po4519, po4520, po4521, po4522, po4523, po4524, po4525, po4526, po4527, po4528, po4529, po4530, po4531, po4532, po4533, po4534, po4535, po4536, po4537, po4538, po4539, po4540, po4541, po4542, po4543, po4544, po4545, po4546, po4547, po4548, po4549, po4550, po4551, po4552, po4553, po4554, po4555, po4556, po4557, po4558, po4559, po4560, po4561, po4562, po4563, po4564, po4565, po4566, po4567, po4568, po4569, po4570, po4571, po4572, po4573, po4574, po4575, po4576, po4577, po4578, po4579, po4580, po4581, po4582, po4583, po4584, po4585, po4586, po4587, po4588, po4589, po4590, po4591, po4592, po4593, po4594, po4595, po4596, po4597, po4598, po4599, po4600, po4601, po4602, po4603, po4604, po4605, po4606, po4607, po4608, po4609, po4610, po4611, po4612, po4613, po4614, po4615, po4616, po4617, po4618, po4619, po4620, po4621, po4622, po4623, po4624, po4625, po4626, po4627, po4628, po4629, po4630, po4631, po4632, po4633, po4634, po4635, po4636, po4637, po4638, po4639, po4640, po4641, po4642, po4643, po4644, po4645, po4646, po4647, po4648, po4649, po4650, po4651, po4652, po4653, po4654, po4655, po4656, po4657, po4658, po4659, po4660, po4661, po4662, po4663, po4664, po4665, po4666, po4667, po4668, po4669, po4670, po4671, po4672, po4673, po4674, po4675, po4676, po4677, po4678, po4679, po4680, po4681, po4682, po4683, po4684, po4685, po4686, po4687, po4688, po4689, po4690, po4691, po4692, po4693, po4694, po4695, po4696, po4697, po4698, po4699, po4700, po4701, po4702, po4703, po4704, po4705, po4706, po4707, po4708, po4709, po4710, po4711, po4712, po4713, po4714, po4715, po4716, po4717, po4718, po4719, po4720, po4721, po4722, po4723, po4724, po4725, po4726, po4727, po4728, po4729, po4730, po4731, po4732, po4733, po4734, po4735, po4736, po4737, po4738, po4739, po4740, po4741, po4742, po4743, po4744, po4745, po4746, po4747, po4748, po4749, po4750, po4751, po4752, po4753, po4754, po4755, po4756, po4757, po4758, po4759, po4760, po4761, po4762, po4763, po4764, po4765, po4766, po4767, po4768, po4769, po4770, po4771, po4772, po4773, po4774, po4775, po4776, po4777, po4778, po4779, po4780, po4781, po4782, po4783, po4784, po4785, po4786, po4787, po4788, po4789, po4790, po4791, po4792, po4793, po4794, po4795, po4796, po4797, po4798, po4799, po4800, po4801, po4802, po4803, po4804, po4805, po4806, po4807, po4808, po4809, po4810, po4811, po4812, po4813, po4814, po4815, po4816, po4817, po4818, po4819, po4820, po4821, po4822, po4823, po4824, po4825, po4826, po4827, po4828, po4829, po4830, po4831, po4832, po4833, po4834, po4835, po4836, po4837, po4838, po4839, po4840, po4841, po4842, po4843, po4844, po4845, po4846, po4847, po4848, po4849, po4850, po4851, po4852, po4853, po4854, po4855, po4856, po4857, po4858, po4859, po4860, po4861, po4862, po4863, po4864, po4865, po4866, po4867, po4868, po4869, po4870, po4871, po4872, po4873, po4874, po4875, po4876, po4877, po4878, po4879, po4880, po4881, po4882, po4883, po4884, po4885, po4886, po4887, po4888, po4889, po4890, po4891, po4892, po4893, po4894, po4895, po4896, po4897, po4898, po4899, po4900, po4901, po4902, po4903, po4904, po4905, po4906, po4907, po4908, po4909, po4910, po4911, po4912, po4913, po4914, po4915, po4916, po4917, po4918, po4919, po4920, po4921, po4922, po4923, po4924, po4925, po4926, po4927, po4928, po4929, po4930, po4931, po4932, po4933, po4934, po4935, po4936, po4937, po4938, po4939, po4940, po4941, po4942, po4943, po4944, po4945, po4946, po4947, po4948, po4949, po4950, po4951, po4952, po4953, po4954, po4955, po4956, po4957, po4958, po4959, po4960, po4961, po4962, po4963, po4964, po4965, po4966, po4967, po4968, po4969, po4970, po4971, po4972, po4973, po4974, po4975, po4976, po4977, po4978, po4979, po4980, po4981, po4982, po4983, po4984, po4985, po4986, po4987, po4988, po4989, po4990, po4991, po4992, po4993, po4994, po4995, po4996, po4997, po4998, po4999, po5000, po5001, po5002, po5003, po5004, po5005, po5006, po5007, po5008, po5009, po5010, po5011, po5012, po5013, po5014, po5015, po5016, po5017, po5018, po5019, po5020, po5021, po5022, po5023, po5024, po5025, po5026, po5027, po5028, po5029, po5030, po5031, po5032, po5033, po5034, po5035, po5036, po5037, po5038, po5039, po5040, po5041, po5042, po5043, po5044, po5045, po5046, po5047, po5048, po5049, po5050, po5051, po5052, po5053, po5054, po5055, po5056, po5057, po5058, po5059, po5060, po5061, po5062, po5063, po5064, po5065, po5066, po5067, po5068, po5069, po5070, po5071, po5072, po5073, po5074, po5075, po5076, po5077, po5078, po5079, po5080, po5081, po5082, po5083, po5084, po5085, po5086, po5087, po5088, po5089, po5090, po5091, po5092, po5093, po5094, po5095, po5096, po5097, po5098, po5099, po5100, po5101, po5102, po5103, po5104, po5105, po5106, po5107, po5108, po5109, po5110, po5111, po5112, po5113, po5114, po5115, po5116, po5117, po5118, po5119, po5120, po5121, po5122, po5123, po5124, po5125, po5126, po5127, po5128, po5129, po5130, po5131, po5132, po5133, po5134, po5135, po5136, po5137, po5138, po5139, po5140, po5141, po5142, po5143, po5144, po5145, po5146, po5147, po5148, po5149, po5150, po5151, po5152, po5153, po5154, po5155, po5156, po5157, po5158, po5159, po5160, po5161, po5162, po5163, po5164, po5165, po5166, po5167, po5168, po5169, po5170, po5171, po5172, po5173, po5174, po5175, po5176, po5177, po5178, po5179, po5180, po5181, po5182, po5183, po5184, po5185, po5186, po5187, po5188, po5189, po5190, po5191, po5192, po5193, po5194, po5195, po5196, po5197, po5198, po5199, po5200, po5201, po5202, po5203, po5204, po5205, po5206, po5207, po5208, po5209, po5210, po5211, po5212, po5213, po5214, po5215, po5216, po5217, po5218, po5219, po5220, po5221, po5222, po5223, po5224, po5225, po5226, po5227, po5228, po5229, po5230, po5231, po5232, po5233, po5234, po5235, po5236, po5237, po5238, po5239, po5240, po5241, po5242, po5243, po5244, po5245, po5246, po5247, po5248, po5249, po5250, po5251, po5252, po5253, po5254, po5255, po5256, po5257, po5258, po5259, po5260, po5261, po5262, po5263, po5264, po5265, po5266, po5267, po5268, po5269, po5270, po5271, po5272, po5273, po5274, po5275, po5276, po5277, po5278, po5279, po5280, po5281, po5282, po5283, po5284, po5285, po5286, po5287, po5288, po5289, po5290, po5291, po5292, po5293, po5294, po5295, po5296, po5297, po5298, po5299, po5300, po5301, po5302, po5303, po5304, po5305, po5306, po5307, po5308, po5309, po5310, po5311, po5312, po5313, po5314, po5315, po5316, po5317, po5318, po5319, po5320, po5321, po5322, po5323, po5324, po5325, po5326, po5327, po5328, po5329, po5330, po5331, po5332, po5333, po5334, po5335, po5336, po5337, po5338, po5339, po5340, po5341, po5342, po5343, po5344, po5345, po5346, po5347, po5348, po5349, po5350, po5351, po5352, po5353, po5354, po5355, po5356, po5357, po5358, po5359, po5360, po5361, po5362, po5363, po5364, po5365, po5366, po5367, po5368, po5369, po5370, po5371, po5372, po5373, po5374, po5375, po5376, po5377, po5378, po5379, po5380, po5381, po5382, po5383, po5384, po5385, po5386, po5387, po5388, po5389, po5390, po5391, po5392, po5393, po5394, po5395, po5396, po5397, po5398, po5399, po5400, po5401, po5402, po5403, po5404, po5405, po5406, po5407, po5408, po5409, po5410, po5411, po5412, po5413, po5414, po5415, po5416, po5417, po5418, po5419, po5420, po5421, po5422, po5423, po5424, po5425, po5426, po5427, po5428, po5429, po5430, po5431, po5432, po5433, po5434, po5435, po5436, po5437, po5438, po5439, po5440, po5441, po5442, po5443, po5444, po5445, po5446, po5447, po5448, po5449, po5450, po5451, po5452, po5453, po5454, po5455, po5456, po5457, po5458, po5459, po5460, po5461, po5462, po5463, po5464, po5465, po5466, po5467, po5468, po5469, po5470, po5471, po5472, po5473, po5474, po5475, po5476, po5477, po5478, po5479, po5480, po5481, po5482, po5483, po5484, po5485, po5486, po5487, po5488, po5489, po5490, po5491, po5492, po5493, po5494, po5495, po5496, po5497, po5498, po5499, po5500, po5501, po5502, po5503, po5504, po5505, po5506, po5507, po5508, po5509, po5510, po5511, po5512, po5513, po5514, po5515, po5516, po5517, po5518, po5519, po5520, po5521, po5522, po5523, po5524, po5525, po5526, po5527, po5528, po5529, po5530, po5531, po5532, po5533, po5534, po5535, po5536, po5537, po5538, po5539, po5540, po5541, po5542, po5543, po5544, po5545, po5546, po5547, po5548, po5549, po5550, po5551, po5552, po5553, po5554, po5555, po5556, po5557, po5558, po5559, po5560, po5561, po5562, po5563, po5564, po5565, po5566, po5567, po5568, po5569, po5570, po5571, po5572, po5573, po5574, po5575, po5576, po5577, po5578, po5579, po5580, po5581, po5582, po5583, po5584, po5585, po5586, po5587, po5588, po5589, po5590, po5591, po5592, po5593, po5594, po5595, po5596, po5597, po5598, po5599, po5600, po5601, po5602, po5603, po5604, po5605, po5606, po5607, po5608, po5609, po5610, po5611, po5612, po5613, po5614, po5615, po5616, po5617, po5618, po5619, po5620, po5621, po5622, po5623, po5624, po5625, po5626, po5627, po5628, po5629, po5630, po5631, po5632, po5633, po5634, po5635, po5636, po5637, po5638, po5639, po5640, po5641, po5642, po5643, po5644, po5645, po5646, po5647, po5648, po5649, po5650, po5651, po5652, po5653, po5654, po5655, po5656, po5657, po5658, po5659, po5660, po5661, po5662, po5663, po5664, po5665, po5666, po5667, po5668, po5669, po5670, po5671, po5672, po5673, po5674, po5675, po5676, po5677, po5678, po5679, po5680, po5681, po5682, po5683, po5684, po5685, po5686, po5687, po5688, po5689, po5690, po5691, po5692, po5693, po5694, po5695, po5696, po5697, po5698, po5699, po5700, po5701, po5702, po5703, po5704, po5705, po5706, po5707, po5708, po5709, po5710, po5711, po5712, po5713, po5714, po5715, po5716, po5717, po5718, po5719, po5720, po5721, po5722, po5723, po5724, po5725, po5726, po5727, po5728, po5729, po5730, po5731, po5732, po5733, po5734, po5735, po5736, po5737, po5738, po5739, po5740, po5741, po5742, po5743, po5744, po5745, po5746, po5747, po5748, po5749, po5750, po5751, po5752, po5753, po5754, po5755, po5756, po5757, po5758, po5759, po5760, po5761, po5762, po5763, po5764, po5765, po5766, po5767, po5768, po5769, po5770, po5771, po5772, po5773, po5774, po5775, po5776, po5777, po5778, po5779, po5780, po5781, po5782, po5783, po5784, po5785, po5786, po5787, po5788, po5789, po5790, po5791, po5792, po5793, po5794, po5795, po5796, po5797, po5798, po5799, po5800, po5801, po5802, po5803, po5804, po5805, po5806, po5807, po5808, po5809, po5810, po5811, po5812, po5813, po5814, po5815, po5816, po5817, po5818, po5819, po5820, po5821, po5822, po5823, po5824, po5825, po5826, po5827, po5828, po5829, po5830, po5831, po5832, po5833, po5834, po5835, po5836, po5837, po5838, po5839, po5840, po5841, po5842, po5843, po5844, po5845, po5846, po5847, po5848, po5849, po5850, po5851, po5852, po5853, po5854, po5855, po5856, po5857, po5858, po5859, po5860, po5861, po5862, po5863, po5864, po5865, po5866, po5867, po5868, po5869, po5870, po5871, po5872, po5873, po5874, po5875, po5876, po5877, po5878, po5879, po5880, po5881, po5882, po5883, po5884, po5885, po5886, po5887, po5888, po5889, po5890, po5891, po5892, po5893, po5894, po5895, po5896, po5897, po5898, po5899, po5900, po5901, po5902, po5903, po5904, po5905, po5906, po5907, po5908, po5909, po5910, po5911, po5912, po5913, po5914, po5915, po5916, po5917, po5918, po5919, po5920, po5921, po5922, po5923, po5924, po5925, po5926, po5927, po5928, po5929, po5930, po5931, po5932, po5933, po5934, po5935, po5936, po5937, po5938, po5939, po5940, po5941, po5942, po5943, po5944, po5945, po5946, po5947, po5948, po5949, po5950, po5951, po5952, po5953, po5954, po5955, po5956, po5957, po5958, po5959, po5960, po5961, po5962, po5963, po5964, po5965, po5966, po5967, po5968, po5969, po5970, po5971, po5972, po5973, po5974, po5975, po5976, po5977, po5978, po5979, po5980, po5981, po5982, po5983, po5984, po5985, po5986, po5987, po5988, po5989, po5990, po5991, po5992, po5993, po5994, po5995, po5996, po5997, po5998, po5999, po6000, po6001, po6002, po6003, po6004, po6005, po6006, po6007, po6008, po6009, po6010, po6011, po6012, po6013, po6014, po6015, po6016, po6017, po6018, po6019, po6020, po6021, po6022, po6023, po6024, po6025, po6026, po6027, po6028, po6029, po6030, po6031, po6032, po6033, po6034, po6035, po6036, po6037, po6038, po6039, po6040, po6041, po6042, po6043, po6044, po6045, po6046, po6047, po6048, po6049, po6050, po6051, po6052, po6053, po6054, po6055, po6056, po6057, po6058, po6059, po6060, po6061, po6062, po6063, po6064, po6065, po6066, po6067, po6068, po6069, po6070, po6071, po6072, po6073, po6074, po6075, po6076, po6077, po6078, po6079, po6080, po6081, po6082, po6083, po6084, po6085, po6086, po6087, po6088, po6089, po6090, po6091, po6092, po6093, po6094, po6095, po6096, po6097, po6098, po6099, po6100, po6101, po6102, po6103, po6104, po6105, po6106, po6107, po6108, po6109, po6110, po6111, po6112, po6113, po6114, po6115, po6116, po6117, po6118, po6119, po6120, po6121, po6122, po6123, po6124, po6125, po6126, po6127, po6128, po6129, po6130, po6131, po6132, po6133, po6134, po6135, po6136, po6137, po6138, po6139, po6140, po6141, po6142, po6143, po6144, po6145, po6146, po6147, po6148, po6149, po6150, po6151, po6152, po6153, po6154, po6155, po6156, po6157, po6158, po6159, po6160, po6161, po6162, po6163, po6164, po6165, po6166, po6167, po6168, po6169, po6170, po6171, po6172, po6173, po6174, po6175, po6176, po6177, po6178, po6179, po6180, po6181, po6182, po6183, po6184, po6185, po6186, po6187, po6188, po6189, po6190, po6191, po6192, po6193, po6194, po6195, po6196, po6197, po6198, po6199, po6200, po6201, po6202, po6203, po6204, po6205, po6206, po6207, po6208, po6209, po6210, po6211, po6212, po6213, po6214, po6215, po6216, po6217, po6218, po6219, po6220, po6221, po6222, po6223, po6224, po6225, po6226, po6227, po6228, po6229, po6230, po6231, po6232, po6233, po6234, po6235, po6236, po6237, po6238, po6239, po6240, po6241, po6242, po6243, po6244, po6245, po6246, po6247, po6248, po6249, po6250, po6251, po6252, po6253, po6254, po6255, po6256, po6257, po6258, po6259, po6260, po6261, po6262, po6263, po6264, po6265, po6266, po6267, po6268, po6269, po6270, po6271, po6272, po6273, po6274, po6275, po6276, po6277, po6278, po6279, po6280, po6281, po6282, po6283, po6284, po6285, po6286, po6287, po6288, po6289, po6290, po6291, po6292, po6293, po6294, po6295, po6296, po6297, po6298, po6299, po6300, po6301, po6302, po6303, po6304, po6305, po6306, po6307, po6308, po6309, po6310, po6311, po6312, po6313, po6314, po6315, po6316, po6317, po6318, po6319, po6320, po6321, po6322, po6323, po6324, po6325, po6326, po6327, po6328, po6329, po6330, po6331, po6332, po6333, po6334, po6335, po6336, po6337, po6338, po6339, po6340, po6341, po6342, po6343, po6344, po6345, po6346, po6347, po6348, po6349, po6350, po6351, po6352, po6353, po6354, po6355, po6356, po6357, po6358, po6359, po6360, po6361, po6362, po6363, po6364, po6365, po6366, po6367, po6368, po6369, po6370, po6371, po6372, po6373, po6374, po6375, po6376, po6377, po6378, po6379, po6380, po6381, po6382, po6383, po6384, po6385, po6386, po6387, po6388, po6389, po6390, po6391, po6392, po6393, po6394, po6395, po6396, po6397, po6398, po6399, po6400, po6401, po6402, po6403, po6404, po6405, po6406, po6407, po6408, po6409, po6410, po6411, po6412, po6413, po6414, po6415, po6416, po6417, po6418, po6419, po6420, po6421, po6422, po6423, po6424, po6425, po6426, po6427, po6428, po6429, po6430, po6431, po6432, po6433, po6434, po6435, po6436, po6437, po6438, po6439, po6440, po6441, po6442, po6443, po6444, po6445, po6446, po6447, po6448, po6449, po6450, po6451, po6452, po6453, po6454, po6455, po6456, po6457, po6458, po6459, po6460, po6461, po6462, po6463, po6464, po6465, po6466, po6467, po6468, po6469, po6470, po6471, po6472, po6473, po6474, po6475, po6476, po6477, po6478, po6479, po6480, po6481, po6482, po6483, po6484, po6485, po6486, po6487, po6488, po6489, po6490, po6491, po6492, po6493, po6494, po6495, po6496, po6497, po6498, po6499, po6500, po6501, po6502, po6503, po6504, po6505, po6506, po6507, po6508, po6509, po6510, po6511, po6512, po6513, po6514, po6515, po6516, po6517, po6518, po6519, po6520, po6521, po6522, po6523, po6524, po6525, po6526, po6527, po6528, po6529, po6530, po6531, po6532, po6533, po6534, po6535, po6536, po6537, po6538, po6539, po6540, po6541, po6542, po6543, po6544, po6545, po6546, po6547, po6548, po6549, po6550, po6551, po6552, po6553, po6554, po6555, po6556, po6557, po6558, po6559, po6560, po6561, po6562, po6563, po6564, po6565, po6566, po6567, po6568, po6569, po6570, po6571, po6572, po6573, po6574, po6575, po6576, po6577, po6578, po6579, po6580, po6581, po6582, po6583, po6584, po6585, po6586, po6587, po6588, po6589, po6590, po6591, po6592, po6593, po6594, po6595, po6596, po6597, po6598, po6599, po6600, po6601, po6602, po6603, po6604, po6605, po6606, po6607, po6608, po6609, po6610, po6611, po6612, po6613, po6614, po6615, po6616, po6617, po6618, po6619, po6620, po6621, po6622, po6623, po6624, po6625, po6626, po6627, po6628, po6629, po6630, po6631, po6632, po6633, po6634, po6635, po6636, po6637, po6638, po6639, po6640, po6641, po6642, po6643, po6644, po6645, po6646, po6647, po6648, po6649, po6650, po6651, po6652, po6653, po6654, po6655, po6656, po6657, po6658, po6659, po6660, po6661, po6662, po6663, po6664, po6665, po6666, po6667, po6668, po6669, po6670, po6671, po6672, po6673, po6674, po6675, po6676, po6677, po6678, po6679, po6680, po6681, po6682, po6683, po6684, po6685, po6686, po6687, po6688, po6689, po6690, po6691, po6692, po6693, po6694, po6695, po6696, po6697, po6698, po6699, po6700, po6701, po6702, po6703, po6704, po6705, po6706, po6707, po6708, po6709, po6710, po6711, po6712, po6713, po6714, po6715, po6716, po6717, po6718, po6719, po6720, po6721, po6722, po6723, po6724, po6725, po6726, po6727, po6728, po6729, po6730, po6731, po6732, po6733, po6734, po6735, po6736, po6737, po6738, po6739, po6740, po6741, po6742, po6743, po6744, po6745, po6746, po6747, po6748, po6749, po6750, po6751, po6752, po6753, po6754, po6755, po6756, po6757, po6758, po6759, po6760, po6761, po6762, po6763, po6764, po6765, po6766, po6767, po6768, po6769, po6770, po6771, po6772, po6773, po6774, po6775, po6776, po6777, po6778, po6779, po6780, po6781, po6782, po6783, po6784, po6785, po6786, po6787, po6788, po6789, po6790, po6791, po6792, po6793, po6794, po6795, po6796, po6797, po6798, po6799, po6800, po6801, po6802, po6803, po6804, po6805, po6806, po6807, po6808, po6809, po6810, po6811, po6812, po6813, po6814, po6815, po6816, po6817, po6818, po6819, po6820, po6821, po6822, po6823, po6824, po6825, po6826, po6827, po6828, po6829, po6830, po6831, po6832, po6833, po6834, po6835, po6836, po6837, po6838, po6839, po6840, po6841, po6842, po6843, po6844, po6845, po6846, po6847, po6848, po6849, po6850, po6851, po6852, po6853, po6854, po6855, po6856, po6857, po6858, po6859, po6860, po6861, po6862, po6863, po6864, po6865, po6866, po6867, po6868, po6869, po6870, po6871, po6872, po6873, po6874, po6875, po6876, po6877, po6878, po6879, po6880, po6881, po6882, po6883, po6884, po6885, po6886, po6887, po6888, po6889, po6890, po6891, po6892, po6893, po6894, po6895, po6896, po6897, po6898, po6899, po6900, po6901, po6902, po6903, po6904, po6905, po6906, po6907, po6908, po6909, po6910, po6911, po6912, po6913, po6914, po6915, po6916, po6917, po6918, po6919, po6920, po6921, po6922, po6923, po6924, po6925, po6926, po6927, po6928, po6929, po6930, po6931, po6932, po6933, po6934, po6935, po6936, po6937, po6938, po6939, po6940, po6941, po6942, po6943, po6944, po6945, po6946, po6947, po6948, po6949, po6950, po6951, po6952, po6953, po6954, po6955, po6956, po6957, po6958, po6959, po6960, po6961, po6962, po6963, po6964, po6965, po6966, po6967, po6968, po6969, po6970, po6971, po6972, po6973, po6974, po6975, po6976, po6977, po6978, po6979, po6980, po6981, po6982, po6983, po6984, po6985, po6986, po6987, po6988, po6989, po6990, po6991, po6992, po6993, po6994, po6995, po6996, po6997, po6998, po6999, po7000, po7001, po7002, po7003, po7004, po7005, po7006, po7007, po7008, po7009, po7010, po7011, po7012, po7013, po7014, po7015, po7016, po7017, po7018, po7019, po7020, po7021, po7022, po7023, po7024, po7025, po7026, po7027, po7028, po7029, po7030, po7031, po7032, po7033, po7034, po7035, po7036, po7037, po7038, po7039, po7040, po7041, po7042, po7043, po7044, po7045, po7046, po7047, po7048, po7049, po7050, po7051, po7052, po7053, po7054, po7055, po7056, po7057, po7058, po7059, po7060, po7061, po7062, po7063, po7064, po7065, po7066, po7067, po7068, po7069, po7070, po7071, po7072, po7073, po7074, po7075, po7076, po7077, po7078, po7079, po7080, po7081, po7082, po7083, po7084, po7085, po7086, po7087, po7088, po7089, po7090, po7091, po7092, po7093, po7094, po7095, po7096, po7097, po7098, po7099, po7100, po7101, po7102, po7103, po7104, po7105, po7106, po7107, po7108, po7109, po7110, po7111, po7112, po7113, po7114, po7115, po7116, po7117, po7118, po7119, po7120, po7121, po7122, po7123, po7124, po7125, po7126, po7127, po7128, po7129, po7130, po7131, po7132, po7133, po7134, po7135, po7136, po7137, po7138, po7139, po7140, po7141, po7142, po7143, po7144, po7145, po7146, po7147, po7148, po7149, po7150, po7151, po7152, po7153, po7154, po7155, po7156, po7157, po7158, po7159, po7160, po7161, po7162, po7163, po7164, po7165, po7166, po7167, po7168, po7169, po7170, po7171, po7172, po7173, po7174, po7175, po7176, po7177, po7178, po7179, po7180, po7181, po7182, po7183, po7184, po7185, po7186, po7187, po7188, po7189, po7190, po7191, po7192, po7193, po7194, po7195, po7196, po7197, po7198, po7199, po7200, po7201, po7202, po7203, po7204, po7205, po7206, po7207, po7208, po7209, po7210, po7211, po7212, po7213, po7214, po7215, po7216, po7217, po7218, po7219, po7220, po7221, po7222, po7223, po7224, po7225, po7226, po7227, po7228, po7229, po7230, po7231, po7232, po7233, po7234, po7235, po7236, po7237, po7238, po7239, po7240, po7241, po7242, po7243, po7244, po7245, po7246, po7247, po7248, po7249, po7250, po7251, po7252, po7253, po7254, po7255, po7256, po7257, po7258, po7259, po7260, po7261, po7262, po7263, po7264, po7265, po7266, po7267, po7268, po7269, po7270, po7271, po7272, po7273, po7274, po7275, po7276, po7277, po7278, po7279, po7280, po7281, po7282, po7283, po7284, po7285, po7286, po7287, po7288, po7289, po7290, po7291, po7292, po7293, po7294, po7295, po7296, po7297, po7298, po7299, po7300, po7301, po7302, po7303, po7304, po7305, po7306, po7307, po7308, po7309, po7310, po7311, po7312, po7313, po7314, po7315, po7316, po7317, po7318, po7319, po7320, po7321, po7322, po7323, po7324, po7325, po7326, po7327, po7328, po7329, po7330, po7331, po7332, po7333, po7334, po7335, po7336, po7337, po7338, po7339, po7340, po7341, po7342, po7343, po7344, po7345, po7346, po7347, po7348, po7349, po7350, po7351, po7352, po7353, po7354, po7355, po7356, po7357, po7358, po7359, po7360, po7361, po7362, po7363, po7364, po7365, po7366, po7367, po7368, po7369, po7370, po7371, po7372, po7373, po7374, po7375, po7376, po7377, po7378, po7379, po7380, po7381, po7382, po7383, po7384, po7385, po7386, po7387, po7388, po7389, po7390, po7391, po7392, po7393, po7394, po7395, po7396, po7397, po7398, po7399, po7400, po7401, po7402, po7403, po7404, po7405, po7406, po7407, po7408, po7409, po7410, po7411, po7412, po7413, po7414, po7415, po7416, po7417, po7418, po7419, po7420, po7421, po7422, po7423, po7424, po7425, po7426, po7427, po7428, po7429, po7430, po7431, po7432, po7433, po7434, po7435, po7436, po7437, po7438, po7439, po7440, po7441, po7442, po7443, po7444, po7445, po7446, po7447, po7448, po7449, po7450, po7451, po7452, po7453, po7454, po7455, po7456, po7457, po7458, po7459, po7460, po7461, po7462, po7463, po7464, po7465, po7466, po7467, po7468, po7469, po7470, po7471, po7472, po7473, po7474, po7475, po7476, po7477, po7478, po7479, po7480, po7481, po7482, po7483, po7484, po7485, po7486, po7487, po7488, po7489, po7490, po7491, po7492, po7493, po7494, po7495, po7496, po7497, po7498, po7499, po7500, po7501, po7502, po7503, po7504, po7505, po7506, po7507, po7508, po7509, po7510, po7511, po7512, po7513, po7514, po7515, po7516, po7517, po7518, po7519, po7520, po7521, po7522, po7523, po7524, po7525, po7526, po7527, po7528, po7529, po7530, po7531, po7532, po7533, po7534, po7535, po7536, po7537, po7538, po7539, po7540, po7541, po7542, po7543, po7544, po7545, po7546, po7547, po7548, po7549, po7550, po7551, po7552, po7553, po7554, po7555, po7556, po7557, po7558, po7559, po7560, po7561, po7562, po7563, po7564, po7565, po7566, po7567, po7568, po7569, po7570, po7571, po7572, po7573, po7574, po7575, po7576, po7577, po7578, po7579, po7580, po7581, po7582, po7583, po7584, po7585, po7586, po7587, po7588, po7589, po7590, po7591, po7592, po7593, po7594, po7595, po7596, po7597, po7598, po7599, po7600, po7601, po7602, po7603, po7604, po7605, po7606, po7607, po7608, po7609, po7610, po7611, po7612, po7613, po7614, po7615, po7616, po7617, po7618, po7619, po7620, po7621, po7622, po7623, po7624, po7625, po7626, po7627, po7628, po7629, po7630, po7631, po7632, po7633, po7634, po7635, po7636, po7637, po7638, po7639, po7640, po7641, po7642, po7643, po7644, po7645, po7646, po7647, po7648, po7649, po7650, po7651, po7652, po7653, po7654, po7655, po7656, po7657, po7658, po7659, po7660, po7661, po7662, po7663, po7664, po7665, po7666, po7667, po7668, po7669, po7670, po7671, po7672, po7673, po7674, po7675, po7676, po7677, po7678, po7679, po7680, po7681, po7682, po7683, po7684, po7685, po7686, po7687, po7688, po7689, po7690, po7691, po7692, po7693, po7694, po7695, po7696, po7697, po7698, po7699, po7700, po7701, po7702, po7703, po7704, po7705, po7706, po7707, po7708, po7709, po7710, po7711, po7712, po7713, po7714, po7715, po7716, po7717, po7718, po7719, po7720, po7721, po7722, po7723, po7724, po7725, po7726, po7727, po7728, po7729, po7730, po7731, po7732, po7733, po7734, po7735, po7736, po7737, po7738, po7739, po7740, po7741, po7742, po7743, po7744, po7745, po7746, po7747, po7748, po7749, po7750, po7751, po7752, po7753, po7754, po7755, po7756, po7757, po7758, po7759, po7760, po7761, po7762, po7763, po7764, po7765, po7766, po7767, po7768, po7769, po7770, po7771, po7772, po7773, po7774, po7775, po7776, po7777, po7778, po7779, po7780, po7781, po7782, po7783, po7784, po7785, po7786, po7787, po7788, po7789, po7790, po7791, po7792, po7793, po7794, po7795, po7796, po7797, po7798, po7799, po7800, po7801, po7802, po7803, po7804, po7805, po7806, po7807, po7808, po7809, po7810, po7811, po7812, po7813, po7814, po7815, po7816, po7817, po7818, po7819, po7820, po7821, po7822, po7823, po7824, po7825, po7826, po7827, po7828, po7829, po7830, po7831, po7832, po7833, po7834, po7835, po7836, po7837, po7838, po7839, po7840, po7841, po7842, po7843, po7844, po7845, po7846, po7847, po7848, po7849, po7850, po7851, po7852, po7853, po7854, po7855, po7856, po7857, po7858, po7859, po7860, po7861, po7862, po7863, po7864, po7865, po7866, po7867, po7868, po7869, po7870, po7871, po7872, po7873, po7874, po7875, po7876, po7877, po7878, po7879, po7880, po7881, po7882, po7883, po7884, po7885, po7886, po7887, po7888, po7889, po7890, po7891, po7892, po7893, po7894, po7895, po7896, po7897, po7898, po7899, po7900, po7901, po7902, po7903, po7904, po7905, po7906, po7907, po7908, po7909, po7910, po7911, po7912, po7913, po7914, po7915, po7916, po7917, po7918, po7919, po7920, po7921, po7922, po7923, po7924, po7925, po7926, po7927, po7928, po7929, po7930, po7931, po7932, po7933, po7934, po7935, po7936, po7937, po7938, po7939, po7940, po7941, po7942, po7943, po7944, po7945, po7946, po7947, po7948, po7949, po7950, po7951, po7952, po7953, po7954, po7955, po7956, po7957, po7958, po7959, po7960, po7961, po7962, po7963, po7964, po7965, po7966, po7967, po7968, po7969, po7970, po7971, po7972, po7973, po7974, po7975, po7976, po7977, po7978, po7979, po7980, po7981, po7982, po7983, po7984, po7985, po7986, po7987, po7988, po7989, po7990, po7991, po7992, po7993, po7994, po7995, po7996, po7997, po7998, po7999, po8000, po8001, po8002, po8003, po8004, po8005, po8006, po8007, po8008, po8009, po8010, po8011, po8012, po8013, po8014, po8015, po8016, po8017, po8018, po8019, po8020, po8021, po8022, po8023, po8024, po8025, po8026, po8027, po8028, po8029, po8030, po8031, po8032, po8033, po8034, po8035, po8036, po8037, po8038, po8039, po8040, po8041, po8042, po8043, po8044, po8045, po8046, po8047, po8048, po8049, po8050, po8051, po8052, po8053, po8054, po8055, po8056, po8057, po8058, po8059, po8060, po8061, po8062, po8063, po8064, po8065, po8066, po8067, po8068, po8069, po8070, po8071, po8072, po8073, po8074, po8075, po8076, po8077, po8078, po8079, po8080, po8081, po8082, po8083, po8084, po8085, po8086, po8087, po8088, po8089, po8090, po8091, po8092, po8093, po8094, po8095, po8096, po8097, po8098, po8099, po8100, po8101, po8102, po8103, po8104, po8105, po8106, po8107, po8108, po8109, po8110, po8111, po8112, po8113, po8114, po8115, po8116, po8117, po8118, po8119, po8120, po8121, po8122, po8123, po8124, po8125, po8126, po8127, po8128, po8129, po8130, po8131, po8132, po8133, po8134, po8135, po8136, po8137, po8138, po8139, po8140, po8141, po8142, po8143, po8144, po8145, po8146, po8147, po8148, po8149, po8150, po8151, po8152, po8153, po8154, po8155, po8156, po8157, po8158, po8159, po8160, po8161, po8162, po8163, po8164, po8165, po8166, po8167, po8168, po8169, po8170, po8171, po8172, po8173, po8174, po8175, po8176, po8177, po8178, po8179, po8180, po8181, po8182, po8183, po8184, po8185, po8186, po8187, po8188, po8189, po8190, po8191, po8192, po8193, po8194, po8195, po8196, po8197, po8198, po8199, po8200, po8201, po8202, po8203, po8204, po8205, po8206, po8207, po8208, po8209, po8210, po8211, po8212, po8213, po8214, po8215, po8216, po8217, po8218, po8219, po8220, po8221, po8222, po8223, po8224, po8225, po8226, po8227, po8228, po8229, po8230, po8231, po8232, po8233, po8234, po8235, po8236, po8237, po8238, po8239, po8240, po8241, po8242, po8243, po8244, po8245, po8246, po8247, po8248, po8249, po8250, po8251, po8252, po8253, po8254, po8255, po8256, po8257, po8258, po8259, po8260, po8261, po8262, po8263, po8264, po8265, po8266, po8267, po8268, po8269, po8270, po8271, po8272, po8273, po8274, po8275, po8276, po8277, po8278, po8279, po8280, po8281, po8282, po8283, po8284, po8285, po8286, po8287, po8288, po8289, po8290, po8291, po8292, po8293, po8294, po8295, po8296, po8297, po8298, po8299, po8300, po8301, po8302, po8303, po8304, po8305, po8306, po8307, po8308, po8309, po8310, po8311, po8312, po8313, po8314, po8315, po8316, po8317, po8318, po8319, po8320, po8321, po8322, po8323, po8324, po8325, po8326, po8327, po8328, po8329, po8330, po8331, po8332, po8333, po8334, po8335, po8336, po8337, po8338, po8339, po8340, po8341, po8342, po8343, po8344, po8345, po8346, po8347, po8348, po8349, po8350, po8351, po8352, po8353, po8354, po8355, po8356, po8357, po8358, po8359, po8360, po8361, po8362, po8363, po8364, po8365, po8366, po8367, po8368, po8369, po8370, po8371, po8372, po8373, po8374, po8375, po8376, po8377, po8378, po8379, po8380, po8381, po8382, po8383, po8384, po8385, po8386, po8387, po8388, po8389, po8390, po8391, po8392, po8393, po8394, po8395, po8396, po8397, po8398, po8399, po8400, po8401, po8402, po8403, po8404, po8405, po8406, po8407, po8408, po8409, po8410, po8411, po8412, po8413, po8414, po8415, po8416, po8417, po8418, po8419, po8420, po8421, po8422, po8423, po8424, po8425, po8426, po8427, po8428, po8429, po8430, po8431, po8432, po8433, po8434, po8435, po8436, po8437, po8438, po8439, po8440, po8441, po8442, po8443, po8444, po8445, po8446, po8447, po8448, po8449, po8450, po8451, po8452, po8453, po8454, po8455, po8456, po8457, po8458, po8459, po8460, po8461, po8462, po8463, po8464, po8465, po8466, po8467, po8468, po8469, po8470, po8471, po8472, po8473, po8474, po8475, po8476, po8477, po8478, po8479, po8480, po8481, po8482, po8483, po8484, po8485, po8486, po8487, po8488, po8489, po8490, po8491, po8492, po8493, po8494, po8495, po8496, po8497, po8498, po8499, po8500, po8501, po8502, po8503, po8504, po8505, po8506, po8507, po8508, po8509, po8510, po8511, po8512, po8513, po8514, po8515, po8516, po8517, po8518, po8519, po8520, po8521, po8522, po8523, po8524, po8525, po8526, po8527, po8528, po8529, po8530, po8531, po8532, po8533, po8534, po8535, po8536, po8537, po8538, po8539, po8540, po8541, po8542, po8543, po8544, po8545, po8546, po8547, po8548, po8549, po8550, po8551, po8552, po8553, po8554, po8555, po8556, po8557, po8558, po8559, po8560, po8561, po8562, po8563, po8564, po8565, po8566, po8567, po8568, po8569, po8570, po8571, po8572, po8573, po8574, po8575, po8576, po8577, po8578, po8579, po8580, po8581, po8582, po8583, po8584, po8585, po8586, po8587, po8588, po8589, po8590, po8591, po8592, po8593, po8594, po8595, po8596, po8597, po8598, po8599, po8600, po8601, po8602, po8603, po8604, po8605, po8606, po8607, po8608, po8609, po8610, po8611, po8612, po8613, po8614, po8615, po8616, po8617, po8618, po8619, po8620, po8621, po8622, po8623, po8624, po8625, po8626, po8627, po8628, po8629, po8630, po8631, po8632, po8633, po8634, po8635, po8636, po8637, po8638, po8639, po8640, po8641, po8642, po8643, po8644, po8645, po8646, po8647, po8648, po8649, po8650, po8651, po8652, po8653, po8654, po8655, po8656, po8657, po8658, po8659, po8660, po8661, po8662, po8663, po8664, po8665, po8666, po8667, po8668, po8669, po8670, po8671, po8672, po8673, po8674, po8675, po8676, po8677, po8678, po8679, po8680, po8681, po8682, po8683, po8684, po8685, po8686, po8687, po8688, po8689, po8690, po8691, po8692, po8693, po8694, po8695, po8696, po8697, po8698, po8699, po8700, po8701, po8702, po8703, po8704, po8705, po8706, po8707, po8708, po8709, po8710, po8711, po8712, po8713, po8714, po8715, po8716, po8717, po8718, po8719, po8720, po8721, po8722, po8723, po8724, po8725, po8726, po8727, po8728, po8729, po8730, po8731, po8732, po8733, po8734, po8735, po8736, po8737, po8738, po8739, po8740, po8741, po8742, po8743, po8744, po8745, po8746, po8747, po8748, po8749, po8750, po8751, po8752, po8753, po8754, po8755, po8756, po8757, po8758, po8759, po8760, po8761, po8762, po8763, po8764, po8765, po8766, po8767, po8768, po8769, po8770, po8771, po8772, po8773, po8774, po8775, po8776, po8777, po8778, po8779, po8780, po8781, po8782, po8783, po8784, po8785, po8786, po8787, po8788, po8789, po8790, po8791, po8792, po8793, po8794, po8795, po8796, po8797, po8798, po8799, po8800, po8801, po8802, po8803, po8804, po8805, po8806, po8807, po8808, po8809, po8810, po8811, po8812, po8813, po8814, po8815, po8816, po8817, po8818, po8819, po8820, po8821, po8822, po8823, po8824, po8825, po8826, po8827, po8828, po8829, po8830, po8831, po8832, po8833, po8834, po8835, po8836, po8837, po8838, po8839, po8840, po8841, po8842, po8843, po8844, po8845, po8846, po8847, po8848, po8849, po8850, po8851, po8852, po8853, po8854, po8855, po8856, po8857, po8858, po8859, po8860, po8861, po8862, po8863, po8864, po8865, po8866, po8867, po8868, po8869, po8870, po8871, po8872, po8873, po8874, po8875, po8876, po8877, po8878, po8879, po8880, po8881, po8882, po8883, po8884, po8885, po8886, po8887, po8888, po8889, po8890, po8891, po8892, po8893, po8894, po8895, po8896, po8897, po8898, po8899, po8900, po8901, po8902, po8903, po8904, po8905, po8906, po8907, po8908, po8909, po8910, po8911, po8912, po8913, po8914, po8915, po8916, po8917, po8918, po8919, po8920, po8921, po8922, po8923, po8924, po8925, po8926, po8927, po8928, po8929, po8930, po8931, po8932, po8933, po8934, po8935, po8936, po8937, po8938, po8939, po8940, po8941, po8942, po8943, po8944, po8945, po8946, po8947, po8948, po8949, po8950, po8951, po8952, po8953, po8954, po8955, po8956, po8957, po8958, po8959, po8960, po8961, po8962, po8963, po8964, po8965, po8966, po8967, po8968, po8969, po8970, po8971, po8972, po8973, po8974, po8975, po8976, po8977, po8978, po8979, po8980, po8981, po8982, po8983, po8984, po8985, po8986, po8987, po8988, po8989, po8990, po8991, po8992, po8993, po8994, po8995, po8996, po8997, po8998, po8999, po9000, po9001, po9002, po9003, po9004, po9005, po9006, po9007, po9008, po9009, po9010, po9011, po9012, po9013, po9014, po9015, po9016, po9017, po9018, po9019, po9020, po9021, po9022, po9023, po9024, po9025, po9026, po9027, po9028, po9029, po9030, po9031, po9032, po9033, po9034, po9035, po9036, po9037;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211, w40212, w40213, w40214, w40215, w40216, w40217, w40218, w40219, w40220, w40221, w40222, w40223, w40224, w40225, w40226, w40227, w40228, w40229, w40230, w40231, w40232, w40233, w40234, w40235, w40236, w40237, w40238, w40239, w40240, w40241, w40242, w40243, w40244, w40245, w40246, w40247, w40248, w40249, w40250, w40251, w40252, w40253, w40254, w40255, w40256, w40257, w40258, w40259, w40260, w40261, w40262, w40263, w40264, w40265, w40266, w40267, w40268, w40269, w40270, w40271, w40272, w40273, w40274, w40275, w40276, w40277, w40278, w40279, w40280, w40281, w40282, w40283, w40284, w40285, w40286, w40287, w40288, w40289, w40290, w40291, w40292, w40293, w40294, w40295, w40296, w40297, w40298, w40299, w40300, w40301, w40302, w40303, w40304, w40305, w40306, w40307, w40308, w40309, w40310, w40311, w40312, w40313, w40314, w40315, w40316, w40317, w40318, w40319, w40320, w40321, w40322, w40323, w40324, w40325, w40326, w40327, w40328, w40329, w40330, w40331, w40332, w40333, w40334, w40335, w40336, w40337, w40338, w40339, w40340, w40341, w40342, w40343, w40344, w40345, w40346, w40347, w40348, w40349, w40350, w40351, w40352, w40353, w40354, w40355, w40356, w40357, w40358, w40359, w40360, w40361, w40362, w40363, w40364, w40365, w40366, w40367, w40368, w40369, w40370, w40371, w40372, w40373, w40374, w40375, w40376, w40377, w40378, w40379, w40380, w40381, w40382, w40383, w40384, w40385, w40386, w40387, w40388, w40389, w40390, w40391, w40392, w40393, w40394, w40395, w40396, w40397, w40398, w40399, w40400, w40401, w40402, w40403, w40404, w40405, w40406, w40407, w40408, w40409, w40410, w40411, w40412, w40413, w40414, w40415, w40416, w40417, w40418, w40419, w40420, w40421, w40422, w40423, w40424, w40425, w40426, w40427, w40428, w40429, w40430, w40431, w40432, w40433, w40434, w40435, w40436, w40437, w40438, w40439, w40440, w40441, w40442, w40443, w40444, w40445, w40446, w40447, w40448, w40449, w40450, w40451, w40452, w40453, w40454, w40455, w40456, w40457, w40458, w40459, w40460, w40461, w40462, w40463, w40464, w40465, w40466, w40467, w40468, w40469, w40470, w40471, w40472, w40473, w40474, w40475, w40476, w40477, w40478, w40479, w40480, w40481, w40482, w40483, w40484, w40485, w40486, w40487, w40488, w40489, w40490, w40491, w40492, w40493, w40494, w40495, w40496, w40497, w40498, w40499, w40500, w40501, w40502, w40503, w40504, w40505, w40506, w40507, w40508, w40509, w40510, w40511, w40512, w40513, w40514, w40515, w40516, w40517, w40518, w40519, w40520, w40521, w40522, w40523, w40524, w40525, w40526, w40527, w40528, w40529, w40530, w40531, w40532, w40533, w40534, w40535, w40536, w40537, w40538, w40539, w40540, w40541, w40542, w40543, w40544, w40545, w40546, w40547, w40548, w40549, w40550, w40551, w40552, w40553, w40554, w40555, w40556, w40557, w40558, w40559, w40560, w40561, w40562, w40563, w40564, w40565, w40566, w40567, w40568, w40569, w40570, w40571, w40572, w40573, w40574, w40575, w40576, w40577, w40578, w40579, w40580, w40581, w40582, w40583, w40584, w40585, w40586, w40587, w40588, w40589, w40590, w40591, w40592, w40593, w40594, w40595, w40596, w40597, w40598, w40599, w40600, w40601, w40602, w40603, w40604, w40605, w40606, w40607, w40608, w40609, w40610, w40611, w40612, w40613, w40614, w40615, w40616, w40617, w40618, w40619, w40620, w40621, w40622, w40623, w40624, w40625, w40626, w40627, w40628, w40629, w40630, w40631, w40632, w40633, w40634, w40635, w40636, w40637, w40638, w40639, w40640, w40641, w40642, w40643, w40644, w40645, w40646, w40647, w40648, w40649, w40650, w40651, w40652, w40653, w40654, w40655, w40656, w40657, w40658, w40659, w40660, w40661, w40662, w40663, w40664, w40665, w40666, w40667, w40668, w40669, w40670, w40671, w40672, w40673, w40674, w40675, w40676, w40677, w40678, w40679, w40680, w40681, w40682, w40683, w40684, w40685, w40686, w40687, w40688, w40689, w40690, w40691, w40692, w40693, w40694, w40695, w40696, w40697, w40698, w40699, w40700, w40701, w40702, w40703, w40704, w40705, w40706, w40707, w40708, w40709, w40710, w40711, w40712, w40713, w40714, w40715, w40716, w40717, w40718, w40719, w40720, w40721, w40722, w40723, w40724, w40725, w40726, w40727, w40728, w40729, w40730, w40731, w40732, w40733, w40734, w40735, w40736, w40737, w40738, w40739, w40740, w40741, w40742, w40743, w40744, w40745, w40746, w40747, w40748, w40749, w40750, w40751, w40752, w40753, w40754, w40755, w40756, w40757, w40758, w40759, w40760, w40761, w40762, w40763, w40764, w40765, w40766, w40767, w40768, w40769, w40770, w40771, w40772, w40773, w40774, w40775, w40776, w40777, w40778, w40779, w40780, w40781, w40782, w40783, w40784, w40785, w40786, w40787, w40788, w40789, w40790, w40791, w40792, w40793, w40794, w40795, w40796, w40797, w40798, w40799, w40800, w40801, w40802, w40803, w40804, w40805, w40806, w40807, w40808, w40809, w40810, w40811, w40812, w40813, w40814, w40815, w40816, w40817, w40818, w40819, w40820, w40821, w40822, w40823, w40824, w40825, w40826, w40827, w40828, w40829, w40830, w40831, w40832, w40833, w40834, w40835, w40836, w40837, w40838, w40839, w40840, w40841, w40842, w40843, w40844, w40845, w40846, w40847, w40848, w40849, w40850, w40851, w40852, w40853, w40854, w40855, w40856, w40857, w40858, w40859, w40860, w40861, w40862, w40863, w40864, w40865, w40866, w40867, w40868, w40869, w40870, w40871, w40872, w40873, w40874, w40875, w40876, w40877, w40878, w40879, w40880, w40881, w40882, w40883, w40884, w40885, w40886, w40887, w40888, w40889, w40890, w40891, w40892, w40893, w40894, w40895, w40896, w40897, w40898, w40899, w40900, w40901, w40902, w40903, w40904, w40905, w40906, w40907, w40908, w40909, w40910, w40911, w40912, w40913, w40914, w40915, w40916, w40917, w40918, w40919, w40920, w40921, w40922, w40923, w40924, w40925, w40926, w40927, w40928, w40929, w40930, w40931, w40932, w40933, w40934, w40935, w40936, w40937, w40938, w40939, w40940, w40941, w40942, w40943, w40944, w40945, w40946, w40947, w40948, w40949, w40950, w40951, w40952, w40953, w40954, w40955, w40956, w40957, w40958, w40959, w40960, w40961, w40962, w40963, w40964, w40965, w40966, w40967, w40968, w40969, w40970, w40971, w40972, w40973, w40974, w40975, w40976, w40977, w40978, w40979, w40980, w40981, w40982, w40983, w40984, w40985, w40986, w40987, w40988, w40989, w40990, w40991, w40992, w40993, w40994, w40995, w40996, w40997, w40998, w40999, w41000, w41001, w41002, w41003, w41004, w41005, w41006, w41007, w41008, w41009, w41010, w41011, w41012, w41013, w41014, w41015, w41016, w41017, w41018, w41019, w41020, w41021, w41022, w41023, w41024, w41025, w41026, w41027, w41028, w41029, w41030, w41031, w41032, w41033, w41034, w41035, w41036, w41037, w41038, w41039, w41040, w41041, w41042, w41043, w41044, w41045, w41046, w41047, w41048, w41049, w41050, w41051, w41052, w41053, w41054, w41055, w41056, w41057, w41058, w41059, w41060, w41061, w41062, w41063, w41064, w41065, w41066, w41067, w41068, w41069, w41070, w41071, w41072, w41073, w41074, w41075, w41076, w41077, w41078, w41079, w41080, w41081, w41082, w41083, w41084, w41085, w41086, w41087, w41088, w41089, w41090, w41091, w41092, w41093, w41094, w41095, w41096, w41097, w41098, w41099, w41100, w41101, w41102, w41103, w41104, w41105, w41106, w41107, w41108, w41109, w41110, w41111, w41112, w41113, w41114, w41115, w41116, w41117, w41118, w41119, w41120, w41121, w41122, w41123, w41124, w41125, w41126, w41127, w41128, w41129, w41130, w41131, w41132, w41133, w41134, w41135, w41136, w41137, w41138, w41139, w41140, w41141, w41142, w41143, w41144, w41145, w41146, w41147, w41148, w41149, w41150, w41151, w41152, w41153, w41154, w41155, w41156, w41157, w41158, w41159, w41160, w41161, w41162, w41163, w41164, w41165, w41166, w41167, w41168, w41169, w41170, w41171, w41172, w41173, w41174, w41175, w41176, w41177, w41178, w41179, w41180, w41181, w41182, w41183, w41184, w41185, w41186, w41187, w41188, w41189, w41190, w41191, w41192, w41193, w41194, w41195, w41196, w41197, w41198, w41199, w41200, w41201, w41202, w41203, w41204, w41205, w41206, w41207, w41208, w41209, w41210, w41211, w41212, w41213, w41214, w41215, w41216, w41217, w41218, w41219, w41220, w41221, w41222, w41223, w41224, w41225, w41226, w41227, w41228, w41229, w41230, w41231, w41232, w41233, w41234, w41235, w41236, w41237, w41238, w41239, w41240, w41241, w41242, w41243, w41244, w41245, w41246, w41247, w41248, w41249, w41250, w41251, w41252, w41253, w41254, w41255, w41256, w41257, w41258, w41259, w41260, w41261, w41262, w41263, w41264, w41265, w41266, w41267, w41268, w41269, w41270, w41271, w41272, w41273, w41274, w41275, w41276, w41277, w41278, w41279, w41280, w41281, w41282, w41283, w41284, w41285, w41286, w41287, w41288, w41289, w41290, w41291, w41292, w41293, w41294, w41295, w41296, w41297, w41298, w41299, w41300, w41301, w41302, w41303, w41304, w41305, w41306, w41307, w41308, w41309, w41310, w41311, w41312, w41313, w41314, w41315, w41316, w41317, w41318, w41319, w41320, w41321, w41322, w41323, w41324, w41325, w41326, w41327, w41328, w41329, w41330, w41331, w41332, w41333, w41334, w41335, w41336, w41337, w41338, w41339, w41340, w41341, w41342, w41343, w41344, w41345, w41346, w41347, w41348, w41349, w41350, w41351, w41352, w41353, w41354, w41355, w41356, w41357, w41358, w41359, w41360, w41361, w41362, w41363, w41364, w41365, w41366, w41367, w41368, w41369, w41370, w41371, w41372, w41373, w41374, w41375, w41376, w41377, w41378, w41379, w41380, w41381, w41382, w41383, w41384, w41385, w41386, w41387, w41388, w41389, w41390, w41391, w41392, w41393, w41394, w41395, w41396, w41397, w41398, w41399, w41400, w41401, w41402, w41403, w41404, w41405, w41406, w41407, w41408, w41409, w41410, w41411, w41412, w41413, w41414, w41415, w41416, w41417, w41418, w41419, w41420, w41421, w41422, w41423, w41424, w41425, w41426, w41427, w41428, w41429, w41430, w41431, w41432, w41433, w41434, w41435, w41436, w41437, w41438, w41439, w41440, w41441, w41442, w41443, w41444, w41445, w41446, w41447, w41448, w41449, w41450, w41451, w41452, w41453, w41454, w41455, w41456, w41457, w41458, w41459, w41460, w41461, w41462, w41463, w41464, w41465, w41466, w41467, w41468, w41469, w41470, w41471, w41472, w41473, w41474, w41475, w41476, w41477, w41478, w41479, w41480, w41481, w41482, w41483, w41484, w41485, w41486, w41487, w41488, w41489, w41490, w41491, w41492, w41493, w41494, w41495, w41496, w41497, w41498, w41499, w41500, w41501, w41502, w41503, w41504, w41505, w41506, w41507, w41508, w41509, w41510, w41511, w41512, w41513, w41514, w41515, w41516, w41517, w41518, w41519, w41520, w41521, w41522, w41523, w41524, w41525, w41526, w41527, w41528, w41529, w41530, w41531, w41532, w41533, w41534, w41535, w41536, w41537, w41538, w41539, w41540, w41541, w41542, w41543, w41544, w41545, w41546, w41547, w41548, w41549, w41550, w41551, w41552, w41553, w41554, w41555, w41556, w41557, w41558, w41559, w41560, w41561, w41562, w41563, w41564, w41565, w41566, w41567, w41568, w41569, w41570, w41571, w41572, w41573, w41574, w41575, w41576, w41577, w41578, w41579, w41580, w41581, w41582, w41583, w41584, w41585, w41586, w41587, w41588, w41589, w41590, w41591, w41592, w41593, w41594, w41595, w41596, w41597, w41598, w41599, w41600, w41601, w41602, w41603, w41604, w41605, w41606, w41607, w41608, w41609, w41610, w41611, w41612, w41613, w41614, w41615, w41616, w41617, w41618, w41619, w41620, w41621, w41622, w41623, w41624, w41625, w41626, w41627, w41628, w41629, w41630, w41631, w41632, w41633, w41634, w41635, w41636, w41637, w41638, w41639, w41640, w41641, w41642, w41643, w41644, w41645, w41646, w41647, w41648, w41649, w41650, w41651, w41652, w41653, w41654, w41655, w41656, w41657, w41658, w41659, w41660, w41661, w41662, w41663, w41664, w41665, w41666, w41667, w41668, w41669, w41670, w41671, w41672, w41673, w41674, w41675, w41676, w41677, w41678, w41679, w41680, w41681, w41682, w41683, w41684, w41685, w41686, w41687, w41688, w41689, w41690, w41691, w41692, w41693, w41694, w41695, w41696, w41697, w41698, w41699, w41700, w41701, w41702, w41703, w41704, w41705, w41706, w41707, w41708, w41709, w41710, w41711, w41712, w41713, w41714, w41715, w41716, w41717, w41718, w41719, w41720, w41721, w41722, w41723, w41724, w41725, w41726, w41727, w41728, w41729, w41730, w41731, w41732, w41733, w41734, w41735, w41736, w41737, w41738, w41739, w41740, w41741, w41742, w41743, w41744, w41745, w41746, w41747, w41748, w41749, w41750, w41751, w41752, w41753, w41754, w41755, w41756, w41757, w41758, w41759, w41760, w41761, w41762, w41763, w41764, w41765, w41766, w41767, w41768, w41769, w41770, w41771, w41772, w41773, w41774, w41775, w41776, w41777, w41778, w41779, w41780, w41781, w41782, w41783, w41784, w41785, w41786, w41787, w41788, w41789, w41790, w41791, w41792, w41793, w41794, w41795, w41796, w41797, w41798, w41799, w41800, w41801, w41802, w41803, w41804, w41805, w41806, w41807, w41808, w41809, w41810, w41811, w41812, w41813, w41814, w41815, w41816, w41817, w41818, w41819, w41820, w41821, w41822, w41823, w41824, w41825, w41826, w41827, w41828, w41829, w41830, w41831, w41832, w41833, w41834, w41835, w41836, w41837, w41838, w41839, w41840, w41841, w41842, w41843, w41844, w41845, w41846, w41847, w41848, w41849, w41850, w41851, w41852, w41853, w41854, w41855, w41856, w41857, w41858, w41859, w41860, w41861, w41862, w41863, w41864, w41865, w41866, w41867, w41868, w41869, w41870, w41871, w41872, w41873, w41874, w41875, w41876, w41877, w41878, w41879, w41880, w41881, w41882, w41883, w41884, w41885, w41886, w41887, w41888, w41889, w41890, w41891, w41892, w41893, w41894, w41895, w41896, w41897, w41898, w41899, w41900, w41901, w41902, w41903, w41904, w41905, w41906, w41907, w41908, w41909, w41910, w41911, w41912, w41913, w41914, w41915, w41916, w41917, w41918, w41919, w41920, w41921, w41922, w41923, w41924, w41925, w41926, w41927, w41928, w41929, w41930, w41931, w41932, w41933, w41934, w41935, w41936, w41937, w41938, w41939, w41940, w41941, w41942, w41943, w41944, w41945, w41946, w41947, w41948, w41949, w41950, w41951, w41952, w41953, w41954, w41955, w41956, w41957, w41958, w41959, w41960, w41961, w41962, w41963, w41964, w41965, w41966, w41967, w41968, w41969, w41970, w41971, w41972, w41973, w41974, w41975, w41976, w41977, w41978, w41979, w41980, w41981, w41982, w41983, w41984, w41985, w41986, w41987, w41988, w41989, w41990, w41991, w41992, w41993, w41994, w41995, w41996, w41997, w41998, w41999, w42000, w42001, w42002, w42003, w42004, w42005, w42006, w42007, w42008, w42009, w42010, w42011, w42012, w42013, w42014, w42015, w42016, w42017, w42018, w42019, w42020, w42021, w42022, w42023, w42024, w42025, w42026, w42027, w42028, w42029, w42030, w42031, w42032, w42033, w42034, w42035, w42036, w42037, w42038, w42039, w42040, w42041, w42042, w42043, w42044, w42045, w42046, w42047, w42048, w42049, w42050, w42051, w42052, w42053, w42054, w42055, w42056, w42057, w42058, w42059, w42060, w42061, w42062, w42063, w42064, w42065, w42066, w42067, w42068, w42069, w42070, w42071, w42072, w42073, w42074, w42075, w42076, w42077, w42078, w42079, w42080, w42081, w42082, w42083, w42084, w42085, w42086, w42087, w42088, w42089, w42090, w42091, w42092, w42093, w42094, w42095, w42096, w42097, w42098, w42099, w42100, w42101, w42102, w42103, w42104, w42105, w42106, w42107, w42108, w42109, w42110, w42111, w42112, w42113, w42114, w42115, w42116, w42117, w42118, w42119, w42120, w42121, w42122, w42123, w42124, w42125, w42126, w42127, w42128, w42129, w42130, w42131, w42132, w42133, w42134, w42135, w42136, w42137, w42138, w42139, w42140, w42141, w42142, w42143, w42144, w42145, w42146, w42147, w42148, w42149, w42150, w42151, w42152, w42153, w42154, w42155, w42156, w42157, w42158, w42159, w42160, w42161, w42162, w42163, w42164, w42165, w42166, w42167, w42168, w42169, w42170, w42171, w42172, w42173, w42174, w42175, w42176, w42177, w42178, w42179, w42180, w42181, w42182, w42183, w42184, w42185, w42186, w42187, w42188, w42189, w42190, w42191, w42192, w42193, w42194, w42195, w42196, w42197, w42198, w42199, w42200, w42201, w42202, w42203, w42204, w42205, w42206, w42207, w42208, w42209, w42210, w42211, w42212, w42213, w42214, w42215, w42216, w42217, w42218, w42219, w42220, w42221, w42222, w42223, w42224, w42225, w42226, w42227, w42228, w42229, w42230, w42231, w42232, w42233, w42234, w42235, w42236, w42237, w42238, w42239, w42240, w42241, w42242, w42243, w42244, w42245, w42246, w42247, w42248, w42249, w42250, w42251, w42252, w42253, w42254, w42255, w42256, w42257, w42258, w42259, w42260, w42261, w42262, w42263, w42264, w42265, w42266, w42267, w42268, w42269, w42270, w42271, w42272, w42273, w42274, w42275, w42276, w42277, w42278, w42279, w42280, w42281, w42282, w42283, w42284, w42285, w42286, w42287, w42288, w42289, w42290, w42291, w42292, w42293, w42294, w42295, w42296, w42297, w42298, w42299, w42300, w42301, w42302, w42303, w42304, w42305, w42306, w42307, w42308, w42309, w42310, w42311, w42312, w42313, w42314, w42315, w42316, w42317, w42318, w42319, w42320, w42321, w42322, w42323, w42324, w42325, w42326, w42327, w42328, w42329, w42330, w42331, w42332, w42333, w42334, w42335, w42336, w42337, w42338, w42339, w42340, w42341, w42342, w42343, w42344, w42345, w42346, w42347, w42348, w42349, w42350, w42351, w42352, w42353, w42354, w42355, w42356, w42357, w42358, w42359, w42360, w42361, w42362, w42363, w42364, w42365, w42366, w42367, w42368, w42369, w42370, w42371, w42372, w42373, w42374, w42375, w42376, w42377, w42378, w42379, w42380, w42381, w42382, w42383, w42384, w42385, w42386, w42387, w42388, w42389, w42390, w42391, w42392, w42393, w42394, w42395, w42396, w42397, w42398, w42399, w42400, w42401, w42402, w42403, w42404, w42405, w42406, w42407, w42408, w42409, w42410, w42411, w42412, w42413, w42414, w42415, w42416, w42417, w42418, w42419, w42420, w42421, w42422, w42423, w42424, w42425, w42426, w42427, w42428, w42429, w42430, w42431, w42432, w42433, w42434, w42435, w42436, w42437, w42438, w42439, w42440, w42441, w42442, w42443, w42444, w42445, w42446, w42447, w42448, w42449, w42450, w42451, w42452, w42453, w42454, w42455, w42456, w42457, w42458, w42459, w42460, w42461, w42462, w42463, w42464, w42465, w42466, w42467, w42468, w42469, w42470, w42471, w42472, w42473, w42474, w42475, w42476, w42477, w42478, w42479, w42480, w42481, w42482, w42483, w42484, w42485, w42486, w42487, w42488, w42489, w42490, w42491, w42492, w42493, w42494, w42495, w42496, w42497, w42498, w42499, w42500, w42501, w42502, w42503, w42504, w42505, w42506, w42507, w42508, w42509, w42510, w42511, w42512, w42513, w42514, w42515, w42516, w42517, w42518, w42519, w42520, w42521, w42522, w42523, w42524, w42525, w42526, w42527, w42528, w42529, w42530, w42531, w42532, w42533, w42534, w42535, w42536, w42537, w42538, w42539, w42540, w42541, w42542, w42543, w42544, w42545, w42546, w42547, w42548, w42549, w42550, w42551, w42552, w42553, w42554, w42555, w42556, w42557, w42558, w42559, w42560, w42561, w42562, w42563, w42564, w42565, w42566, w42567, w42568, w42569, w42570, w42571, w42572, w42573, w42574, w42575, w42576, w42577, w42578, w42579, w42580, w42581, w42582, w42583, w42584, w42585, w42586, w42587, w42588, w42589, w42590, w42591, w42592, w42593, w42594, w42595, w42596, w42597, w42598, w42599, w42600, w42601, w42602, w42603, w42604, w42605, w42606, w42607, w42608, w42609, w42610, w42611, w42612, w42613, w42614, w42615, w42616, w42617, w42618, w42619, w42620, w42621, w42622, w42623, w42624, w42625, w42626, w42627, w42628, w42629, w42630, w42631, w42632, w42633, w42634, w42635, w42636, w42637, w42638, w42639, w42640, w42641, w42642, w42643, w42644, w42645, w42646, w42647, w42648, w42649, w42650, w42651, w42652, w42653, w42654, w42655, w42656, w42657, w42658, w42659, w42660, w42661, w42662, w42663, w42664, w42665, w42666, w42667, w42668, w42669, w42670, w42671, w42672, w42673, w42674, w42675, w42676, w42677, w42678, w42679, w42680, w42681, w42682, w42683, w42684, w42685, w42686, w42687, w42688, w42689, w42690, w42691, w42692, w42693, w42694, w42695, w42696, w42697, w42698, w42699, w42700, w42701, w42702, w42703, w42704, w42705, w42706, w42707, w42708, w42709, w42710, w42711, w42712, w42713, w42714, w42715, w42716, w42717, w42718, w42719, w42720, w42721, w42722, w42723, w42724, w42725, w42726, w42727, w42728, w42729, w42730, w42731, w42732, w42733, w42734, w42735, w42736, w42737, w42738, w42739, w42740, w42741, w42742, w42743, w42744, w42745, w42746, w42747, w42748, w42749, w42750, w42751, w42752, w42753, w42754, w42755, w42756, w42757, w42758, w42759, w42760, w42761, w42762, w42763, w42764, w42765, w42766, w42767, w42768, w42769, w42770, w42771, w42772, w42773, w42774, w42775, w42776, w42777, w42778, w42779, w42780, w42781, w42782, w42783, w42784, w42785, w42786, w42787, w42788, w42789, w42790, w42791, w42792, w42793, w42794, w42795, w42796, w42797, w42798, w42799, w42800, w42801, w42802, w42803, w42804, w42805, w42806, w42807, w42808, w42809, w42810, w42811, w42812, w42813, w42814, w42815, w42816, w42817, w42818, w42819, w42820, w42821, w42822, w42823, w42824, w42825, w42826, w42827, w42828, w42829, w42830, w42831, w42832, w42833, w42834, w42835, w42836, w42837, w42838, w42839, w42840, w42841, w42842, w42843, w42844, w42845, w42846, w42847, w42848, w42849, w42850, w42851, w42852, w42853, w42854, w42855, w42856, w42857, w42858, w42859, w42860, w42861, w42862, w42863, w42864, w42865, w42866, w42867, w42868, w42869, w42870, w42871, w42872, w42873, w42874, w42875, w42876, w42877, w42878, w42879, w42880, w42881, w42882, w42883, w42884, w42885, w42886, w42887, w42888, w42889, w42890, w42891, w42892, w42893, w42894, w42895, w42896, w42897, w42898, w42899, w42900, w42901, w42902, w42903, w42904, w42905, w42906, w42907, w42908, w42909, w42910, w42911, w42912, w42913, w42914, w42915, w42916, w42917, w42918, w42919, w42920, w42921, w42922, w42923, w42924, w42925, w42926, w42927, w42928, w42929, w42930, w42931, w42932, w42933, w42934, w42935, w42936, w42937, w42938, w42939, w42940, w42941, w42942, w42943, w42944, w42945, w42946, w42947, w42948, w42949, w42950, w42951, w42952, w42953, w42954, w42955, w42956, w42957, w42958, w42959, w42960, w42961, w42962, w42963, w42964, w42965, w42966, w42967, w42968, w42969, w42970, w42971, w42972, w42973, w42974, w42975, w42976, w42977, w42978, w42979, w42980, w42981, w42982, w42983, w42984, w42985, w42986, w42987, w42988, w42989, w42990, w42991, w42992, w42993, w42994, w42995, w42996, w42997, w42998, w42999, w43000, w43001, w43002, w43003, w43004, w43005, w43006, w43007, w43008, w43009, w43010, w43011, w43012, w43013, w43014, w43015, w43016, w43017, w43018, w43019, w43020, w43021, w43022, w43023, w43024, w43025, w43026, w43027, w43028, w43029, w43030, w43031, w43032, w43033, w43034, w43035, w43036, w43037, w43038, w43039, w43040, w43041, w43042, w43043, w43044, w43045, w43046, w43047, w43048, w43049, w43050, w43051, w43052, w43053, w43054, w43055, w43056, w43057, w43058, w43059, w43060, w43061, w43062, w43063, w43064, w43065, w43066, w43067, w43068, w43069, w43070, w43071, w43072, w43073, w43074, w43075, w43076, w43077, w43078, w43079, w43080, w43081, w43082, w43083, w43084, w43085, w43086, w43087, w43088, w43089, w43090, w43091, w43092, w43093, w43094, w43095, w43096, w43097, w43098, w43099, w43100, w43101, w43102, w43103, w43104, w43105, w43106, w43107, w43108, w43109, w43110, w43111, w43112, w43113, w43114, w43115, w43116, w43117, w43118, w43119, w43120, w43121, w43122, w43123, w43124, w43125, w43126, w43127, w43128, w43129, w43130, w43131, w43132, w43133, w43134, w43135, w43136, w43137, w43138, w43139, w43140, w43141, w43142, w43143, w43144, w43145, w43146, w43147, w43148, w43149, w43150, w43151, w43152, w43153, w43154, w43155, w43156, w43157, w43158, w43159, w43160, w43161, w43162, w43163, w43164, w43165, w43166, w43167, w43168, w43169, w43170, w43171, w43172, w43173, w43174, w43175, w43176, w43177, w43178, w43179, w43180, w43181, w43182, w43183, w43184, w43185, w43186, w43187, w43188, w43189, w43190, w43191, w43192, w43193, w43194, w43195, w43196, w43197, w43198, w43199, w43200, w43201, w43202, w43203, w43204, w43205, w43206, w43207, w43208, w43209, w43210, w43211, w43212, w43213, w43214, w43215, w43216, w43217, w43218, w43219, w43220, w43221, w43222, w43223, w43224, w43225, w43226, w43227, w43228, w43229, w43230, w43231, w43232, w43233, w43234, w43235, w43236, w43237, w43238, w43239, w43240, w43241, w43242, w43243, w43244, w43245, w43246, w43247, w43248, w43249, w43250, w43251, w43252, w43253, w43254, w43255, w43256, w43257, w43258, w43259, w43260, w43261, w43262, w43263, w43264, w43265, w43266, w43267, w43268, w43269, w43270, w43271, w43272, w43273, w43274, w43275, w43276, w43277, w43278, w43279, w43280, w43281, w43282, w43283, w43284, w43285, w43286, w43287, w43288, w43289, w43290, w43291, w43292, w43293, w43294, w43295, w43296, w43297, w43298, w43299, w43300, w43301, w43302, w43303, w43304, w43305, w43306, w43307, w43308, w43309, w43310, w43311, w43312, w43313, w43314, w43315, w43316, w43317, w43318, w43319, w43320, w43321, w43322, w43323, w43324, w43325, w43326, w43327, w43328, w43329, w43330, w43331, w43332, w43333, w43334, w43335, w43336, w43337, w43338, w43339, w43340, w43341, w43342, w43343, w43344, w43345, w43346, w43347, w43348, w43349, w43350, w43351, w43352, w43353, w43354, w43355, w43356, w43357, w43358, w43359, w43360, w43361, w43362, w43363, w43364, w43365, w43366, w43367, w43368, w43369, w43370, w43371, w43372, w43373, w43374, w43375, w43376, w43377, w43378, w43379, w43380, w43381, w43382, w43383, w43384, w43385, w43386, w43387, w43388, w43389, w43390, w43391, w43392, w43393, w43394, w43395, w43396, w43397, w43398, w43399, w43400, w43401, w43402, w43403, w43404, w43405, w43406, w43407, w43408, w43409, w43410, w43411, w43412, w43413, w43414, w43415, w43416, w43417, w43418, w43419, w43420, w43421, w43422, w43423, w43424, w43425, w43426, w43427, w43428, w43429, w43430, w43431, w43432, w43433, w43434, w43435, w43436, w43437, w43438, w43439, w43440, w43441, w43442, w43443, w43444, w43445, w43446, w43447, w43448, w43449, w43450, w43451, w43452, w43453, w43454, w43455, w43456, w43457, w43458, w43459, w43460, w43461, w43462, w43463, w43464, w43465, w43466, w43467, w43468, w43469, w43470, w43471, w43472, w43473, w43474, w43475, w43476, w43477, w43478, w43479, w43480, w43481, w43482, w43483, w43484, w43485, w43486, w43487, w43488, w43489, w43490, w43491, w43492, w43493, w43494, w43495, w43496, w43497, w43498, w43499, w43500, w43501, w43502, w43503, w43504, w43505, w43506, w43507, w43508, w43509, w43510, w43511, w43512, w43513, w43514, w43515, w43516, w43517, w43518, w43519, w43520, w43521, w43522, w43523, w43524, w43525, w43526, w43527, w43528, w43529, w43530, w43531, w43532, w43533, w43534, w43535, w43536, w43537, w43538, w43539, w43540, w43541, w43542, w43543, w43544, w43545, w43546, w43547, w43548, w43549, w43550, w43551, w43552, w43553, w43554, w43555, w43556, w43557, w43558, w43559, w43560, w43561, w43562, w43563, w43564, w43565, w43566, w43567, w43568, w43569, w43570, w43571, w43572, w43573, w43574, w43575, w43576, w43577, w43578, w43579, w43580, w43581, w43582, w43583, w43584, w43585, w43586, w43587, w43588, w43589, w43590, w43591, w43592, w43593, w43594, w43595, w43596, w43597, w43598, w43599, w43600, w43601, w43602, w43603, w43604, w43605, w43606, w43607, w43608, w43609, w43610, w43611, w43612, w43613, w43614, w43615, w43616, w43617, w43618, w43619, w43620, w43621, w43622, w43623, w43624, w43625, w43626, w43627, w43628, w43629, w43630, w43631, w43632, w43633, w43634, w43635, w43636, w43637, w43638, w43639, w43640, w43641, w43642, w43643, w43644, w43645, w43646, w43647, w43648, w43649, w43650, w43651, w43652, w43653, w43654, w43655, w43656, w43657, w43658, w43659, w43660, w43661, w43662, w43663, w43664, w43665, w43666, w43667, w43668, w43669, w43670, w43671, w43672, w43673, w43674, w43675, w43676, w43677, w43678, w43679, w43680, w43681, w43682, w43683, w43684, w43685, w43686, w43687, w43688, w43689, w43690, w43691, w43692, w43693, w43694, w43695, w43696, w43697, w43698, w43699, w43700, w43701, w43702, w43703, w43704, w43705, w43706, w43707, w43708, w43709, w43710, w43711, w43712, w43713, w43714, w43715, w43716, w43717, w43718, w43719, w43720, w43721, w43722, w43723, w43724, w43725, w43726, w43727, w43728, w43729, w43730, w43731, w43732, w43733, w43734, w43735, w43736, w43737, w43738, w43739, w43740, w43741, w43742, w43743, w43744, w43745, w43746, w43747, w43748, w43749, w43750, w43751, w43752, w43753, w43754, w43755, w43756, w43757, w43758, w43759, w43760, w43761, w43762, w43763, w43764, w43765, w43766, w43767, w43768, w43769, w43770, w43771, w43772, w43773, w43774, w43775, w43776, w43777, w43778, w43779, w43780, w43781, w43782, w43783, w43784, w43785, w43786, w43787, w43788, w43789, w43790, w43791, w43792, w43793, w43794, w43795, w43796, w43797, w43798, w43799, w43800, w43801, w43802, w43803, w43804, w43805, w43806, w43807, w43808, w43809, w43810, w43811, w43812, w43813, w43814, w43815, w43816, w43817, w43818, w43819, w43820, w43821, w43822, w43823, w43824, w43825, w43826, w43827, w43828, w43829, w43830, w43831, w43832, w43833, w43834, w43835, w43836, w43837, w43838, w43839, w43840, w43841, w43842, w43843, w43844, w43845, w43846, w43847, w43848, w43849, w43850, w43851, w43852, w43853, w43854, w43855, w43856, w43857, w43858, w43859, w43860, w43861, w43862, w43863, w43864, w43865, w43866, w43867, w43868, w43869, w43870, w43871, w43872, w43873, w43874, w43875, w43876, w43877, w43878, w43879, w43880, w43881, w43882, w43883, w43884, w43885, w43886, w43887, w43888, w43889, w43890, w43891, w43892, w43893, w43894, w43895, w43896, w43897, w43898, w43899, w43900, w43901, w43902, w43903, w43904, w43905, w43906, w43907, w43908, w43909, w43910, w43911, w43912, w43913, w43914, w43915, w43916, w43917, w43918, w43919, w43920, w43921, w43922, w43923, w43924, w43925, w43926, w43927, w43928, w43929, w43930, w43931, w43932, w43933, w43934, w43935, w43936, w43937, w43938, w43939, w43940, w43941, w43942, w43943, w43944, w43945, w43946, w43947, w43948, w43949, w43950, w43951, w43952, w43953, w43954, w43955, w43956, w43957, w43958, w43959, w43960, w43961, w43962, w43963, w43964, w43965, w43966, w43967, w43968, w43969, w43970, w43971, w43972, w43973, w43974, w43975, w43976, w43977, w43978, w43979, w43980, w43981, w43982, w43983, w43984, w43985, w43986, w43987, w43988, w43989, w43990, w43991, w43992, w43993, w43994, w43995, w43996, w43997, w43998, w43999, w44000, w44001, w44002, w44003, w44004, w44005, w44006, w44007, w44008, w44009, w44010, w44011, w44012, w44013, w44014, w44015, w44016, w44017, w44018, w44019, w44020, w44021, w44022, w44023, w44024, w44025, w44026, w44027, w44028, w44029, w44030, w44031, w44032, w44033, w44034, w44035, w44036, w44037, w44038, w44039, w44040, w44041, w44042, w44043, w44044, w44045, w44046, w44047, w44048, w44049, w44050, w44051, w44052, w44053, w44054, w44055, w44056, w44057, w44058, w44059, w44060, w44061, w44062, w44063, w44064, w44065, w44066, w44067, w44068, w44069, w44070, w44071, w44072, w44073, w44074, w44075, w44076, w44077, w44078, w44079, w44080, w44081, w44082, w44083, w44084, w44085, w44086, w44087, w44088, w44089, w44090, w44091, w44092, w44093, w44094, w44095, w44096, w44097, w44098, w44099, w44100, w44101, w44102, w44103, w44104, w44105, w44106, w44107, w44108, w44109, w44110, w44111, w44112, w44113, w44114, w44115, w44116, w44117, w44118, w44119, w44120, w44121, w44122, w44123, w44124, w44125, w44126, w44127, w44128, w44129, w44130, w44131, w44132, w44133, w44134, w44135, w44136, w44137, w44138, w44139, w44140, w44141, w44142, w44143, w44144, w44145, w44146, w44147, w44148, w44149, w44150, w44151, w44152, w44153, w44154, w44155, w44156, w44157, w44158, w44159, w44160, w44161, w44162, w44163, w44164, w44165, w44166, w44167, w44168, w44169, w44170, w44171, w44172, w44173, w44174, w44175, w44176, w44177, w44178, w44179, w44180, w44181, w44182, w44183, w44184, w44185, w44186, w44187, w44188, w44189, w44190, w44191, w44192, w44193, w44194, w44195, w44196, w44197, w44198, w44199, w44200, w44201, w44202, w44203, w44204, w44205, w44206, w44207, w44208, w44209, w44210, w44211, w44212, w44213, w44214, w44215, w44216, w44217, w44218, w44219, w44220, w44221, w44222, w44223, w44224, w44225, w44226, w44227, w44228, w44229, w44230, w44231, w44232, w44233, w44234, w44235, w44236, w44237, w44238, w44239, w44240, w44241, w44242, w44243, w44244, w44245, w44246, w44247, w44248, w44249, w44250, w44251, w44252, w44253, w44254, w44255, w44256, w44257, w44258, w44259, w44260, w44261, w44262, w44263, w44264, w44265, w44266, w44267, w44268, w44269, w44270, w44271, w44272, w44273, w44274, w44275, w44276, w44277, w44278, w44279, w44280, w44281, w44282, w44283, w44284, w44285, w44286, w44287, w44288, w44289, w44290, w44291, w44292, w44293, w44294, w44295, w44296, w44297, w44298, w44299, w44300, w44301, w44302, w44303, w44304, w44305, w44306, w44307, w44308, w44309, w44310, w44311, w44312, w44313, w44314, w44315, w44316, w44317, w44318, w44319, w44320, w44321, w44322, w44323, w44324, w44325, w44326, w44327, w44328, w44329, w44330, w44331, w44332, w44333, w44334, w44335, w44336, w44337, w44338, w44339, w44340, w44341, w44342, w44343, w44344, w44345, w44346, w44347, w44348, w44349, w44350, w44351, w44352, w44353, w44354, w44355, w44356, w44357, w44358, w44359, w44360, w44361, w44362, w44363, w44364, w44365, w44366, w44367, w44368, w44369, w44370, w44371, w44372, w44373, w44374, w44375, w44376, w44377, w44378, w44379, w44380, w44381, w44382, w44383, w44384, w44385, w44386, w44387, w44388, w44389, w44390, w44391, w44392, w44393, w44394, w44395, w44396, w44397, w44398, w44399, w44400, w44401, w44402, w44403, w44404, w44405, w44406, w44407, w44408, w44409, w44410, w44411, w44412, w44413, w44414, w44415, w44416, w44417, w44418, w44419, w44420, w44421, w44422, w44423, w44424, w44425, w44426, w44427, w44428, w44429, w44430, w44431, w44432, w44433, w44434, w44435, w44436, w44437, w44438, w44439, w44440, w44441, w44442, w44443, w44444, w44445, w44446, w44447, w44448, w44449, w44450, w44451, w44452, w44453, w44454, w44455, w44456, w44457, w44458, w44459, w44460, w44461, w44462, w44463, w44464, w44465, w44466, w44467, w44468, w44469, w44470, w44471, w44472, w44473, w44474, w44475, w44476, w44477, w44478, w44479, w44480, w44481, w44482, w44483, w44484, w44485, w44486, w44487, w44488, w44489, w44490, w44491, w44492, w44493, w44494, w44495, w44496, w44497, w44498, w44499, w44500, w44501, w44502, w44503, w44504, w44505, w44506, w44507, w44508, w44509, w44510, w44511, w44512, w44513, w44514, w44515, w44516, w44517, w44518, w44519, w44520, w44521, w44522, w44523, w44524, w44525, w44526, w44527, w44528, w44529, w44530, w44531, w44532, w44533, w44534, w44535, w44536, w44537, w44538, w44539, w44540, w44541, w44542, w44543, w44544, w44545, w44546, w44547, w44548, w44549, w44550, w44551, w44552, w44553, w44554, w44555, w44556, w44557, w44558, w44559, w44560, w44561, w44562, w44563, w44564, w44565, w44566, w44567, w44568, w44569, w44570, w44571, w44572, w44573, w44574, w44575, w44576, w44577, w44578, w44579, w44580, w44581, w44582, w44583, w44584, w44585, w44586, w44587, w44588, w44589, w44590, w44591, w44592, w44593, w44594, w44595, w44596, w44597, w44598, w44599, w44600, w44601, w44602, w44603, w44604, w44605, w44606, w44607, w44608, w44609, w44610, w44611, w44612, w44613, w44614, w44615, w44616, w44617, w44618, w44619, w44620, w44621, w44622, w44623, w44624, w44625, w44626, w44627, w44628, w44629, w44630, w44631, w44632, w44633, w44634, w44635, w44636, w44637, w44638, w44639, w44640, w44641, w44642, w44643, w44644, w44645, w44646, w44647, w44648, w44649, w44650, w44651, w44652, w44653, w44654, w44655, w44656, w44657, w44658, w44659, w44660, w44661, w44662, w44663, w44664, w44665, w44666, w44667, w44668, w44669, w44670, w44671, w44672, w44673, w44674, w44675, w44676, w44677, w44678, w44679, w44680, w44681, w44682, w44683, w44684, w44685, w44686, w44687, w44688, w44689, w44690, w44691, w44692, w44693, w44694, w44695, w44696, w44697, w44698, w44699, w44700, w44701, w44702, w44703, w44704, w44705, w44706, w44707, w44708, w44709, w44710, w44711, w44712, w44713, w44714, w44715, w44716, w44717, w44718, w44719, w44720, w44721, w44722, w44723, w44724, w44725, w44726, w44727, w44728, w44729, w44730, w44731, w44732, w44733, w44734, w44735, w44736, w44737, w44738, w44739, w44740, w44741, w44742, w44743, w44744, w44745, w44746, w44747, w44748, w44749, w44750, w44751, w44752, w44753, w44754, w44755, w44756, w44757, w44758, w44759, w44760, w44761, w44762, w44763, w44764, w44765, w44766, w44767, w44768, w44769, w44770, w44771, w44772, w44773, w44774, w44775, w44776, w44777, w44778, w44779, w44780, w44781, w44782, w44783, w44784, w44785, w44786, w44787, w44788, w44789, w44790, w44791, w44792, w44793, w44794, w44795, w44796, w44797, w44798, w44799, w44800, w44801, w44802, w44803, w44804, w44805, w44806, w44807, w44808, w44809, w44810, w44811, w44812, w44813, w44814, w44815, w44816, w44817, w44818, w44819, w44820, w44821, w44822, w44823, w44824, w44825, w44826, w44827, w44828, w44829, w44830, w44831, w44832, w44833, w44834, w44835, w44836, w44837, w44838, w44839, w44840, w44841, w44842, w44843, w44844, w44845, w44846, w44847, w44848, w44849, w44850, w44851, w44852, w44853, w44854, w44855, w44856, w44857, w44858, w44859, w44860, w44861, w44862, w44863, w44864, w44865, w44866, w44867, w44868, w44869, w44870, w44871, w44872, w44873, w44874, w44875, w44876, w44877, w44878, w44879, w44880, w44881, w44882, w44883, w44884, w44885, w44886, w44887, w44888, w44889, w44890, w44891, w44892, w44893, w44894, w44895, w44896, w44897, w44898, w44899, w44900, w44901, w44902, w44903, w44904, w44905, w44906, w44907, w44908, w44909, w44910, w44911, w44912, w44913, w44914, w44915, w44916, w44917, w44918, w44919, w44920, w44921, w44922, w44923, w44924, w44925, w44926, w44927, w44928, w44929, w44930, w44931, w44932, w44933, w44934, w44935, w44936, w44937, w44938, w44939, w44940, w44941, w44942, w44943, w44944, w44945, w44946, w44947, w44948, w44949, w44950, w44951, w44952, w44953, w44954, w44955, w44956, w44957, w44958, w44959, w44960, w44961, w44962, w44963, w44964, w44965, w44966, w44967, w44968, w44969, w44970, w44971, w44972, w44973, w44974, w44975, w44976, w44977, w44978, w44979, w44980, w44981, w44982, w44983, w44984, w44985, w44986, w44987, w44988, w44989, w44990, w44991, w44992, w44993, w44994, w44995, w44996, w44997, w44998, w44999, w45000, w45001, w45002, w45003, w45004, w45005, w45006, w45007, w45008, w45009, w45010, w45011, w45012, w45013, w45014, w45015, w45016, w45017, w45018, w45019, w45020, w45021, w45022, w45023, w45024, w45025, w45026, w45027, w45028, w45029, w45030, w45031, w45032, w45033, w45034, w45035, w45036, w45037, w45038, w45039, w45040, w45041, w45042, w45043, w45044, w45045, w45046, w45047, w45048, w45049, w45050, w45051, w45052, w45053, w45054, w45055, w45056, w45057, w45058, w45059, w45060, w45061, w45062, w45063, w45064, w45065, w45066, w45067, w45068, w45069, w45070, w45071, w45072, w45073, w45074, w45075, w45076, w45077, w45078, w45079, w45080, w45081, w45082, w45083, w45084, w45085, w45086, w45087, w45088, w45089, w45090, w45091, w45092, w45093, w45094, w45095, w45096, w45097, w45098, w45099, w45100, w45101, w45102, w45103, w45104, w45105, w45106, w45107, w45108, w45109, w45110, w45111, w45112, w45113, w45114, w45115, w45116, w45117, w45118, w45119, w45120, w45121, w45122, w45123, w45124, w45125, w45126, w45127, w45128, w45129, w45130, w45131, w45132, w45133, w45134, w45135, w45136, w45137, w45138, w45139, w45140, w45141, w45142, w45143, w45144, w45145, w45146, w45147, w45148, w45149, w45150, w45151, w45152, w45153, w45154, w45155, w45156, w45157, w45158, w45159, w45160, w45161, w45162, w45163, w45164, w45165, w45166, w45167, w45168, w45169, w45170, w45171, w45172, w45173, w45174, w45175, w45176, w45177, w45178, w45179, w45180, w45181, w45182, w45183, w45184, w45185, w45186, w45187, w45188, w45189, w45190, w45191, w45192, w45193, w45194, w45195, w45196, w45197, w45198, w45199, w45200, w45201, w45202, w45203, w45204, w45205, w45206, w45207, w45208, w45209, w45210, w45211, w45212, w45213, w45214, w45215, w45216, w45217, w45218, w45219, w45220, w45221, w45222, w45223, w45224, w45225, w45226, w45227, w45228, w45229, w45230, w45231, w45232, w45233, w45234, w45235, w45236, w45237, w45238, w45239, w45240, w45241, w45242, w45243, w45244, w45245, w45246, w45247, w45248, w45249, w45250, w45251, w45252, w45253, w45254, w45255, w45256, w45257, w45258, w45259, w45260, w45261, w45262, w45263, w45264, w45265, w45266, w45267, w45268, w45269, w45270, w45271, w45272, w45273, w45274, w45275, w45276, w45277, w45278, w45279, w45280, w45281, w45282, w45283, w45284, w45285, w45286, w45287, w45288, w45289, w45290, w45291, w45292, w45293, w45294, w45295, w45296, w45297, w45298, w45299, w45300, w45301, w45302, w45303, w45304, w45305, w45306, w45307, w45308, w45309, w45310, w45311, w45312, w45313, w45314, w45315, w45316, w45317, w45318, w45319, w45320, w45321, w45322, w45323, w45324, w45325, w45326, w45327, w45328, w45329, w45330, w45331, w45332, w45333, w45334, w45335, w45336, w45337, w45338, w45339, w45340, w45341, w45342, w45343, w45344, w45345, w45346, w45347, w45348, w45349, w45350, w45351, w45352, w45353, w45354, w45355, w45356, w45357, w45358, w45359, w45360, w45361, w45362, w45363, w45364, w45365, w45366, w45367, w45368, w45369, w45370, w45371, w45372, w45373, w45374, w45375, w45376, w45377, w45378, w45379, w45380, w45381, w45382, w45383, w45384, w45385, w45386, w45387, w45388, w45389, w45390, w45391, w45392, w45393, w45394, w45395, w45396, w45397, w45398, w45399, w45400, w45401, w45402, w45403, w45404, w45405, w45406, w45407, w45408, w45409, w45410, w45411, w45412, w45413, w45414, w45415, w45416, w45417, w45418, w45419, w45420, w45421, w45422, w45423, w45424, w45425, w45426, w45427, w45428, w45429, w45430, w45431, w45432, w45433, w45434, w45435, w45436, w45437, w45438, w45439, w45440, w45441, w45442, w45443, w45444, w45445, w45446, w45447, w45448, w45449, w45450, w45451, w45452, w45453, w45454, w45455, w45456, w45457, w45458, w45459, w45460, w45461, w45462, w45463, w45464, w45465, w45466, w45467, w45468, w45469, w45470, w45471, w45472, w45473, w45474, w45475, w45476, w45477, w45478, w45479, w45480, w45481, w45482, w45483, w45484, w45485, w45486, w45487, w45488, w45489, w45490, w45491, w45492, w45493, w45494, w45495, w45496, w45497, w45498, w45499, w45500, w45501, w45502, w45503, w45504, w45505, w45506, w45507, w45508, w45509, w45510, w45511, w45512, w45513, w45514, w45515, w45516, w45517, w45518, w45519, w45520, w45521, w45522, w45523, w45524, w45525, w45526, w45527, w45528, w45529, w45530, w45531, w45532, w45533, w45534, w45535, w45536, w45537, w45538, w45539, w45540, w45541, w45542, w45543, w45544, w45545, w45546, w45547, w45548, w45549, w45550, w45551, w45552, w45553, w45554, w45555, w45556, w45557, w45558, w45559, w45560, w45561, w45562, w45563, w45564, w45565, w45566, w45567, w45568, w45569, w45570, w45571, w45572, w45573, w45574, w45575, w45576, w45577, w45578, w45579, w45580, w45581, w45582, w45583, w45584, w45585, w45586, w45587, w45588, w45589, w45590, w45591, w45592, w45593, w45594, w45595, w45596, w45597, w45598, w45599, w45600, w45601, w45602, w45603, w45604, w45605, w45606, w45607, w45608, w45609, w45610, w45611, w45612, w45613, w45614, w45615, w45616, w45617, w45618, w45619, w45620, w45621, w45622, w45623, w45624, w45625, w45626, w45627, w45628, w45629, w45630, w45631, w45632, w45633, w45634, w45635, w45636, w45637, w45638, w45639, w45640, w45641, w45642, w45643, w45644, w45645, w45646, w45647, w45648, w45649, w45650, w45651, w45652, w45653, w45654, w45655, w45656, w45657, w45658, w45659, w45660, w45661, w45662, w45663, w45664, w45665, w45666, w45667, w45668, w45669, w45670, w45671, w45672, w45673, w45674, w45675, w45676, w45677, w45678, w45679, w45680, w45681, w45682, w45683, w45684, w45685, w45686, w45687, w45688, w45689, w45690, w45691, w45692, w45693, w45694, w45695, w45696, w45697, w45698, w45699, w45700, w45701, w45702, w45703, w45704, w45705, w45706, w45707, w45708, w45709, w45710, w45711, w45712, w45713, w45714, w45715, w45716, w45717, w45718, w45719, w45720, w45721, w45722, w45723, w45724, w45725, w45726, w45727, w45728, w45729, w45730, w45731, w45732, w45733, w45734, w45735, w45736, w45737, w45738, w45739, w45740, w45741, w45742, w45743, w45744, w45745, w45746, w45747, w45748, w45749, w45750, w45751, w45752, w45753, w45754, w45755, w45756, w45757, w45758, w45759, w45760, w45761, w45762, w45763, w45764, w45765, w45766, w45767, w45768, w45769, w45770, w45771, w45772, w45773, w45774, w45775, w45776, w45777, w45778, w45779, w45780, w45781, w45782, w45783, w45784, w45785, w45786, w45787, w45788, w45789, w45790, w45791, w45792, w45793, w45794, w45795, w45796, w45797, w45798, w45799, w45800, w45801, w45802, w45803, w45804, w45805, w45806, w45807, w45808, w45809, w45810, w45811, w45812, w45813, w45814, w45815, w45816, w45817, w45818, w45819, w45820, w45821, w45822, w45823, w45824, w45825, w45826, w45827, w45828, w45829, w45830, w45831, w45832, w45833, w45834, w45835, w45836, w45837, w45838, w45839, w45840, w45841, w45842, w45843, w45844, w45845, w45846, w45847, w45848, w45849, w45850, w45851, w45852, w45853, w45854, w45855, w45856, w45857, w45858, w45859, w45860, w45861, w45862, w45863, w45864, w45865, w45866, w45867, w45868, w45869, w45870, w45871, w45872, w45873, w45874, w45875, w45876, w45877, w45878, w45879, w45880, w45881, w45882, w45883, w45884, w45885, w45886, w45887, w45888, w45889, w45890, w45891, w45892, w45893, w45894, w45895, w45896, w45897, w45898, w45899, w45900, w45901, w45902, w45903, w45904, w45905, w45906, w45907, w45908, w45909, w45910, w45911, w45912, w45913, w45914, w45915, w45916, w45917, w45918, w45919, w45920, w45921, w45922, w45923, w45924, w45925, w45926, w45927, w45928, w45929, w45930, w45931, w45932, w45933, w45934, w45935, w45936, w45937, w45938, w45939, w45940, w45941, w45942, w45943, w45944, w45945, w45946, w45947, w45948, w45949, w45950, w45951, w45952, w45953, w45954, w45955, w45956, w45957, w45958, w45959, w45960, w45961, w45962, w45963, w45964, w45965, w45966, w45967, w45968, w45969, w45970, w45971, w45972, w45973, w45974, w45975, w45976, w45977, w45978, w45979, w45980, w45981, w45982, w45983, w45984, w45985, w45986, w45987, w45988, w45989, w45990, w45991, w45992, w45993, w45994, w45995, w45996, w45997, w45998, w45999, w46000, w46001, w46002, w46003, w46004, w46005, w46006, w46007, w46008, w46009, w46010, w46011, w46012, w46013, w46014, w46015, w46016, w46017, w46018, w46019, w46020, w46021, w46022, w46023, w46024, w46025, w46026, w46027, w46028, w46029, w46030, w46031, w46032, w46033, w46034, w46035, w46036, w46037, w46038, w46039, w46040, w46041, w46042, w46043, w46044, w46045, w46046, w46047, w46048, w46049, w46050, w46051, w46052, w46053, w46054, w46055, w46056, w46057, w46058, w46059, w46060, w46061, w46062, w46063, w46064, w46065, w46066, w46067, w46068, w46069, w46070, w46071, w46072, w46073, w46074, w46075, w46076, w46077, w46078, w46079, w46080, w46081, w46082, w46083, w46084, w46085, w46086, w46087, w46088, w46089, w46090, w46091, w46092, w46093, w46094, w46095, w46096, w46097, w46098, w46099, w46100, w46101, w46102, w46103, w46104, w46105, w46106, w46107, w46108, w46109, w46110, w46111, w46112, w46113, w46114, w46115, w46116, w46117, w46118, w46119, w46120, w46121, w46122, w46123, w46124, w46125, w46126, w46127, w46128, w46129, w46130, w46131, w46132, w46133, w46134, w46135, w46136, w46137, w46138, w46139, w46140, w46141, w46142, w46143, w46144, w46145, w46146, w46147, w46148, w46149, w46150, w46151, w46152, w46153, w46154, w46155, w46156, w46157, w46158, w46159, w46160, w46161, w46162, w46163, w46164, w46165, w46166, w46167, w46168, w46169, w46170, w46171, w46172, w46173, w46174, w46175, w46176, w46177, w46178, w46179, w46180, w46181, w46182, w46183, w46184, w46185, w46186, w46187, w46188, w46189, w46190, w46191, w46192, w46193, w46194, w46195, w46196, w46197, w46198, w46199, w46200, w46201, w46202, w46203, w46204, w46205, w46206, w46207, w46208, w46209, w46210, w46211, w46212, w46213, w46214, w46215, w46216, w46217, w46218, w46219, w46220, w46221, w46222, w46223, w46224, w46225, w46226, w46227, w46228, w46229, w46230, w46231, w46232, w46233, w46234, w46235, w46236, w46237, w46238, w46239, w46240, w46241, w46242, w46243, w46244, w46245, w46246, w46247, w46248, w46249, w46250, w46251, w46252, w46253, w46254, w46255, w46256, w46257, w46258, w46259, w46260, w46261, w46262, w46263, w46264, w46265, w46266, w46267, w46268, w46269, w46270, w46271, w46272, w46273, w46274, w46275, w46276, w46277, w46278, w46279, w46280, w46281, w46282, w46283, w46284, w46285, w46286, w46287, w46288, w46289, w46290, w46291, w46292, w46293, w46294, w46295, w46296, w46297, w46298, w46299, w46300, w46301, w46302, w46303, w46304, w46305, w46306, w46307, w46308, w46309, w46310, w46311, w46312, w46313, w46314, w46315, w46316, w46317, w46318, w46319, w46320, w46321, w46322, w46323, w46324, w46325, w46326, w46327, w46328, w46329, w46330, w46331, w46332, w46333, w46334, w46335, w46336, w46337, w46338, w46339, w46340, w46341, w46342, w46343, w46344, w46345, w46346, w46347, w46348, w46349, w46350, w46351, w46352, w46353, w46354, w46355, w46356, w46357, w46358, w46359, w46360, w46361, w46362, w46363, w46364, w46365, w46366, w46367, w46368, w46369, w46370, w46371, w46372, w46373, w46374, w46375, w46376, w46377, w46378, w46379, w46380, w46381, w46382, w46383, w46384, w46385, w46386, w46387, w46388, w46389, w46390, w46391, w46392, w46393, w46394, w46395, w46396, w46397, w46398, w46399, w46400, w46401, w46402, w46403, w46404, w46405, w46406, w46407, w46408, w46409, w46410, w46411, w46412, w46413, w46414, w46415, w46416, w46417, w46418, w46419, w46420, w46421, w46422, w46423, w46424, w46425, w46426, w46427, w46428, w46429, w46430, w46431, w46432, w46433, w46434, w46435, w46436, w46437, w46438, w46439, w46440, w46441, w46442, w46443, w46444, w46445, w46446, w46447, w46448, w46449, w46450, w46451, w46452, w46453, w46454, w46455, w46456, w46457, w46458, w46459, w46460, w46461, w46462, w46463, w46464, w46465, w46466, w46467, w46468, w46469, w46470, w46471, w46472, w46473, w46474, w46475, w46476, w46477, w46478, w46479, w46480, w46481, w46482, w46483, w46484, w46485, w46486, w46487, w46488, w46489, w46490, w46491, w46492, w46493, w46494, w46495, w46496, w46497, w46498, w46499, w46500, w46501, w46502, w46503, w46504, w46505, w46506, w46507, w46508, w46509, w46510, w46511, w46512, w46513, w46514, w46515, w46516, w46517, w46518, w46519, w46520, w46521, w46522, w46523, w46524, w46525, w46526, w46527, w46528, w46529, w46530, w46531, w46532, w46533, w46534, w46535, w46536, w46537, w46538, w46539, w46540, w46541, w46542, w46543, w46544, w46545, w46546, w46547, w46548, w46549, w46550, w46551, w46552, w46553, w46554, w46555, w46556, w46557, w46558, w46559, w46560, w46561, w46562, w46563, w46564, w46565, w46566, w46567, w46568, w46569, w46570, w46571, w46572, w46573, w46574, w46575, w46576, w46577, w46578, w46579, w46580, w46581, w46582, w46583, w46584, w46585, w46586, w46587, w46588, w46589, w46590, w46591, w46592, w46593, w46594, w46595, w46596, w46597, w46598, w46599, w46600, w46601, w46602, w46603, w46604, w46605, w46606, w46607, w46608, w46609, w46610, w46611, w46612, w46613, w46614, w46615, w46616, w46617, w46618, w46619, w46620, w46621, w46622, w46623, w46624, w46625, w46626, w46627, w46628, w46629, w46630, w46631, w46632, w46633, w46634, w46635, w46636, w46637, w46638, w46639, w46640, w46641, w46642, w46643, w46644, w46645, w46646, w46647, w46648, w46649, w46650, w46651, w46652, w46653, w46654, w46655, w46656, w46657, w46658, w46659, w46660, w46661, w46662, w46663, w46664, w46665, w46666, w46667, w46668, w46669, w46670, w46671, w46672, w46673, w46674, w46675, w46676, w46677, w46678, w46679, w46680, w46681, w46682, w46683, w46684, w46685, w46686, w46687, w46688, w46689, w46690, w46691, w46692, w46693, w46694, w46695, w46696, w46697, w46698, w46699, w46700, w46701, w46702, w46703, w46704, w46705, w46706, w46707, w46708, w46709, w46710, w46711, w46712, w46713, w46714, w46715, w46716, w46717, w46718, w46719, w46720, w46721, w46722, w46723, w46724, w46725, w46726, w46727, w46728, w46729, w46730, w46731, w46732, w46733, w46734, w46735, w46736, w46737, w46738, w46739, w46740, w46741, w46742, w46743, w46744, w46745, w46746, w46747, w46748, w46749, w46750, w46751, w46752, w46753, w46754, w46755, w46756, w46757, w46758, w46759, w46760, w46761, w46762, w46763, w46764, w46765, w46766, w46767, w46768, w46769, w46770, w46771, w46772, w46773, w46774, w46775, w46776, w46777, w46778, w46779, w46780, w46781, w46782, w46783, w46784, w46785, w46786, w46787, w46788, w46789, w46790, w46791, w46792, w46793, w46794, w46795, w46796, w46797, w46798, w46799, w46800, w46801, w46802, w46803, w46804, w46805, w46806, w46807, w46808, w46809, w46810, w46811, w46812, w46813, w46814, w46815, w46816, w46817, w46818, w46819, w46820, w46821, w46822, w46823, w46824, w46825, w46826, w46827, w46828, w46829, w46830, w46831, w46832, w46833, w46834, w46835, w46836, w46837, w46838, w46839, w46840, w46841, w46842, w46843, w46844, w46845, w46846, w46847, w46848, w46849, w46850, w46851, w46852, w46853, w46854, w46855, w46856, w46857, w46858, w46859, w46860, w46861, w46862, w46863, w46864, w46865, w46866, w46867, w46868, w46869, w46870, w46871, w46872, w46873, w46874, w46875, w46876, w46877, w46878, w46879, w46880, w46881, w46882, w46883, w46884, w46885, w46886, w46887, w46888, w46889, w46890, w46891, w46892, w46893, w46894, w46895, w46896, w46897, w46898, w46899, w46900, w46901, w46902, w46903, w46904, w46905, w46906, w46907, w46908, w46909, w46910, w46911, w46912, w46913, w46914, w46915, w46916, w46917, w46918, w46919, w46920, w46921, w46922, w46923, w46924, w46925, w46926, w46927, w46928, w46929, w46930, w46931, w46932, w46933, w46934, w46935, w46936, w46937, w46938, w46939, w46940, w46941, w46942, w46943, w46944, w46945, w46946, w46947, w46948, w46949, w46950, w46951, w46952, w46953, w46954, w46955, w46956, w46957, w46958, w46959, w46960, w46961, w46962, w46963, w46964, w46965, w46966, w46967, w46968, w46969, w46970, w46971, w46972, w46973, w46974, w46975, w46976, w46977, w46978, w46979, w46980, w46981, w46982, w46983, w46984, w46985, w46986, w46987, w46988, w46989, w46990, w46991, w46992, w46993, w46994, w46995, w46996, w46997, w46998, w46999, w47000, w47001, w47002, w47003, w47004, w47005, w47006, w47007, w47008, w47009, w47010, w47011, w47012, w47013, w47014, w47015, w47016, w47017, w47018, w47019, w47020, w47021, w47022, w47023, w47024, w47025, w47026, w47027, w47028, w47029, w47030, w47031, w47032, w47033, w47034, w47035, w47036, w47037, w47038, w47039, w47040, w47041, w47042, w47043, w47044, w47045, w47046, w47047, w47048, w47049, w47050, w47051, w47052, w47053, w47054, w47055, w47056, w47057, w47058, w47059, w47060, w47061, w47062, w47063, w47064, w47065, w47066, w47067, w47068, w47069, w47070, w47071, w47072, w47073, w47074, w47075, w47076, w47077, w47078, w47079, w47080, w47081, w47082, w47083, w47084, w47085, w47086, w47087, w47088, w47089, w47090, w47091, w47092, w47093, w47094, w47095, w47096, w47097, w47098, w47099, w47100, w47101, w47102, w47103, w47104, w47105, w47106, w47107, w47108, w47109, w47110, w47111, w47112, w47113, w47114, w47115, w47116, w47117, w47118, w47119, w47120, w47121, w47122, w47123, w47124, w47125, w47126, w47127, w47128, w47129, w47130, w47131, w47132, w47133, w47134, w47135, w47136, w47137, w47138, w47139, w47140, w47141, w47142, w47143, w47144, w47145, w47146, w47147, w47148, w47149, w47150, w47151, w47152, w47153, w47154, w47155, w47156, w47157, w47158, w47159, w47160, w47161, w47162, w47163, w47164, w47165, w47166, w47167, w47168, w47169, w47170, w47171, w47172, w47173, w47174, w47175, w47176, w47177, w47178, w47179, w47180, w47181, w47182, w47183, w47184, w47185, w47186, w47187, w47188, w47189, w47190, w47191, w47192, w47193, w47194, w47195, w47196, w47197, w47198, w47199, w47200, w47201, w47202, w47203, w47204, w47205, w47206, w47207, w47208, w47209, w47210, w47211, w47212, w47213, w47214, w47215, w47216, w47217, w47218, w47219, w47220, w47221, w47222, w47223, w47224, w47225, w47226, w47227, w47228, w47229, w47230, w47231, w47232, w47233, w47234, w47235, w47236, w47237, w47238, w47239, w47240, w47241, w47242, w47243, w47244, w47245, w47246, w47247, w47248, w47249, w47250, w47251, w47252, w47253, w47254, w47255, w47256, w47257, w47258, w47259, w47260, w47261, w47262, w47263, w47264, w47265, w47266, w47267, w47268, w47269, w47270, w47271, w47272, w47273, w47274, w47275, w47276, w47277, w47278, w47279, w47280, w47281, w47282, w47283, w47284, w47285, w47286, w47287, w47288, w47289, w47290, w47291, w47292, w47293, w47294, w47295, w47296, w47297, w47298, w47299, w47300, w47301, w47302, w47303, w47304, w47305, w47306, w47307, w47308, w47309, w47310, w47311, w47312, w47313, w47314, w47315, w47316, w47317, w47318, w47319, w47320, w47321, w47322, w47323, w47324, w47325, w47326, w47327, w47328, w47329, w47330, w47331, w47332, w47333, w47334, w47335, w47336, w47337, w47338, w47339, w47340, w47341, w47342, w47343, w47344, w47345, w47346, w47347, w47348, w47349, w47350, w47351, w47352, w47353, w47354, w47355, w47356, w47357, w47358, w47359, w47360, w47361, w47362, w47363, w47364, w47365, w47366, w47367, w47368, w47369, w47370, w47371, w47372, w47373, w47374, w47375, w47376, w47377, w47378, w47379, w47380, w47381, w47382, w47383, w47384, w47385, w47386, w47387, w47388, w47389, w47390, w47391, w47392, w47393, w47394, w47395, w47396, w47397, w47398, w47399, w47400, w47401, w47402, w47403, w47404, w47405, w47406, w47407, w47408, w47409, w47410, w47411, w47412, w47413, w47414, w47415, w47416, w47417, w47418, w47419, w47420, w47421, w47422, w47423, w47424, w47425, w47426, w47427, w47428, w47429, w47430, w47431, w47432, w47433, w47434, w47435, w47436, w47437, w47438, w47439, w47440, w47441, w47442, w47443, w47444, w47445, w47446, w47447, w47448, w47449, w47450, w47451, w47452, w47453, w47454, w47455, w47456, w47457, w47458, w47459, w47460, w47461, w47462, w47463, w47464, w47465, w47466, w47467, w47468, w47469, w47470, w47471, w47472, w47473, w47474, w47475, w47476, w47477, w47478, w47479, w47480, w47481, w47482, w47483, w47484, w47485, w47486, w47487, w47488, w47489, w47490, w47491, w47492, w47493, w47494, w47495, w47496, w47497, w47498, w47499, w47500, w47501, w47502, w47503, w47504, w47505, w47506, w47507, w47508, w47509, w47510, w47511, w47512, w47513, w47514, w47515, w47516, w47517, w47518, w47519, w47520, w47521, w47522, w47523, w47524, w47525, w47526, w47527, w47528, w47529, w47530, w47531, w47532, w47533, w47534, w47535, w47536, w47537, w47538, w47539, w47540, w47541, w47542, w47543, w47544, w47545, w47546, w47547, w47548, w47549, w47550, w47551, w47552, w47553, w47554, w47555, w47556, w47557, w47558, w47559, w47560, w47561, w47562, w47563, w47564, w47565, w47566, w47567, w47568, w47569, w47570, w47571, w47572, w47573, w47574, w47575, w47576, w47577, w47578, w47579, w47580, w47581, w47582, w47583, w47584, w47585, w47586, w47587, w47588, w47589, w47590, w47591, w47592, w47593, w47594, w47595, w47596, w47597, w47598, w47599, w47600, w47601, w47602, w47603, w47604, w47605, w47606, w47607, w47608, w47609, w47610, w47611, w47612, w47613, w47614, w47615, w47616, w47617, w47618, w47619, w47620, w47621, w47622, w47623, w47624, w47625, w47626, w47627, w47628, w47629, w47630, w47631, w47632, w47633, w47634, w47635, w47636, w47637, w47638, w47639, w47640, w47641, w47642, w47643, w47644, w47645, w47646, w47647, w47648, w47649, w47650, w47651, w47652, w47653, w47654, w47655, w47656, w47657, w47658, w47659, w47660, w47661, w47662, w47663, w47664, w47665, w47666, w47667, w47668, w47669, w47670, w47671, w47672, w47673, w47674, w47675, w47676, w47677, w47678, w47679, w47680, w47681, w47682, w47683, w47684, w47685, w47686, w47687, w47688, w47689, w47690, w47691, w47692, w47693, w47694, w47695, w47696, w47697, w47698, w47699, w47700, w47701, w47702, w47703, w47704, w47705, w47706, w47707, w47708, w47709, w47710, w47711, w47712, w47713, w47714, w47715, w47716, w47717, w47718, w47719, w47720, w47721, w47722, w47723, w47724, w47725, w47726, w47727, w47728, w47729, w47730, w47731, w47732, w47733, w47734, w47735, w47736, w47737, w47738, w47739, w47740, w47741, w47742, w47743, w47744, w47745, w47746, w47747, w47748, w47749, w47750, w47751, w47752, w47753, w47754, w47755, w47756, w47757, w47758, w47759, w47760, w47761, w47762, w47763, w47764, w47765, w47766, w47767, w47768, w47769, w47770, w47771, w47772, w47773, w47774, w47775, w47776, w47777, w47778, w47779, w47780, w47781, w47782, w47783, w47784, w47785, w47786, w47787, w47788, w47789, w47790, w47791, w47792, w47793, w47794, w47795, w47796, w47797, w47798, w47799, w47800, w47801, w47802, w47803, w47804, w47805, w47806, w47807, w47808, w47809, w47810, w47811, w47812, w47813, w47814, w47815, w47816, w47817, w47818, w47819, w47820, w47821, w47822, w47823, w47824, w47825, w47826, w47827, w47828, w47829, w47830, w47831, w47832, w47833, w47834, w47835, w47836, w47837, w47838, w47839, w47840, w47841, w47842, w47843, w47844, w47845, w47846, w47847, w47848, w47849, w47850, w47851, w47852, w47853, w47854, w47855, w47856, w47857, w47858, w47859, w47860, w47861, w47862, w47863, w47864, w47865, w47866, w47867, w47868, w47869, w47870, w47871, w47872, w47873, w47874, w47875, w47876, w47877, w47878, w47879, w47880, w47881, w47882, w47883, w47884, w47885, w47886, w47887, w47888, w47889, w47890, w47891, w47892, w47893, w47894, w47895, w47896, w47897, w47898, w47899, w47900, w47901, w47902, w47903, w47904, w47905, w47906, w47907, w47908, w47909, w47910, w47911, w47912, w47913, w47914, w47915, w47916, w47917, w47918, w47919, w47920, w47921, w47922, w47923, w47924, w47925, w47926, w47927, w47928, w47929, w47930, w47931, w47932, w47933, w47934, w47935, w47936, w47937, w47938, w47939, w47940, w47941, w47942, w47943, w47944, w47945, w47946, w47947, w47948, w47949, w47950, w47951, w47952, w47953, w47954, w47955, w47956, w47957, w47958, w47959, w47960, w47961, w47962, w47963, w47964, w47965, w47966, w47967, w47968, w47969, w47970, w47971, w47972, w47973, w47974, w47975, w47976, w47977, w47978, w47979, w47980, w47981, w47982, w47983, w47984, w47985, w47986, w47987, w47988, w47989, w47990, w47991, w47992, w47993, w47994, w47995, w47996, w47997, w47998, w47999, w48000, w48001, w48002, w48003, w48004, w48005, w48006, w48007, w48008, w48009, w48010, w48011, w48012, w48013, w48014, w48015, w48016, w48017, w48018, w48019, w48020, w48021, w48022, w48023, w48024, w48025, w48026, w48027, w48028, w48029, w48030, w48031, w48032, w48033, w48034, w48035, w48036, w48037, w48038, w48039, w48040, w48041, w48042, w48043, w48044, w48045, w48046, w48047, w48048, w48049, w48050, w48051, w48052, w48053, w48054, w48055, w48056, w48057, w48058, w48059, w48060, w48061, w48062, w48063, w48064, w48065, w48066, w48067, w48068, w48069, w48070, w48071, w48072, w48073, w48074, w48075, w48076, w48077, w48078, w48079, w48080, w48081, w48082, w48083, w48084, w48085, w48086, w48087, w48088, w48089, w48090, w48091, w48092, w48093, w48094, w48095, w48096, w48097, w48098, w48099, w48100, w48101, w48102, w48103, w48104, w48105, w48106, w48107, w48108, w48109, w48110, w48111, w48112, w48113, w48114, w48115, w48116, w48117, w48118, w48119, w48120, w48121, w48122, w48123, w48124, w48125, w48126, w48127, w48128, w48129, w48130, w48131, w48132, w48133, w48134, w48135, w48136, w48137, w48138, w48139, w48140, w48141, w48142, w48143, w48144, w48145, w48146, w48147, w48148, w48149, w48150, w48151, w48152, w48153, w48154, w48155, w48156, w48157, w48158, w48159, w48160, w48161, w48162, w48163, w48164, w48165, w48166, w48167, w48168, w48169, w48170, w48171, w48172, w48173, w48174, w48175, w48176, w48177, w48178, w48179, w48180, w48181, w48182, w48183, w48184, w48185, w48186, w48187, w48188, w48189, w48190, w48191, w48192, w48193, w48194, w48195, w48196, w48197, w48198, w48199, w48200, w48201, w48202, w48203, w48204, w48205, w48206, w48207, w48208, w48209, w48210, w48211, w48212, w48213, w48214, w48215, w48216, w48217, w48218, w48219, w48220, w48221, w48222, w48223, w48224, w48225, w48226, w48227, w48228, w48229, w48230, w48231, w48232, w48233, w48234, w48235, w48236, w48237, w48238, w48239, w48240, w48241, w48242, w48243, w48244, w48245, w48246, w48247, w48248, w48249, w48250, w48251, w48252, w48253, w48254, w48255, w48256, w48257, w48258, w48259, w48260, w48261, w48262, w48263, w48264, w48265, w48266, w48267, w48268, w48269, w48270, w48271, w48272, w48273, w48274, w48275, w48276, w48277, w48278, w48279, w48280, w48281, w48282, w48283, w48284, w48285, w48286, w48287, w48288, w48289, w48290, w48291, w48292, w48293, w48294, w48295, w48296, w48297, w48298, w48299, w48300, w48301, w48302, w48303, w48304, w48305, w48306, w48307, w48308, w48309, w48310, w48311, w48312, w48313, w48314, w48315, w48316, w48317, w48318, w48319, w48320, w48321, w48322, w48323, w48324, w48325, w48326, w48327, w48328, w48329, w48330, w48331, w48332, w48333, w48334, w48335, w48336, w48337, w48338, w48339, w48340, w48341, w48342, w48343, w48344, w48345, w48346, w48347, w48348, w48349, w48350, w48351, w48352, w48353, w48354, w48355, w48356, w48357, w48358, w48359, w48360, w48361, w48362, w48363, w48364, w48365, w48366, w48367, w48368, w48369, w48370, w48371, w48372, w48373, w48374, w48375, w48376, w48377, w48378, w48379, w48380, w48381, w48382, w48383, w48384, w48385, w48386, w48387, w48388, w48389, w48390, w48391, w48392, w48393, w48394, w48395, w48396, w48397, w48398, w48399, w48400, w48401, w48402, w48403, w48404, w48405, w48406, w48407, w48408, w48409, w48410, w48411, w48412, w48413, w48414, w48415, w48416, w48417, w48418, w48419, w48420, w48421, w48422, w48423, w48424, w48425, w48426, w48427, w48428, w48429, w48430, w48431, w48432, w48433, w48434, w48435, w48436, w48437, w48438, w48439, w48440, w48441, w48442, w48443, w48444, w48445, w48446, w48447, w48448, w48449, w48450, w48451, w48452, w48453, w48454, w48455, w48456, w48457, w48458, w48459, w48460, w48461, w48462, w48463, w48464, w48465, w48466, w48467, w48468, w48469, w48470, w48471, w48472, w48473, w48474, w48475, w48476, w48477, w48478, w48479, w48480, w48481, w48482, w48483, w48484, w48485, w48486, w48487, w48488, w48489, w48490, w48491, w48492, w48493, w48494, w48495, w48496, w48497, w48498, w48499, w48500, w48501, w48502, w48503, w48504, w48505, w48506, w48507, w48508, w48509, w48510, w48511, w48512, w48513, w48514, w48515, w48516, w48517, w48518, w48519, w48520, w48521, w48522, w48523, w48524, w48525, w48526, w48527, w48528, w48529, w48530, w48531, w48532, w48533, w48534, w48535, w48536, w48537, w48538, w48539, w48540, w48541, w48542, w48543, w48544, w48545, w48546, w48547, w48548, w48549, w48550, w48551, w48552, w48553, w48554, w48555, w48556, w48557, w48558, w48559, w48560, w48561, w48562, w48563, w48564, w48565, w48566, w48567, w48568, w48569, w48570, w48571, w48572, w48573, w48574, w48575, w48576, w48577, w48578, w48579, w48580, w48581, w48582, w48583, w48584, w48585, w48586, w48587, w48588, w48589, w48590, w48591, w48592, w48593, w48594, w48595, w48596, w48597, w48598, w48599, w48600, w48601, w48602, w48603, w48604, w48605, w48606, w48607, w48608, w48609, w48610, w48611, w48612, w48613, w48614, w48615, w48616, w48617, w48618, w48619, w48620, w48621, w48622, w48623, w48624, w48625, w48626, w48627, w48628, w48629, w48630, w48631, w48632, w48633, w48634, w48635, w48636, w48637, w48638, w48639, w48640, w48641, w48642, w48643, w48644, w48645, w48646, w48647, w48648, w48649, w48650, w48651, w48652, w48653, w48654, w48655, w48656, w48657, w48658, w48659, w48660, w48661, w48662, w48663, w48664, w48665, w48666, w48667, w48668, w48669, w48670, w48671, w48672, w48673, w48674, w48675, w48676, w48677, w48678, w48679, w48680, w48681, w48682, w48683, w48684, w48685, w48686, w48687, w48688, w48689, w48690, w48691, w48692, w48693, w48694, w48695, w48696, w48697, w48698, w48699, w48700, w48701, w48702, w48703, w48704, w48705, w48706, w48707, w48708, w48709, w48710, w48711, w48712, w48713, w48714, w48715, w48716, w48717, w48718, w48719, w48720, w48721, w48722, w48723, w48724, w48725, w48726, w48727, w48728, w48729, w48730, w48731, w48732, w48733, w48734, w48735, w48736, w48737, w48738, w48739, w48740, w48741, w48742, w48743, w48744, w48745, w48746, w48747, w48748, w48749, w48750, w48751, w48752, w48753, w48754, w48755, w48756, w48757, w48758, w48759, w48760, w48761, w48762, w48763, w48764, w48765, w48766, w48767, w48768, w48769, w48770, w48771, w48772, w48773, w48774, w48775, w48776, w48777, w48778, w48779, w48780, w48781, w48782, w48783, w48784, w48785, w48786, w48787, w48788, w48789, w48790, w48791, w48792, w48793, w48794, w48795, w48796, w48797, w48798, w48799, w48800, w48801, w48802, w48803, w48804, w48805, w48806, w48807, w48808, w48809, w48810, w48811, w48812, w48813, w48814, w48815, w48816, w48817, w48818, w48819, w48820, w48821, w48822, w48823, w48824, w48825, w48826, w48827, w48828, w48829, w48830, w48831, w48832, w48833, w48834, w48835, w48836, w48837, w48838, w48839, w48840, w48841, w48842, w48843, w48844, w48845, w48846, w48847, w48848, w48849, w48850, w48851, w48852, w48853, w48854, w48855, w48856, w48857, w48858, w48859, w48860, w48861, w48862, w48863, w48864, w48865, w48866, w48867, w48868, w48869, w48870, w48871, w48872, w48873, w48874, w48875, w48876, w48877, w48878, w48879, w48880, w48881, w48882, w48883, w48884, w48885, w48886, w48887, w48888, w48889, w48890, w48891, w48892, w48893, w48894, w48895, w48896, w48897, w48898, w48899, w48900, w48901, w48902, w48903, w48904, w48905, w48906, w48907, w48908, w48909, w48910, w48911, w48912, w48913, w48914, w48915, w48916, w48917, w48918, w48919, w48920, w48921, w48922, w48923, w48924, w48925, w48926, w48927, w48928, w48929, w48930, w48931, w48932, w48933, w48934, w48935, w48936, w48937, w48938, w48939, w48940, w48941, w48942, w48943, w48944, w48945, w48946, w48947, w48948, w48949, w48950, w48951, w48952, w48953, w48954, w48955, w48956, w48957, w48958, w48959, w48960, w48961, w48962, w48963, w48964, w48965, w48966, w48967, w48968, w48969, w48970, w48971, w48972, w48973, w48974, w48975, w48976, w48977, w48978, w48979, w48980, w48981, w48982, w48983, w48984, w48985, w48986, w48987, w48988, w48989, w48990, w48991, w48992, w48993, w48994, w48995, w48996, w48997, w48998, w48999, w49000, w49001, w49002, w49003, w49004, w49005, w49006, w49007, w49008, w49009, w49010, w49011, w49012, w49013, w49014, w49015, w49016, w49017, w49018, w49019, w49020, w49021, w49022, w49023, w49024, w49025, w49026, w49027, w49028, w49029, w49030, w49031, w49032, w49033, w49034, w49035, w49036, w49037, w49038, w49039, w49040, w49041, w49042, w49043, w49044, w49045, w49046, w49047, w49048, w49049, w49050, w49051, w49052, w49053, w49054, w49055, w49056, w49057, w49058, w49059, w49060, w49061, w49062, w49063, w49064, w49065, w49066, w49067, w49068, w49069, w49070, w49071, w49072, w49073, w49074, w49075, w49076, w49077, w49078, w49079, w49080, w49081, w49082, w49083, w49084, w49085, w49086, w49087, w49088, w49089, w49090, w49091, w49092, w49093, w49094, w49095, w49096, w49097, w49098, w49099, w49100, w49101, w49102, w49103, w49104, w49105, w49106, w49107, w49108, w49109, w49110, w49111, w49112, w49113, w49114, w49115, w49116, w49117, w49118, w49119, w49120, w49121, w49122, w49123, w49124, w49125, w49126, w49127, w49128, w49129, w49130, w49131, w49132, w49133, w49134, w49135, w49136, w49137, w49138, w49139, w49140, w49141, w49142, w49143, w49144, w49145, w49146, w49147, w49148, w49149, w49150, w49151, w49152, w49153, w49154, w49155, w49156, w49157, w49158, w49159, w49160, w49161, w49162, w49163, w49164, w49165, w49166, w49167, w49168, w49169, w49170, w49171, w49172, w49173, w49174, w49175, w49176, w49177, w49178, w49179, w49180, w49181, w49182, w49183, w49184, w49185, w49186, w49187, w49188, w49189, w49190, w49191, w49192, w49193, w49194, w49195, w49196, w49197, w49198, w49199, w49200, w49201, w49202, w49203, w49204, w49205, w49206, w49207, w49208, w49209, w49210, w49211, w49212, w49213, w49214, w49215, w49216, w49217, w49218, w49219, w49220, w49221, w49222, w49223, w49224, w49225, w49226, w49227, w49228, w49229, w49230, w49231, w49232, w49233, w49234, w49235, w49236, w49237, w49238, w49239, w49240, w49241, w49242, w49243, w49244, w49245, w49246, w49247, w49248, w49249, w49250, w49251, w49252, w49253, w49254, w49255, w49256, w49257, w49258, w49259, w49260, w49261, w49262, w49263, w49264, w49265, w49266, w49267, w49268, w49269, w49270, w49271, w49272, w49273, w49274, w49275, w49276, w49277, w49278, w49279, w49280, w49281, w49282, w49283, w49284, w49285, w49286, w49287, w49288, w49289, w49290, w49291, w49292, w49293, w49294, w49295, w49296, w49297, w49298, w49299, w49300, w49301, w49302, w49303, w49304, w49305, w49306, w49307, w49308, w49309, w49310, w49311, w49312, w49313, w49314, w49315, w49316, w49317, w49318, w49319, w49320, w49321, w49322, w49323, w49324, w49325, w49326, w49327, w49328, w49329, w49330, w49331, w49332, w49333, w49334, w49335, w49336, w49337, w49338, w49339, w49340, w49341, w49342, w49343, w49344, w49345, w49346, w49347, w49348, w49349, w49350, w49351, w49352, w49353, w49354, w49355, w49356, w49357, w49358, w49359, w49360, w49361, w49362, w49363, w49364, w49365, w49366, w49367, w49368, w49369, w49370, w49371, w49372, w49373, w49374, w49375, w49376, w49377, w49378, w49379, w49380, w49381, w49382, w49383, w49384, w49385, w49386, w49387, w49388, w49389, w49390, w49391, w49392, w49393, w49394, w49395, w49396, w49397, w49398, w49399, w49400, w49401, w49402, w49403, w49404, w49405, w49406, w49407, w49408, w49409, w49410, w49411, w49412, w49413, w49414, w49415, w49416, w49417, w49418, w49419, w49420, w49421, w49422, w49423, w49424, w49425, w49426, w49427, w49428, w49429, w49430, w49431, w49432, w49433, w49434, w49435, w49436, w49437, w49438, w49439, w49440, w49441, w49442, w49443, w49444, w49445, w49446, w49447, w49448, w49449, w49450, w49451, w49452, w49453, w49454, w49455, w49456, w49457, w49458, w49459, w49460, w49461, w49462, w49463, w49464, w49465, w49466, w49467, w49468, w49469, w49470, w49471, w49472, w49473, w49474, w49475, w49476, w49477, w49478, w49479, w49480, w49481, w49482, w49483, w49484, w49485, w49486, w49487, w49488, w49489, w49490, w49491, w49492, w49493, w49494, w49495, w49496, w49497, w49498, w49499, w49500, w49501, w49502, w49503, w49504, w49505, w49506, w49507, w49508, w49509, w49510, w49511, w49512, w49513, w49514, w49515, w49516, w49517, w49518, w49519, w49520, w49521, w49522, w49523, w49524, w49525, w49526, w49527, w49528, w49529, w49530, w49531, w49532, w49533, w49534, w49535, w49536, w49537, w49538, w49539, w49540, w49541, w49542, w49543, w49544, w49545, w49546, w49547, w49548, w49549, w49550, w49551, w49552, w49553, w49554, w49555, w49556, w49557, w49558, w49559, w49560, w49561, w49562, w49563, w49564, w49565, w49566, w49567, w49568, w49569, w49570, w49571, w49572, w49573, w49574, w49575, w49576, w49577, w49578, w49579, w49580, w49581, w49582, w49583, w49584, w49585, w49586, w49587, w49588, w49589, w49590, w49591, w49592, w49593, w49594, w49595, w49596, w49597, w49598, w49599, w49600, w49601, w49602, w49603, w49604, w49605, w49606, w49607, w49608, w49609, w49610, w49611, w49612, w49613, w49614, w49615, w49616, w49617, w49618, w49619, w49620, w49621, w49622, w49623, w49624, w49625, w49626, w49627, w49628, w49629, w49630, w49631, w49632, w49633, w49634, w49635, w49636, w49637, w49638, w49639, w49640, w49641, w49642, w49643, w49644, w49645, w49646, w49647, w49648, w49649, w49650, w49651, w49652, w49653, w49654, w49655, w49656, w49657, w49658, w49659, w49660, w49661, w49662, w49663, w49664, w49665, w49666, w49667, w49668, w49669, w49670, w49671, w49672, w49673, w49674, w49675, w49676, w49677, w49678, w49679, w49680, w49681, w49682, w49683, w49684, w49685, w49686, w49687, w49688, w49689, w49690, w49691, w49692, w49693, w49694, w49695, w49696, w49697, w49698, w49699, w49700, w49701, w49702, w49703, w49704, w49705, w49706, w49707, w49708, w49709, w49710, w49711, w49712, w49713, w49714, w49715, w49716, w49717, w49718, w49719, w49720, w49721, w49722, w49723, w49724, w49725, w49726, w49727, w49728, w49729, w49730, w49731, w49732, w49733, w49734, w49735, w49736, w49737, w49738, w49739, w49740, w49741, w49742, w49743, w49744, w49745, w49746, w49747, w49748, w49749, w49750, w49751, w49752, w49753, w49754, w49755, w49756, w49757, w49758, w49759, w49760, w49761, w49762, w49763, w49764, w49765, w49766, w49767, w49768, w49769, w49770, w49771, w49772, w49773, w49774, w49775, w49776, w49777, w49778, w49779, w49780, w49781, w49782, w49783, w49784, w49785, w49786, w49787, w49788, w49789, w49790, w49791, w49792, w49793, w49794, w49795, w49796, w49797, w49798, w49799, w49800, w49801, w49802, w49803, w49804, w49805, w49806, w49807, w49808, w49809, w49810, w49811, w49812, w49813, w49814, w49815, w49816, w49817, w49818, w49819, w49820, w49821, w49822, w49823, w49824, w49825, w49826, w49827, w49828, w49829, w49830, w49831, w49832, w49833, w49834, w49835, w49836, w49837, w49838, w49839, w49840, w49841, w49842, w49843, w49844, w49845, w49846, w49847, w49848, w49849, w49850, w49851, w49852, w49853, w49854, w49855, w49856, w49857, w49858, w49859, w49860, w49861, w49862, w49863, w49864, w49865, w49866, w49867, w49868, w49869, w49870, w49871, w49872, w49873, w49874, w49875, w49876, w49877, w49878, w49879, w49880, w49881, w49882, w49883, w49884, w49885, w49886, w49887, w49888, w49889, w49890, w49891, w49892, w49893, w49894, w49895, w49896, w49897, w49898, w49899, w49900, w49901, w49902, w49903, w49904, w49905, w49906, w49907, w49908, w49909, w49910, w49911, w49912, w49913, w49914, w49915, w49916, w49917, w49918, w49919, w49920, w49921, w49922, w49923, w49924, w49925, w49926, w49927, w49928, w49929, w49930, w49931, w49932, w49933, w49934, w49935, w49936, w49937, w49938, w49939, w49940, w49941, w49942, w49943, w49944, w49945, w49946, w49947, w49948, w49949, w49950, w49951, w49952, w49953, w49954, w49955, w49956, w49957, w49958, w49959, w49960, w49961, w49962, w49963, w49964, w49965, w49966, w49967, w49968, w49969, w49970, w49971, w49972, w49973, w49974, w49975, w49976, w49977, w49978, w49979, w49980, w49981, w49982, w49983, w49984, w49985, w49986, w49987, w49988, w49989, w49990, w49991, w49992, w49993, w49994, w49995, w49996, w49997, w49998, w49999, w50000, w50001, w50002, w50003, w50004, w50005, w50006, w50007, w50008, w50009, w50010, w50011, w50012, w50013, w50014, w50015, w50016, w50017, w50018, w50019, w50020, w50021, w50022, w50023, w50024, w50025, w50026, w50027, w50028, w50029, w50030, w50031, w50032, w50033, w50034, w50035, w50036, w50037, w50038, w50039, w50040, w50041, w50042, w50043, w50044, w50045, w50046, w50047, w50048, w50049, w50050, w50051, w50052, w50053, w50054, w50055, w50056, w50057, w50058, w50059, w50060, w50061, w50062, w50063, w50064, w50065, w50066, w50067, w50068, w50069, w50070, w50071, w50072, w50073, w50074, w50075, w50076, w50077, w50078, w50079, w50080, w50081, w50082, w50083, w50084, w50085, w50086, w50087, w50088, w50089, w50090, w50091, w50092, w50093, w50094, w50095, w50096, w50097, w50098, w50099, w50100, w50101, w50102, w50103, w50104, w50105, w50106, w50107, w50108, w50109, w50110, w50111, w50112, w50113, w50114, w50115, w50116, w50117, w50118, w50119, w50120, w50121, w50122, w50123, w50124, w50125, w50126, w50127, w50128, w50129, w50130, w50131, w50132, w50133, w50134, w50135, w50136, w50137, w50138, w50139, w50140, w50141, w50142, w50143, w50144, w50145, w50146, w50147, w50148, w50149, w50150, w50151, w50152, w50153, w50154, w50155, w50156, w50157, w50158, w50159, w50160, w50161, w50162, w50163, w50164, w50165, w50166, w50167, w50168, w50169, w50170, w50171, w50172, w50173, w50174, w50175, w50176, w50177, w50178, w50179, w50180, w50181, w50182, w50183, w50184, w50185, w50186, w50187, w50188, w50189, w50190, w50191, w50192, w50193, w50194, w50195, w50196, w50197, w50198, w50199, w50200, w50201, w50202, w50203, w50204, w50205, w50206, w50207, w50208, w50209, w50210, w50211, w50212, w50213, w50214, w50215, w50216, w50217, w50218, w50219, w50220, w50221, w50222, w50223, w50224, w50225, w50226, w50227, w50228, w50229, w50230, w50231, w50232, w50233, w50234, w50235, w50236, w50237, w50238, w50239, w50240, w50241, w50242, w50243, w50244, w50245, w50246, w50247, w50248, w50249, w50250, w50251, w50252, w50253, w50254, w50255, w50256, w50257, w50258, w50259, w50260, w50261, w50262, w50263, w50264, w50265, w50266, w50267, w50268, w50269, w50270, w50271, w50272, w50273, w50274, w50275, w50276, w50277, w50278, w50279, w50280, w50281, w50282, w50283, w50284, w50285, w50286, w50287, w50288, w50289, w50290, w50291, w50292, w50293, w50294, w50295, w50296, w50297, w50298, w50299, w50300, w50301, w50302, w50303, w50304, w50305, w50306, w50307, w50308, w50309, w50310, w50311, w50312, w50313, w50314, w50315, w50316, w50317, w50318, w50319, w50320, w50321, w50322, w50323, w50324, w50325, w50326, w50327, w50328, w50329, w50330, w50331, w50332, w50333, w50334, w50335, w50336, w50337, w50338, w50339, w50340, w50341, w50342, w50343, w50344, w50345, w50346, w50347, w50348, w50349, w50350, w50351, w50352, w50353, w50354, w50355, w50356, w50357, w50358, w50359, w50360, w50361, w50362, w50363, w50364, w50365, w50366, w50367, w50368, w50369, w50370, w50371, w50372, w50373, w50374, w50375, w50376, w50377, w50378, w50379, w50380, w50381, w50382, w50383, w50384, w50385, w50386, w50387, w50388, w50389, w50390, w50391, w50392, w50393, w50394, w50395, w50396, w50397, w50398, w50399, w50400, w50401, w50402, w50403, w50404, w50405, w50406, w50407, w50408, w50409, w50410, w50411, w50412, w50413, w50414, w50415, w50416, w50417, w50418, w50419, w50420, w50421, w50422, w50423, w50424, w50425, w50426, w50427, w50428, w50429, w50430, w50431, w50432, w50433, w50434, w50435, w50436, w50437, w50438, w50439, w50440, w50441, w50442, w50443, w50444, w50445, w50446, w50447, w50448, w50449, w50450, w50451, w50452, w50453, w50454, w50455, w50456, w50457, w50458, w50459, w50460, w50461, w50462, w50463, w50464, w50465, w50466, w50467, w50468, w50469, w50470, w50471, w50472, w50473, w50474, w50475, w50476, w50477, w50478, w50479, w50480, w50481, w50482, w50483, w50484, w50485, w50486, w50487, w50488, w50489, w50490, w50491, w50492, w50493, w50494, w50495, w50496, w50497, w50498, w50499, w50500, w50501, w50502, w50503, w50504, w50505, w50506, w50507, w50508, w50509, w50510, w50511, w50512, w50513, w50514, w50515, w50516, w50517, w50518, w50519, w50520, w50521, w50522, w50523, w50524, w50525, w50526, w50527, w50528, w50529, w50530, w50531, w50532, w50533, w50534, w50535, w50536, w50537, w50538, w50539, w50540, w50541, w50542, w50543, w50544, w50545, w50546, w50547, w50548, w50549, w50550, w50551, w50552, w50553, w50554, w50555, w50556, w50557, w50558, w50559, w50560, w50561, w50562, w50563, w50564, w50565, w50566, w50567, w50568, w50569, w50570, w50571, w50572, w50573, w50574, w50575, w50576, w50577, w50578, w50579, w50580, w50581, w50582, w50583, w50584, w50585, w50586, w50587, w50588, w50589, w50590, w50591, w50592, w50593, w50594, w50595, w50596, w50597, w50598, w50599, w50600, w50601, w50602, w50603, w50604, w50605, w50606, w50607, w50608, w50609, w50610, w50611, w50612, w50613, w50614, w50615, w50616, w50617, w50618, w50619, w50620, w50621, w50622, w50623, w50624, w50625, w50626, w50627, w50628, w50629, w50630, w50631, w50632, w50633, w50634, w50635, w50636, w50637, w50638, w50639, w50640, w50641, w50642, w50643, w50644, w50645, w50646, w50647, w50648, w50649, w50650, w50651, w50652, w50653, w50654, w50655, w50656, w50657, w50658, w50659, w50660, w50661, w50662, w50663, w50664, w50665, w50666, w50667, w50668, w50669, w50670, w50671, w50672, w50673, w50674, w50675, w50676, w50677, w50678, w50679, w50680, w50681, w50682, w50683, w50684, w50685, w50686, w50687, w50688, w50689, w50690, w50691, w50692, w50693, w50694, w50695, w50696, w50697, w50698, w50699, w50700, w50701, w50702, w50703, w50704, w50705, w50706, w50707, w50708, w50709, w50710, w50711, w50712, w50713, w50714, w50715, w50716, w50717, w50718, w50719, w50720, w50721, w50722, w50723, w50724, w50725, w50726, w50727, w50728, w50729, w50730, w50731, w50732, w50733, w50734, w50735, w50736, w50737, w50738, w50739, w50740, w50741, w50742, w50743, w50744, w50745, w50746, w50747, w50748, w50749, w50750, w50751, w50752, w50753, w50754, w50755, w50756, w50757, w50758, w50759, w50760, w50761, w50762, w50763, w50764, w50765, w50766, w50767, w50768, w50769, w50770, w50771, w50772, w50773, w50774, w50775, w50776, w50777, w50778, w50779, w50780, w50781, w50782, w50783, w50784, w50785, w50786, w50787, w50788, w50789, w50790, w50791, w50792, w50793, w50794, w50795, w50796, w50797, w50798, w50799, w50800, w50801, w50802, w50803, w50804, w50805, w50806, w50807, w50808, w50809, w50810, w50811, w50812, w50813, w50814, w50815, w50816, w50817, w50818, w50819, w50820, w50821, w50822, w50823, w50824, w50825, w50826, w50827, w50828, w50829, w50830, w50831, w50832, w50833, w50834, w50835, w50836, w50837, w50838, w50839, w50840, w50841, w50842, w50843, w50844, w50845, w50846, w50847, w50848, w50849, w50850, w50851, w50852, w50853, w50854, w50855, w50856, w50857, w50858, w50859, w50860, w50861, w50862, w50863, w50864, w50865, w50866, w50867, w50868, w50869, w50870, w50871, w50872, w50873, w50874, w50875, w50876, w50877, w50878, w50879, w50880, w50881, w50882, w50883, w50884, w50885, w50886, w50887, w50888, w50889, w50890, w50891, w50892, w50893, w50894, w50895, w50896, w50897, w50898, w50899, w50900, w50901, w50902, w50903, w50904, w50905, w50906, w50907, w50908, w50909, w50910, w50911, w50912, w50913, w50914, w50915, w50916, w50917, w50918, w50919, w50920, w50921, w50922, w50923, w50924, w50925, w50926, w50927, w50928, w50929, w50930, w50931, w50932, w50933, w50934, w50935, w50936, w50937, w50938, w50939, w50940, w50941, w50942, w50943, w50944, w50945, w50946, w50947, w50948, w50949, w50950, w50951, w50952, w50953, w50954, w50955, w50956, w50957, w50958, w50959, w50960, w50961, w50962, w50963, w50964, w50965, w50966, w50967, w50968, w50969, w50970, w50971, w50972, w50973, w50974, w50975, w50976, w50977, w50978, w50979, w50980, w50981, w50982, w50983, w50984, w50985, w50986, w50987, w50988, w50989, w50990, w50991, w50992, w50993, w50994, w50995, w50996, w50997, w50998, w50999, w51000, w51001, w51002, w51003, w51004, w51005, w51006, w51007, w51008, w51009, w51010, w51011, w51012, w51013, w51014, w51015, w51016, w51017, w51018, w51019, w51020, w51021, w51022, w51023, w51024, w51025, w51026, w51027, w51028, w51029, w51030, w51031, w51032, w51033, w51034, w51035, w51036, w51037, w51038, w51039, w51040, w51041, w51042, w51043, w51044, w51045, w51046, w51047, w51048, w51049, w51050, w51051, w51052, w51053, w51054, w51055, w51056, w51057, w51058, w51059, w51060, w51061, w51062, w51063, w51064, w51065, w51066, w51067, w51068, w51069, w51070, w51071, w51072, w51073, w51074, w51075, w51076, w51077, w51078, w51079, w51080, w51081, w51082, w51083, w51084, w51085, w51086, w51087, w51088, w51089, w51090, w51091, w51092, w51093, w51094, w51095, w51096, w51097, w51098, w51099, w51100, w51101, w51102, w51103, w51104, w51105, w51106, w51107, w51108, w51109, w51110, w51111, w51112, w51113, w51114, w51115, w51116, w51117, w51118, w51119, w51120, w51121, w51122, w51123, w51124, w51125, w51126, w51127, w51128, w51129, w51130, w51131, w51132, w51133, w51134, w51135, w51136, w51137, w51138, w51139, w51140, w51141, w51142, w51143, w51144, w51145, w51146, w51147, w51148, w51149, w51150, w51151, w51152, w51153, w51154, w51155, w51156, w51157, w51158, w51159, w51160, w51161, w51162, w51163, w51164, w51165, w51166, w51167, w51168, w51169, w51170, w51171, w51172, w51173, w51174, w51175, w51176, w51177, w51178, w51179, w51180, w51181, w51182, w51183, w51184, w51185, w51186, w51187, w51188, w51189, w51190, w51191, w51192, w51193, w51194, w51195, w51196, w51197, w51198, w51199, w51200, w51201, w51202, w51203, w51204, w51205, w51206, w51207, w51208, w51209, w51210, w51211, w51212, w51213, w51214, w51215, w51216, w51217, w51218, w51219, w51220, w51221, w51222, w51223, w51224, w51225, w51226, w51227, w51228, w51229, w51230, w51231, w51232, w51233, w51234, w51235, w51236, w51237, w51238, w51239, w51240, w51241, w51242, w51243, w51244, w51245, w51246, w51247, w51248, w51249, w51250, w51251, w51252, w51253, w51254, w51255, w51256, w51257, w51258, w51259, w51260, w51261, w51262, w51263, w51264, w51265, w51266, w51267, w51268, w51269, w51270, w51271, w51272, w51273, w51274, w51275, w51276, w51277, w51278, w51279, w51280, w51281, w51282, w51283, w51284, w51285, w51286, w51287, w51288, w51289, w51290, w51291, w51292, w51293, w51294, w51295, w51296, w51297, w51298, w51299, w51300, w51301, w51302, w51303, w51304, w51305, w51306, w51307, w51308, w51309, w51310, w51311, w51312, w51313, w51314, w51315, w51316, w51317, w51318, w51319, w51320, w51321, w51322, w51323, w51324, w51325, w51326, w51327, w51328, w51329, w51330, w51331, w51332, w51333, w51334, w51335, w51336, w51337, w51338, w51339, w51340, w51341, w51342, w51343, w51344, w51345, w51346, w51347, w51348, w51349, w51350, w51351, w51352, w51353, w51354, w51355, w51356, w51357, w51358, w51359, w51360, w51361, w51362, w51363, w51364, w51365, w51366, w51367, w51368, w51369, w51370, w51371, w51372, w51373, w51374, w51375, w51376, w51377, w51378, w51379, w51380, w51381, w51382, w51383, w51384, w51385, w51386, w51387, w51388, w51389, w51390, w51391, w51392, w51393, w51394, w51395, w51396, w51397, w51398, w51399, w51400, w51401, w51402, w51403, w51404, w51405, w51406, w51407, w51408, w51409, w51410, w51411, w51412, w51413, w51414, w51415, w51416, w51417, w51418, w51419, w51420, w51421, w51422, w51423, w51424, w51425, w51426, w51427, w51428, w51429, w51430, w51431, w51432, w51433, w51434, w51435, w51436, w51437, w51438, w51439, w51440, w51441, w51442, w51443, w51444, w51445, w51446, w51447, w51448, w51449, w51450, w51451, w51452, w51453, w51454, w51455, w51456, w51457, w51458, w51459, w51460, w51461, w51462, w51463, w51464, w51465, w51466, w51467, w51468, w51469, w51470, w51471, w51472, w51473, w51474, w51475, w51476, w51477, w51478, w51479, w51480, w51481, w51482, w51483, w51484, w51485, w51486, w51487, w51488, w51489, w51490, w51491, w51492, w51493, w51494, w51495, w51496, w51497, w51498, w51499, w51500, w51501, w51502, w51503, w51504, w51505, w51506, w51507, w51508, w51509, w51510, w51511, w51512, w51513, w51514, w51515, w51516, w51517, w51518, w51519, w51520, w51521, w51522, w51523, w51524, w51525, w51526, w51527, w51528, w51529, w51530, w51531, w51532, w51533, w51534, w51535, w51536, w51537, w51538, w51539, w51540, w51541, w51542, w51543, w51544, w51545, w51546, w51547, w51548, w51549, w51550, w51551, w51552, w51553, w51554, w51555, w51556, w51557, w51558, w51559, w51560, w51561, w51562, w51563, w51564, w51565, w51566, w51567, w51568, w51569, w51570, w51571, w51572, w51573, w51574, w51575, w51576, w51577, w51578, w51579, w51580, w51581, w51582, w51583, w51584, w51585, w51586, w51587, w51588, w51589, w51590, w51591, w51592, w51593, w51594, w51595, w51596, w51597, w51598, w51599, w51600, w51601, w51602, w51603, w51604, w51605, w51606, w51607, w51608, w51609, w51610, w51611, w51612, w51613, w51614, w51615, w51616, w51617, w51618, w51619, w51620, w51621, w51622, w51623, w51624, w51625, w51626, w51627, w51628, w51629, w51630, w51631, w51632, w51633, w51634, w51635, w51636, w51637, w51638, w51639, w51640, w51641, w51642, w51643, w51644, w51645, w51646, w51647, w51648, w51649, w51650, w51651, w51652, w51653, w51654, w51655, w51656, w51657, w51658, w51659, w51660, w51661, w51662, w51663, w51664, w51665, w51666, w51667, w51668, w51669, w51670, w51671, w51672, w51673, w51674, w51675, w51676, w51677, w51678, w51679, w51680, w51681, w51682, w51683, w51684, w51685, w51686, w51687, w51688, w51689, w51690, w51691, w51692, w51693, w51694, w51695, w51696, w51697, w51698, w51699, w51700, w51701, w51702, w51703, w51704, w51705, w51706, w51707, w51708, w51709, w51710, w51711, w51712, w51713, w51714, w51715, w51716, w51717, w51718, w51719, w51720, w51721, w51722, w51723, w51724, w51725, w51726, w51727, w51728, w51729, w51730, w51731, w51732, w51733, w51734, w51735, w51736, w51737, w51738, w51739, w51740, w51741, w51742, w51743, w51744, w51745, w51746, w51747, w51748, w51749, w51750, w51751, w51752, w51753, w51754, w51755, w51756, w51757, w51758, w51759, w51760, w51761, w51762, w51763, w51764, w51765, w51766, w51767, w51768, w51769, w51770, w51771, w51772, w51773, w51774, w51775, w51776, w51777, w51778, w51779, w51780, w51781, w51782, w51783, w51784, w51785, w51786, w51787, w51788, w51789, w51790, w51791, w51792, w51793, w51794, w51795, w51796, w51797, w51798, w51799, w51800, w51801, w51802, w51803, w51804, w51805, w51806, w51807, w51808, w51809, w51810, w51811, w51812, w51813, w51814, w51815, w51816, w51817, w51818, w51819, w51820, w51821, w51822, w51823, w51824, w51825, w51826, w51827, w51828, w51829, w51830, w51831, w51832, w51833, w51834, w51835, w51836, w51837, w51838, w51839, w51840, w51841, w51842, w51843, w51844, w51845, w51846, w51847, w51848, w51849, w51850, w51851, w51852, w51853, w51854, w51855, w51856, w51857, w51858, w51859, w51860, w51861, w51862, w51863, w51864, w51865, w51866, w51867, w51868, w51869, w51870, w51871, w51872, w51873, w51874, w51875, w51876, w51877, w51878, w51879, w51880, w51881, w51882, w51883, w51884, w51885, w51886, w51887, w51888, w51889, w51890, w51891, w51892, w51893, w51894, w51895, w51896, w51897, w51898, w51899, w51900, w51901, w51902, w51903, w51904, w51905, w51906, w51907, w51908, w51909, w51910, w51911, w51912, w51913, w51914, w51915, w51916, w51917, w51918, w51919, w51920, w51921, w51922, w51923, w51924, w51925, w51926, w51927, w51928, w51929, w51930, w51931, w51932, w51933, w51934, w51935, w51936, w51937, w51938, w51939, w51940, w51941, w51942, w51943, w51944, w51945, w51946, w51947, w51948, w51949, w51950, w51951, w51952, w51953, w51954, w51955, w51956, w51957, w51958, w51959, w51960, w51961, w51962, w51963, w51964, w51965, w51966, w51967, w51968, w51969, w51970, w51971, w51972, w51973, w51974, w51975, w51976, w51977, w51978, w51979, w51980, w51981, w51982, w51983, w51984, w51985, w51986, w51987, w51988, w51989, w51990, w51991, w51992, w51993, w51994, w51995, w51996, w51997, w51998, w51999, w52000, w52001, w52002, w52003, w52004, w52005, w52006, w52007, w52008, w52009, w52010, w52011, w52012, w52013, w52014, w52015, w52016, w52017, w52018, w52019, w52020, w52021, w52022, w52023, w52024, w52025, w52026, w52027, w52028, w52029, w52030, w52031, w52032, w52033, w52034, w52035, w52036, w52037, w52038, w52039, w52040, w52041, w52042, w52043, w52044, w52045, w52046, w52047, w52048, w52049, w52050, w52051, w52052, w52053, w52054, w52055, w52056, w52057, w52058, w52059, w52060, w52061, w52062, w52063, w52064, w52065, w52066, w52067, w52068, w52069, w52070, w52071, w52072, w52073, w52074, w52075, w52076, w52077, w52078, w52079, w52080, w52081, w52082, w52083, w52084, w52085, w52086, w52087, w52088, w52089, w52090, w52091, w52092, w52093, w52094, w52095, w52096, w52097, w52098, w52099, w52100, w52101, w52102, w52103, w52104, w52105, w52106, w52107, w52108, w52109, w52110, w52111, w52112, w52113, w52114, w52115, w52116, w52117, w52118, w52119, w52120, w52121, w52122, w52123, w52124, w52125, w52126, w52127, w52128, w52129, w52130, w52131, w52132, w52133, w52134, w52135, w52136, w52137, w52138, w52139, w52140, w52141, w52142, w52143, w52144, w52145, w52146, w52147, w52148, w52149, w52150, w52151, w52152, w52153, w52154, w52155, w52156, w52157, w52158, w52159, w52160, w52161, w52162, w52163, w52164, w52165, w52166, w52167, w52168, w52169, w52170, w52171, w52172, w52173, w52174, w52175, w52176, w52177, w52178, w52179, w52180, w52181, w52182, w52183, w52184, w52185, w52186, w52187, w52188, w52189, w52190, w52191, w52192, w52193, w52194, w52195, w52196, w52197, w52198, w52199, w52200, w52201, w52202, w52203, w52204, w52205, w52206, w52207, w52208, w52209, w52210, w52211, w52212, w52213, w52214, w52215, w52216, w52217, w52218, w52219, w52220, w52221, w52222, w52223, w52224, w52225, w52226, w52227, w52228, w52229, w52230, w52231, w52232, w52233, w52234, w52235, w52236, w52237, w52238, w52239, w52240, w52241, w52242, w52243, w52244, w52245, w52246, w52247, w52248, w52249, w52250, w52251, w52252, w52253, w52254, w52255, w52256, w52257, w52258, w52259, w52260, w52261, w52262, w52263, w52264, w52265, w52266, w52267, w52268, w52269, w52270, w52271, w52272, w52273, w52274, w52275, w52276, w52277, w52278, w52279, w52280, w52281, w52282, w52283, w52284, w52285, w52286, w52287, w52288, w52289, w52290, w52291, w52292, w52293, w52294, w52295, w52296, w52297, w52298, w52299, w52300, w52301, w52302, w52303, w52304, w52305, w52306, w52307, w52308, w52309, w52310, w52311, w52312, w52313, w52314, w52315, w52316, w52317, w52318, w52319, w52320, w52321, w52322, w52323, w52324, w52325, w52326, w52327, w52328, w52329, w52330, w52331, w52332, w52333, w52334, w52335, w52336, w52337, w52338, w52339, w52340, w52341, w52342, w52343, w52344, w52345, w52346, w52347, w52348, w52349, w52350, w52351, w52352, w52353, w52354, w52355, w52356, w52357, w52358, w52359, w52360, w52361, w52362, w52363, w52364, w52365, w52366, w52367, w52368, w52369, w52370, w52371, w52372, w52373, w52374, w52375, w52376, w52377, w52378, w52379, w52380, w52381, w52382, w52383, w52384, w52385, w52386, w52387, w52388, w52389, w52390, w52391, w52392, w52393, w52394, w52395, w52396, w52397, w52398, w52399, w52400, w52401, w52402, w52403, w52404, w52405, w52406, w52407, w52408, w52409, w52410, w52411, w52412, w52413, w52414, w52415, w52416, w52417, w52418, w52419, w52420, w52421, w52422, w52423, w52424, w52425, w52426, w52427, w52428, w52429, w52430, w52431, w52432, w52433, w52434, w52435, w52436, w52437, w52438, w52439, w52440, w52441, w52442, w52443, w52444, w52445, w52446, w52447, w52448, w52449, w52450, w52451, w52452, w52453, w52454, w52455, w52456, w52457, w52458, w52459, w52460, w52461, w52462, w52463, w52464, w52465, w52466, w52467, w52468, w52469, w52470, w52471, w52472, w52473, w52474, w52475, w52476, w52477, w52478, w52479, w52480, w52481, w52482, w52483, w52484, w52485, w52486, w52487, w52488, w52489, w52490, w52491, w52492, w52493, w52494, w52495, w52496, w52497, w52498, w52499, w52500, w52501, w52502, w52503, w52504, w52505, w52506, w52507, w52508, w52509, w52510, w52511, w52512, w52513, w52514, w52515, w52516, w52517, w52518, w52519, w52520, w52521, w52522, w52523, w52524, w52525, w52526, w52527, w52528, w52529, w52530, w52531, w52532, w52533, w52534, w52535, w52536, w52537, w52538, w52539, w52540, w52541, w52542, w52543, w52544, w52545, w52546, w52547, w52548, w52549, w52550, w52551, w52552, w52553, w52554, w52555, w52556, w52557, w52558, w52559, w52560, w52561, w52562, w52563, w52564, w52565, w52566, w52567, w52568, w52569, w52570, w52571, w52572, w52573, w52574, w52575, w52576, w52577, w52578, w52579, w52580, w52581, w52582, w52583, w52584, w52585, w52586, w52587, w52588, w52589, w52590, w52591, w52592, w52593, w52594, w52595, w52596, w52597, w52598, w52599, w52600, w52601, w52602, w52603, w52604, w52605, w52606, w52607, w52608, w52609, w52610, w52611, w52612, w52613, w52614, w52615, w52616, w52617, w52618, w52619, w52620, w52621, w52622, w52623, w52624, w52625, w52626, w52627, w52628, w52629, w52630, w52631, w52632, w52633, w52634, w52635, w52636, w52637, w52638, w52639, w52640, w52641, w52642, w52643, w52644, w52645, w52646, w52647, w52648, w52649, w52650, w52651, w52652, w52653, w52654, w52655, w52656, w52657, w52658, w52659, w52660, w52661, w52662, w52663, w52664, w52665, w52666, w52667, w52668, w52669, w52670, w52671, w52672, w52673, w52674, w52675, w52676, w52677, w52678, w52679, w52680, w52681, w52682, w52683, w52684, w52685, w52686, w52687, w52688, w52689, w52690, w52691, w52692, w52693, w52694, w52695, w52696, w52697, w52698, w52699, w52700, w52701, w52702, w52703, w52704, w52705, w52706, w52707, w52708, w52709, w52710, w52711, w52712, w52713, w52714, w52715, w52716, w52717, w52718, w52719, w52720, w52721, w52722, w52723, w52724, w52725, w52726, w52727, w52728, w52729, w52730, w52731, w52732, w52733, w52734, w52735, w52736, w52737, w52738, w52739, w52740, w52741, w52742, w52743, w52744, w52745, w52746, w52747, w52748, w52749, w52750, w52751, w52752, w52753, w52754, w52755, w52756, w52757, w52758, w52759, w52760, w52761, w52762, w52763, w52764, w52765, w52766, w52767, w52768, w52769, w52770, w52771, w52772, w52773, w52774, w52775, w52776, w52777, w52778, w52779, w52780, w52781, w52782, w52783, w52784, w52785, w52786, w52787, w52788, w52789, w52790, w52791, w52792, w52793, w52794, w52795, w52796, w52797, w52798, w52799, w52800, w52801, w52802, w52803, w52804, w52805, w52806, w52807, w52808, w52809, w52810, w52811, w52812, w52813, w52814, w52815, w52816, w52817, w52818, w52819, w52820, w52821, w52822, w52823, w52824, w52825, w52826, w52827, w52828, w52829, w52830, w52831, w52832, w52833, w52834, w52835, w52836, w52837, w52838, w52839, w52840, w52841, w52842, w52843, w52844, w52845, w52846, w52847, w52848, w52849, w52850, w52851, w52852, w52853, w52854, w52855, w52856, w52857, w52858, w52859, w52860, w52861, w52862, w52863, w52864, w52865, w52866, w52867, w52868, w52869, w52870, w52871, w52872, w52873, w52874, w52875, w52876, w52877, w52878, w52879, w52880, w52881, w52882, w52883, w52884, w52885, w52886, w52887, w52888, w52889, w52890, w52891, w52892, w52893, w52894, w52895, w52896, w52897, w52898, w52899, w52900, w52901, w52902, w52903, w52904, w52905, w52906, w52907, w52908, w52909, w52910, w52911, w52912, w52913, w52914, w52915, w52916, w52917, w52918, w52919, w52920, w52921, w52922, w52923, w52924, w52925, w52926, w52927, w52928, w52929, w52930, w52931, w52932, w52933, w52934, w52935, w52936, w52937, w52938, w52939, w52940, w52941, w52942, w52943, w52944, w52945, w52946, w52947, w52948, w52949, w52950, w52951, w52952, w52953, w52954, w52955, w52956, w52957, w52958, w52959, w52960, w52961, w52962, w52963, w52964, w52965, w52966, w52967, w52968, w52969, w52970, w52971, w52972, w52973, w52974, w52975, w52976, w52977, w52978, w52979, w52980, w52981, w52982, w52983, w52984, w52985, w52986, w52987, w52988, w52989, w52990, w52991, w52992, w52993, w52994, w52995, w52996, w52997, w52998, w52999, w53000, w53001, w53002, w53003, w53004, w53005, w53006, w53007, w53008, w53009, w53010, w53011, w53012, w53013, w53014, w53015, w53016, w53017, w53018, w53019, w53020, w53021, w53022, w53023, w53024, w53025, w53026, w53027, w53028, w53029, w53030, w53031, w53032, w53033, w53034, w53035, w53036, w53037, w53038, w53039, w53040, w53041, w53042, w53043, w53044, w53045, w53046, w53047, w53048, w53049, w53050, w53051, w53052, w53053, w53054, w53055, w53056, w53057, w53058, w53059, w53060, w53061, w53062, w53063, w53064, w53065, w53066, w53067, w53068, w53069, w53070, w53071, w53072, w53073, w53074, w53075, w53076, w53077, w53078, w53079, w53080, w53081, w53082, w53083, w53084, w53085, w53086, w53087, w53088, w53089, w53090, w53091, w53092, w53093, w53094, w53095, w53096, w53097, w53098, w53099, w53100, w53101, w53102, w53103, w53104, w53105, w53106, w53107, w53108, w53109, w53110, w53111, w53112, w53113, w53114, w53115, w53116, w53117, w53118, w53119, w53120, w53121, w53122, w53123, w53124, w53125, w53126, w53127, w53128, w53129, w53130, w53131, w53132, w53133, w53134, w53135, w53136, w53137, w53138, w53139, w53140, w53141, w53142, w53143, w53144, w53145, w53146, w53147, w53148, w53149, w53150, w53151, w53152, w53153, w53154, w53155, w53156, w53157, w53158, w53159, w53160, w53161, w53162, w53163, w53164, w53165, w53166, w53167, w53168, w53169, w53170, w53171, w53172, w53173, w53174, w53175, w53176, w53177, w53178, w53179, w53180, w53181, w53182, w53183, w53184, w53185, w53186, w53187, w53188, w53189, w53190, w53191, w53192, w53193, w53194, w53195, w53196, w53197, w53198, w53199, w53200, w53201, w53202, w53203, w53204, w53205, w53206, w53207, w53208, w53209, w53210, w53211, w53212, w53213, w53214, w53215, w53216, w53217, w53218, w53219, w53220, w53221, w53222, w53223, w53224, w53225, w53226, w53227, w53228, w53229, w53230, w53231, w53232, w53233, w53234, w53235, w53236, w53237, w53238, w53239, w53240, w53241, w53242, w53243, w53244, w53245, w53246, w53247, w53248, w53249, w53250, w53251, w53252, w53253, w53254, w53255, w53256, w53257, w53258, w53259, w53260, w53261, w53262, w53263, w53264, w53265, w53266, w53267, w53268, w53269, w53270, w53271, w53272, w53273, w53274, w53275, w53276, w53277, w53278, w53279, w53280, w53281, w53282, w53283, w53284, w53285, w53286, w53287, w53288, w53289, w53290, w53291, w53292, w53293, w53294, w53295, w53296, w53297, w53298, w53299, w53300, w53301, w53302, w53303, w53304, w53305, w53306, w53307, w53308, w53309, w53310, w53311, w53312, w53313, w53314, w53315, w53316, w53317, w53318, w53319, w53320, w53321, w53322, w53323, w53324, w53325, w53326, w53327, w53328, w53329, w53330, w53331, w53332, w53333, w53334, w53335, w53336, w53337, w53338, w53339, w53340, w53341, w53342, w53343, w53344, w53345, w53346, w53347, w53348, w53349, w53350, w53351, w53352, w53353, w53354, w53355, w53356, w53357, w53358, w53359, w53360, w53361, w53362, w53363, w53364, w53365, w53366, w53367, w53368, w53369, w53370, w53371, w53372, w53373, w53374, w53375, w53376, w53377, w53378, w53379, w53380, w53381, w53382, w53383, w53384, w53385, w53386, w53387, w53388, w53389, w53390, w53391, w53392, w53393, w53394, w53395, w53396, w53397, w53398, w53399, w53400, w53401, w53402, w53403, w53404, w53405, w53406, w53407, w53408, w53409, w53410, w53411, w53412, w53413, w53414, w53415, w53416, w53417, w53418, w53419, w53420, w53421, w53422, w53423, w53424, w53425, w53426, w53427, w53428, w53429, w53430, w53431, w53432, w53433, w53434, w53435, w53436, w53437, w53438, w53439, w53440, w53441, w53442, w53443, w53444, w53445, w53446, w53447, w53448, w53449, w53450, w53451, w53452, w53453, w53454, w53455, w53456, w53457, w53458, w53459, w53460, w53461, w53462, w53463, w53464, w53465, w53466, w53467, w53468, w53469, w53470, w53471, w53472, w53473, w53474, w53475, w53476, w53477, w53478, w53479, w53480, w53481, w53482, w53483, w53484, w53485, w53486, w53487, w53488, w53489, w53490, w53491, w53492, w53493, w53494, w53495, w53496, w53497, w53498, w53499, w53500, w53501, w53502, w53503, w53504, w53505, w53506, w53507, w53508, w53509, w53510, w53511, w53512, w53513, w53514, w53515, w53516, w53517, w53518, w53519, w53520, w53521, w53522, w53523, w53524, w53525, w53526, w53527, w53528, w53529, w53530, w53531, w53532, w53533, w53534, w53535, w53536, w53537, w53538, w53539, w53540, w53541, w53542, w53543, w53544, w53545, w53546, w53547, w53548, w53549, w53550, w53551, w53552, w53553, w53554, w53555, w53556, w53557, w53558, w53559, w53560, w53561, w53562, w53563, w53564, w53565, w53566, w53567, w53568, w53569, w53570, w53571, w53572, w53573, w53574, w53575, w53576, w53577, w53578, w53579, w53580, w53581, w53582, w53583, w53584, w53585, w53586, w53587, w53588, w53589, w53590, w53591, w53592, w53593, w53594, w53595, w53596, w53597, w53598, w53599, w53600, w53601, w53602, w53603, w53604, w53605, w53606, w53607, w53608, w53609, w53610, w53611, w53612, w53613, w53614, w53615, w53616, w53617, w53618, w53619, w53620, w53621, w53622, w53623, w53624, w53625, w53626, w53627, w53628, w53629, w53630, w53631, w53632, w53633, w53634, w53635, w53636, w53637, w53638, w53639, w53640, w53641, w53642, w53643, w53644, w53645, w53646, w53647, w53648, w53649, w53650, w53651, w53652, w53653, w53654, w53655, w53656, w53657, w53658, w53659, w53660, w53661, w53662, w53663, w53664, w53665, w53666, w53667, w53668, w53669, w53670, w53671, w53672, w53673, w53674, w53675, w53676, w53677, w53678, w53679, w53680, w53681, w53682, w53683, w53684, w53685, w53686, w53687, w53688, w53689, w53690, w53691, w53692, w53693, w53694, w53695, w53696, w53697, w53698, w53699, w53700, w53701, w53702, w53703, w53704, w53705, w53706, w53707, w53708, w53709, w53710, w53711, w53712, w53713, w53714, w53715, w53716, w53717, w53718, w53719, w53720, w53721, w53722, w53723, w53724, w53725, w53726, w53727, w53728, w53729, w53730, w53731, w53732, w53733, w53734, w53735, w53736, w53737, w53738, w53739, w53740, w53741, w53742, w53743, w53744, w53745, w53746, w53747, w53748, w53749, w53750, w53751, w53752, w53753, w53754, w53755, w53756, w53757, w53758, w53759, w53760, w53761, w53762, w53763, w53764, w53765, w53766, w53767, w53768, w53769, w53770, w53771, w53772, w53773, w53774, w53775, w53776, w53777, w53778, w53779, w53780, w53781, w53782, w53783, w53784, w53785, w53786, w53787, w53788, w53789, w53790, w53791, w53792, w53793, w53794, w53795, w53796, w53797, w53798, w53799, w53800, w53801, w53802, w53803, w53804, w53805, w53806, w53807, w53808, w53809, w53810, w53811, w53812, w53813, w53814, w53815, w53816, w53817, w53818, w53819, w53820, w53821, w53822, w53823, w53824, w53825, w53826, w53827, w53828, w53829, w53830, w53831, w53832, w53833, w53834, w53835, w53836, w53837, w53838, w53839, w53840, w53841, w53842, w53843, w53844, w53845, w53846, w53847, w53848, w53849, w53850, w53851, w53852, w53853, w53854, w53855, w53856, w53857, w53858, w53859, w53860, w53861, w53862, w53863, w53864, w53865, w53866, w53867, w53868, w53869, w53870, w53871, w53872, w53873, w53874, w53875, w53876, w53877, w53878, w53879, w53880, w53881, w53882, w53883, w53884, w53885, w53886, w53887, w53888, w53889, w53890, w53891, w53892, w53893, w53894, w53895, w53896, w53897, w53898, w53899, w53900, w53901, w53902, w53903, w53904, w53905, w53906, w53907, w53908, w53909, w53910, w53911, w53912, w53913, w53914, w53915, w53916, w53917, w53918, w53919, w53920, w53921, w53922, w53923, w53924, w53925, w53926, w53927, w53928, w53929, w53930, w53931, w53932, w53933, w53934, w53935, w53936, w53937, w53938, w53939, w53940, w53941, w53942, w53943, w53944, w53945, w53946, w53947, w53948, w53949, w53950, w53951, w53952, w53953, w53954, w53955, w53956, w53957, w53958, w53959, w53960, w53961, w53962, w53963, w53964, w53965, w53966, w53967, w53968, w53969, w53970, w53971, w53972, w53973, w53974, w53975, w53976, w53977, w53978, w53979, w53980, w53981, w53982, w53983, w53984, w53985, w53986, w53987, w53988, w53989, w53990, w53991, w53992, w53993, w53994, w53995, w53996, w53997, w53998, w53999, w54000, w54001, w54002, w54003, w54004, w54005, w54006, w54007, w54008, w54009, w54010, w54011, w54012, w54013, w54014, w54015, w54016, w54017, w54018, w54019, w54020, w54021, w54022, w54023, w54024, w54025, w54026, w54027, w54028, w54029, w54030, w54031, w54032, w54033, w54034, w54035, w54036, w54037, w54038, w54039, w54040, w54041, w54042, w54043, w54044, w54045, w54046, w54047, w54048, w54049, w54050, w54051, w54052, w54053, w54054, w54055, w54056, w54057, w54058, w54059, w54060, w54061, w54062, w54063, w54064, w54065, w54066, w54067, w54068, w54069, w54070, w54071, w54072, w54073, w54074, w54075, w54076, w54077, w54078, w54079, w54080, w54081, w54082, w54083, w54084, w54085, w54086, w54087, w54088, w54089, w54090, w54091, w54092, w54093, w54094, w54095, w54096, w54097, w54098, w54099, w54100, w54101, w54102, w54103, w54104, w54105, w54106, w54107, w54108, w54109, w54110, w54111, w54112, w54113, w54114, w54115, w54116, w54117, w54118, w54119, w54120, w54121, w54122, w54123, w54124, w54125, w54126, w54127, w54128, w54129, w54130, w54131, w54132, w54133, w54134, w54135, w54136, w54137, w54138, w54139, w54140, w54141, w54142, w54143, w54144, w54145, w54146, w54147, w54148, w54149, w54150, w54151, w54152, w54153, w54154, w54155, w54156, w54157, w54158, w54159, w54160, w54161, w54162, w54163, w54164, w54165, w54166, w54167, w54168, w54169, w54170, w54171, w54172, w54173, w54174, w54175, w54176, w54177, w54178, w54179, w54180, w54181, w54182, w54183, w54184, w54185, w54186, w54187, w54188, w54189, w54190, w54191, w54192, w54193, w54194, w54195, w54196, w54197, w54198, w54199, w54200, w54201, w54202, w54203, w54204, w54205, w54206, w54207, w54208, w54209, w54210, w54211, w54212, w54213, w54214, w54215, w54216, w54217, w54218, w54219, w54220, w54221, w54222, w54223, w54224, w54225, w54226, w54227, w54228, w54229, w54230, w54231, w54232, w54233, w54234, w54235, w54236, w54237, w54238, w54239, w54240, w54241, w54242, w54243, w54244, w54245, w54246, w54247, w54248, w54249, w54250, w54251, w54252, w54253, w54254, w54255, w54256, w54257, w54258, w54259, w54260, w54261, w54262, w54263, w54264, w54265, w54266, w54267, w54268, w54269, w54270, w54271, w54272, w54273, w54274, w54275, w54276, w54277, w54278, w54279, w54280, w54281, w54282, w54283, w54284, w54285, w54286, w54287, w54288, w54289, w54290, w54291, w54292, w54293, w54294, w54295, w54296, w54297, w54298, w54299, w54300, w54301, w54302, w54303, w54304, w54305, w54306, w54307, w54308, w54309, w54310, w54311, w54312, w54313, w54314, w54315, w54316, w54317, w54318, w54319, w54320, w54321, w54322, w54323, w54324, w54325, w54326, w54327, w54328, w54329, w54330, w54331, w54332, w54333, w54334, w54335, w54336, w54337, w54338, w54339, w54340, w54341, w54342, w54343, w54344, w54345, w54346, w54347, w54348, w54349, w54350, w54351, w54352, w54353, w54354, w54355, w54356, w54357, w54358, w54359, w54360, w54361, w54362, w54363, w54364, w54365, w54366, w54367, w54368, w54369, w54370, w54371, w54372, w54373, w54374, w54375, w54376, w54377, w54378, w54379, w54380, w54381, w54382, w54383, w54384, w54385, w54386, w54387, w54388, w54389, w54390, w54391, w54392, w54393, w54394, w54395, w54396, w54397, w54398, w54399, w54400, w54401, w54402, w54403, w54404, w54405, w54406, w54407, w54408, w54409, w54410, w54411, w54412, w54413, w54414, w54415, w54416, w54417, w54418, w54419, w54420, w54421, w54422, w54423, w54424, w54425, w54426, w54427, w54428, w54429, w54430, w54431, w54432, w54433, w54434, w54435, w54436, w54437, w54438, w54439, w54440, w54441, w54442, w54443, w54444, w54445, w54446, w54447, w54448, w54449, w54450, w54451, w54452, w54453, w54454, w54455, w54456, w54457, w54458, w54459, w54460, w54461, w54462, w54463, w54464, w54465, w54466, w54467, w54468, w54469, w54470, w54471, w54472, w54473, w54474, w54475, w54476, w54477, w54478, w54479, w54480, w54481, w54482, w54483, w54484, w54485, w54486, w54487, w54488, w54489, w54490, w54491, w54492, w54493, w54494, w54495, w54496, w54497, w54498, w54499, w54500, w54501, w54502, w54503, w54504, w54505, w54506, w54507, w54508, w54509, w54510, w54511, w54512, w54513, w54514, w54515, w54516, w54517, w54518, w54519, w54520, w54521, w54522, w54523, w54524, w54525, w54526, w54527, w54528, w54529, w54530, w54531, w54532, w54533, w54534, w54535, w54536, w54537, w54538, w54539, w54540, w54541, w54542, w54543, w54544, w54545, w54546, w54547, w54548, w54549, w54550, w54551, w54552, w54553, w54554, w54555, w54556, w54557, w54558, w54559, w54560, w54561, w54562, w54563, w54564, w54565, w54566, w54567, w54568, w54569, w54570, w54571, w54572, w54573, w54574, w54575, w54576, w54577, w54578, w54579, w54580, w54581, w54582, w54583, w54584, w54585, w54586, w54587, w54588, w54589, w54590, w54591, w54592, w54593, w54594, w54595, w54596, w54597, w54598, w54599, w54600, w54601, w54602, w54603, w54604, w54605, w54606, w54607, w54608, w54609, w54610, w54611, w54612, w54613, w54614, w54615, w54616, w54617, w54618, w54619, w54620, w54621, w54622, w54623, w54624, w54625, w54626, w54627, w54628, w54629, w54630, w54631, w54632, w54633, w54634, w54635, w54636, w54637, w54638, w54639, w54640, w54641, w54642, w54643, w54644, w54645, w54646, w54647, w54648, w54649, w54650, w54651, w54652, w54653, w54654, w54655, w54656, w54657, w54658, w54659, w54660, w54661, w54662, w54663, w54664, w54665, w54666, w54667, w54668, w54669, w54670, w54671, w54672, w54673, w54674, w54675, w54676, w54677, w54678, w54679, w54680, w54681, w54682, w54683, w54684, w54685, w54686, w54687, w54688, w54689, w54690, w54691, w54692, w54693, w54694, w54695, w54696, w54697, w54698, w54699, w54700, w54701, w54702, w54703, w54704, w54705, w54706, w54707, w54708, w54709, w54710, w54711, w54712, w54713, w54714, w54715, w54716, w54717, w54718, w54719, w54720, w54721, w54722, w54723, w54724, w54725, w54726, w54727, w54728, w54729, w54730, w54731, w54732, w54733, w54734, w54735, w54736, w54737, w54738, w54739, w54740, w54741, w54742, w54743, w54744, w54745, w54746, w54747, w54748, w54749, w54750, w54751, w54752, w54753, w54754, w54755, w54756, w54757, w54758, w54759, w54760, w54761, w54762, w54763, w54764, w54765, w54766, w54767, w54768, w54769, w54770, w54771, w54772, w54773, w54774, w54775, w54776, w54777, w54778, w54779, w54780, w54781, w54782, w54783, w54784, w54785, w54786, w54787, w54788, w54789, w54790, w54791, w54792, w54793, w54794, w54795, w54796, w54797, w54798, w54799, w54800, w54801, w54802, w54803, w54804, w54805, w54806, w54807, w54808, w54809, w54810, w54811, w54812, w54813, w54814, w54815, w54816, w54817, w54818, w54819, w54820, w54821, w54822, w54823, w54824, w54825, w54826, w54827, w54828, w54829, w54830, w54831, w54832, w54833, w54834, w54835, w54836, w54837, w54838, w54839, w54840, w54841, w54842, w54843, w54844, w54845, w54846, w54847, w54848, w54849, w54850, w54851, w54852, w54853, w54854, w54855, w54856, w54857, w54858, w54859, w54860, w54861, w54862, w54863, w54864, w54865, w54866, w54867, w54868, w54869, w54870, w54871, w54872, w54873, w54874, w54875, w54876, w54877, w54878, w54879, w54880, w54881, w54882, w54883, w54884, w54885, w54886, w54887, w54888, w54889, w54890, w54891, w54892, w54893, w54894, w54895, w54896, w54897, w54898, w54899, w54900, w54901, w54902, w54903, w54904, w54905, w54906, w54907, w54908, w54909, w54910, w54911, w54912, w54913, w54914, w54915, w54916, w54917, w54918, w54919, w54920, w54921, w54922, w54923, w54924, w54925, w54926, w54927, w54928, w54929, w54930, w54931, w54932, w54933, w54934, w54935, w54936, w54937, w54938, w54939, w54940, w54941, w54942, w54943, w54944, w54945, w54946, w54947, w54948, w54949, w54950, w54951, w54952, w54953, w54954, w54955, w54956, w54957, w54958, w54959, w54960, w54961, w54962, w54963, w54964, w54965, w54966, w54967, w54968, w54969, w54970, w54971, w54972, w54973, w54974, w54975, w54976, w54977, w54978, w54979, w54980, w54981, w54982, w54983, w54984, w54985, w54986, w54987, w54988, w54989, w54990, w54991, w54992, w54993, w54994, w54995, w54996, w54997, w54998, w54999, w55000, w55001, w55002, w55003, w55004, w55005, w55006, w55007, w55008, w55009, w55010, w55011, w55012, w55013, w55014, w55015, w55016, w55017, w55018, w55019, w55020, w55021, w55022, w55023, w55024, w55025, w55026, w55027, w55028, w55029, w55030, w55031, w55032, w55033, w55034, w55035, w55036, w55037, w55038, w55039, w55040, w55041, w55042, w55043, w55044, w55045, w55046, w55047, w55048, w55049, w55050, w55051, w55052, w55053, w55054, w55055, w55056, w55057, w55058, w55059, w55060, w55061, w55062, w55063, w55064, w55065, w55066, w55067, w55068, w55069, w55070, w55071, w55072, w55073, w55074, w55075, w55076, w55077, w55078, w55079, w55080, w55081, w55082, w55083, w55084, w55085, w55086, w55087, w55088, w55089, w55090, w55091, w55092, w55093, w55094, w55095, w55096, w55097, w55098, w55099, w55100, w55101, w55102, w55103, w55104, w55105, w55106, w55107, w55108, w55109, w55110, w55111, w55112, w55113, w55114, w55115, w55116, w55117, w55118, w55119, w55120, w55121, w55122, w55123, w55124, w55125, w55126, w55127, w55128, w55129, w55130, w55131, w55132, w55133, w55134, w55135, w55136, w55137, w55138, w55139, w55140, w55141, w55142, w55143, w55144, w55145, w55146, w55147, w55148, w55149, w55150, w55151, w55152, w55153, w55154, w55155, w55156, w55157, w55158, w55159, w55160, w55161, w55162, w55163, w55164, w55165, w55166, w55167, w55168, w55169, w55170, w55171, w55172, w55173, w55174, w55175, w55176, w55177, w55178, w55179, w55180, w55181, w55182, w55183, w55184, w55185, w55186, w55187, w55188, w55189, w55190, w55191, w55192, w55193, w55194, w55195, w55196, w55197, w55198, w55199, w55200, w55201, w55202, w55203, w55204, w55205, w55206, w55207, w55208, w55209, w55210, w55211, w55212, w55213, w55214, w55215, w55216, w55217, w55218, w55219, w55220, w55221, w55222, w55223, w55224, w55225, w55226, w55227, w55228, w55229, w55230, w55231, w55232, w55233, w55234, w55235, w55236, w55237, w55238, w55239, w55240, w55241, w55242, w55243, w55244, w55245, w55246, w55247, w55248, w55249, w55250, w55251, w55252, w55253, w55254, w55255, w55256, w55257, w55258, w55259, w55260, w55261, w55262, w55263, w55264, w55265, w55266, w55267, w55268, w55269, w55270, w55271, w55272, w55273, w55274, w55275, w55276, w55277, w55278, w55279, w55280, w55281, w55282, w55283, w55284, w55285, w55286, w55287, w55288, w55289, w55290, w55291, w55292, w55293, w55294, w55295, w55296, w55297, w55298, w55299, w55300, w55301, w55302, w55303, w55304, w55305, w55306, w55307, w55308, w55309, w55310, w55311, w55312, w55313, w55314, w55315, w55316, w55317, w55318, w55319, w55320, w55321, w55322, w55323, w55324, w55325, w55326, w55327, w55328, w55329, w55330, w55331, w55332, w55333, w55334, w55335, w55336, w55337, w55338, w55339, w55340, w55341, w55342, w55343, w55344, w55345, w55346, w55347, w55348, w55349, w55350, w55351, w55352, w55353, w55354, w55355, w55356, w55357, w55358, w55359, w55360, w55361, w55362, w55363, w55364, w55365, w55366, w55367, w55368, w55369, w55370, w55371, w55372, w55373, w55374, w55375, w55376, w55377, w55378, w55379, w55380, w55381, w55382, w55383, w55384, w55385, w55386, w55387, w55388, w55389, w55390, w55391, w55392, w55393, w55394, w55395, w55396, w55397, w55398, w55399, w55400, w55401, w55402, w55403, w55404, w55405, w55406, w55407, w55408, w55409, w55410, w55411, w55412, w55413, w55414, w55415, w55416, w55417, w55418, w55419, w55420, w55421, w55422, w55423, w55424, w55425, w55426, w55427, w55428, w55429, w55430, w55431, w55432, w55433, w55434, w55435, w55436, w55437, w55438, w55439, w55440, w55441, w55442, w55443, w55444, w55445, w55446, w55447, w55448, w55449, w55450, w55451, w55452, w55453, w55454, w55455, w55456, w55457, w55458, w55459, w55460, w55461, w55462, w55463, w55464, w55465, w55466, w55467, w55468, w55469, w55470, w55471, w55472, w55473, w55474, w55475, w55476, w55477, w55478, w55479, w55480, w55481, w55482, w55483, w55484, w55485, w55486, w55487, w55488, w55489, w55490, w55491, w55492, w55493, w55494, w55495, w55496, w55497, w55498, w55499, w55500, w55501, w55502, w55503, w55504, w55505, w55506, w55507, w55508, w55509, w55510, w55511, w55512, w55513, w55514, w55515, w55516, w55517, w55518, w55519, w55520, w55521, w55522, w55523, w55524, w55525, w55526, w55527, w55528, w55529, w55530, w55531, w55532, w55533, w55534, w55535, w55536, w55537, w55538, w55539, w55540, w55541, w55542, w55543, w55544, w55545, w55546, w55547, w55548, w55549, w55550, w55551, w55552, w55553, w55554, w55555, w55556, w55557, w55558, w55559, w55560, w55561, w55562, w55563, w55564, w55565, w55566, w55567, w55568, w55569, w55570, w55571, w55572, w55573, w55574, w55575, w55576, w55577, w55578, w55579, w55580, w55581, w55582, w55583, w55584, w55585, w55586, w55587, w55588, w55589, w55590, w55591, w55592, w55593, w55594, w55595, w55596, w55597, w55598, w55599, w55600, w55601, w55602, w55603, w55604, w55605, w55606, w55607, w55608, w55609, w55610, w55611, w55612, w55613, w55614, w55615, w55616, w55617, w55618, w55619, w55620, w55621, w55622, w55623, w55624, w55625, w55626, w55627, w55628, w55629, w55630, w55631, w55632, w55633, w55634, w55635, w55636, w55637, w55638, w55639, w55640, w55641, w55642, w55643, w55644, w55645, w55646, w55647, w55648, w55649, w55650, w55651, w55652, w55653, w55654, w55655, w55656, w55657, w55658, w55659, w55660, w55661, w55662, w55663, w55664, w55665, w55666, w55667, w55668, w55669, w55670, w55671, w55672, w55673, w55674, w55675, w55676, w55677, w55678, w55679, w55680, w55681, w55682, w55683, w55684, w55685, w55686, w55687, w55688, w55689, w55690, w55691, w55692, w55693, w55694, w55695, w55696, w55697, w55698, w55699, w55700, w55701, w55702, w55703, w55704, w55705, w55706, w55707, w55708, w55709, w55710, w55711, w55712, w55713, w55714, w55715, w55716, w55717, w55718, w55719, w55720, w55721, w55722, w55723, w55724, w55725, w55726, w55727, w55728, w55729, w55730, w55731, w55732, w55733, w55734, w55735, w55736, w55737, w55738, w55739, w55740, w55741, w55742, w55743, w55744, w55745, w55746, w55747, w55748, w55749, w55750, w55751, w55752, w55753, w55754, w55755, w55756, w55757, w55758, w55759, w55760, w55761, w55762, w55763, w55764, w55765, w55766, w55767, w55768, w55769, w55770, w55771, w55772, w55773, w55774, w55775, w55776, w55777, w55778, w55779, w55780, w55781, w55782, w55783, w55784, w55785, w55786, w55787, w55788, w55789, w55790, w55791, w55792, w55793, w55794, w55795, w55796, w55797, w55798, w55799, w55800, w55801, w55802, w55803, w55804, w55805, w55806, w55807, w55808, w55809, w55810, w55811, w55812, w55813, w55814, w55815, w55816, w55817, w55818, w55819, w55820, w55821, w55822, w55823, w55824, w55825, w55826, w55827, w55828, w55829, w55830, w55831, w55832, w55833, w55834, w55835, w55836, w55837, w55838, w55839, w55840, w55841, w55842, w55843, w55844, w55845, w55846, w55847, w55848, w55849, w55850, w55851, w55852, w55853, w55854, w55855, w55856, w55857, w55858, w55859, w55860, w55861, w55862, w55863, w55864, w55865, w55866, w55867, w55868, w55869, w55870, w55871, w55872, w55873, w55874, w55875, w55876, w55877, w55878, w55879, w55880, w55881, w55882, w55883, w55884, w55885, w55886, w55887, w55888, w55889, w55890, w55891, w55892, w55893, w55894, w55895, w55896, w55897, w55898, w55899, w55900, w55901, w55902, w55903, w55904, w55905, w55906, w55907, w55908, w55909, w55910, w55911, w55912, w55913, w55914, w55915, w55916, w55917, w55918, w55919, w55920, w55921, w55922, w55923, w55924, w55925, w55926, w55927, w55928, w55929, w55930, w55931, w55932, w55933, w55934, w55935, w55936, w55937, w55938, w55939, w55940, w55941, w55942, w55943, w55944, w55945, w55946, w55947, w55948, w55949, w55950, w55951, w55952, w55953, w55954, w55955, w55956, w55957, w55958, w55959, w55960, w55961, w55962, w55963, w55964, w55965, w55966, w55967, w55968, w55969, w55970, w55971, w55972, w55973, w55974, w55975, w55976, w55977, w55978, w55979, w55980, w55981, w55982, w55983, w55984, w55985, w55986, w55987, w55988, w55989, w55990, w55991, w55992, w55993, w55994, w55995, w55996, w55997, w55998, w55999, w56000, w56001, w56002, w56003, w56004, w56005, w56006, w56007, w56008, w56009, w56010, w56011, w56012, w56013, w56014, w56015, w56016, w56017, w56018, w56019, w56020, w56021, w56022, w56023, w56024, w56025, w56026, w56027, w56028, w56029, w56030, w56031, w56032, w56033, w56034, w56035, w56036, w56037, w56038, w56039, w56040, w56041, w56042, w56043, w56044, w56045, w56046, w56047, w56048, w56049, w56050, w56051, w56052, w56053, w56054, w56055, w56056, w56057, w56058, w56059, w56060, w56061, w56062, w56063, w56064, w56065, w56066, w56067, w56068, w56069, w56070, w56071, w56072, w56073, w56074, w56075, w56076, w56077, w56078, w56079, w56080, w56081, w56082, w56083, w56084, w56085, w56086, w56087, w56088, w56089, w56090, w56091, w56092, w56093, w56094, w56095, w56096, w56097, w56098, w56099, w56100, w56101, w56102, w56103, w56104, w56105, w56106, w56107, w56108, w56109, w56110, w56111, w56112, w56113, w56114, w56115, w56116, w56117, w56118, w56119, w56120, w56121, w56122, w56123, w56124, w56125, w56126, w56127, w56128, w56129, w56130, w56131, w56132, w56133, w56134, w56135, w56136, w56137, w56138, w56139, w56140, w56141, w56142, w56143, w56144, w56145, w56146, w56147, w56148, w56149, w56150, w56151, w56152, w56153, w56154, w56155, w56156, w56157, w56158, w56159, w56160, w56161, w56162, w56163, w56164, w56165, w56166, w56167, w56168, w56169, w56170, w56171, w56172, w56173, w56174, w56175, w56176, w56177, w56178, w56179, w56180, w56181, w56182, w56183, w56184, w56185, w56186, w56187, w56188, w56189, w56190, w56191, w56192, w56193, w56194, w56195, w56196, w56197, w56198, w56199, w56200, w56201, w56202, w56203, w56204, w56205, w56206, w56207, w56208, w56209, w56210, w56211, w56212, w56213, w56214, w56215, w56216, w56217, w56218, w56219, w56220, w56221, w56222, w56223, w56224, w56225, w56226, w56227, w56228, w56229, w56230, w56231, w56232, w56233, w56234, w56235, w56236, w56237, w56238, w56239, w56240, w56241, w56242, w56243, w56244, w56245, w56246, w56247, w56248, w56249, w56250, w56251, w56252, w56253, w56254, w56255, w56256, w56257, w56258, w56259, w56260, w56261, w56262, w56263, w56264, w56265, w56266, w56267, w56268, w56269, w56270, w56271, w56272, w56273, w56274, w56275, w56276, w56277, w56278, w56279, w56280, w56281, w56282, w56283, w56284, w56285, w56286, w56287, w56288, w56289, w56290, w56291, w56292, w56293, w56294, w56295, w56296, w56297, w56298, w56299, w56300, w56301, w56302, w56303, w56304, w56305, w56306, w56307, w56308, w56309, w56310, w56311, w56312, w56313, w56314, w56315, w56316, w56317, w56318, w56319, w56320, w56321, w56322, w56323, w56324, w56325, w56326, w56327, w56328, w56329, w56330, w56331, w56332, w56333, w56334, w56335, w56336, w56337, w56338, w56339, w56340, w56341, w56342, w56343, w56344, w56345, w56346, w56347, w56348, w56349, w56350, w56351, w56352, w56353, w56354, w56355, w56356, w56357, w56358, w56359, w56360, w56361, w56362, w56363, w56364, w56365, w56366, w56367, w56368, w56369, w56370, w56371, w56372, w56373, w56374, w56375, w56376, w56377, w56378, w56379, w56380, w56381, w56382, w56383, w56384, w56385, w56386, w56387, w56388, w56389, w56390, w56391, w56392, w56393, w56394, w56395, w56396, w56397, w56398, w56399, w56400, w56401, w56402, w56403, w56404, w56405, w56406, w56407, w56408, w56409, w56410, w56411, w56412, w56413, w56414, w56415, w56416, w56417, w56418, w56419, w56420, w56421, w56422, w56423, w56424, w56425, w56426, w56427, w56428, w56429, w56430, w56431, w56432, w56433, w56434, w56435, w56436, w56437, w56438, w56439, w56440, w56441, w56442, w56443, w56444, w56445, w56446, w56447, w56448, w56449, w56450, w56451, w56452, w56453, w56454, w56455, w56456, w56457, w56458, w56459, w56460, w56461, w56462, w56463, w56464, w56465, w56466, w56467, w56468, w56469, w56470, w56471, w56472, w56473, w56474, w56475, w56476, w56477, w56478, w56479, w56480, w56481, w56482, w56483, w56484, w56485, w56486, w56487, w56488, w56489, w56490, w56491, w56492, w56493, w56494, w56495, w56496, w56497, w56498, w56499, w56500, w56501, w56502, w56503, w56504, w56505, w56506, w56507, w56508, w56509, w56510, w56511, w56512, w56513, w56514, w56515, w56516, w56517, w56518, w56519, w56520, w56521, w56522, w56523, w56524, w56525, w56526, w56527, w56528, w56529, w56530, w56531, w56532, w56533, w56534, w56535, w56536, w56537, w56538, w56539, w56540, w56541, w56542, w56543, w56544, w56545, w56546, w56547, w56548, w56549, w56550, w56551, w56552, w56553, w56554, w56555, w56556, w56557, w56558, w56559, w56560, w56561, w56562, w56563, w56564, w56565, w56566, w56567, w56568, w56569, w56570, w56571, w56572, w56573, w56574, w56575, w56576, w56577, w56578, w56579, w56580, w56581, w56582, w56583, w56584, w56585, w56586, w56587, w56588, w56589, w56590, w56591, w56592, w56593, w56594, w56595, w56596, w56597, w56598, w56599, w56600, w56601, w56602, w56603, w56604, w56605, w56606, w56607, w56608, w56609, w56610, w56611, w56612, w56613, w56614, w56615, w56616, w56617, w56618, w56619, w56620, w56621, w56622, w56623, w56624, w56625, w56626, w56627, w56628, w56629, w56630, w56631, w56632, w56633, w56634, w56635, w56636, w56637, w56638, w56639, w56640, w56641, w56642, w56643, w56644, w56645, w56646, w56647, w56648, w56649, w56650, w56651, w56652, w56653, w56654, w56655, w56656, w56657, w56658, w56659, w56660, w56661, w56662, w56663, w56664, w56665, w56666, w56667, w56668, w56669, w56670, w56671, w56672, w56673, w56674, w56675, w56676, w56677, w56678, w56679, w56680, w56681, w56682, w56683, w56684, w56685, w56686, w56687, w56688, w56689, w56690, w56691, w56692, w56693, w56694, w56695, w56696, w56697, w56698, w56699, w56700, w56701, w56702, w56703, w56704, w56705, w56706, w56707, w56708, w56709, w56710, w56711, w56712, w56713, w56714, w56715, w56716, w56717, w56718, w56719, w56720, w56721, w56722, w56723, w56724, w56725, w56726, w56727, w56728, w56729, w56730, w56731, w56732, w56733, w56734, w56735, w56736, w56737, w56738, w56739, w56740, w56741, w56742, w56743, w56744, w56745, w56746, w56747, w56748, w56749, w56750, w56751, w56752, w56753, w56754, w56755, w56756, w56757, w56758, w56759, w56760, w56761, w56762, w56763, w56764, w56765, w56766, w56767, w56768, w56769, w56770, w56771, w56772, w56773, w56774, w56775, w56776, w56777, w56778, w56779, w56780, w56781, w56782, w56783, w56784, w56785, w56786, w56787, w56788, w56789, w56790, w56791, w56792, w56793, w56794, w56795, w56796, w56797, w56798, w56799, w56800, w56801, w56802, w56803, w56804, w56805, w56806, w56807, w56808, w56809, w56810, w56811, w56812, w56813, w56814, w56815, w56816, w56817, w56818, w56819, w56820, w56821, w56822, w56823, w56824, w56825, w56826, w56827, w56828, w56829, w56830, w56831, w56832, w56833, w56834, w56835, w56836, w56837, w56838, w56839, w56840, w56841, w56842, w56843, w56844, w56845, w56846, w56847, w56848, w56849, w56850, w56851, w56852, w56853, w56854, w56855, w56856, w56857, w56858, w56859, w56860, w56861, w56862, w56863, w56864, w56865, w56866, w56867, w56868, w56869, w56870, w56871, w56872, w56873, w56874, w56875, w56876, w56877, w56878, w56879, w56880, w56881, w56882, w56883, w56884, w56885, w56886, w56887, w56888, w56889, w56890, w56891, w56892, w56893, w56894, w56895, w56896, w56897, w56898, w56899, w56900, w56901, w56902, w56903, w56904, w56905, w56906, w56907, w56908, w56909, w56910, w56911, w56912, w56913, w56914, w56915, w56916, w56917, w56918, w56919, w56920, w56921, w56922, w56923, w56924, w56925, w56926, w56927, w56928, w56929, w56930, w56931, w56932, w56933, w56934, w56935, w56936, w56937, w56938, w56939, w56940, w56941, w56942, w56943, w56944, w56945, w56946, w56947, w56948, w56949, w56950, w56951, w56952, w56953, w56954, w56955, w56956, w56957, w56958, w56959, w56960, w56961, w56962, w56963, w56964, w56965, w56966, w56967, w56968, w56969, w56970, w56971, w56972, w56973, w56974, w56975, w56976, w56977, w56978, w56979, w56980, w56981, w56982, w56983, w56984, w56985, w56986, w56987, w56988, w56989, w56990, w56991, w56992, w56993, w56994, w56995, w56996, w56997, w56998, w56999, w57000, w57001, w57002, w57003, w57004, w57005, w57006, w57007, w57008, w57009, w57010, w57011, w57012, w57013, w57014, w57015, w57016, w57017, w57018, w57019, w57020, w57021, w57022, w57023, w57024, w57025, w57026, w57027, w57028, w57029, w57030, w57031, w57032, w57033, w57034, w57035, w57036, w57037, w57038, w57039, w57040, w57041, w57042, w57043, w57044, w57045, w57046, w57047, w57048, w57049, w57050, w57051, w57052, w57053, w57054, w57055, w57056, w57057, w57058, w57059, w57060, w57061, w57062, w57063, w57064, w57065, w57066, w57067, w57068, w57069, w57070, w57071, w57072, w57073, w57074, w57075, w57076, w57077, w57078, w57079, w57080, w57081, w57082, w57083, w57084, w57085, w57086, w57087, w57088, w57089, w57090, w57091, w57092, w57093, w57094, w57095, w57096, w57097, w57098, w57099, w57100, w57101, w57102, w57103, w57104, w57105, w57106, w57107, w57108, w57109, w57110, w57111, w57112, w57113, w57114, w57115, w57116, w57117, w57118, w57119, w57120, w57121, w57122, w57123, w57124, w57125, w57126, w57127, w57128, w57129, w57130, w57131, w57132, w57133, w57134, w57135, w57136, w57137, w57138, w57139, w57140, w57141, w57142, w57143, w57144, w57145, w57146, w57147, w57148, w57149, w57150, w57151, w57152, w57153, w57154, w57155, w57156, w57157, w57158, w57159, w57160, w57161, w57162, w57163, w57164, w57165, w57166, w57167, w57168, w57169, w57170, w57171, w57172, w57173, w57174, w57175, w57176, w57177, w57178, w57179, w57180, w57181, w57182, w57183, w57184, w57185, w57186, w57187, w57188, w57189, w57190, w57191, w57192, w57193, w57194, w57195, w57196, w57197, w57198, w57199, w57200, w57201, w57202, w57203, w57204, w57205, w57206, w57207, w57208, w57209, w57210, w57211, w57212, w57213, w57214, w57215, w57216, w57217, w57218, w57219, w57220, w57221, w57222, w57223, w57224, w57225, w57226, w57227, w57228, w57229, w57230, w57231, w57232, w57233, w57234, w57235, w57236, w57237, w57238, w57239, w57240, w57241, w57242, w57243, w57244, w57245, w57246, w57247, w57248, w57249, w57250, w57251, w57252, w57253, w57254, w57255, w57256, w57257, w57258, w57259, w57260, w57261, w57262, w57263, w57264, w57265, w57266, w57267, w57268, w57269, w57270, w57271, w57272, w57273, w57274, w57275, w57276, w57277, w57278, w57279, w57280, w57281, w57282, w57283, w57284, w57285, w57286, w57287, w57288, w57289, w57290, w57291, w57292, w57293, w57294, w57295, w57296, w57297, w57298, w57299, w57300, w57301, w57302, w57303, w57304, w57305, w57306, w57307, w57308, w57309, w57310, w57311, w57312, w57313, w57314, w57315, w57316, w57317, w57318, w57319, w57320, w57321, w57322, w57323, w57324, w57325, w57326, w57327, w57328, w57329, w57330, w57331, w57332, w57333, w57334, w57335, w57336, w57337, w57338, w57339, w57340, w57341, w57342, w57343, w57344, w57345, w57346, w57347, w57348, w57349, w57350, w57351, w57352, w57353, w57354, w57355, w57356, w57357, w57358, w57359, w57360, w57361, w57362, w57363, w57364, w57365, w57366, w57367, w57368, w57369, w57370, w57371, w57372, w57373, w57374, w57375, w57376, w57377, w57378, w57379, w57380, w57381, w57382, w57383, w57384, w57385, w57386, w57387, w57388, w57389, w57390, w57391, w57392, w57393, w57394, w57395, w57396, w57397, w57398, w57399, w57400, w57401, w57402, w57403, w57404, w57405, w57406, w57407, w57408, w57409, w57410, w57411, w57412, w57413, w57414, w57415, w57416, w57417, w57418, w57419, w57420, w57421, w57422, w57423, w57424, w57425, w57426, w57427, w57428, w57429, w57430, w57431, w57432, w57433, w57434, w57435, w57436, w57437, w57438, w57439, w57440, w57441, w57442, w57443, w57444, w57445, w57446, w57447, w57448, w57449, w57450, w57451, w57452, w57453, w57454, w57455, w57456, w57457, w57458, w57459, w57460, w57461, w57462, w57463, w57464, w57465, w57466, w57467, w57468, w57469, w57470, w57471, w57472, w57473, w57474, w57475, w57476, w57477, w57478, w57479, w57480, w57481, w57482, w57483, w57484, w57485, w57486, w57487, w57488, w57489, w57490, w57491, w57492, w57493, w57494, w57495, w57496, w57497, w57498, w57499, w57500, w57501, w57502, w57503, w57504, w57505, w57506, w57507, w57508, w57509, w57510, w57511, w57512, w57513, w57514, w57515, w57516, w57517, w57518, w57519, w57520, w57521, w57522, w57523, w57524, w57525, w57526, w57527, w57528, w57529, w57530, w57531, w57532, w57533, w57534, w57535, w57536, w57537, w57538, w57539, w57540, w57541, w57542, w57543, w57544, w57545, w57546, w57547, w57548, w57549, w57550, w57551, w57552, w57553, w57554, w57555, w57556, w57557, w57558, w57559, w57560, w57561, w57562, w57563, w57564, w57565, w57566, w57567, w57568, w57569, w57570, w57571, w57572, w57573, w57574, w57575, w57576, w57577, w57578, w57579, w57580, w57581, w57582, w57583, w57584, w57585, w57586, w57587, w57588, w57589, w57590, w57591, w57592, w57593, w57594, w57595, w57596, w57597, w57598, w57599, w57600, w57601, w57602, w57603, w57604, w57605, w57606, w57607, w57608, w57609, w57610, w57611, w57612, w57613, w57614, w57615, w57616, w57617, w57618, w57619, w57620, w57621, w57622, w57623, w57624, w57625, w57626, w57627, w57628, w57629, w57630, w57631, w57632, w57633, w57634, w57635, w57636, w57637, w57638, w57639, w57640, w57641, w57642, w57643, w57644, w57645, w57646, w57647, w57648, w57649, w57650, w57651, w57652, w57653, w57654, w57655, w57656, w57657, w57658, w57659, w57660, w57661, w57662, w57663, w57664, w57665, w57666, w57667, w57668, w57669, w57670, w57671, w57672, w57673, w57674, w57675, w57676, w57677, w57678, w57679, w57680, w57681, w57682, w57683, w57684, w57685, w57686, w57687, w57688, w57689, w57690, w57691, w57692, w57693, w57694, w57695, w57696, w57697, w57698, w57699, w57700, w57701, w57702, w57703, w57704, w57705, w57706, w57707, w57708, w57709, w57710, w57711, w57712, w57713, w57714, w57715, w57716, w57717, w57718, w57719, w57720, w57721, w57722, w57723, w57724, w57725, w57726, w57727, w57728, w57729, w57730, w57731, w57732, w57733, w57734, w57735, w57736, w57737, w57738, w57739, w57740, w57741, w57742, w57743, w57744, w57745, w57746, w57747, w57748, w57749, w57750, w57751, w57752, w57753, w57754, w57755, w57756, w57757, w57758, w57759, w57760, w57761, w57762, w57763, w57764, w57765, w57766, w57767, w57768, w57769, w57770, w57771, w57772, w57773, w57774, w57775, w57776, w57777, w57778, w57779, w57780, w57781, w57782, w57783, w57784, w57785, w57786, w57787, w57788, w57789, w57790, w57791, w57792, w57793, w57794, w57795, w57796, w57797, w57798, w57799, w57800, w57801, w57802, w57803, w57804, w57805, w57806, w57807, w57808, w57809, w57810, w57811, w57812, w57813, w57814, w57815, w57816, w57817, w57818, w57819, w57820, w57821, w57822, w57823, w57824, w57825, w57826, w57827, w57828, w57829, w57830, w57831, w57832, w57833, w57834, w57835, w57836, w57837, w57838, w57839, w57840, w57841, w57842, w57843, w57844, w57845, w57846, w57847, w57848, w57849, w57850, w57851, w57852, w57853, w57854, w57855, w57856, w57857, w57858, w57859, w57860, w57861, w57862, w57863, w57864, w57865, w57866, w57867, w57868, w57869, w57870, w57871, w57872, w57873, w57874, w57875, w57876, w57877, w57878, w57879, w57880, w57881, w57882, w57883, w57884, w57885, w57886, w57887, w57888, w57889, w57890, w57891, w57892, w57893, w57894, w57895, w57896, w57897, w57898, w57899, w57900, w57901, w57902, w57903, w57904, w57905, w57906, w57907, w57908, w57909, w57910, w57911, w57912, w57913, w57914, w57915, w57916, w57917, w57918, w57919, w57920, w57921, w57922, w57923, w57924, w57925, w57926, w57927, w57928, w57929, w57930, w57931, w57932, w57933, w57934, w57935, w57936, w57937, w57938, w57939, w57940, w57941, w57942, w57943, w57944, w57945, w57946, w57947, w57948, w57949, w57950, w57951, w57952, w57953, w57954, w57955, w57956, w57957, w57958, w57959, w57960, w57961, w57962, w57963, w57964, w57965, w57966, w57967, w57968, w57969, w57970, w57971, w57972, w57973, w57974, w57975, w57976, w57977, w57978, w57979, w57980, w57981, w57982, w57983, w57984, w57985, w57986, w57987, w57988, w57989, w57990, w57991, w57992, w57993, w57994, w57995, w57996, w57997, w57998, w57999, w58000, w58001, w58002, w58003, w58004, w58005, w58006, w58007, w58008, w58009, w58010, w58011, w58012, w58013, w58014, w58015, w58016, w58017, w58018, w58019, w58020, w58021, w58022, w58023, w58024, w58025, w58026, w58027, w58028, w58029, w58030, w58031, w58032, w58033, w58034, w58035, w58036, w58037, w58038, w58039, w58040, w58041, w58042, w58043, w58044, w58045, w58046, w58047, w58048, w58049, w58050, w58051, w58052, w58053, w58054, w58055, w58056, w58057, w58058, w58059, w58060, w58061, w58062, w58063, w58064, w58065, w58066, w58067, w58068, w58069, w58070, w58071, w58072, w58073, w58074, w58075, w58076, w58077, w58078, w58079, w58080, w58081, w58082, w58083, w58084, w58085, w58086, w58087, w58088, w58089, w58090, w58091, w58092, w58093, w58094, w58095, w58096, w58097, w58098, w58099, w58100, w58101, w58102, w58103, w58104, w58105, w58106, w58107, w58108, w58109, w58110, w58111, w58112, w58113, w58114, w58115, w58116, w58117, w58118, w58119, w58120, w58121, w58122, w58123, w58124, w58125, w58126, w58127, w58128, w58129, w58130, w58131, w58132, w58133, w58134, w58135, w58136, w58137, w58138, w58139, w58140, w58141, w58142, w58143, w58144, w58145, w58146, w58147, w58148, w58149, w58150, w58151, w58152, w58153, w58154, w58155, w58156, w58157, w58158, w58159, w58160, w58161, w58162, w58163, w58164, w58165, w58166, w58167, w58168, w58169, w58170, w58171, w58172, w58173, w58174, w58175, w58176, w58177, w58178, w58179, w58180, w58181, w58182, w58183, w58184, w58185, w58186, w58187, w58188, w58189, w58190, w58191, w58192, w58193, w58194, w58195, w58196, w58197, w58198, w58199, w58200, w58201, w58202, w58203, w58204, w58205, w58206, w58207, w58208, w58209, w58210, w58211, w58212, w58213, w58214, w58215, w58216, w58217, w58218, w58219, w58220, w58221, w58222, w58223, w58224, w58225, w58226, w58227, w58228, w58229, w58230, w58231, w58232, w58233, w58234, w58235, w58236, w58237, w58238, w58239, w58240, w58241, w58242, w58243, w58244, w58245, w58246, w58247, w58248, w58249, w58250, w58251, w58252, w58253, w58254, w58255, w58256, w58257, w58258, w58259, w58260, w58261, w58262, w58263, w58264, w58265, w58266, w58267, w58268, w58269, w58270, w58271, w58272, w58273, w58274, w58275, w58276, w58277, w58278, w58279, w58280, w58281, w58282, w58283, w58284, w58285, w58286, w58287, w58288, w58289, w58290, w58291, w58292, w58293, w58294, w58295, w58296, w58297, w58298, w58299, w58300, w58301, w58302, w58303, w58304, w58305, w58306, w58307, w58308, w58309, w58310, w58311, w58312, w58313, w58314, w58315, w58316, w58317, w58318, w58319, w58320, w58321, w58322, w58323, w58324, w58325, w58326, w58327, w58328, w58329, w58330, w58331, w58332, w58333, w58334, w58335, w58336, w58337, w58338, w58339, w58340, w58341, w58342, w58343, w58344, w58345, w58346, w58347, w58348, w58349, w58350, w58351, w58352, w58353, w58354, w58355, w58356, w58357, w58358, w58359, w58360, w58361, w58362, w58363, w58364, w58365, w58366, w58367, w58368, w58369, w58370, w58371, w58372, w58373, w58374, w58375, w58376, w58377, w58378, w58379, w58380, w58381, w58382, w58383, w58384, w58385, w58386, w58387, w58388, w58389, w58390, w58391, w58392, w58393, w58394, w58395, w58396, w58397, w58398, w58399, w58400, w58401, w58402, w58403, w58404, w58405, w58406, w58407, w58408, w58409, w58410, w58411, w58412, w58413, w58414, w58415, w58416, w58417, w58418, w58419, w58420, w58421, w58422, w58423, w58424, w58425, w58426, w58427, w58428, w58429, w58430, w58431, w58432, w58433, w58434, w58435, w58436, w58437, w58438, w58439, w58440, w58441, w58442, w58443, w58444, w58445, w58446, w58447, w58448, w58449, w58450, w58451, w58452, w58453, w58454, w58455, w58456, w58457, w58458, w58459, w58460, w58461, w58462, w58463, w58464, w58465, w58466, w58467, w58468, w58469, w58470, w58471, w58472, w58473, w58474, w58475, w58476, w58477, w58478, w58479, w58480, w58481, w58482, w58483, w58484, w58485, w58486, w58487, w58488, w58489, w58490, w58491, w58492, w58493, w58494, w58495, w58496, w58497, w58498, w58499, w58500, w58501, w58502, w58503, w58504, w58505, w58506, w58507, w58508, w58509, w58510, w58511, w58512, w58513, w58514, w58515, w58516, w58517, w58518, w58519, w58520, w58521, w58522, w58523, w58524, w58525, w58526, w58527, w58528, w58529, w58530, w58531, w58532, w58533, w58534, w58535, w58536, w58537, w58538, w58539, w58540, w58541, w58542, w58543, w58544, w58545, w58546, w58547, w58548, w58549, w58550, w58551, w58552, w58553, w58554, w58555, w58556, w58557, w58558, w58559, w58560, w58561, w58562, w58563, w58564, w58565, w58566, w58567, w58568, w58569, w58570, w58571, w58572, w58573, w58574, w58575, w58576, w58577, w58578, w58579, w58580, w58581, w58582, w58583, w58584, w58585, w58586, w58587, w58588, w58589, w58590, w58591, w58592, w58593, w58594, w58595, w58596, w58597, w58598, w58599, w58600, w58601, w58602, w58603, w58604, w58605, w58606, w58607, w58608, w58609, w58610, w58611, w58612, w58613, w58614, w58615, w58616, w58617, w58618, w58619, w58620, w58621, w58622, w58623, w58624, w58625, w58626, w58627, w58628, w58629, w58630, w58631, w58632, w58633, w58634, w58635, w58636, w58637, w58638, w58639, w58640, w58641, w58642, w58643, w58644, w58645, w58646, w58647, w58648, w58649, w58650, w58651, w58652, w58653, w58654, w58655, w58656, w58657, w58658, w58659, w58660, w58661, w58662, w58663, w58664, w58665, w58666, w58667, w58668, w58669, w58670, w58671, w58672, w58673, w58674, w58675, w58676, w58677, w58678, w58679, w58680, w58681, w58682, w58683, w58684, w58685, w58686, w58687, w58688, w58689, w58690, w58691, w58692, w58693, w58694, w58695, w58696, w58697, w58698, w58699, w58700, w58701, w58702, w58703, w58704, w58705, w58706, w58707, w58708, w58709, w58710, w58711, w58712, w58713, w58714, w58715, w58716, w58717, w58718, w58719, w58720, w58721, w58722, w58723, w58724, w58725, w58726, w58727, w58728, w58729, w58730, w58731, w58732, w58733, w58734, w58735, w58736, w58737, w58738, w58739, w58740, w58741, w58742, w58743, w58744, w58745, w58746, w58747, w58748, w58749, w58750, w58751, w58752, w58753, w58754, w58755, w58756, w58757, w58758, w58759, w58760, w58761, w58762, w58763, w58764, w58765, w58766, w58767, w58768, w58769, w58770, w58771, w58772, w58773, w58774, w58775, w58776, w58777, w58778, w58779, w58780, w58781, w58782, w58783, w58784, w58785, w58786, w58787, w58788, w58789, w58790, w58791, w58792, w58793, w58794, w58795, w58796, w58797, w58798, w58799, w58800, w58801, w58802, w58803, w58804, w58805, w58806, w58807, w58808, w58809, w58810, w58811, w58812, w58813, w58814, w58815, w58816, w58817, w58818, w58819, w58820, w58821, w58822, w58823, w58824, w58825, w58826, w58827, w58828, w58829, w58830, w58831, w58832, w58833, w58834, w58835, w58836, w58837, w58838, w58839, w58840, w58841, w58842, w58843, w58844, w58845, w58846, w58847, w58848, w58849, w58850, w58851, w58852, w58853, w58854, w58855, w58856, w58857, w58858, w58859, w58860, w58861, w58862, w58863, w58864, w58865, w58866, w58867, w58868, w58869, w58870, w58871, w58872, w58873, w58874, w58875, w58876, w58877, w58878, w58879, w58880, w58881, w58882, w58883, w58884, w58885, w58886, w58887, w58888, w58889, w58890, w58891, w58892, w58893, w58894, w58895, w58896, w58897, w58898, w58899, w58900, w58901, w58902, w58903, w58904, w58905, w58906, w58907, w58908, w58909, w58910, w58911, w58912, w58913, w58914, w58915, w58916, w58917, w58918, w58919, w58920, w58921, w58922, w58923, w58924, w58925, w58926, w58927, w58928, w58929, w58930, w58931, w58932, w58933, w58934, w58935, w58936, w58937, w58938, w58939, w58940, w58941, w58942, w58943, w58944, w58945, w58946, w58947, w58948, w58949, w58950, w58951, w58952, w58953, w58954, w58955, w58956, w58957, w58958, w58959, w58960, w58961, w58962, w58963, w58964, w58965, w58966, w58967, w58968, w58969, w58970, w58971, w58972, w58973, w58974, w58975, w58976, w58977, w58978, w58979, w58980, w58981, w58982, w58983, w58984, w58985, w58986, w58987, w58988, w58989, w58990, w58991, w58992, w58993, w58994, w58995, w58996, w58997, w58998, w58999, w59000, w59001, w59002, w59003, w59004, w59005, w59006, w59007, w59008, w59009, w59010, w59011, w59012, w59013, w59014, w59015, w59016, w59017, w59018, w59019, w59020, w59021, w59022, w59023, w59024, w59025, w59026, w59027, w59028, w59029, w59030, w59031, w59032, w59033, w59034, w59035, w59036, w59037, w59038, w59039, w59040, w59041, w59042, w59043, w59044, w59045, w59046, w59047, w59048, w59049, w59050, w59051, w59052, w59053, w59054, w59055, w59056, w59057, w59058, w59059, w59060, w59061, w59062, w59063, w59064, w59065, w59066, w59067, w59068, w59069, w59070, w59071, w59072, w59073, w59074, w59075, w59076, w59077, w59078, w59079, w59080, w59081, w59082, w59083, w59084, w59085, w59086, w59087, w59088, w59089, w59090, w59091, w59092, w59093, w59094, w59095, w59096, w59097, w59098, w59099, w59100, w59101, w59102, w59103, w59104, w59105, w59106, w59107, w59108, w59109, w59110, w59111, w59112, w59113, w59114, w59115, w59116, w59117, w59118, w59119, w59120, w59121, w59122, w59123, w59124, w59125, w59126, w59127, w59128, w59129, w59130, w59131, w59132, w59133, w59134, w59135, w59136, w59137, w59138, w59139, w59140, w59141, w59142, w59143, w59144, w59145, w59146, w59147, w59148, w59149, w59150, w59151, w59152, w59153, w59154, w59155, w59156, w59157, w59158, w59159, w59160, w59161, w59162, w59163, w59164, w59165, w59166, w59167, w59168, w59169, w59170, w59171, w59172, w59173, w59174, w59175, w59176, w59177, w59178, w59179, w59180, w59181, w59182, w59183, w59184, w59185, w59186, w59187, w59188, w59189, w59190, w59191, w59192, w59193, w59194, w59195, w59196, w59197, w59198, w59199, w59200, w59201, w59202, w59203, w59204, w59205, w59206, w59207, w59208, w59209, w59210, w59211, w59212, w59213, w59214, w59215, w59216, w59217, w59218, w59219, w59220, w59221, w59222, w59223, w59224, w59225, w59226, w59227, w59228, w59229, w59230, w59231, w59232, w59233, w59234, w59235, w59236, w59237, w59238, w59239, w59240, w59241, w59242, w59243, w59244, w59245, w59246, w59247, w59248, w59249, w59250, w59251, w59252, w59253, w59254, w59255, w59256, w59257, w59258, w59259, w59260, w59261, w59262, w59263, w59264, w59265, w59266, w59267, w59268, w59269, w59270, w59271, w59272, w59273, w59274, w59275, w59276, w59277, w59278, w59279, w59280, w59281, w59282, w59283, w59284, w59285, w59286, w59287, w59288, w59289, w59290, w59291, w59292, w59293, w59294, w59295, w59296, w59297, w59298, w59299, w59300, w59301, w59302, w59303, w59304, w59305, w59306, w59307, w59308, w59309, w59310, w59311, w59312, w59313, w59314, w59315, w59316, w59317, w59318, w59319, w59320, w59321, w59322, w59323, w59324, w59325, w59326, w59327, w59328, w59329, w59330, w59331, w59332, w59333, w59334, w59335, w59336, w59337, w59338, w59339, w59340, w59341, w59342, w59343, w59344, w59345, w59346, w59347, w59348, w59349, w59350, w59351, w59352, w59353, w59354, w59355, w59356, w59357, w59358, w59359, w59360, w59361, w59362, w59363, w59364, w59365, w59366, w59367, w59368, w59369, w59370, w59371, w59372, w59373, w59374, w59375, w59376, w59377, w59378, w59379, w59380, w59381, w59382, w59383, w59384, w59385, w59386, w59387, w59388, w59389, w59390, w59391, w59392, w59393, w59394, w59395, w59396, w59397, w59398, w59399, w59400, w59401, w59402, w59403, w59404, w59405, w59406, w59407, w59408, w59409, w59410, w59411, w59412, w59413, w59414, w59415, w59416, w59417, w59418, w59419, w59420, w59421, w59422, w59423, w59424, w59425, w59426, w59427, w59428, w59429, w59430, w59431, w59432, w59433, w59434, w59435, w59436, w59437, w59438, w59439, w59440, w59441, w59442, w59443, w59444, w59445, w59446, w59447, w59448, w59449, w59450, w59451, w59452, w59453, w59454, w59455, w59456, w59457, w59458, w59459, w59460, w59461, w59462, w59463, w59464, w59465, w59466, w59467, w59468, w59469, w59470, w59471, w59472, w59473, w59474, w59475, w59476, w59477, w59478, w59479, w59480, w59481, w59482, w59483, w59484, w59485, w59486, w59487, w59488, w59489, w59490, w59491, w59492, w59493, w59494, w59495, w59496, w59497, w59498, w59499, w59500, w59501, w59502, w59503, w59504, w59505, w59506, w59507, w59508, w59509, w59510, w59511, w59512, w59513, w59514, w59515, w59516, w59517, w59518, w59519, w59520, w59521, w59522, w59523, w59524, w59525, w59526, w59527, w59528, w59529, w59530, w59531, w59532, w59533, w59534, w59535, w59536, w59537, w59538, w59539, w59540, w59541, w59542, w59543, w59544, w59545, w59546, w59547, w59548, w59549, w59550, w59551, w59552, w59553, w59554, w59555, w59556, w59557, w59558, w59559, w59560, w59561, w59562, w59563, w59564, w59565, w59566, w59567, w59568, w59569, w59570, w59571, w59572, w59573, w59574, w59575, w59576, w59577, w59578, w59579, w59580, w59581, w59582, w59583, w59584, w59585, w59586, w59587, w59588, w59589, w59590, w59591, w59592, w59593, w59594, w59595, w59596, w59597, w59598, w59599, w59600, w59601, w59602, w59603, w59604, w59605, w59606, w59607, w59608, w59609, w59610, w59611, w59612, w59613, w59614, w59615, w59616, w59617, w59618, w59619, w59620, w59621, w59622, w59623, w59624, w59625, w59626, w59627, w59628, w59629, w59630, w59631, w59632, w59633, w59634, w59635, w59636, w59637, w59638, w59639, w59640, w59641, w59642, w59643, w59644, w59645, w59646, w59647, w59648, w59649, w59650, w59651, w59652, w59653, w59654, w59655, w59656, w59657, w59658, w59659, w59660, w59661, w59662, w59663, w59664, w59665, w59666, w59667, w59668, w59669, w59670, w59671, w59672, w59673, w59674, w59675, w59676, w59677, w59678, w59679, w59680, w59681, w59682, w59683, w59684, w59685, w59686, w59687, w59688, w59689, w59690, w59691, w59692, w59693, w59694, w59695, w59696, w59697, w59698, w59699, w59700, w59701, w59702, w59703, w59704, w59705, w59706, w59707, w59708, w59709, w59710, w59711, w59712, w59713, w59714, w59715, w59716, w59717, w59718, w59719, w59720, w59721, w59722, w59723, w59724, w59725, w59726, w59727, w59728, w59729, w59730, w59731, w59732, w59733, w59734, w59735, w59736, w59737, w59738, w59739, w59740, w59741, w59742, w59743, w59744, w59745, w59746, w59747, w59748, w59749, w59750, w59751, w59752, w59753, w59754, w59755, w59756, w59757, w59758, w59759, w59760, w59761, w59762, w59763, w59764, w59765, w59766, w59767, w59768, w59769, w59770, w59771, w59772, w59773, w59774, w59775, w59776, w59777, w59778, w59779, w59780, w59781, w59782, w59783, w59784, w59785, w59786, w59787, w59788, w59789, w59790, w59791, w59792, w59793, w59794, w59795, w59796, w59797, w59798, w59799, w59800, w59801, w59802, w59803, w59804, w59805, w59806, w59807, w59808, w59809, w59810, w59811, w59812, w59813, w59814, w59815, w59816, w59817, w59818, w59819, w59820, w59821, w59822, w59823, w59824, w59825, w59826, w59827, w59828, w59829, w59830, w59831, w59832, w59833, w59834, w59835, w59836, w59837, w59838, w59839, w59840, w59841, w59842, w59843, w59844, w59845, w59846, w59847, w59848, w59849, w59850, w59851, w59852, w59853, w59854, w59855, w59856, w59857, w59858, w59859, w59860, w59861, w59862, w59863, w59864, w59865, w59866, w59867, w59868, w59869, w59870, w59871, w59872, w59873, w59874, w59875, w59876, w59877, w59878, w59879, w59880, w59881, w59882, w59883, w59884, w59885, w59886, w59887, w59888, w59889, w59890, w59891, w59892, w59893, w59894, w59895, w59896, w59897, w59898, w59899, w59900, w59901, w59902, w59903, w59904, w59905, w59906, w59907, w59908, w59909, w59910, w59911, w59912, w59913, w59914, w59915, w59916, w59917, w59918, w59919, w59920, w59921, w59922, w59923, w59924, w59925, w59926, w59927, w59928, w59929, w59930, w59931, w59932, w59933, w59934, w59935, w59936, w59937, w59938, w59939, w59940, w59941, w59942, w59943, w59944, w59945, w59946, w59947, w59948, w59949, w59950, w59951, w59952, w59953, w59954, w59955, w59956, w59957, w59958, w59959, w59960, w59961, w59962, w59963, w59964, w59965, w59966, w59967, w59968, w59969, w59970, w59971, w59972, w59973, w59974, w59975, w59976, w59977, w59978, w59979, w59980, w59981, w59982, w59983, w59984, w59985, w59986, w59987, w59988, w59989, w59990, w59991, w59992, w59993, w59994, w59995, w59996, w59997, w59998, w59999, w60000, w60001, w60002, w60003, w60004, w60005, w60006, w60007, w60008, w60009, w60010, w60011, w60012, w60013, w60014, w60015, w60016, w60017, w60018, w60019, w60020, w60021, w60022, w60023, w60024, w60025, w60026, w60027, w60028, w60029, w60030, w60031, w60032, w60033, w60034, w60035, w60036, w60037, w60038, w60039, w60040, w60041, w60042, w60043, w60044, w60045, w60046, w60047, w60048, w60049, w60050, w60051, w60052, w60053, w60054, w60055, w60056, w60057, w60058, w60059, w60060, w60061, w60062, w60063, w60064, w60065, w60066, w60067, w60068, w60069, w60070, w60071, w60072, w60073, w60074, w60075, w60076, w60077, w60078, w60079, w60080, w60081, w60082, w60083, w60084, w60085, w60086, w60087, w60088, w60089, w60090, w60091, w60092, w60093, w60094, w60095, w60096, w60097, w60098, w60099, w60100, w60101, w60102, w60103, w60104, w60105, w60106, w60107, w60108, w60109, w60110, w60111, w60112, w60113, w60114, w60115, w60116, w60117, w60118, w60119, w60120, w60121, w60122, w60123, w60124, w60125, w60126, w60127, w60128, w60129, w60130, w60131, w60132, w60133, w60134, w60135, w60136, w60137, w60138, w60139, w60140, w60141, w60142, w60143, w60144, w60145, w60146, w60147, w60148, w60149, w60150, w60151, w60152, w60153, w60154, w60155, w60156, w60157, w60158, w60159, w60160, w60161, w60162, w60163, w60164, w60165, w60166, w60167, w60168, w60169, w60170, w60171, w60172, w60173, w60174, w60175, w60176, w60177, w60178, w60179, w60180, w60181, w60182, w60183, w60184, w60185, w60186, w60187, w60188, w60189, w60190, w60191, w60192, w60193, w60194, w60195, w60196, w60197, w60198, w60199, w60200, w60201, w60202, w60203, w60204, w60205, w60206, w60207, w60208, w60209, w60210, w60211, w60212, w60213, w60214, w60215, w60216, w60217, w60218, w60219, w60220, w60221, w60222, w60223, w60224, w60225, w60226, w60227, w60228, w60229, w60230, w60231, w60232, w60233, w60234, w60235, w60236, w60237, w60238, w60239, w60240, w60241, w60242, w60243, w60244, w60245, w60246, w60247, w60248, w60249, w60250, w60251, w60252, w60253, w60254, w60255, w60256, w60257, w60258, w60259, w60260, w60261, w60262, w60263, w60264, w60265, w60266, w60267, w60268, w60269, w60270, w60271, w60272, w60273, w60274, w60275, w60276, w60277, w60278, w60279, w60280, w60281, w60282, w60283, w60284, w60285, w60286, w60287, w60288, w60289, w60290, w60291, w60292, w60293, w60294, w60295, w60296, w60297, w60298, w60299, w60300, w60301, w60302, w60303, w60304, w60305, w60306, w60307, w60308, w60309, w60310, w60311, w60312, w60313, w60314, w60315, w60316, w60317, w60318, w60319, w60320, w60321, w60322, w60323, w60324, w60325, w60326, w60327, w60328, w60329, w60330, w60331, w60332, w60333, w60334, w60335, w60336, w60337, w60338, w60339, w60340, w60341, w60342, w60343, w60344, w60345, w60346, w60347, w60348, w60349, w60350, w60351, w60352, w60353, w60354, w60355, w60356, w60357, w60358, w60359, w60360, w60361, w60362, w60363, w60364, w60365, w60366, w60367, w60368, w60369, w60370, w60371, w60372, w60373, w60374, w60375, w60376, w60377, w60378, w60379, w60380, w60381, w60382, w60383, w60384, w60385, w60386, w60387, w60388, w60389, w60390, w60391, w60392, w60393, w60394, w60395, w60396, w60397, w60398, w60399, w60400, w60401, w60402, w60403, w60404, w60405, w60406, w60407, w60408, w60409, w60410, w60411, w60412, w60413, w60414, w60415, w60416, w60417, w60418, w60419, w60420, w60421, w60422, w60423, w60424, w60425, w60426, w60427, w60428, w60429, w60430, w60431, w60432, w60433, w60434, w60435, w60436, w60437, w60438, w60439, w60440, w60441, w60442, w60443, w60444, w60445, w60446, w60447, w60448, w60449, w60450, w60451, w60452, w60453, w60454, w60455, w60456, w60457, w60458, w60459, w60460, w60461, w60462, w60463, w60464, w60465, w60466, w60467, w60468, w60469, w60470, w60471, w60472, w60473, w60474, w60475, w60476, w60477, w60478, w60479, w60480, w60481, w60482, w60483, w60484, w60485, w60486, w60487, w60488, w60489, w60490, w60491, w60492, w60493, w60494, w60495, w60496, w60497, w60498, w60499, w60500, w60501, w60502, w60503, w60504, w60505, w60506, w60507, w60508, w60509, w60510, w60511, w60512, w60513, w60514, w60515, w60516, w60517, w60518, w60519, w60520, w60521, w60522, w60523, w60524, w60525, w60526, w60527, w60528, w60529, w60530, w60531, w60532, w60533, w60534, w60535, w60536, w60537, w60538, w60539, w60540, w60541, w60542, w60543, w60544, w60545, w60546, w60547, w60548, w60549, w60550, w60551, w60552, w60553, w60554, w60555, w60556, w60557, w60558, w60559, w60560, w60561, w60562, w60563, w60564, w60565, w60566, w60567, w60568, w60569, w60570, w60571, w60572, w60573, w60574, w60575, w60576, w60577, w60578, w60579, w60580, w60581, w60582, w60583, w60584, w60585, w60586, w60587, w60588, w60589, w60590, w60591, w60592, w60593, w60594, w60595, w60596, w60597, w60598, w60599, w60600, w60601, w60602, w60603, w60604, w60605, w60606, w60607, w60608, w60609, w60610, w60611, w60612, w60613, w60614, w60615, w60616, w60617, w60618, w60619, w60620, w60621, w60622, w60623, w60624, w60625, w60626, w60627, w60628, w60629, w60630, w60631, w60632, w60633, w60634, w60635, w60636, w60637, w60638, w60639, w60640, w60641, w60642, w60643, w60644, w60645, w60646, w60647, w60648, w60649, w60650, w60651, w60652, w60653, w60654, w60655, w60656, w60657, w60658, w60659, w60660, w60661, w60662, w60663, w60664, w60665, w60666, w60667, w60668, w60669, w60670, w60671, w60672, w60673, w60674, w60675, w60676, w60677, w60678, w60679, w60680, w60681, w60682, w60683, w60684, w60685, w60686, w60687, w60688, w60689, w60690, w60691, w60692, w60693, w60694, w60695, w60696, w60697, w60698, w60699, w60700, w60701, w60702, w60703, w60704, w60705, w60706, w60707, w60708, w60709, w60710, w60711, w60712, w60713, w60714, w60715, w60716, w60717, w60718, w60719, w60720, w60721, w60722, w60723, w60724, w60725, w60726, w60727, w60728, w60729, w60730, w60731, w60732, w60733, w60734, w60735, w60736, w60737, w60738, w60739, w60740, w60741, w60742, w60743, w60744, w60745, w60746, w60747, w60748, w60749, w60750, w60751, w60752, w60753, w60754, w60755, w60756, w60757, w60758, w60759, w60760, w60761, w60762, w60763, w60764, w60765, w60766, w60767, w60768, w60769, w60770, w60771, w60772, w60773, w60774, w60775, w60776, w60777, w60778, w60779, w60780, w60781, w60782, w60783, w60784, w60785, w60786, w60787, w60788, w60789, w60790, w60791, w60792, w60793, w60794, w60795, w60796, w60797, w60798, w60799, w60800, w60801, w60802, w60803, w60804, w60805, w60806, w60807, w60808, w60809, w60810, w60811, w60812, w60813, w60814, w60815, w60816, w60817, w60818, w60819, w60820, w60821, w60822, w60823, w60824, w60825, w60826, w60827, w60828, w60829, w60830, w60831, w60832, w60833, w60834, w60835, w60836, w60837, w60838, w60839, w60840, w60841, w60842, w60843, w60844, w60845, w60846, w60847, w60848, w60849, w60850, w60851, w60852, w60853, w60854, w60855, w60856, w60857, w60858, w60859, w60860, w60861, w60862, w60863, w60864, w60865, w60866, w60867, w60868, w60869, w60870, w60871, w60872, w60873, w60874, w60875, w60876, w60877, w60878, w60879, w60880, w60881, w60882, w60883, w60884, w60885, w60886, w60887, w60888, w60889, w60890, w60891, w60892, w60893, w60894, w60895, w60896, w60897, w60898, w60899, w60900, w60901, w60902, w60903, w60904, w60905, w60906, w60907, w60908, w60909, w60910, w60911, w60912, w60913, w60914, w60915, w60916, w60917, w60918, w60919, w60920, w60921, w60922, w60923, w60924, w60925, w60926, w60927, w60928, w60929, w60930, w60931, w60932, w60933, w60934, w60935, w60936, w60937, w60938, w60939, w60940, w60941, w60942, w60943, w60944, w60945, w60946, w60947, w60948, w60949, w60950, w60951, w60952, w60953, w60954, w60955, w60956, w60957, w60958, w60959, w60960, w60961, w60962, w60963, w60964, w60965, w60966, w60967, w60968, w60969, w60970, w60971, w60972, w60973, w60974, w60975, w60976, w60977, w60978, w60979, w60980, w60981, w60982, w60983, w60984, w60985, w60986, w60987, w60988, w60989, w60990, w60991, w60992, w60993, w60994, w60995, w60996, w60997, w60998, w60999, w61000, w61001, w61002, w61003, w61004, w61005, w61006, w61007, w61008, w61009, w61010, w61011, w61012, w61013, w61014, w61015, w61016, w61017, w61018, w61019, w61020, w61021, w61022, w61023, w61024, w61025, w61026, w61027, w61028, w61029, w61030, w61031, w61032, w61033, w61034, w61035, w61036, w61037, w61038, w61039, w61040, w61041, w61042, w61043, w61044, w61045, w61046, w61047, w61048, w61049, w61050, w61051, w61052, w61053, w61054, w61055, w61056, w61057, w61058, w61059, w61060, w61061, w61062, w61063, w61064, w61065, w61066, w61067, w61068, w61069, w61070, w61071, w61072, w61073, w61074, w61075, w61076, w61077, w61078, w61079, w61080, w61081, w61082, w61083, w61084, w61085, w61086, w61087, w61088, w61089, w61090, w61091, w61092, w61093, w61094, w61095, w61096, w61097, w61098, w61099, w61100, w61101, w61102, w61103, w61104, w61105, w61106, w61107, w61108, w61109, w61110, w61111, w61112, w61113, w61114, w61115, w61116, w61117, w61118, w61119, w61120, w61121, w61122, w61123, w61124, w61125, w61126, w61127, w61128, w61129, w61130, w61131, w61132, w61133, w61134, w61135, w61136, w61137, w61138, w61139, w61140, w61141, w61142, w61143, w61144, w61145, w61146, w61147, w61148, w61149, w61150, w61151, w61152, w61153, w61154, w61155, w61156, w61157, w61158, w61159, w61160, w61161, w61162, w61163, w61164, w61165, w61166, w61167, w61168, w61169, w61170, w61171, w61172, w61173, w61174, w61175, w61176, w61177, w61178, w61179, w61180, w61181, w61182, w61183, w61184, w61185, w61186, w61187, w61188, w61189, w61190, w61191, w61192, w61193, w61194, w61195, w61196, w61197, w61198, w61199, w61200, w61201, w61202, w61203, w61204, w61205, w61206, w61207, w61208, w61209, w61210, w61211, w61212, w61213, w61214, w61215, w61216, w61217, w61218, w61219, w61220, w61221, w61222, w61223, w61224, w61225, w61226, w61227, w61228, w61229, w61230, w61231, w61232, w61233, w61234, w61235, w61236, w61237, w61238, w61239, w61240, w61241, w61242, w61243, w61244, w61245, w61246, w61247, w61248, w61249, w61250, w61251, w61252, w61253, w61254, w61255, w61256, w61257, w61258, w61259, w61260, w61261, w61262, w61263, w61264, w61265, w61266, w61267, w61268, w61269, w61270, w61271, w61272, w61273, w61274, w61275, w61276, w61277, w61278, w61279, w61280, w61281, w61282, w61283, w61284, w61285, w61286, w61287, w61288, w61289, w61290, w61291, w61292, w61293, w61294, w61295, w61296, w61297, w61298, w61299, w61300, w61301, w61302, w61303, w61304, w61305, w61306, w61307, w61308, w61309, w61310, w61311, w61312, w61313, w61314, w61315, w61316, w61317, w61318, w61319, w61320, w61321, w61322, w61323, w61324, w61325, w61326, w61327, w61328, w61329, w61330, w61331, w61332, w61333, w61334, w61335, w61336, w61337, w61338, w61339, w61340, w61341, w61342, w61343, w61344, w61345, w61346, w61347, w61348, w61349, w61350, w61351, w61352, w61353, w61354, w61355, w61356, w61357, w61358, w61359, w61360, w61361, w61362, w61363, w61364, w61365, w61366, w61367, w61368, w61369, w61370, w61371, w61372, w61373, w61374, w61375, w61376, w61377, w61378, w61379, w61380, w61381, w61382, w61383, w61384, w61385, w61386, w61387, w61388, w61389, w61390, w61391, w61392, w61393, w61394, w61395, w61396, w61397, w61398, w61399, w61400, w61401, w61402, w61403, w61404, w61405, w61406, w61407, w61408, w61409, w61410, w61411, w61412, w61413, w61414, w61415, w61416, w61417, w61418, w61419, w61420, w61421, w61422, w61423, w61424, w61425, w61426, w61427, w61428, w61429, w61430, w61431, w61432, w61433, w61434, w61435, w61436, w61437, w61438, w61439, w61440, w61441, w61442, w61443, w61444, w61445, w61446, w61447, w61448, w61449, w61450, w61451, w61452, w61453, w61454, w61455, w61456, w61457, w61458, w61459, w61460, w61461, w61462, w61463, w61464, w61465, w61466, w61467, w61468, w61469, w61470, w61471, w61472, w61473, w61474, w61475, w61476, w61477, w61478, w61479, w61480, w61481, w61482, w61483, w61484, w61485, w61486, w61487, w61488, w61489, w61490, w61491, w61492, w61493, w61494, w61495, w61496, w61497, w61498, w61499, w61500, w61501, w61502, w61503, w61504, w61505, w61506, w61507, w61508, w61509, w61510, w61511, w61512, w61513, w61514, w61515, w61516, w61517, w61518, w61519, w61520, w61521, w61522, w61523, w61524, w61525, w61526, w61527, w61528, w61529, w61530, w61531, w61532, w61533, w61534, w61535, w61536, w61537, w61538, w61539, w61540, w61541, w61542, w61543, w61544, w61545, w61546, w61547, w61548, w61549, w61550, w61551, w61552, w61553, w61554, w61555, w61556, w61557, w61558, w61559, w61560, w61561, w61562, w61563, w61564, w61565, w61566, w61567, w61568, w61569, w61570, w61571, w61572, w61573, w61574, w61575, w61576, w61577, w61578, w61579, w61580, w61581, w61582, w61583, w61584, w61585, w61586, w61587, w61588, w61589, w61590, w61591, w61592, w61593, w61594, w61595, w61596, w61597, w61598, w61599, w61600, w61601, w61602, w61603, w61604, w61605, w61606, w61607, w61608, w61609, w61610, w61611, w61612, w61613, w61614, w61615, w61616, w61617, w61618, w61619, w61620, w61621, w61622, w61623, w61624, w61625, w61626, w61627, w61628, w61629, w61630, w61631, w61632, w61633, w61634, w61635, w61636, w61637, w61638, w61639, w61640, w61641, w61642, w61643, w61644, w61645, w61646, w61647, w61648, w61649, w61650, w61651, w61652, w61653, w61654, w61655, w61656, w61657, w61658, w61659, w61660, w61661, w61662, w61663, w61664, w61665, w61666, w61667, w61668, w61669, w61670, w61671, w61672, w61673, w61674, w61675, w61676, w61677, w61678, w61679, w61680, w61681, w61682, w61683, w61684, w61685, w61686, w61687, w61688, w61689, w61690, w61691, w61692, w61693, w61694, w61695, w61696, w61697, w61698, w61699, w61700, w61701, w61702, w61703, w61704, w61705, w61706, w61707, w61708, w61709, w61710, w61711, w61712, w61713, w61714, w61715, w61716, w61717, w61718, w61719, w61720, w61721, w61722, w61723, w61724, w61725, w61726, w61727, w61728, w61729, w61730, w61731, w61732, w61733, w61734, w61735, w61736, w61737, w61738, w61739, w61740, w61741, w61742, w61743, w61744, w61745, w61746, w61747, w61748, w61749, w61750, w61751, w61752, w61753, w61754, w61755, w61756, w61757, w61758, w61759, w61760, w61761, w61762, w61763, w61764, w61765, w61766, w61767, w61768, w61769, w61770, w61771, w61772, w61773, w61774, w61775, w61776, w61777, w61778, w61779, w61780, w61781, w61782, w61783, w61784, w61785, w61786, w61787, w61788, w61789, w61790, w61791, w61792, w61793, w61794, w61795, w61796, w61797, w61798, w61799, w61800, w61801, w61802, w61803, w61804, w61805, w61806, w61807, w61808, w61809, w61810, w61811, w61812, w61813, w61814, w61815, w61816, w61817, w61818, w61819, w61820, w61821, w61822, w61823, w61824, w61825, w61826, w61827, w61828, w61829, w61830, w61831, w61832, w61833, w61834, w61835, w61836, w61837, w61838, w61839, w61840, w61841, w61842, w61843, w61844, w61845, w61846, w61847, w61848, w61849, w61850, w61851, w61852, w61853, w61854, w61855, w61856, w61857, w61858, w61859, w61860, w61861, w61862, w61863, w61864, w61865, w61866, w61867, w61868, w61869, w61870, w61871, w61872, w61873, w61874, w61875, w61876, w61877, w61878, w61879, w61880, w61881, w61882, w61883, w61884, w61885, w61886, w61887, w61888, w61889, w61890, w61891, w61892, w61893, w61894, w61895, w61896, w61897, w61898, w61899, w61900, w61901, w61902, w61903, w61904, w61905, w61906, w61907, w61908, w61909, w61910, w61911, w61912, w61913, w61914, w61915, w61916, w61917, w61918, w61919, w61920, w61921, w61922, w61923, w61924, w61925, w61926, w61927, w61928, w61929, w61930, w61931, w61932, w61933, w61934, w61935, w61936, w61937, w61938, w61939, w61940, w61941, w61942, w61943, w61944, w61945, w61946, w61947, w61948, w61949, w61950, w61951, w61952, w61953, w61954, w61955, w61956, w61957, w61958, w61959, w61960, w61961, w61962, w61963, w61964, w61965, w61966, w61967, w61968, w61969, w61970, w61971, w61972, w61973, w61974, w61975, w61976, w61977, w61978, w61979, w61980, w61981, w61982, w61983, w61984, w61985, w61986, w61987, w61988, w61989, w61990, w61991, w61992, w61993, w61994, w61995, w61996, w61997, w61998, w61999, w62000, w62001, w62002, w62003, w62004, w62005, w62006, w62007, w62008, w62009, w62010, w62011, w62012, w62013, w62014, w62015, w62016, w62017, w62018, w62019, w62020, w62021, w62022, w62023, w62024, w62025, w62026, w62027, w62028, w62029, w62030, w62031, w62032, w62033, w62034, w62035, w62036, w62037, w62038, w62039, w62040, w62041, w62042, w62043, w62044, w62045, w62046, w62047, w62048, w62049, w62050, w62051, w62052, w62053, w62054, w62055, w62056, w62057, w62058, w62059, w62060, w62061, w62062, w62063, w62064, w62065, w62066, w62067, w62068, w62069, w62070, w62071, w62072, w62073, w62074, w62075, w62076, w62077, w62078, w62079, w62080, w62081, w62082, w62083, w62084, w62085, w62086, w62087, w62088, w62089, w62090, w62091, w62092, w62093, w62094, w62095, w62096, w62097, w62098, w62099, w62100, w62101, w62102, w62103, w62104, w62105, w62106, w62107, w62108, w62109, w62110, w62111, w62112, w62113, w62114, w62115, w62116, w62117, w62118, w62119, w62120, w62121, w62122, w62123, w62124, w62125, w62126, w62127, w62128, w62129, w62130, w62131, w62132, w62133, w62134, w62135, w62136, w62137, w62138, w62139, w62140, w62141, w62142, w62143, w62144, w62145, w62146, w62147, w62148, w62149, w62150, w62151, w62152, w62153, w62154, w62155, w62156, w62157, w62158, w62159, w62160, w62161, w62162, w62163, w62164, w62165, w62166, w62167, w62168, w62169, w62170, w62171, w62172, w62173, w62174, w62175, w62176, w62177, w62178, w62179, w62180, w62181, w62182, w62183, w62184, w62185, w62186, w62187, w62188, w62189, w62190, w62191, w62192, w62193, w62194, w62195, w62196, w62197, w62198, w62199, w62200, w62201, w62202, w62203, w62204, w62205, w62206, w62207, w62208, w62209, w62210, w62211, w62212, w62213, w62214, w62215, w62216, w62217, w62218, w62219, w62220, w62221, w62222, w62223, w62224, w62225, w62226, w62227, w62228, w62229, w62230, w62231, w62232, w62233, w62234, w62235, w62236, w62237, w62238, w62239, w62240, w62241, w62242, w62243, w62244, w62245, w62246, w62247, w62248, w62249, w62250, w62251, w62252, w62253, w62254, w62255, w62256, w62257, w62258, w62259, w62260, w62261, w62262, w62263, w62264, w62265, w62266, w62267, w62268, w62269, w62270, w62271, w62272, w62273, w62274, w62275, w62276, w62277, w62278, w62279, w62280, w62281, w62282, w62283, w62284, w62285, w62286, w62287, w62288, w62289, w62290, w62291, w62292, w62293, w62294, w62295, w62296, w62297, w62298, w62299, w62300, w62301, w62302, w62303, w62304, w62305, w62306, w62307, w62308, w62309, w62310, w62311, w62312, w62313, w62314, w62315, w62316, w62317, w62318, w62319, w62320, w62321, w62322, w62323, w62324, w62325, w62326, w62327, w62328, w62329, w62330, w62331, w62332, w62333, w62334, w62335, w62336, w62337, w62338, w62339, w62340, w62341, w62342, w62343, w62344, w62345, w62346, w62347, w62348, w62349, w62350, w62351, w62352, w62353, w62354, w62355, w62356, w62357, w62358, w62359, w62360, w62361, w62362, w62363, w62364, w62365, w62366, w62367, w62368, w62369, w62370, w62371, w62372, w62373, w62374, w62375, w62376, w62377, w62378, w62379, w62380, w62381, w62382, w62383, w62384, w62385, w62386, w62387, w62388, w62389, w62390, w62391, w62392, w62393, w62394, w62395, w62396, w62397, w62398, w62399, w62400, w62401, w62402, w62403, w62404, w62405, w62406, w62407, w62408, w62409, w62410, w62411, w62412, w62413, w62414, w62415, w62416, w62417, w62418, w62419, w62420, w62421, w62422, w62423, w62424, w62425, w62426, w62427, w62428, w62429, w62430, w62431, w62432, w62433, w62434, w62435, w62436, w62437, w62438, w62439, w62440, w62441, w62442, w62443, w62444, w62445, w62446, w62447, w62448, w62449, w62450, w62451, w62452, w62453, w62454, w62455, w62456, w62457, w62458, w62459, w62460, w62461, w62462, w62463, w62464, w62465, w62466, w62467, w62468, w62469, w62470, w62471, w62472, w62473, w62474, w62475, w62476, w62477, w62478, w62479, w62480, w62481, w62482, w62483, w62484, w62485, w62486, w62487, w62488, w62489, w62490, w62491, w62492, w62493, w62494, w62495, w62496, w62497, w62498, w62499, w62500, w62501, w62502, w62503, w62504, w62505, w62506, w62507, w62508, w62509, w62510, w62511, w62512, w62513, w62514, w62515, w62516, w62517, w62518, w62519, w62520, w62521, w62522, w62523, w62524, w62525, w62526, w62527, w62528, w62529, w62530, w62531, w62532, w62533, w62534, w62535, w62536, w62537, w62538, w62539, w62540, w62541, w62542, w62543, w62544, w62545, w62546, w62547, w62548, w62549, w62550, w62551, w62552, w62553, w62554, w62555, w62556, w62557, w62558, w62559, w62560, w62561, w62562, w62563, w62564, w62565, w62566, w62567, w62568, w62569, w62570, w62571, w62572, w62573, w62574, w62575, w62576, w62577, w62578, w62579, w62580, w62581, w62582, w62583, w62584, w62585, w62586, w62587, w62588, w62589, w62590, w62591, w62592, w62593, w62594, w62595, w62596, w62597, w62598, w62599, w62600, w62601, w62602, w62603, w62604, w62605, w62606, w62607, w62608, w62609, w62610, w62611, w62612, w62613, w62614, w62615, w62616, w62617, w62618, w62619, w62620, w62621, w62622, w62623, w62624, w62625, w62626, w62627, w62628, w62629, w62630, w62631, w62632, w62633, w62634, w62635, w62636, w62637, w62638, w62639, w62640, w62641, w62642, w62643, w62644, w62645, w62646, w62647, w62648, w62649, w62650, w62651, w62652, w62653, w62654, w62655, w62656, w62657, w62658, w62659, w62660, w62661, w62662, w62663, w62664, w62665, w62666, w62667, w62668, w62669, w62670, w62671, w62672, w62673, w62674, w62675, w62676, w62677, w62678, w62679, w62680, w62681, w62682, w62683, w62684, w62685, w62686, w62687, w62688, w62689, w62690, w62691, w62692, w62693, w62694, w62695, w62696, w62697, w62698, w62699, w62700, w62701, w62702, w62703, w62704, w62705, w62706, w62707, w62708, w62709, w62710, w62711, w62712, w62713, w62714, w62715, w62716, w62717, w62718, w62719, w62720, w62721, w62722, w62723, w62724, w62725, w62726, w62727, w62728, w62729, w62730, w62731, w62732, w62733, w62734, w62735, w62736, w62737, w62738, w62739, w62740, w62741, w62742, w62743, w62744, w62745, w62746, w62747, w62748, w62749, w62750, w62751, w62752, w62753, w62754, w62755, w62756, w62757, w62758, w62759, w62760, w62761, w62762, w62763, w62764, w62765, w62766, w62767, w62768, w62769, w62770, w62771, w62772, w62773, w62774, w62775, w62776, w62777, w62778, w62779, w62780, w62781, w62782, w62783, w62784, w62785, w62786, w62787, w62788, w62789, w62790, w62791, w62792, w62793, w62794, w62795, w62796, w62797, w62798, w62799, w62800, w62801, w62802, w62803, w62804, w62805, w62806, w62807, w62808, w62809, w62810, w62811, w62812, w62813, w62814, w62815, w62816, w62817, w62818, w62819, w62820, w62821, w62822, w62823, w62824, w62825, w62826, w62827, w62828, w62829, w62830, w62831, w62832, w62833, w62834, w62835, w62836, w62837, w62838, w62839, w62840, w62841, w62842, w62843, w62844, w62845, w62846, w62847, w62848, w62849, w62850, w62851, w62852, w62853, w62854, w62855, w62856, w62857, w62858, w62859, w62860, w62861, w62862, w62863, w62864, w62865, w62866, w62867, w62868, w62869, w62870, w62871, w62872, w62873, w62874, w62875, w62876, w62877, w62878, w62879, w62880, w62881, w62882, w62883, w62884, w62885, w62886, w62887, w62888, w62889, w62890, w62891, w62892, w62893, w62894, w62895, w62896, w62897, w62898, w62899, w62900, w62901, w62902, w62903, w62904, w62905, w62906, w62907, w62908, w62909, w62910, w62911, w62912, w62913, w62914, w62915, w62916, w62917, w62918, w62919, w62920, w62921, w62922, w62923, w62924, w62925, w62926, w62927, w62928, w62929, w62930, w62931, w62932, w62933, w62934, w62935, w62936, w62937, w62938, w62939, w62940, w62941, w62942, w62943, w62944, w62945, w62946, w62947, w62948, w62949, w62950, w62951, w62952, w62953, w62954, w62955, w62956, w62957, w62958, w62959, w62960, w62961, w62962, w62963, w62964, w62965, w62966, w62967, w62968, w62969, w62970, w62971, w62972, w62973, w62974, w62975, w62976, w62977, w62978, w62979, w62980, w62981, w62982, w62983, w62984, w62985, w62986, w62987, w62988, w62989, w62990, w62991, w62992, w62993, w62994, w62995, w62996, w62997, w62998, w62999, w63000, w63001, w63002, w63003, w63004, w63005, w63006, w63007, w63008, w63009, w63010, w63011, w63012, w63013, w63014, w63015, w63016, w63017, w63018, w63019, w63020, w63021, w63022, w63023, w63024, w63025, w63026, w63027, w63028, w63029, w63030, w63031, w63032, w63033, w63034, w63035, w63036, w63037, w63038, w63039, w63040, w63041, w63042, w63043, w63044, w63045, w63046, w63047, w63048, w63049, w63050, w63051, w63052, w63053, w63054, w63055, w63056, w63057, w63058, w63059, w63060, w63061, w63062, w63063, w63064, w63065, w63066, w63067, w63068, w63069, w63070, w63071, w63072, w63073, w63074, w63075, w63076, w63077, w63078, w63079, w63080, w63081, w63082, w63083, w63084, w63085, w63086, w63087, w63088, w63089, w63090, w63091, w63092, w63093, w63094, w63095, w63096, w63097, w63098, w63099, w63100, w63101, w63102, w63103, w63104, w63105, w63106, w63107, w63108, w63109, w63110, w63111, w63112, w63113, w63114, w63115, w63116, w63117, w63118, w63119, w63120, w63121, w63122, w63123, w63124, w63125, w63126, w63127, w63128, w63129, w63130, w63131, w63132, w63133, w63134, w63135, w63136, w63137, w63138, w63139, w63140, w63141, w63142, w63143, w63144, w63145, w63146, w63147, w63148, w63149, w63150, w63151, w63152, w63153, w63154, w63155, w63156, w63157, w63158, w63159, w63160, w63161, w63162, w63163, w63164, w63165, w63166, w63167, w63168, w63169, w63170, w63171, w63172, w63173, w63174, w63175, w63176, w63177, w63178, w63179, w63180, w63181, w63182, w63183, w63184, w63185, w63186, w63187, w63188, w63189, w63190, w63191, w63192, w63193, w63194, w63195, w63196, w63197, w63198, w63199, w63200, w63201, w63202, w63203, w63204, w63205, w63206, w63207, w63208, w63209, w63210, w63211, w63212, w63213, w63214, w63215, w63216, w63217, w63218, w63219, w63220, w63221, w63222, w63223, w63224, w63225, w63226, w63227, w63228, w63229, w63230, w63231, w63232, w63233, w63234, w63235, w63236, w63237, w63238, w63239, w63240, w63241, w63242, w63243, w63244, w63245, w63246, w63247, w63248, w63249, w63250, w63251, w63252, w63253, w63254, w63255, w63256, w63257, w63258, w63259, w63260, w63261, w63262, w63263, w63264, w63265, w63266, w63267, w63268, w63269, w63270, w63271, w63272, w63273, w63274, w63275, w63276, w63277, w63278, w63279, w63280, w63281, w63282, w63283, w63284, w63285, w63286, w63287, w63288, w63289, w63290, w63291, w63292, w63293, w63294, w63295, w63296, w63297, w63298, w63299, w63300, w63301, w63302, w63303, w63304, w63305, w63306, w63307, w63308, w63309, w63310, w63311, w63312, w63313, w63314, w63315, w63316, w63317, w63318, w63319, w63320, w63321, w63322, w63323, w63324, w63325, w63326, w63327, w63328, w63329, w63330, w63331, w63332, w63333, w63334, w63335, w63336, w63337, w63338, w63339, w63340, w63341, w63342, w63343, w63344, w63345, w63346, w63347, w63348, w63349, w63350, w63351, w63352, w63353, w63354, w63355, w63356, w63357, w63358, w63359, w63360, w63361, w63362, w63363, w63364, w63365, w63366, w63367, w63368, w63369, w63370, w63371, w63372, w63373, w63374, w63375, w63376, w63377, w63378, w63379, w63380, w63381, w63382, w63383, w63384, w63385, w63386, w63387, w63388, w63389, w63390, w63391, w63392, w63393, w63394, w63395, w63396, w63397, w63398, w63399, w63400, w63401, w63402, w63403, w63404, w63405, w63406, w63407, w63408, w63409, w63410, w63411, w63412, w63413, w63414, w63415, w63416, w63417, w63418, w63419, w63420, w63421, w63422, w63423, w63424, w63425, w63426, w63427, w63428, w63429, w63430, w63431, w63432, w63433, w63434, w63435, w63436, w63437, w63438, w63439, w63440, w63441, w63442, w63443, w63444, w63445, w63446, w63447, w63448, w63449, w63450, w63451, w63452, w63453, w63454, w63455, w63456, w63457, w63458, w63459, w63460, w63461, w63462, w63463, w63464, w63465, w63466, w63467, w63468, w63469, w63470, w63471, w63472, w63473, w63474, w63475, w63476, w63477, w63478, w63479, w63480, w63481, w63482, w63483, w63484, w63485, w63486, w63487, w63488, w63489, w63490, w63491, w63492, w63493, w63494, w63495, w63496, w63497, w63498, w63499, w63500, w63501, w63502, w63503, w63504, w63505, w63506, w63507, w63508, w63509, w63510, w63511, w63512, w63513, w63514, w63515, w63516, w63517, w63518, w63519, w63520, w63521, w63522, w63523, w63524, w63525, w63526, w63527, w63528, w63529, w63530, w63531, w63532, w63533, w63534, w63535, w63536, w63537, w63538, w63539, w63540, w63541, w63542, w63543, w63544, w63545, w63546, w63547, w63548, w63549, w63550, w63551, w63552, w63553, w63554, w63555, w63556, w63557, w63558, w63559, w63560, w63561, w63562, w63563, w63564, w63565, w63566, w63567, w63568, w63569, w63570, w63571, w63572, w63573, w63574, w63575, w63576, w63577, w63578, w63579, w63580, w63581, w63582, w63583, w63584, w63585, w63586, w63587, w63588, w63589, w63590, w63591, w63592, w63593, w63594, w63595, w63596, w63597, w63598, w63599, w63600, w63601, w63602, w63603, w63604, w63605, w63606, w63607, w63608, w63609, w63610, w63611, w63612, w63613, w63614, w63615, w63616, w63617, w63618, w63619, w63620, w63621, w63622, w63623, w63624, w63625, w63626, w63627, w63628, w63629, w63630, w63631, w63632, w63633, w63634, w63635, w63636, w63637, w63638, w63639, w63640, w63641, w63642, w63643, w63644, w63645, w63646, w63647, w63648, w63649, w63650, w63651, w63652, w63653, w63654, w63655, w63656, w63657, w63658, w63659, w63660, w63661, w63662, w63663, w63664, w63665, w63666, w63667, w63668, w63669, w63670, w63671, w63672, w63673, w63674, w63675, w63676, w63677, w63678, w63679, w63680, w63681, w63682, w63683, w63684, w63685, w63686, w63687, w63688, w63689, w63690, w63691, w63692, w63693, w63694, w63695, w63696, w63697, w63698, w63699, w63700, w63701, w63702, w63703, w63704, w63705, w63706, w63707, w63708, w63709, w63710, w63711, w63712, w63713, w63714, w63715, w63716, w63717, w63718, w63719, w63720, w63721, w63722, w63723, w63724, w63725, w63726, w63727, w63728, w63729, w63730, w63731, w63732, w63733, w63734, w63735, w63736, w63737, w63738, w63739, w63740, w63741, w63742, w63743, w63744, w63745, w63746, w63747, w63748, w63749, w63750, w63751, w63752, w63753, w63754, w63755, w63756, w63757, w63758, w63759, w63760, w63761, w63762, w63763, w63764, w63765, w63766, w63767, w63768, w63769, w63770, w63771, w63772, w63773, w63774, w63775, w63776, w63777, w63778, w63779, w63780, w63781, w63782, w63783, w63784, w63785, w63786, w63787, w63788, w63789, w63790, w63791, w63792, w63793, w63794, w63795, w63796, w63797, w63798, w63799, w63800, w63801, w63802, w63803, w63804, w63805, w63806, w63807, w63808, w63809, w63810, w63811, w63812, w63813, w63814, w63815, w63816, w63817, w63818, w63819, w63820, w63821, w63822, w63823, w63824, w63825, w63826, w63827, w63828, w63829, w63830, w63831, w63832, w63833, w63834, w63835, w63836, w63837, w63838, w63839, w63840, w63841, w63842, w63843, w63844, w63845, w63846, w63847, w63848, w63849, w63850, w63851, w63852, w63853, w63854, w63855, w63856, w63857, w63858, w63859, w63860, w63861, w63862, w63863, w63864, w63865, w63866, w63867, w63868, w63869, w63870, w63871, w63872, w63873, w63874, w63875, w63876, w63877, w63878, w63879, w63880, w63881, w63882, w63883, w63884, w63885, w63886, w63887, w63888, w63889, w63890, w63891, w63892, w63893, w63894, w63895, w63896, w63897, w63898, w63899, w63900, w63901, w63902, w63903, w63904, w63905, w63906, w63907, w63908, w63909, w63910, w63911, w63912, w63913, w63914, w63915, w63916, w63917, w63918, w63919, w63920, w63921, w63922, w63923, w63924, w63925, w63926, w63927, w63928, w63929, w63930, w63931, w63932, w63933, w63934, w63935, w63936, w63937, w63938, w63939, w63940, w63941, w63942, w63943, w63944, w63945, w63946, w63947, w63948, w63949, w63950, w63951, w63952, w63953, w63954, w63955, w63956, w63957, w63958, w63959, w63960, w63961, w63962, w63963, w63964, w63965, w63966, w63967, w63968, w63969, w63970, w63971, w63972, w63973, w63974, w63975, w63976, w63977, w63978, w63979, w63980, w63981, w63982, w63983, w63984, w63985, w63986, w63987, w63988, w63989, w63990, w63991, w63992, w63993, w63994, w63995, w63996, w63997, w63998, w63999, w64000, w64001, w64002, w64003, w64004, w64005, w64006, w64007, w64008, w64009, w64010, w64011, w64012, w64013, w64014, w64015, w64016, w64017, w64018, w64019, w64020, w64021, w64022, w64023, w64024, w64025, w64026, w64027, w64028, w64029, w64030, w64031, w64032, w64033, w64034, w64035, w64036, w64037, w64038, w64039, w64040, w64041, w64042, w64043, w64044, w64045, w64046, w64047, w64048, w64049, w64050, w64051, w64052, w64053, w64054, w64055, w64056, w64057, w64058, w64059, w64060, w64061, w64062, w64063, w64064, w64065, w64066, w64067, w64068, w64069, w64070, w64071, w64072, w64073, w64074, w64075, w64076, w64077, w64078, w64079, w64080, w64081, w64082, w64083, w64084, w64085, w64086, w64087, w64088, w64089, w64090, w64091, w64092, w64093, w64094, w64095, w64096, w64097, w64098, w64099, w64100, w64101, w64102, w64103, w64104, w64105, w64106, w64107, w64108, w64109, w64110, w64111, w64112, w64113, w64114, w64115, w64116, w64117, w64118, w64119, w64120, w64121, w64122, w64123, w64124, w64125, w64126, w64127, w64128, w64129, w64130, w64131, w64132, w64133, w64134, w64135, w64136, w64137, w64138, w64139, w64140, w64141, w64142, w64143, w64144, w64145, w64146, w64147, w64148, w64149, w64150, w64151, w64152, w64153, w64154, w64155, w64156, w64157, w64158, w64159, w64160, w64161, w64162, w64163, w64164, w64165, w64166, w64167, w64168, w64169, w64170, w64171, w64172, w64173, w64174, w64175, w64176, w64177, w64178, w64179, w64180, w64181, w64182, w64183, w64184, w64185, w64186, w64187, w64188, w64189, w64190, w64191, w64192, w64193, w64194, w64195, w64196, w64197, w64198, w64199, w64200, w64201, w64202, w64203, w64204, w64205, w64206, w64207, w64208, w64209, w64210, w64211, w64212, w64213, w64214, w64215, w64216, w64217, w64218, w64219, w64220, w64221, w64222, w64223, w64224, w64225, w64226, w64227, w64228, w64229, w64230, w64231, w64232, w64233, w64234, w64235, w64236, w64237, w64238, w64239, w64240, w64241, w64242, w64243, w64244, w64245, w64246, w64247, w64248, w64249, w64250, w64251, w64252, w64253, w64254, w64255, w64256, w64257, w64258, w64259, w64260, w64261, w64262, w64263, w64264, w64265, w64266, w64267, w64268, w64269, w64270, w64271, w64272, w64273, w64274, w64275, w64276, w64277, w64278, w64279, w64280, w64281, w64282, w64283, w64284, w64285, w64286, w64287, w64288, w64289, w64290, w64291, w64292, w64293, w64294, w64295, w64296, w64297, w64298, w64299, w64300, w64301, w64302, w64303, w64304, w64305, w64306, w64307, w64308, w64309, w64310, w64311, w64312, w64313, w64314, w64315, w64316, w64317, w64318, w64319, w64320, w64321, w64322, w64323, w64324, w64325, w64326, w64327, w64328, w64329, w64330, w64331, w64332, w64333, w64334, w64335, w64336, w64337, w64338, w64339, w64340, w64341, w64342, w64343, w64344, w64345, w64346, w64347, w64348, w64349, w64350, w64351, w64352, w64353, w64354, w64355, w64356, w64357, w64358, w64359, w64360, w64361, w64362, w64363, w64364, w64365, w64366, w64367, w64368, w64369, w64370, w64371, w64372, w64373, w64374, w64375, w64376, w64377, w64378, w64379, w64380, w64381, w64382, w64383, w64384, w64385, w64386, w64387, w64388, w64389, w64390, w64391, w64392, w64393, w64394, w64395, w64396, w64397, w64398, w64399, w64400, w64401, w64402, w64403, w64404, w64405, w64406, w64407, w64408, w64409, w64410, w64411, w64412, w64413, w64414, w64415, w64416, w64417, w64418, w64419, w64420, w64421, w64422, w64423, w64424, w64425, w64426, w64427, w64428, w64429, w64430, w64431, w64432, w64433, w64434, w64435, w64436, w64437, w64438, w64439, w64440, w64441, w64442, w64443, w64444, w64445, w64446, w64447, w64448, w64449, w64450, w64451, w64452, w64453, w64454, w64455, w64456, w64457, w64458, w64459, w64460, w64461, w64462, w64463, w64464, w64465, w64466, w64467, w64468, w64469, w64470, w64471, w64472, w64473, w64474, w64475, w64476, w64477, w64478, w64479, w64480, w64481, w64482, w64483, w64484, w64485, w64486, w64487, w64488, w64489, w64490, w64491, w64492, w64493, w64494, w64495, w64496, w64497, w64498, w64499, w64500, w64501, w64502, w64503, w64504, w64505, w64506, w64507, w64508, w64509, w64510, w64511, w64512, w64513, w64514, w64515, w64516, w64517, w64518, w64519, w64520, w64521, w64522, w64523, w64524, w64525, w64526, w64527, w64528, w64529, w64530, w64531, w64532, w64533, w64534, w64535, w64536, w64537, w64538, w64539, w64540, w64541, w64542, w64543, w64544, w64545, w64546, w64547, w64548, w64549, w64550, w64551, w64552, w64553, w64554, w64555, w64556, w64557, w64558, w64559, w64560, w64561, w64562, w64563, w64564, w64565, w64566, w64567, w64568, w64569, w64570, w64571, w64572, w64573, w64574, w64575, w64576, w64577, w64578, w64579, w64580, w64581, w64582, w64583, w64584, w64585, w64586, w64587, w64588, w64589, w64590, w64591, w64592, w64593, w64594, w64595, w64596, w64597, w64598, w64599, w64600, w64601, w64602, w64603, w64604, w64605, w64606, w64607, w64608, w64609, w64610, w64611, w64612, w64613, w64614, w64615, w64616, w64617, w64618, w64619, w64620, w64621, w64622, w64623, w64624, w64625, w64626, w64627, w64628, w64629, w64630, w64631, w64632, w64633, w64634, w64635, w64636, w64637, w64638, w64639, w64640, w64641, w64642, w64643, w64644, w64645, w64646, w64647, w64648, w64649, w64650, w64651, w64652, w64653, w64654, w64655, w64656, w64657, w64658, w64659, w64660, w64661, w64662, w64663, w64664, w64665, w64666, w64667, w64668, w64669, w64670, w64671, w64672, w64673, w64674, w64675, w64676, w64677, w64678, w64679, w64680, w64681, w64682, w64683, w64684, w64685, w64686, w64687, w64688, w64689, w64690, w64691, w64692, w64693, w64694, w64695, w64696, w64697, w64698, w64699, w64700, w64701, w64702, w64703, w64704, w64705, w64706, w64707, w64708, w64709, w64710, w64711, w64712, w64713, w64714, w64715, w64716, w64717, w64718, w64719, w64720, w64721, w64722, w64723, w64724, w64725, w64726, w64727, w64728, w64729, w64730, w64731, w64732, w64733, w64734, w64735, w64736, w64737, w64738, w64739, w64740, w64741, w64742, w64743, w64744, w64745, w64746, w64747, w64748, w64749, w64750, w64751, w64752, w64753, w64754, w64755, w64756, w64757, w64758, w64759, w64760, w64761, w64762, w64763, w64764, w64765, w64766, w64767, w64768, w64769, w64770, w64771, w64772, w64773, w64774, w64775, w64776, w64777, w64778, w64779, w64780, w64781, w64782, w64783, w64784, w64785, w64786, w64787, w64788, w64789, w64790, w64791, w64792, w64793, w64794, w64795, w64796, w64797, w64798, w64799, w64800, w64801, w64802, w64803, w64804, w64805, w64806, w64807, w64808, w64809, w64810, w64811, w64812, w64813, w64814, w64815, w64816, w64817, w64818, w64819, w64820, w64821, w64822, w64823, w64824, w64825, w64826, w64827, w64828, w64829, w64830, w64831, w64832, w64833, w64834, w64835, w64836, w64837, w64838, w64839, w64840, w64841, w64842, w64843, w64844, w64845, w64846, w64847, w64848, w64849, w64850, w64851, w64852, w64853, w64854, w64855, w64856, w64857, w64858, w64859, w64860, w64861, w64862, w64863, w64864, w64865, w64866, w64867, w64868, w64869, w64870, w64871, w64872, w64873, w64874, w64875, w64876, w64877, w64878, w64879, w64880, w64881, w64882, w64883, w64884, w64885, w64886, w64887, w64888, w64889, w64890, w64891, w64892, w64893, w64894, w64895, w64896, w64897, w64898, w64899, w64900, w64901, w64902, w64903, w64904, w64905, w64906, w64907, w64908, w64909, w64910, w64911, w64912, w64913, w64914, w64915, w64916, w64917, w64918, w64919, w64920, w64921, w64922, w64923, w64924, w64925, w64926, w64927, w64928, w64929, w64930, w64931, w64932, w64933, w64934, w64935, w64936, w64937, w64938, w64939, w64940, w64941, w64942, w64943, w64944, w64945, w64946, w64947, w64948, w64949, w64950, w64951, w64952, w64953, w64954, w64955, w64956, w64957, w64958, w64959, w64960, w64961, w64962, w64963, w64964, w64965, w64966, w64967, w64968, w64969, w64970, w64971, w64972, w64973, w64974, w64975, w64976, w64977, w64978, w64979, w64980, w64981, w64982, w64983, w64984, w64985, w64986, w64987, w64988, w64989, w64990, w64991, w64992, w64993, w64994, w64995, w64996, w64997, w64998, w64999, w65000, w65001, w65002, w65003, w65004, w65005, w65006, w65007, w65008, w65009, w65010, w65011, w65012, w65013, w65014, w65015, w65016, w65017, w65018, w65019, w65020, w65021, w65022, w65023, w65024, w65025, w65026, w65027, w65028, w65029, w65030, w65031, w65032, w65033, w65034, w65035, w65036, w65037, w65038, w65039, w65040, w65041, w65042, w65043, w65044, w65045, w65046, w65047, w65048, w65049, w65050, w65051, w65052, w65053, w65054, w65055, w65056, w65057, w65058, w65059, w65060, w65061, w65062, w65063, w65064, w65065, w65066, w65067, w65068, w65069, w65070, w65071, w65072, w65073, w65074, w65075, w65076, w65077, w65078, w65079, w65080, w65081, w65082, w65083, w65084, w65085, w65086, w65087, w65088, w65089, w65090, w65091, w65092, w65093, w65094, w65095, w65096, w65097, w65098, w65099, w65100, w65101, w65102, w65103, w65104, w65105, w65106, w65107, w65108, w65109, w65110, w65111, w65112, w65113, w65114, w65115, w65116, w65117, w65118, w65119, w65120, w65121, w65122, w65123, w65124, w65125, w65126, w65127, w65128, w65129, w65130, w65131, w65132, w65133, w65134, w65135, w65136, w65137, w65138, w65139, w65140, w65141, w65142, w65143, w65144, w65145, w65146, w65147, w65148, w65149, w65150, w65151, w65152, w65153, w65154, w65155, w65156, w65157, w65158, w65159, w65160, w65161, w65162, w65163, w65164, w65165, w65166, w65167, w65168, w65169, w65170, w65171, w65172, w65173, w65174, w65175, w65176, w65177, w65178, w65179, w65180, w65181, w65182, w65183, w65184, w65185, w65186, w65187, w65188, w65189, w65190, w65191, w65192, w65193, w65194, w65195, w65196, w65197, w65198, w65199, w65200, w65201, w65202, w65203, w65204, w65205, w65206, w65207, w65208, w65209, w65210, w65211, w65212, w65213, w65214, w65215, w65216, w65217, w65218, w65219, w65220, w65221, w65222, w65223, w65224, w65225, w65226, w65227, w65228, w65229, w65230, w65231, w65232, w65233, w65234, w65235, w65236, w65237, w65238, w65239, w65240, w65241, w65242, w65243, w65244, w65245, w65246, w65247, w65248, w65249, w65250, w65251, w65252, w65253, w65254, w65255, w65256, w65257, w65258, w65259, w65260, w65261, w65262, w65263, w65264, w65265, w65266, w65267, w65268, w65269, w65270, w65271, w65272, w65273, w65274, w65275, w65276, w65277, w65278, w65279, w65280, w65281, w65282, w65283, w65284, w65285, w65286, w65287, w65288, w65289, w65290, w65291, w65292, w65293, w65294, w65295, w65296, w65297, w65298, w65299, w65300, w65301, w65302, w65303, w65304, w65305, w65306, w65307, w65308, w65309, w65310, w65311, w65312, w65313, w65314, w65315, w65316, w65317, w65318, w65319, w65320, w65321, w65322, w65323, w65324, w65325, w65326, w65327, w65328, w65329, w65330, w65331, w65332, w65333, w65334, w65335, w65336, w65337, w65338, w65339, w65340, w65341, w65342, w65343, w65344, w65345, w65346, w65347, w65348, w65349, w65350, w65351, w65352, w65353, w65354, w65355, w65356, w65357, w65358, w65359, w65360, w65361, w65362, w65363, w65364, w65365, w65366, w65367, w65368, w65369, w65370, w65371, w65372, w65373, w65374, w65375, w65376, w65377, w65378, w65379, w65380, w65381, w65382, w65383, w65384, w65385, w65386, w65387, w65388, w65389, w65390, w65391, w65392, w65393, w65394, w65395, w65396, w65397, w65398, w65399, w65400, w65401, w65402, w65403, w65404, w65405, w65406, w65407, w65408, w65409, w65410, w65411, w65412, w65413, w65414, w65415, w65416, w65417, w65418, w65419, w65420, w65421, w65422, w65423, w65424, w65425, w65426, w65427, w65428, w65429, w65430, w65431, w65432, w65433, w65434, w65435, w65436, w65437, w65438, w65439, w65440, w65441, w65442, w65443, w65444, w65445, w65446, w65447, w65448, w65449, w65450, w65451, w65452, w65453, w65454, w65455, w65456, w65457, w65458, w65459, w65460, w65461, w65462, w65463, w65464, w65465, w65466, w65467, w65468, w65469, w65470, w65471, w65472, w65473, w65474, w65475, w65476, w65477, w65478, w65479, w65480, w65481, w65482, w65483, w65484, w65485, w65486, w65487, w65488, w65489, w65490, w65491, w65492, w65493, w65494, w65495, w65496, w65497, w65498, w65499, w65500, w65501, w65502, w65503, w65504, w65505, w65506, w65507, w65508, w65509, w65510, w65511, w65512, w65513, w65514, w65515, w65516, w65517, w65518, w65519, w65520, w65521, w65522, w65523, w65524, w65525, w65526, w65527, w65528, w65529, w65530, w65531, w65532, w65533, w65534, w65535, w65536, w65537, w65538, w65539, w65540, w65541, w65542, w65543, w65544, w65545, w65546, w65547, w65548, w65549, w65550, w65551, w65552, w65553, w65554, w65555, w65556, w65557, w65558, w65559, w65560, w65561, w65562, w65563, w65564, w65565, w65566, w65567, w65568, w65569, w65570, w65571, w65572, w65573, w65574, w65575, w65576, w65577, w65578, w65579, w65580, w65581, w65582, w65583, w65584, w65585, w65586, w65587, w65588, w65589, w65590, w65591, w65592, w65593, w65594, w65595, w65596, w65597, w65598, w65599, w65600, w65601, w65602, w65603, w65604, w65605, w65606, w65607, w65608, w65609, w65610, w65611, w65612, w65613, w65614, w65615, w65616, w65617, w65618, w65619, w65620, w65621, w65622, w65623, w65624, w65625, w65626, w65627, w65628, w65629, w65630, w65631, w65632, w65633, w65634, w65635, w65636, w65637, w65638, w65639, w65640, w65641, w65642, w65643, w65644, w65645, w65646, w65647, w65648, w65649, w65650, w65651, w65652, w65653, w65654, w65655, w65656, w65657, w65658, w65659, w65660, w65661, w65662, w65663, w65664, w65665, w65666, w65667, w65668, w65669, w65670, w65671, w65672, w65673, w65674, w65675, w65676, w65677, w65678, w65679, w65680, w65681, w65682, w65683, w65684, w65685, w65686, w65687, w65688, w65689, w65690, w65691, w65692, w65693, w65694, w65695, w65696, w65697, w65698, w65699, w65700, w65701, w65702, w65703, w65704, w65705, w65706, w65707, w65708, w65709, w65710, w65711, w65712, w65713, w65714, w65715, w65716, w65717, w65718, w65719, w65720, w65721, w65722, w65723, w65724, w65725, w65726, w65727, w65728, w65729, w65730, w65731, w65732, w65733, w65734, w65735, w65736, w65737, w65738, w65739, w65740, w65741, w65742, w65743, w65744, w65745, w65746, w65747, w65748, w65749, w65750, w65751, w65752, w65753, w65754, w65755, w65756, w65757, w65758, w65759, w65760, w65761, w65762, w65763, w65764, w65765, w65766, w65767, w65768, w65769, w65770, w65771, w65772, w65773, w65774, w65775, w65776, w65777, w65778, w65779, w65780, w65781, w65782, w65783, w65784, w65785, w65786, w65787, w65788, w65789, w65790, w65791, w65792, w65793, w65794, w65795, w65796, w65797, w65798, w65799, w65800, w65801, w65802, w65803, w65804, w65805, w65806, w65807, w65808, w65809, w65810, w65811, w65812, w65813, w65814, w65815, w65816, w65817, w65818, w65819, w65820, w65821, w65822, w65823, w65824, w65825, w65826, w65827, w65828, w65829, w65830, w65831, w65832, w65833, w65834, w65835, w65836, w65837, w65838, w65839, w65840, w65841, w65842, w65843, w65844, w65845, w65846, w65847, w65848, w65849, w65850, w65851, w65852, w65853, w65854, w65855, w65856, w65857, w65858, w65859, w65860, w65861, w65862, w65863, w65864, w65865, w65866, w65867, w65868, w65869, w65870, w65871, w65872, w65873, w65874, w65875, w65876, w65877, w65878, w65879, w65880, w65881, w65882, w65883, w65884, w65885, w65886, w65887, w65888, w65889, w65890, w65891, w65892, w65893, w65894, w65895, w65896, w65897, w65898, w65899, w65900, w65901, w65902, w65903, w65904, w65905, w65906, w65907, w65908, w65909, w65910, w65911, w65912, w65913, w65914, w65915, w65916, w65917, w65918, w65919, w65920, w65921, w65922, w65923, w65924, w65925, w65926, w65927, w65928, w65929, w65930, w65931, w65932, w65933, w65934, w65935, w65936, w65937, w65938, w65939, w65940, w65941, w65942, w65943, w65944, w65945, w65946, w65947, w65948, w65949, w65950, w65951, w65952, w65953, w65954, w65955, w65956, w65957, w65958, w65959, w65960, w65961, w65962, w65963, w65964, w65965, w65966, w65967, w65968, w65969, w65970, w65971, w65972, w65973, w65974, w65975, w65976, w65977, w65978, w65979, w65980, w65981, w65982, w65983, w65984, w65985, w65986, w65987, w65988, w65989, w65990, w65991, w65992, w65993, w65994, w65995, w65996, w65997, w65998, w65999, w66000, w66001, w66002, w66003, w66004, w66005, w66006, w66007, w66008, w66009, w66010, w66011, w66012, w66013, w66014, w66015, w66016, w66017, w66018, w66019, w66020, w66021, w66022, w66023, w66024, w66025, w66026, w66027, w66028, w66029, w66030, w66031, w66032, w66033, w66034, w66035, w66036, w66037, w66038, w66039, w66040, w66041, w66042, w66043, w66044, w66045, w66046, w66047, w66048, w66049, w66050, w66051, w66052, w66053, w66054, w66055, w66056, w66057, w66058, w66059, w66060, w66061, w66062, w66063, w66064, w66065, w66066, w66067, w66068, w66069, w66070, w66071, w66072, w66073, w66074, w66075, w66076, w66077, w66078, w66079, w66080, w66081, w66082, w66083, w66084, w66085, w66086, w66087, w66088, w66089, w66090, w66091, w66092, w66093, w66094, w66095, w66096, w66097, w66098, w66099, w66100, w66101, w66102, w66103, w66104, w66105, w66106, w66107, w66108, w66109, w66110, w66111, w66112, w66113, w66114, w66115, w66116, w66117, w66118, w66119, w66120, w66121, w66122, w66123, w66124, w66125, w66126, w66127, w66128, w66129, w66130, w66131, w66132, w66133, w66134, w66135, w66136, w66137, w66138, w66139, w66140, w66141, w66142, w66143, w66144, w66145, w66146, w66147, w66148, w66149, w66150, w66151, w66152, w66153, w66154, w66155, w66156, w66157, w66158, w66159, w66160, w66161, w66162, w66163, w66164, w66165, w66166, w66167, w66168, w66169, w66170, w66171, w66172, w66173, w66174, w66175, w66176, w66177, w66178, w66179, w66180, w66181, w66182, w66183, w66184, w66185, w66186, w66187, w66188, w66189, w66190, w66191, w66192, w66193, w66194, w66195, w66196, w66197, w66198, w66199, w66200, w66201, w66202, w66203, w66204, w66205, w66206, w66207, w66208, w66209, w66210, w66211, w66212, w66213, w66214, w66215, w66216, w66217, w66218, w66219, w66220, w66221, w66222, w66223, w66224, w66225, w66226, w66227, w66228, w66229, w66230, w66231, w66232, w66233, w66234, w66235, w66236, w66237, w66238, w66239, w66240, w66241, w66242, w66243, w66244, w66245, w66246, w66247, w66248, w66249, w66250, w66251, w66252, w66253, w66254, w66255, w66256, w66257, w66258, w66259, w66260, w66261, w66262, w66263, w66264, w66265, w66266, w66267, w66268, w66269, w66270, w66271, w66272, w66273, w66274, w66275, w66276, w66277, w66278, w66279, w66280, w66281, w66282, w66283, w66284, w66285, w66286, w66287, w66288, w66289, w66290, w66291, w66292, w66293, w66294, w66295, w66296, w66297, w66298, w66299, w66300, w66301, w66302, w66303, w66304, w66305, w66306, w66307, w66308, w66309, w66310, w66311, w66312, w66313, w66314, w66315, w66316, w66317, w66318, w66319, w66320, w66321, w66322, w66323, w66324, w66325, w66326, w66327, w66328, w66329, w66330, w66331, w66332, w66333, w66334, w66335, w66336, w66337, w66338, w66339, w66340, w66341, w66342, w66343, w66344, w66345, w66346, w66347, w66348, w66349, w66350, w66351, w66352, w66353, w66354, w66355, w66356, w66357, w66358, w66359, w66360, w66361, w66362, w66363, w66364, w66365, w66366, w66367, w66368, w66369, w66370, w66371, w66372, w66373, w66374, w66375, w66376, w66377, w66378, w66379, w66380, w66381, w66382, w66383, w66384, w66385, w66386, w66387, w66388, w66389, w66390, w66391, w66392, w66393, w66394, w66395, w66396, w66397, w66398, w66399, w66400, w66401, w66402, w66403, w66404, w66405, w66406, w66407, w66408, w66409, w66410, w66411, w66412, w66413, w66414, w66415, w66416, w66417, w66418, w66419, w66420, w66421, w66422, w66423, w66424, w66425, w66426, w66427, w66428, w66429, w66430, w66431, w66432, w66433, w66434, w66435, w66436, w66437, w66438, w66439, w66440, w66441, w66442, w66443, w66444, w66445, w66446, w66447, w66448, w66449, w66450, w66451, w66452, w66453, w66454, w66455, w66456, w66457, w66458, w66459, w66460, w66461, w66462, w66463, w66464, w66465, w66466, w66467, w66468, w66469, w66470, w66471, w66472, w66473, w66474, w66475, w66476, w66477, w66478, w66479, w66480, w66481, w66482, w66483, w66484, w66485, w66486, w66487, w66488, w66489, w66490, w66491, w66492, w66493, w66494, w66495, w66496, w66497, w66498, w66499, w66500, w66501, w66502, w66503, w66504, w66505, w66506, w66507, w66508, w66509, w66510, w66511, w66512, w66513, w66514, w66515, w66516, w66517, w66518, w66519, w66520, w66521, w66522, w66523, w66524, w66525, w66526, w66527, w66528, w66529, w66530, w66531, w66532, w66533, w66534, w66535, w66536, w66537, w66538, w66539, w66540, w66541, w66542, w66543, w66544, w66545, w66546, w66547, w66548, w66549, w66550, w66551, w66552, w66553, w66554, w66555, w66556, w66557, w66558, w66559, w66560, w66561, w66562, w66563, w66564, w66565, w66566, w66567, w66568, w66569, w66570, w66571, w66572, w66573, w66574, w66575, w66576, w66577, w66578, w66579, w66580, w66581, w66582, w66583, w66584, w66585, w66586, w66587, w66588, w66589, w66590, w66591, w66592, w66593, w66594, w66595, w66596, w66597, w66598, w66599, w66600, w66601, w66602, w66603, w66604, w66605, w66606, w66607, w66608, w66609, w66610, w66611, w66612, w66613, w66614, w66615, w66616, w66617, w66618, w66619, w66620, w66621, w66622, w66623, w66624, w66625, w66626, w66627, w66628, w66629, w66630, w66631, w66632, w66633, w66634, w66635, w66636, w66637, w66638, w66639, w66640, w66641, w66642, w66643, w66644, w66645, w66646, w66647, w66648, w66649, w66650, w66651, w66652, w66653, w66654, w66655, w66656, w66657, w66658, w66659, w66660, w66661, w66662, w66663, w66664, w66665, w66666, w66667, w66668, w66669, w66670, w66671, w66672, w66673, w66674, w66675, w66676, w66677, w66678, w66679, w66680, w66681, w66682, w66683, w66684, w66685, w66686, w66687, w66688, w66689, w66690, w66691, w66692, w66693, w66694, w66695, w66696, w66697, w66698, w66699, w66700, w66701, w66702, w66703, w66704, w66705, w66706, w66707, w66708, w66709, w66710, w66711, w66712, w66713, w66714, w66715, w66716, w66717, w66718, w66719, w66720, w66721, w66722, w66723, w66724, w66725, w66726, w66727, w66728, w66729, w66730, w66731, w66732, w66733, w66734, w66735, w66736, w66737, w66738, w66739, w66740, w66741, w66742, w66743, w66744, w66745, w66746, w66747, w66748, w66749, w66750, w66751, w66752, w66753, w66754, w66755, w66756, w66757, w66758, w66759, w66760, w66761, w66762, w66763, w66764, w66765, w66766, w66767, w66768, w66769, w66770, w66771, w66772, w66773, w66774, w66775, w66776, w66777, w66778, w66779, w66780, w66781, w66782, w66783, w66784, w66785, w66786, w66787, w66788, w66789, w66790, w66791, w66792, w66793, w66794, w66795, w66796, w66797, w66798, w66799, w66800, w66801, w66802, w66803, w66804, w66805, w66806, w66807, w66808, w66809, w66810, w66811, w66812, w66813, w66814, w66815, w66816, w66817, w66818, w66819, w66820, w66821, w66822, w66823, w66824, w66825, w66826, w66827, w66828, w66829, w66830, w66831, w66832, w66833, w66834, w66835, w66836, w66837, w66838, w66839, w66840, w66841, w66842, w66843, w66844, w66845, w66846, w66847, w66848, w66849, w66850, w66851, w66852, w66853, w66854, w66855, w66856, w66857, w66858, w66859, w66860, w66861, w66862, w66863, w66864, w66865, w66866, w66867, w66868, w66869, w66870, w66871, w66872, w66873, w66874, w66875, w66876, w66877, w66878, w66879, w66880, w66881, w66882, w66883, w66884, w66885, w66886, w66887, w66888, w66889, w66890, w66891, w66892, w66893, w66894, w66895, w66896, w66897, w66898, w66899, w66900, w66901, w66902, w66903, w66904, w66905, w66906, w66907, w66908, w66909, w66910, w66911, w66912, w66913, w66914, w66915, w66916, w66917, w66918, w66919, w66920, w66921, w66922, w66923, w66924, w66925, w66926, w66927, w66928, w66929, w66930, w66931, w66932, w66933, w66934, w66935, w66936, w66937, w66938, w66939, w66940, w66941, w66942, w66943, w66944, w66945, w66946, w66947, w66948, w66949, w66950, w66951, w66952, w66953, w66954, w66955, w66956, w66957, w66958, w66959, w66960, w66961, w66962, w66963, w66964, w66965, w66966, w66967, w66968, w66969, w66970, w66971, w66972, w66973, w66974, w66975, w66976, w66977, w66978, w66979, w66980, w66981, w66982, w66983, w66984, w66985, w66986, w66987, w66988, w66989, w66990, w66991, w66992, w66993, w66994, w66995, w66996, w66997, w66998, w66999, w67000, w67001, w67002, w67003, w67004, w67005, w67006, w67007, w67008, w67009, w67010, w67011, w67012, w67013, w67014, w67015, w67016, w67017, w67018, w67019, w67020, w67021, w67022, w67023, w67024, w67025, w67026, w67027, w67028, w67029, w67030, w67031, w67032, w67033, w67034, w67035, w67036, w67037, w67038, w67039, w67040, w67041, w67042, w67043, w67044, w67045, w67046, w67047, w67048, w67049, w67050, w67051, w67052, w67053, w67054, w67055, w67056, w67057, w67058, w67059, w67060, w67061, w67062, w67063, w67064, w67065, w67066, w67067, w67068, w67069, w67070, w67071, w67072, w67073, w67074, w67075, w67076, w67077, w67078, w67079, w67080, w67081, w67082, w67083, w67084, w67085, w67086, w67087, w67088, w67089, w67090, w67091, w67092, w67093, w67094, w67095, w67096, w67097, w67098, w67099, w67100, w67101, w67102, w67103, w67104, w67105, w67106, w67107, w67108, w67109, w67110, w67111, w67112, w67113, w67114, w67115, w67116, w67117, w67118, w67119, w67120, w67121, w67122, w67123, w67124, w67125, w67126, w67127, w67128, w67129, w67130, w67131, w67132, w67133, w67134, w67135, w67136, w67137, w67138, w67139, w67140, w67141, w67142, w67143, w67144, w67145, w67146, w67147, w67148, w67149, w67150, w67151, w67152, w67153, w67154, w67155, w67156, w67157, w67158, w67159, w67160, w67161, w67162, w67163, w67164, w67165, w67166, w67167, w67168, w67169, w67170, w67171, w67172, w67173, w67174, w67175, w67176, w67177, w67178, w67179, w67180, w67181, w67182, w67183, w67184, w67185, w67186, w67187, w67188, w67189, w67190, w67191, w67192, w67193;
assign w0 = ~pi2998 & pi9040;
assign w1 = ~pi3008 & ~pi9040;
assign w2 = ~w0 & ~w1;
assign w3 = pi0066 & ~w2;
assign w4 = ~pi0066 & w2;
assign w5 = ~w3 & ~w4;
assign w6 = ~pi3003 & pi9040;
assign w7 = ~pi2992 & ~pi9040;
assign w8 = ~w6 & ~w7;
assign w9 = pi0036 & ~w8;
assign w10 = ~pi0036 & w8;
assign w11 = ~w9 & ~w10;
assign w12 = ~w5 & ~w11;
assign w13 = ~pi3010 & pi9040;
assign w14 = ~pi2991 & ~pi9040;
assign w15 = ~w13 & ~w14;
assign w16 = pi0067 & ~w15;
assign w17 = ~pi0067 & w15;
assign w18 = ~w16 & ~w17;
assign w19 = ~w5 & ~w18;
assign w20 = ~pi2984 & pi9040;
assign w21 = ~pi2986 & ~pi9040;
assign w22 = ~w20 & ~w21;
assign w23 = pi0070 & ~w22;
assign w24 = ~pi0070 & w22;
assign w25 = ~w23 & ~w24;
assign w26 = ~w19 & ~w25;
assign w27 = ~w5 & w11;
assign w28 = ~w18 & w25;
assign w29 = w27 & w28;
assign w30 = ~w26 & ~w29;
assign w31 = ~pi2982 & pi9040;
assign w32 = ~pi3103 & ~pi9040;
assign w33 = ~w31 & ~w32;
assign w34 = pi0095 & ~w33;
assign w35 = ~pi0095 & w33;
assign w36 = ~w34 & ~w35;
assign w37 = ~w30 & w36;
assign w38 = w12 & w37;
assign w39 = ~pi3105 & pi9040;
assign w40 = ~pi3001 & ~pi9040;
assign w41 = ~w39 & ~w40;
assign w42 = pi0077 & ~w41;
assign w43 = ~pi0077 & w41;
assign w44 = ~w42 & ~w43;
assign w45 = w5 & w36;
assign w46 = w11 & ~w25;
assign w47 = w5 & w11;
assign w48 = ~w12 & ~w47;
assign w49 = ~w11 & w25;
assign w50 = ~w46 & ~w49;
assign w51 = w48 & ~w50;
assign w52 = w18 & w51;
assign w53 = (~w46 & ~w51) | (~w46 & w64476) | (~w51 & w64476);
assign w54 = w45 & ~w53;
assign w55 = w18 & w54;
assign w56 = w5 & w25;
assign w57 = ~w36 & w56;
assign w58 = ~w11 & w19;
assign w59 = ~w57 & ~w58;
assign w60 = ~w18 & w50;
assign w61 = w59 & w60;
assign w62 = ~w55 & ~w61;
assign w63 = ~w44 & ~w62;
assign w64 = ~w25 & w48;
assign w65 = w25 & ~w48;
assign w66 = ~w64 & ~w65;
assign w67 = w11 & w18;
assign w68 = ~w66 & w67;
assign w69 = ~w11 & ~w18;
assign w70 = w5 & w69;
assign w71 = ~w5 & w18;
assign w72 = w49 & w71;
assign w73 = ~w18 & ~w25;
assign w74 = ~w27 & w73;
assign w75 = ~w72 & ~w74;
assign w76 = ~w44 & ~w75;
assign w77 = ~w70 & ~w76;
assign w78 = ~w68 & w77;
assign w79 = ~w36 & ~w78;
assign w80 = ~w36 & ~w56;
assign w81 = w50 & w80;
assign w82 = w27 & ~w81;
assign w83 = w45 & w64;
assign w84 = w75 & w83;
assign w85 = ~w18 & w36;
assign w86 = ~w56 & w85;
assign w87 = ~w58 & ~w86;
assign w88 = ~w50 & ~w87;
assign w89 = ~w25 & w71;
assign w90 = ~w82 & ~w89;
assign w91 = ~w88 & w90;
assign w92 = ~w84 & w91;
assign w93 = ~w57 & w92;
assign w94 = w44 & ~w93;
assign w95 = w25 & w36;
assign w96 = w19 & w95;
assign w97 = ~w38 & ~w96;
assign w98 = ~w79 & w97;
assign w99 = ~w63 & w98;
assign w100 = ~w94 & w99;
assign w101 = w45 & ~w92;
assign w102 = ~w28 & ~w36;
assign w103 = ~w26 & w102;
assign w104 = w18 & w47;
assign w105 = ~w103 & ~w104;
assign w106 = ~w37 & w105;
assign w107 = w56 & w69;
assign w108 = w44 & ~w107;
assign w109 = w106 & w108;
assign w110 = ~w48 & w95;
assign w111 = w18 & ~w66;
assign w112 = w81 & ~w111;
assign w113 = ~w44 & ~w110;
assign w114 = ~w52 & w113;
assign w115 = ~w112 & w114;
assign w116 = ~w109 & ~w115;
assign w117 = ~w101 & ~w116;
assign w118 = ~pi2991 & pi9040;
assign w119 = ~pi2999 & ~pi9040;
assign w120 = ~w118 & ~w119;
assign w121 = pi0088 & ~w120;
assign w122 = ~pi0088 & w120;
assign w123 = ~w121 & ~w122;
assign w124 = ~pi3001 & pi9040;
assign w125 = ~pi3046 & ~pi9040;
assign w126 = ~w124 & ~w125;
assign w127 = pi0036 & ~w126;
assign w128 = ~pi0036 & w126;
assign w129 = ~w127 & ~w128;
assign w130 = w123 & w129;
assign w131 = ~w123 & ~w129;
assign w132 = ~w130 & ~w131;
assign w133 = ~pi2995 & pi9040;
assign w134 = ~pi3003 & ~pi9040;
assign w135 = ~w133 & ~w134;
assign w136 = pi0071 & ~w135;
assign w137 = ~pi0071 & w135;
assign w138 = ~w136 & ~w137;
assign w139 = ~pi3045 & pi9040;
assign w140 = ~pi2983 & ~pi9040;
assign w141 = ~w139 & ~w140;
assign w142 = pi0077 & ~w141;
assign w143 = ~pi0077 & w141;
assign w144 = ~w142 & ~w143;
assign w145 = ~pi2987 & pi9040;
assign w146 = ~pi2984 & ~pi9040;
assign w147 = ~w145 & ~w146;
assign w148 = pi0091 & ~w147;
assign w149 = ~pi0091 & w147;
assign w150 = ~w148 & ~w149;
assign w151 = w131 & w150;
assign w152 = ~w144 & w151;
assign w153 = w129 & ~w150;
assign w154 = w144 & w153;
assign w155 = ~w152 & ~w154;
assign w156 = w138 & ~w155;
assign w157 = w132 & w156;
assign w158 = w144 & w150;
assign w159 = w132 & w158;
assign w160 = ~w123 & w159;
assign w161 = w144 & ~w150;
assign w162 = ~w132 & w161;
assign w163 = ~w123 & ~w144;
assign w164 = w129 & w163;
assign w165 = ~w162 & ~w164;
assign w166 = ~w129 & w150;
assign w167 = ~w144 & w166;
assign w168 = w123 & w167;
assign w169 = w165 & ~w168;
assign w170 = ~w160 & w169;
assign w171 = ~w138 & ~w170;
assign w172 = ~pi3064 & pi9040;
assign w173 = ~pi3000 & ~pi9040;
assign w174 = ~w172 & ~w173;
assign w175 = pi0086 & ~w174;
assign w176 = ~pi0086 & w174;
assign w177 = ~w175 & ~w176;
assign w178 = w138 & ~w150;
assign w179 = ~w153 & ~w178;
assign w180 = w123 & ~w144;
assign w181 = ~w179 & w180;
assign w182 = w123 & w144;
assign w183 = w132 & ~w182;
assign w184 = w138 & ~w183;
assign w185 = ~w129 & w182;
assign w186 = ~w163 & ~w185;
assign w187 = ~w158 & w186;
assign w188 = w184 & ~w187;
assign w189 = ~w177 & ~w181;
assign w190 = ~w188 & w189;
assign w191 = ~w157 & w190;
assign w192 = ~w171 & w191;
assign w193 = ~w158 & ~w163;
assign w194 = w179 & w193;
assign w195 = w165 & w64477;
assign w196 = w153 & ~w165;
assign w197 = ~w138 & ~w185;
assign w198 = ~w151 & w197;
assign w199 = w131 & ~w150;
assign w200 = w138 & ~w199;
assign w201 = ~w194 & w200;
assign w202 = ~w198 & ~w201;
assign w203 = ~w160 & w177;
assign w204 = ~w196 & w203;
assign w205 = ~w202 & w204;
assign w206 = ~w195 & w205;
assign w207 = ~w192 & ~w206;
assign w208 = ~w48 & w86;
assign w209 = ~w57 & ~w104;
assign w210 = w28 & w47;
assign w211 = ~w48 & w80;
assign w212 = w50 & w71;
assign w213 = w27 & w36;
assign w214 = ~w210 & ~w213;
assign w215 = ~w211 & w214;
assign w216 = ~w212 & w215;
assign w217 = ~w209 & ~w216;
assign w218 = w108 & ~w208;
assign w219 = ~w111 & w218;
assign w220 = ~w217 & w219;
assign w221 = ~w44 & ~w83;
assign w222 = w45 & w52;
assign w223 = w216 & w221;
assign w224 = ~w222 & w223;
assign w225 = ~w220 & ~w224;
assign w226 = ~pi3063 & pi9040;
assign w227 = ~pi3068 & ~pi9040;
assign w228 = ~w226 & ~w227;
assign w229 = pi0076 & ~w228;
assign w230 = ~pi0076 & w228;
assign w231 = ~w229 & ~w230;
assign w232 = ~pi3043 & pi9040;
assign w233 = ~pi3016 & ~pi9040;
assign w234 = ~w232 & ~w233;
assign w235 = pi0069 & ~w234;
assign w236 = ~pi0069 & w234;
assign w237 = ~w235 & ~w236;
assign w238 = ~w231 & ~w237;
assign w239 = ~pi3004 & pi9040;
assign w240 = ~pi3044 & ~pi9040;
assign w241 = ~w239 & ~w240;
assign w242 = pi0068 & ~w241;
assign w243 = ~pi0068 & w241;
assign w244 = ~w242 & ~w243;
assign w245 = ~pi2985 & pi9040;
assign w246 = ~pi3006 & ~pi9040;
assign w247 = ~w245 & ~w246;
assign w248 = pi0050 & ~w247;
assign w249 = ~pi0050 & w247;
assign w250 = ~w248 & ~w249;
assign w251 = ~w244 & ~w250;
assign w252 = w238 & w251;
assign w253 = ~pi3011 & pi9040;
assign w254 = pi3033 & ~pi9040;
assign w255 = ~w253 & ~w254;
assign w256 = pi0061 & ~w255;
assign w257 = ~pi0061 & w255;
assign w258 = ~w256 & ~w257;
assign w259 = ~pi3042 & pi9040;
assign w260 = ~pi2981 & ~pi9040;
assign w261 = ~w259 & ~w260;
assign w262 = pi0087 & ~w261;
assign w263 = ~pi0087 & w261;
assign w264 = ~w262 & ~w263;
assign w265 = w250 & ~w264;
assign w266 = ~w231 & w244;
assign w267 = w265 & w266;
assign w268 = ~w231 & ~w244;
assign w269 = ~w264 & w268;
assign w270 = ~w250 & w269;
assign w271 = w237 & w244;
assign w272 = ~w244 & w264;
assign w273 = w244 & ~w264;
assign w274 = ~w272 & ~w273;
assign w275 = w231 & ~w274;
assign w276 = w264 & w266;
assign w277 = ~w275 & ~w276;
assign w278 = ~w231 & w264;
assign w279 = w250 & w278;
assign w280 = w271 & ~w279;
assign w281 = ~w277 & w280;
assign w282 = ~w267 & ~w270;
assign w283 = ~w281 & w282;
assign w284 = w258 & ~w283;
assign w285 = ~w250 & w264;
assign w286 = ~w231 & w285;
assign w287 = ~w271 & w286;
assign w288 = w250 & w269;
assign w289 = w231 & ~w244;
assign w290 = w264 & w289;
assign w291 = ~w288 & ~w290;
assign w292 = w237 & ~w291;
assign w293 = ~w287 & ~w292;
assign w294 = ~w258 & ~w293;
assign w295 = ~w266 & ~w289;
assign w296 = w265 & ~w295;
assign w297 = w231 & w264;
assign w298 = w244 & ~w250;
assign w299 = w297 & w298;
assign w300 = ~w279 & ~w299;
assign w301 = w258 & ~w300;
assign w302 = ~w244 & w278;
assign w303 = ~w296 & ~w302;
assign w304 = ~w301 & w303;
assign w305 = ~w237 & ~w304;
assign w306 = w231 & w237;
assign w307 = w244 & ~w258;
assign w308 = ~w306 & ~w307;
assign w309 = ~w238 & ~w265;
assign w310 = ~w285 & w309;
assign w311 = ~w308 & w310;
assign w312 = ~w252 & ~w311;
assign w313 = ~w305 & w312;
assign w314 = ~w284 & w313;
assign w315 = ~w294 & w314;
assign w316 = ~w150 & w163;
assign w317 = w130 & ~w144;
assign w318 = ~w316 & ~w317;
assign w319 = w138 & ~w318;
assign w320 = ~w159 & ~w177;
assign w321 = ~w152 & ~w319;
assign w322 = w320 & w321;
assign w323 = w150 & w164;
assign w324 = w131 & w144;
assign w325 = ~w323 & ~w324;
assign w326 = w138 & ~w325;
assign w327 = w161 & ~w197;
assign w328 = ~w138 & ~w318;
assign w329 = w129 & w138;
assign w330 = w182 & w329;
assign w331 = w177 & ~w330;
assign w332 = ~w168 & w331;
assign w333 = ~w327 & w332;
assign w334 = ~w328 & w333;
assign w335 = ~w326 & w334;
assign w336 = ~w322 & ~w335;
assign w337 = w186 & ~w317;
assign w338 = ~w151 & ~w177;
assign w339 = w337 & w338;
assign w340 = ~w160 & ~w167;
assign w341 = ~w339 & w340;
assign w342 = ~w138 & ~w341;
assign w343 = ~w336 & ~w342;
assign w344 = w67 & ~w106;
assign w345 = w59 & w221;
assign w346 = ~w344 & w345;
assign w347 = ~w29 & w44;
assign w348 = ~w38 & w347;
assign w349 = ~w54 & w348;
assign w350 = ~w346 & ~w349;
assign w351 = ~w18 & w83;
assign w352 = ~w64 & ~w72;
assign w353 = w44 & ~w352;
assign w354 = ~w51 & ~w68;
assign w355 = ~w52 & ~w354;
assign w356 = ~w353 & ~w355;
assign w357 = ~w36 & ~w356;
assign w358 = ~w96 & ~w351;
assign w359 = ~w350 & w358;
assign w360 = ~w357 & w359;
assign w361 = ~pi2997 & pi9040;
assign w362 = ~pi3047 & ~pi9040;
assign w363 = ~w361 & ~w362;
assign w364 = pi0064 & ~w363;
assign w365 = ~pi0064 & w363;
assign w366 = ~w364 & ~w365;
assign w367 = ~pi2980 & pi9040;
assign w368 = ~pi3066 & ~pi9040;
assign w369 = ~w367 & ~w368;
assign w370 = pi0058 & ~w369;
assign w371 = ~pi0058 & w369;
assign w372 = ~w370 & ~w371;
assign w373 = ~pi3068 & pi9040;
assign w374 = ~pi3106 & ~pi9040;
assign w375 = ~w373 & ~w374;
assign w376 = pi0076 & ~w375;
assign w377 = ~pi0076 & w375;
assign w378 = ~w376 & ~w377;
assign w379 = w372 & ~w378;
assign w380 = ~pi2990 & pi9040;
assign w381 = ~pi2985 & ~pi9040;
assign w382 = ~w380 & ~w381;
assign w383 = pi0060 & ~w382;
assign w384 = ~pi0060 & w382;
assign w385 = ~w383 & ~w384;
assign w386 = w379 & w385;
assign w387 = w372 & ~w385;
assign w388 = w378 & w387;
assign w389 = ~w386 & ~w388;
assign w390 = w372 & w389;
assign w391 = ~pi3009 & pi9040;
assign w392 = ~pi3042 & ~pi9040;
assign w393 = ~w391 & ~w392;
assign w394 = pi0090 & ~w393;
assign w395 = ~pi0090 & w393;
assign w396 = ~w394 & ~w395;
assign w397 = ~w390 & ~w396;
assign w398 = w378 & w385;
assign w399 = ~w372 & w398;
assign w400 = ~w372 & ~w385;
assign w401 = ~w378 & w400;
assign w402 = ~w399 & ~w401;
assign w403 = ~w386 & w396;
assign w404 = w402 & w403;
assign w405 = w366 & ~w404;
assign w406 = ~w397 & w405;
assign w407 = ~pi3033 & pi9040;
assign w408 = pi2979 & ~pi9040;
assign w409 = ~w407 & ~w408;
assign w410 = pi0087 & ~w409;
assign w411 = ~pi0087 & w409;
assign w412 = ~w410 & ~w411;
assign w413 = w366 & w398;
assign w414 = ~w372 & ~w378;
assign w415 = ~w366 & w385;
assign w416 = w414 & w415;
assign w417 = w396 & ~w416;
assign w418 = ~w366 & ~w388;
assign w419 = ~w390 & w418;
assign w420 = ~w417 & w419;
assign w421 = ~w366 & w378;
assign w422 = w372 & w396;
assign w423 = w421 & w422;
assign w424 = ~w413 & ~w423;
assign w425 = ~w420 & w424;
assign w426 = ~w412 & ~w425;
assign w427 = ~w366 & ~w396;
assign w428 = w414 & w427;
assign w429 = w366 & ~w372;
assign w430 = ~w379 & ~w400;
assign w431 = ~w366 & w430;
assign w432 = ~w429 & ~w431;
assign w433 = w402 & ~w432;
assign w434 = ~w396 & w433;
assign w435 = w387 & w418;
assign w436 = w389 & ~w421;
assign w437 = w396 & ~w436;
assign w438 = ~w433 & w437;
assign w439 = ~w434 & ~w435;
assign w440 = ~w438 & w439;
assign w441 = w412 & ~w440;
assign w442 = ~w406 & ~w428;
assign w443 = ~w426 & w442;
assign w444 = ~w441 & w443;
assign w445 = ~pi3000 & pi9040;
assign w446 = ~pi3038 & ~pi9040;
assign w447 = ~w445 & ~w446;
assign w448 = pi0059 & ~w447;
assign w449 = ~pi0059 & w447;
assign w450 = ~w448 & ~w449;
assign w451 = ~pi3046 & pi9040;
assign w452 = ~pi2996 & ~pi9040;
assign w453 = ~w451 & ~w452;
assign w454 = pi0089 & ~w453;
assign w455 = ~pi0089 & w453;
assign w456 = ~w454 & ~w455;
assign w457 = ~pi3008 & pi9040;
assign w458 = ~pi2987 & ~pi9040;
assign w459 = ~w457 & ~w458;
assign w460 = pi0049 & ~w459;
assign w461 = ~pi0049 & w459;
assign w462 = ~w460 & ~w461;
assign w463 = ~pi3040 & pi9040;
assign w464 = ~pi2995 & ~pi9040;
assign w465 = ~w463 & ~w464;
assign w466 = pi0084 & ~w465;
assign w467 = ~pi0084 & w465;
assign w468 = ~w466 & ~w467;
assign w469 = ~w462 & w468;
assign w470 = ~pi2983 & pi9040;
assign w471 = ~pi3105 & ~pi9040;
assign w472 = ~w470 & ~w471;
assign w473 = pi0083 & ~w472;
assign w474 = ~pi0083 & w472;
assign w475 = ~w473 & ~w474;
assign w476 = w469 & w475;
assign w477 = w469 & w64478;
assign w478 = ~w450 & w477;
assign w479 = ~w462 & ~w475;
assign w480 = w456 & ~w462;
assign w481 = w475 & ~w480;
assign w482 = (~w468 & w480) | (~w468 & w64479) | (w480 & w64479);
assign w483 = ~w479 & ~w482;
assign w484 = w462 & ~w475;
assign w485 = ~w456 & w484;
assign w486 = w450 & ~w480;
assign w487 = ~w485 & w486;
assign w488 = ~w483 & w487;
assign w489 = ~w468 & w488;
assign w490 = ~pi2986 & pi9040;
assign w491 = ~pi2978 & ~pi9040;
assign w492 = ~w490 & ~w491;
assign w493 = pi0092 & ~w492;
assign w494 = ~pi0092 & w492;
assign w495 = ~w493 & ~w494;
assign w496 = w450 & w468;
assign w497 = ~w487 & w496;
assign w498 = w462 & w475;
assign w499 = w462 & ~w468;
assign w500 = ~w456 & w499;
assign w501 = ~w496 & ~w500;
assign w502 = w498 & ~w501;
assign w503 = w450 & ~w468;
assign w504 = w479 & w503;
assign w505 = w456 & ~w475;
assign w506 = w469 & w505;
assign w507 = ~w468 & w479;
assign w508 = ~w456 & w507;
assign w509 = ~w506 & ~w508;
assign w510 = ~w468 & w475;
assign w511 = ~w484 & ~w510;
assign w512 = ~w456 & ~w475;
assign w513 = ~w450 & ~w512;
assign w514 = ~w511 & w513;
assign w515 = ~w504 & ~w514;
assign w516 = ~w497 & w515;
assign w517 = ~w502 & w509;
assign w518 = w516 & w517;
assign w519 = ~w495 & ~w518;
assign w520 = ~w462 & w475;
assign w521 = ~w456 & w520;
assign w522 = ~w469 & ~w499;
assign w523 = w456 & w522;
assign w524 = w475 & w523;
assign w525 = ~w521 & ~w524;
assign w526 = w468 & ~w525;
assign w527 = w479 & w509;
assign w528 = ~w477 & ~w500;
assign w529 = ~w527 & w528;
assign w530 = ~w450 & ~w529;
assign w531 = w450 & ~w499;
assign w532 = ~w511 & w531;
assign w533 = ~w526 & ~w532;
assign w534 = ~w530 & w533;
assign w535 = w495 & ~w534;
assign w536 = ~w478 & ~w489;
assign w537 = ~w519 & w536;
assign w538 = ~w535 & w537;
assign w539 = ~pi2993 & pi9040;
assign w540 = ~pi2990 & ~pi9040;
assign w541 = ~w539 & ~w540;
assign w542 = pi0092 & ~w541;
assign w543 = ~pi0092 & w541;
assign w544 = ~w542 & ~w543;
assign w545 = ~pi3044 & pi9040;
assign w546 = ~pi2997 & ~pi9040;
assign w547 = ~w545 & ~w546;
assign w548 = pi0083 & ~w547;
assign w549 = ~pi0083 & w547;
assign w550 = ~w548 & ~w549;
assign w551 = ~pi3016 & pi9040;
assign w552 = ~pi3058 & ~pi9040;
assign w553 = ~w551 & ~w552;
assign w554 = pi0060 & ~w553;
assign w555 = ~pi0060 & w553;
assign w556 = ~w554 & ~w555;
assign w557 = ~w550 & ~w556;
assign w558 = ~w544 & w557;
assign w559 = ~w544 & w550;
assign w560 = w556 & w559;
assign w561 = ~w558 & ~w560;
assign w562 = ~w544 & w561;
assign w563 = ~pi2988 & pi9040;
assign w564 = ~pi2980 & ~pi9040;
assign w565 = ~w563 & ~w564;
assign w566 = pi0094 & ~w565;
assign w567 = ~pi0094 & w565;
assign w568 = ~w566 & ~w567;
assign w569 = w562 & w568;
assign w570 = ~pi2976 & pi9040;
assign w571 = ~pi3028 & ~pi9040;
assign w572 = ~w570 & ~w571;
assign w573 = pi0085 & ~w572;
assign w574 = ~pi0085 & w572;
assign w575 = ~w573 & ~w574;
assign w576 = w569 & ~w575;
assign w577 = ~pi3106 & pi9040;
assign w578 = ~pi2994 & ~pi9040;
assign w579 = ~w577 & ~w578;
assign w580 = pi0058 & ~w579;
assign w581 = ~pi0058 & w579;
assign w582 = ~w580 & ~w581;
assign w583 = w559 & ~w568;
assign w584 = w544 & w568;
assign w585 = w556 & w584;
assign w586 = ~w583 & ~w585;
assign w587 = ~w558 & w586;
assign w588 = ~w568 & ~w575;
assign w589 = ~w561 & w588;
assign w590 = w544 & w556;
assign w591 = ~w550 & w590;
assign w592 = ~w575 & ~w591;
assign w593 = ~w583 & w592;
assign w594 = ~w587 & ~w589;
assign w595 = ~w593 & w594;
assign w596 = w561 & ~w575;
assign w597 = w586 & w596;
assign w598 = ~w595 & ~w597;
assign w599 = ~w568 & w590;
assign w600 = ~w550 & w599;
assign w601 = w550 & ~w568;
assign w602 = w544 & ~w556;
assign w603 = w601 & w602;
assign w604 = w557 & w584;
assign w605 = ~w603 & ~w604;
assign w606 = ~w600 & w605;
assign w607 = ~w582 & w606;
assign w608 = ~w598 & w607;
assign w609 = w585 & w592;
assign w610 = w550 & ~w556;
assign w611 = ~w544 & w610;
assign w612 = ~w557 & w575;
assign w613 = ~w611 & w612;
assign w614 = w586 & w613;
assign w615 = ~w589 & w606;
assign w616 = ~w609 & ~w614;
assign w617 = w615 & w616;
assign w618 = w582 & ~w617;
assign w619 = w558 & w568;
assign w620 = ~w603 & ~w619;
assign w621 = w575 & ~w620;
assign w622 = ~w576 & ~w621;
assign w623 = ~w618 & w622;
assign w624 = ~w608 & w623;
assign w625 = w398 & w437;
assign w626 = w378 & w400;
assign w627 = w366 & w626;
assign w628 = w379 & w427;
assign w629 = ~w396 & ~w628;
assign w630 = ~w386 & ~w431;
assign w631 = w629 & ~w630;
assign w632 = w366 & w401;
assign w633 = w414 & ~w415;
assign w634 = ~w390 & ~w633;
assign w635 = w396 & ~w632;
assign w636 = ~w634 & w635;
assign w637 = w412 & ~w627;
assign w638 = ~w631 & w637;
assign w639 = ~w636 & w638;
assign w640 = w366 & w372;
assign w641 = w378 & w640;
assign w642 = ~w396 & ~w641;
assign w643 = ~w633 & w642;
assign w644 = w366 & ~w389;
assign w645 = ~w399 & w417;
assign w646 = ~w644 & w645;
assign w647 = ~w643 & ~w646;
assign w648 = ~w366 & w626;
assign w649 = ~w412 & ~w628;
assign w650 = ~w632 & w649;
assign w651 = ~w648 & w650;
assign w652 = ~w647 & w651;
assign w653 = ~w639 & ~w652;
assign w654 = ~w435 & ~w625;
assign w655 = ~w653 & w654;
assign w656 = w396 & ~w402;
assign w657 = ~w387 & ~w396;
assign w658 = w396 & ~w626;
assign w659 = w372 & w415;
assign w660 = w658 & ~w659;
assign w661 = ~w657 & ~w660;
assign w662 = ~w642 & ~w661;
assign w663 = w402 & ~w662;
assign w664 = w412 & ~w656;
assign w665 = ~w663 & w664;
assign w666 = w389 & ~w396;
assign w667 = ~w366 & ~w658;
assign w668 = ~w666 & w667;
assign w669 = ~w399 & w418;
assign w670 = w634 & w669;
assign w671 = w366 & ~w402;
assign w672 = ~w661 & ~w671;
assign w673 = ~w670 & w672;
assign w674 = ~w412 & ~w673;
assign w675 = ~w665 & ~w668;
assign w676 = ~w674 & w675;
assign w677 = w584 & w610;
assign w678 = ~w619 & ~w677;
assign w679 = w575 & ~w678;
assign w680 = ~w601 & ~w610;
assign w681 = ~w556 & ~w584;
assign w682 = ~w680 & ~w681;
assign w683 = w550 & w590;
assign w684 = ~w560 & ~w591;
assign w685 = ~w584 & ~w601;
assign w686 = w684 & w685;
assign w687 = w575 & ~w683;
assign w688 = ~w686 & w687;
assign w689 = ~w593 & ~w688;
assign w690 = ~w682 & ~w689;
assign w691 = ~w544 & ~w568;
assign w692 = ~w602 & ~w691;
assign w693 = w613 & ~w692;
assign w694 = ~w559 & ~w693;
assign w695 = ~w582 & ~w694;
assign w696 = w690 & w695;
assign w697 = w582 & ~w690;
assign w698 = ~w582 & ~w692;
assign w699 = ~w584 & ~w698;
assign w700 = ~w575 & ~w699;
assign w701 = ~w693 & ~w700;
assign w702 = ~w550 & ~w701;
assign w703 = ~w568 & w683;
assign w704 = ~w679 & ~w703;
assign w705 = ~w702 & w704;
assign w706 = ~w696 & w705;
assign w707 = ~w697 & w706;
assign w708 = ~w138 & w150;
assign w709 = ~w186 & w708;
assign w710 = ~w199 & ~w329;
assign w711 = w144 & ~w710;
assign w712 = ~w150 & w182;
assign w713 = ~w138 & ~w712;
assign w714 = ~w324 & w713;
assign w715 = ~w153 & ~w714;
assign w716 = ~w131 & w713;
assign w717 = ~w195 & w716;
assign w718 = ~w715 & ~w717;
assign w719 = w177 & ~w709;
assign w720 = ~w711 & w719;
assign w721 = ~w718 & w720;
assign w722 = w337 & w708;
assign w723 = ~w150 & w183;
assign w724 = ~w190 & ~w320;
assign w725 = ~w722 & ~w723;
assign w726 = ~w195 & w725;
assign w727 = ~w724 & w726;
assign w728 = ~w721 & ~w727;
assign w729 = ~w156 & ~w728;
assign w730 = ~w506 & ~w524;
assign w731 = w450 & ~w730;
assign w732 = ~w456 & w468;
assign w733 = ~w484 & w732;
assign w734 = ~w476 & ~w733;
assign w735 = w495 & ~w734;
assign w736 = w505 & w522;
assign w737 = ~w735 & ~w736;
assign w738 = ~w450 & ~w737;
assign w739 = ~w500 & ~w510;
assign w740 = w450 & ~w739;
assign w741 = ~w498 & w523;
assign w742 = ~w740 & ~w741;
assign w743 = w495 & ~w742;
assign w744 = ~w510 & ~w512;
assign w745 = w462 & ~w503;
assign w746 = ~w744 & w745;
assign w747 = ~w488 & ~w746;
assign w748 = ~w526 & w747;
assign w749 = ~w495 & ~w748;
assign w750 = ~w731 & ~w738;
assign w751 = ~w743 & w750;
assign w752 = ~w749 & w751;
assign w753 = w366 & w430;
assign w754 = ~w669 & ~w753;
assign w755 = ~w412 & w754;
assign w756 = ~w396 & ~w755;
assign w757 = w417 & ~w641;
assign w758 = ~w648 & w757;
assign w759 = ~w756 & ~w758;
assign w760 = ~w386 & ~w401;
assign w761 = w427 & ~w760;
assign w762 = w366 & w387;
assign w763 = w658 & ~w762;
assign w764 = ~w419 & w763;
assign w765 = ~w412 & ~w754;
assign w766 = w764 & w765;
assign w767 = ~w406 & w753;
assign w768 = w629 & ~w659;
assign w769 = ~w767 & w768;
assign w770 = w412 & ~w764;
assign w771 = ~w769 & w770;
assign w772 = ~w761 & ~w766;
assign w773 = ~w759 & w772;
assign w774 = ~w771 & w773;
assign w775 = ~w264 & w289;
assign w776 = ~w302 & ~w775;
assign w777 = w250 & ~w776;
assign w778 = w237 & ~w267;
assign w779 = ~w237 & ~w270;
assign w780 = ~w297 & w779;
assign w781 = ~w778 & ~w780;
assign w782 = ~w277 & w298;
assign w783 = w258 & ~w777;
assign w784 = ~w782 & w783;
assign w785 = ~w781 & w784;
assign w786 = w250 & ~w277;
assign w787 = w237 & w786;
assign w788 = ~w258 & ~w787;
assign w789 = w244 & w279;
assign w790 = ~w250 & ~w776;
assign w791 = ~w237 & ~w265;
assign w792 = w295 & ~w791;
assign w793 = w238 & w273;
assign w794 = ~w789 & ~w793;
assign w795 = ~w792 & w794;
assign w796 = ~w790 & w795;
assign w797 = w788 & w796;
assign w798 = ~w785 & ~w797;
assign w799 = ~w562 & ~w588;
assign w800 = w569 & w614;
assign w801 = ~w582 & ~w800;
assign w802 = ~w691 & ~w799;
assign w803 = ~w801 & w802;
assign w804 = ~w582 & w683;
assign w805 = w556 & w691;
assign w806 = ~w568 & ~w805;
assign w807 = ~w680 & ~w806;
assign w808 = w557 & w691;
assign w809 = ~w591 & ~w808;
assign w810 = w582 & ~w809;
assign w811 = w575 & ~w804;
assign w812 = ~w807 & w811;
assign w813 = ~w810 & w812;
assign w814 = w684 & ~w805;
assign w815 = ~w582 & ~w814;
assign w816 = ~w575 & ~w604;
assign w817 = ~w815 & w816;
assign w818 = ~w813 & ~w817;
assign w819 = w602 & w689;
assign w820 = ~w583 & w678;
assign w821 = ~w819 & w820;
assign w822 = ~w582 & ~w821;
assign w823 = ~w803 & ~w818;
assign w824 = ~w822 & w823;
assign w825 = w450 & w521;
assign w826 = ~w450 & ~w732;
assign w827 = w481 & ~w500;
assign w828 = w483 & w505;
assign w829 = (~w504 & ~w827) | (~w504 & w64480) | (~w827 & w64480);
assign w830 = ~w828 & w829;
assign w831 = w484 & w826;
assign w832 = w502 & w503;
assign w833 = w479 & w496;
assign w834 = ~w831 & ~w833;
assign w835 = ~w478 & w834;
assign w836 = ~w524 & w835;
assign w837 = ~w832 & w836;
assign w838 = w462 & w830;
assign w839 = ~w450 & w507;
assign w840 = ~w825 & ~w839;
assign w841 = w509 & w840;
assign w842 = (w841 & ~w837) | (w841 & w64481) | (~w837 & w64481);
assign w843 = ~w495 & ~w842;
assign w844 = ~w508 & ~w524;
assign w845 = ~w450 & ~w844;
assign w846 = w495 & ~w837;
assign w847 = ~w497 & ~w845;
assign w848 = ~w846 & w847;
assign w849 = ~w843 & w848;
assign w850 = ~pi2994 & pi9040;
assign w851 = ~pi3009 & ~pi9040;
assign w852 = ~w850 & ~w851;
assign w853 = pi0061 & ~w852;
assign w854 = ~pi0061 & w852;
assign w855 = ~w853 & ~w854;
assign w856 = ~pi3047 & pi9040;
assign w857 = ~pi3063 & ~pi9040;
assign w858 = ~w856 & ~w857;
assign w859 = pi0093 & ~w858;
assign w860 = ~pi0093 & w858;
assign w861 = ~w859 & ~w860;
assign w862 = w855 & w861;
assign w863 = ~w855 & ~w861;
assign w864 = ~w862 & ~w863;
assign w865 = ~pi2979 & pi9040;
assign w866 = ~pi2988 & ~pi9040;
assign w867 = ~w865 & ~w866;
assign w868 = pi0066 & ~w867;
assign w869 = ~pi0066 & w867;
assign w870 = ~w868 & ~w869;
assign w871 = ~pi3002 & pi9040;
assign w872 = ~pi2993 & ~pi9040;
assign w873 = ~w871 & ~w872;
assign w874 = pi0068 & ~w873;
assign w875 = ~pi0068 & w873;
assign w876 = ~w874 & ~w875;
assign w877 = ~w870 & ~w876;
assign w878 = ~w864 & w877;
assign w879 = ~w855 & w870;
assign w880 = w864 & ~w879;
assign w881 = w876 & w880;
assign w882 = ~w878 & ~w881;
assign w883 = ~w855 & ~w882;
assign w884 = w870 & ~w876;
assign w885 = w864 & w884;
assign w886 = ~w883 & ~w885;
assign w887 = ~pi3028 & pi9040;
assign w888 = pi2977 & ~pi9040;
assign w889 = ~w887 & ~w888;
assign w890 = pi0074 & ~w889;
assign w891 = ~pi0074 & w889;
assign w892 = ~w890 & ~w891;
assign w893 = ~w886 & w892;
assign w894 = ~w870 & w876;
assign w895 = ~w861 & ~w870;
assign w896 = w861 & w884;
assign w897 = ~w895 & ~w896;
assign w898 = w855 & ~w892;
assign w899 = ~w897 & w898;
assign w900 = w894 & w899;
assign w901 = w855 & ~w870;
assign w902 = w892 & ~w901;
assign w903 = w861 & w870;
assign w904 = ~w862 & w894;
assign w905 = ~w884 & w892;
assign w906 = ~w903 & w905;
assign w907 = ~w904 & w906;
assign w908 = ~w902 & ~w907;
assign w909 = w855 & ~w861;
assign w910 = ~w894 & ~w909;
assign w911 = ~w908 & ~w910;
assign w912 = w876 & w879;
assign w913 = w861 & w912;
assign w914 = ~w864 & ~w892;
assign w915 = ~w876 & w914;
assign w916 = ~pi3066 & pi9040;
assign w917 = ~pi3043 & ~pi9040;
assign w918 = ~w916 & ~w917;
assign w919 = pi0070 & ~w918;
assign w920 = ~pi0070 & w918;
assign w921 = ~w919 & ~w920;
assign w922 = ~w913 & w921;
assign w923 = ~w915 & w922;
assign w924 = ~w911 & w923;
assign w925 = w880 & w908;
assign w926 = w892 & ~w895;
assign w927 = ~w855 & w884;
assign w928 = ~w878 & ~w927;
assign w929 = w926 & ~w928;
assign w930 = w876 & ~w901;
assign w931 = w870 & ~w892;
assign w932 = ~w862 & ~w931;
assign w933 = w930 & ~w932;
assign w934 = ~w921 & ~w933;
assign w935 = ~w929 & w934;
assign w936 = ~w925 & w935;
assign w937 = ~w924 & ~w936;
assign w938 = ~w893 & ~w900;
assign w939 = ~w937 & w938;
assign w940 = ~w485 & w495;
assign w941 = w482 & ~w940;
assign w942 = ~w520 & w733;
assign w943 = ~w941 & ~w942;
assign w944 = ~w450 & ~w943;
assign w945 = ~w487 & w495;
assign w946 = ~w528 & ~w945;
assign w947 = ~w495 & w496;
assign w948 = w734 & w947;
assign w949 = ~w476 & ~w740;
assign w950 = w480 & ~w949;
assign w951 = w469 & w512;
assign w952 = w830 & ~w951;
assign w953 = ~w950 & w952;
assign w954 = w495 & ~w953;
assign w955 = ~w946 & ~w948;
assign w956 = ~w944 & w955;
assign w957 = ~w954 & w956;
assign w958 = w237 & ~w286;
assign w959 = w295 & w958;
assign w960 = ~w251 & ~w266;
assign w961 = w250 & ~w272;
assign w962 = w960 & ~w961;
assign w963 = w297 & ~w962;
assign w964 = ~w237 & w264;
assign w965 = ~w960 & w964;
assign w966 = ~w296 & ~w965;
assign w967 = ~w959 & w966;
assign w968 = ~w963 & w967;
assign w969 = ~w258 & ~w968;
assign w970 = ~w237 & ~w267;
assign w971 = (w237 & ~w265) | (w237 & w64482) | (~w265 & w64482);
assign w972 = ~w299 & w971;
assign w973 = ~w970 & ~w972;
assign w974 = w237 & w258;
assign w975 = ~w231 & ~w250;
assign w976 = ~w274 & w975;
assign w977 = ~w775 & ~w789;
assign w978 = ~w976 & w977;
assign w979 = w974 & ~w978;
assign w980 = ~w269 & ~w962;
assign w981 = w258 & ~w959;
assign w982 = ~w980 & w981;
assign w983 = ~w973 & ~w979;
assign w984 = ~w982 & w983;
assign w985 = ~w969 & w984;
assign w986 = ~w550 & w568;
assign w987 = ~w575 & ~w703;
assign w988 = ~w805 & w987;
assign w989 = ~w986 & ~w988;
assign w990 = ~w602 & ~w989;
assign w991 = ~w693 & ~w990;
assign w992 = ~w582 & ~w991;
assign w993 = ~w599 & ~w611;
assign w994 = ~w987 & ~w993;
assign w995 = ~w604 & ~w994;
assign w996 = w582 & ~w995;
assign w997 = ~w599 & ~w809;
assign w998 = w560 & w582;
assign w999 = ~w603 & ~w998;
assign w1000 = ~w997 & w999;
assign w1001 = ~w575 & ~w1000;
assign w1002 = ~w800 & ~w1001;
assign w1003 = ~w819 & w1002;
assign w1004 = ~w996 & w1003;
assign w1005 = ~w992 & w1004;
assign w1006 = ~w138 & w317;
assign w1007 = ~w184 & ~w714;
assign w1008 = ~w152 & w177;
assign w1009 = ~w1007 & w1008;
assign w1010 = ~w131 & w144;
assign w1011 = w129 & ~w708;
assign w1012 = ~w166 & ~w1010;
assign w1013 = ~w1011 & w1012;
assign w1014 = w320 & ~w330;
assign w1015 = ~w1013 & w1014;
assign w1016 = ~w1009 & ~w1015;
assign w1017 = ~w182 & ~w196;
assign w1018 = w138 & ~w161;
assign w1019 = ~w1017 & w1018;
assign w1020 = ~w1006 & ~w1016;
assign w1021 = ~w1019 & w1020;
assign w1022 = w880 & w933;
assign w1023 = w863 & ~w876;
assign w1024 = ~w881 & w921;
assign w1025 = ~w877 & w897;
assign w1026 = w1024 & w1025;
assign w1027 = ~w1023 & ~w1026;
assign w1028 = w892 & ~w1027;
assign w1029 = ~w855 & ~w892;
assign w1030 = w894 & w1029;
assign w1031 = ~w921 & ~w1030;
assign w1032 = w855 & w894;
assign w1033 = w862 & ~w876;
assign w1034 = ~w1032 & ~w1033;
assign w1035 = w892 & ~w1034;
assign w1036 = ~w930 & ~w931;
assign w1037 = w864 & ~w1036;
assign w1038 = ~w878 & w1031;
assign w1039 = ~w1035 & w1038;
assign w1040 = ~w1037 & w1039;
assign w1041 = w863 & w884;
assign w1042 = ~w855 & w877;
assign w1043 = ~w1032 & ~w1042;
assign w1044 = w861 & ~w1043;
assign w1045 = w921 & ~w1041;
assign w1046 = ~w899 & w1045;
assign w1047 = ~w1044 & w1046;
assign w1048 = ~w1040 & ~w1047;
assign w1049 = ~w1022 & ~w1048;
assign w1050 = ~w1028 & w1049;
assign w1051 = w288 & ~w974;
assign w1052 = ~w250 & ~w268;
assign w1053 = w274 & w1052;
assign w1054 = ~w237 & ~w1053;
assign w1055 = ~w272 & ~w975;
assign w1056 = ~w285 & ~w1055;
assign w1057 = ~w275 & w971;
assign w1058 = ~w1056 & w1057;
assign w1059 = ~w1054 & ~w1058;
assign w1060 = ~w786 & ~w1059;
assign w1061 = ~w1059 & w64483;
assign w1062 = w971 & w1053;
assign w1063 = ~w1061 & ~w1062;
assign w1064 = ~w258 & ~w1063;
assign w1065 = ~w788 & ~w1060;
assign w1066 = ~w1051 & ~w1065;
assign w1067 = ~w1064 & w1066;
assign w1068 = ~w886 & w925;
assign w1069 = w877 & w926;
assign w1070 = ~w855 & ~w895;
assign w1071 = w876 & ~w1070;
assign w1072 = w902 & w1071;
assign w1073 = ~w912 & ~w1023;
assign w1074 = ~w1032 & w1073;
assign w1075 = ~w892 & ~w1074;
assign w1076 = ~w913 & ~w1041;
assign w1077 = w855 & ~w876;
assign w1078 = w897 & w1077;
assign w1079 = w921 & ~w1072;
assign w1080 = w1076 & ~w1078;
assign w1081 = w1079 & w1080;
assign w1082 = ~w1075 & w1081;
assign w1083 = ~w898 & ~w927;
assign w1084 = w903 & ~w1083;
assign w1085 = ~w907 & w1031;
assign w1086 = ~w1084 & w1085;
assign w1087 = ~w1082 & ~w1086;
assign w1088 = ~w900 & ~w1069;
assign w1089 = ~w1068 & w1088;
assign w1090 = ~w1087 & w1089;
assign w1091 = ~pi3103 & pi9040;
assign w1092 = ~pi3005 & ~pi9040;
assign w1093 = ~w1091 & ~w1092;
assign w1094 = pi0086 & ~w1093;
assign w1095 = ~pi0086 & w1093;
assign w1096 = ~w1094 & ~w1095;
assign w1097 = ~pi3007 & pi9040;
assign w1098 = ~pi3040 & ~pi9040;
assign w1099 = ~w1097 & ~w1098;
assign w1100 = pi0084 & ~w1099;
assign w1101 = ~pi0084 & w1099;
assign w1102 = ~w1100 & ~w1101;
assign w1103 = ~w1096 & w1102;
assign w1104 = ~pi3038 & pi9040;
assign w1105 = ~pi2989 & ~pi9040;
assign w1106 = ~w1104 & ~w1105;
assign w1107 = pi0088 & ~w1106;
assign w1108 = ~pi0088 & w1106;
assign w1109 = ~w1107 & ~w1108;
assign w1110 = ~pi2978 & pi9040;
assign w1111 = ~pi3010 & ~pi9040;
assign w1112 = ~w1110 & ~w1111;
assign w1113 = pi0065 & ~w1112;
assign w1114 = ~pi0065 & w1112;
assign w1115 = ~w1113 & ~w1114;
assign w1116 = ~w1109 & ~w1115;
assign w1117 = ~pi2996 & pi9040;
assign w1118 = pi3053 & ~pi9040;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = pi0049 & ~w1119;
assign w1121 = ~pi0049 & w1119;
assign w1122 = ~w1120 & ~w1121;
assign w1123 = ~pi2992 & pi9040;
assign w1124 = ~pi3045 & ~pi9040;
assign w1125 = ~w1123 & ~w1124;
assign w1126 = pi0075 & ~w1125;
assign w1127 = ~pi0075 & w1125;
assign w1128 = ~w1126 & ~w1127;
assign w1129 = w1122 & w1128;
assign w1130 = w1116 & w1129;
assign w1131 = w1109 & w1115;
assign w1132 = w1102 & ~w1128;
assign w1133 = w1131 & w1132;
assign w1134 = ~w1130 & ~w1133;
assign w1135 = ~w1103 & ~w1134;
assign w1136 = w1096 & ~w1102;
assign w1137 = ~w1103 & ~w1136;
assign w1138 = ~w1116 & w1137;
assign w1139 = w1122 & ~w1128;
assign w1140 = w1138 & w1139;
assign w1141 = ~w1096 & ~w1102;
assign w1142 = w1115 & ~w1141;
assign w1143 = ~w1103 & ~w1115;
assign w1144 = ~w1142 & ~w1143;
assign w1145 = w1116 & w1136;
assign w1146 = ~w1144 & ~w1145;
assign w1147 = ~w1096 & ~w1109;
assign w1148 = w1128 & ~w1141;
assign w1149 = ~w1147 & w1148;
assign w1150 = ~w1146 & w1149;
assign w1151 = w1109 & w1141;
assign w1152 = w1128 & w1151;
assign w1153 = w1116 & w1137;
assign w1154 = (~w1128 & ~w1137) | (~w1128 & w64484) | (~w1137 & w64484);
assign w1155 = w1103 & w1115;
assign w1156 = ~w1102 & w1109;
assign w1157 = w1096 & w1156;
assign w1158 = ~w1155 & ~w1157;
assign w1159 = w1154 & w1158;
assign w1160 = w1096 & w1115;
assign w1161 = ~w1109 & w1160;
assign w1162 = w1128 & ~w1161;
assign w1163 = ~w1144 & w1162;
assign w1164 = ~w1159 & ~w1163;
assign w1165 = ~w1102 & w1161;
assign w1166 = ~w1152 & ~w1165;
assign w1167 = ~w1164 & w1166;
assign w1168 = ~w1122 & ~w1167;
assign w1169 = w1142 & w1162;
assign w1170 = ~w1136 & ~w1154;
assign w1171 = w1116 & ~w1170;
assign w1172 = ~w1169 & ~w1171;
assign w1173 = w1122 & ~w1172;
assign w1174 = ~w1135 & ~w1140;
assign w1175 = ~w1150 & w1174;
assign w1176 = ~w1168 & w1175;
assign w1177 = ~w1173 & w1176;
assign w1178 = w892 & ~w1076;
assign w1179 = ~w927 & ~w1071;
assign w1180 = ~w914 & ~w1030;
assign w1181 = w1179 & ~w1180;
assign w1182 = w892 & w1042;
assign w1183 = w892 & ~w1179;
assign w1184 = w896 & ~w1183;
assign w1185 = w1024 & ~w1182;
assign w1186 = ~w1184 & w1185;
assign w1187 = ~w926 & w1077;
assign w1188 = ~w921 & ~w1187;
assign w1189 = ~w1183 & w1188;
assign w1190 = ~w1186 & ~w1189;
assign w1191 = ~w1178 & ~w1181;
assign w1192 = ~w1190 & w1191;
assign w1193 = w1131 & w1136;
assign w1194 = ~w1102 & w1115;
assign w1195 = ~w1136 & ~w1194;
assign w1196 = w1109 & w1195;
assign w1197 = ~w1167 & w1196;
assign w1198 = ~w1131 & w1138;
assign w1199 = ~w1193 & ~w1198;
assign w1200 = ~w1171 & w1199;
assign w1201 = ~w1197 & w1200;
assign w1202 = ~w1122 & ~w1201;
assign w1203 = w1147 & w1163;
assign w1204 = w1102 & ~w1109;
assign w1205 = ~w1156 & ~w1160;
assign w1206 = w1128 & ~w1205;
assign w1207 = w1204 & w1206;
assign w1208 = w1096 & w1102;
assign w1209 = w1122 & w1131;
assign w1210 = ~w1208 & w1209;
assign w1211 = ~w1207 & ~w1210;
assign w1212 = w1137 & ~w1211;
assign w1213 = w1158 & ~w1204;
assign w1214 = w1129 & ~w1213;
assign w1215 = ~w1147 & ~w1156;
assign w1216 = w1139 & w1215;
assign w1217 = w1213 & w1216;
assign w1218 = ~w1203 & ~w1214;
assign w1219 = ~w1217 & w1218;
assign w1220 = ~w1212 & w1219;
assign w1221 = ~w1202 & w1220;
assign w1222 = w1129 & ~w1146;
assign w1223 = ~w1109 & w1155;
assign w1224 = ~w1128 & ~w1160;
assign w1225 = w1215 & w1224;
assign w1226 = ~w1153 & ~w1223;
assign w1227 = ~w1225 & w1226;
assign w1228 = ~w1122 & ~w1227;
assign w1229 = w1109 & w1194;
assign w1230 = ~w1122 & ~w1229;
assign w1231 = w1206 & w1230;
assign w1232 = ~w1151 & ~w1160;
assign w1233 = ~w1128 & ~w1230;
assign w1234 = ~w1232 & w1233;
assign w1235 = w1211 & ~w1231;
assign w1236 = ~w1222 & ~w1234;
assign w1237 = w1235 & w1236;
assign w1238 = ~w1228 & w1237;
assign w1239 = ~w1128 & w1161;
assign w1240 = w1103 & w1209;
assign w1241 = ~w1195 & w1224;
assign w1242 = ~w1109 & ~w1137;
assign w1243 = w1109 & w1208;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = ~w1152 & w1244;
assign w1246 = ~w1115 & ~w1245;
assign w1247 = w1122 & ~w1241;
assign w1248 = ~w1246 & w1247;
assign w1249 = w1102 & w1244;
assign w1250 = ~w1128 & w1195;
assign w1251 = ~w1249 & w1250;
assign w1252 = w1149 & w1244;
assign w1253 = w1116 & w1141;
assign w1254 = ~w1122 & ~w1253;
assign w1255 = ~w1252 & w1254;
assign w1256 = ~w1251 & w1255;
assign w1257 = ~w1248 & ~w1256;
assign w1258 = ~w1151 & w1194;
assign w1259 = w1162 & w1258;
assign w1260 = ~w1239 & ~w1240;
assign w1261 = ~w1259 & w1260;
assign w1262 = ~w1257 & w1261;
assign w1263 = ~pi3031 & pi9040;
assign w1264 = ~pi3013 & ~pi9040;
assign w1265 = ~w1263 & ~w1264;
assign w1266 = pi0107 & ~w1265;
assign w1267 = ~pi0107 & w1265;
assign w1268 = ~w1266 & ~w1267;
assign w1269 = ~pi3062 & pi9040;
assign w1270 = ~pi3029 & ~pi9040;
assign w1271 = ~w1269 & ~w1270;
assign w1272 = pi0146 & ~w1271;
assign w1273 = ~pi0146 & w1271;
assign w1274 = ~w1272 & ~w1273;
assign w1275 = w1268 & w1274;
assign w1276 = ~pi3054 & pi9040;
assign w1277 = ~pi3127 & ~pi9040;
assign w1278 = ~w1276 & ~w1277;
assign w1279 = pi0156 & ~w1278;
assign w1280 = ~pi0156 & w1278;
assign w1281 = ~w1279 & ~w1280;
assign w1282 = ~pi3165 & pi9040;
assign w1283 = ~pi3097 & ~pi9040;
assign w1284 = ~w1282 & ~w1283;
assign w1285 = pi0127 & ~w1284;
assign w1286 = ~pi0127 & w1284;
assign w1287 = ~w1285 & ~w1286;
assign w1288 = w1281 & w1287;
assign w1289 = ~pi3035 & pi9040;
assign w1290 = ~pi3067 & ~pi9040;
assign w1291 = ~w1289 & ~w1290;
assign w1292 = pi0129 & ~w1291;
assign w1293 = ~pi0129 & w1291;
assign w1294 = ~w1292 & ~w1293;
assign w1295 = ~w1288 & w1294;
assign w1296 = w1275 & ~w1295;
assign w1297 = w1274 & w1281;
assign w1298 = w1268 & ~w1274;
assign w1299 = ~w1288 & w1298;
assign w1300 = w1294 & ~w1299;
assign w1301 = w1268 & ~w1287;
assign w1302 = ~w1275 & ~w1301;
assign w1303 = w1294 & ~w1302;
assign w1304 = ~w1300 & ~w1303;
assign w1305 = ~w1281 & ~w1287;
assign w1306 = ~w1288 & ~w1305;
assign w1307 = ~w1297 & w1306;
assign w1308 = w1304 & w1307;
assign w1309 = (~w1296 & ~w1304) | (~w1296 & w64485) | (~w1304 & w64485);
assign w1310 = ~pi3029 & pi9040;
assign w1311 = ~pi3065 & ~pi9040;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = pi0150 & ~w1312;
assign w1314 = ~pi0150 & w1312;
assign w1315 = ~w1313 & ~w1314;
assign w1316 = ~w1309 & ~w1315;
assign w1317 = w1297 & w1301;
assign w1318 = ~w1281 & w1287;
assign w1319 = ~w1298 & ~w1318;
assign w1320 = ~w1304 & ~w1319;
assign w1321 = ~w1268 & w1294;
assign w1322 = w1268 & ~w1318;
assign w1323 = ~w1321 & ~w1322;
assign w1324 = (~w1317 & ~w1323) | (~w1317 & w64486) | (~w1323 & w64486);
assign w1325 = ~w1320 & w1324;
assign w1326 = (w1315 & w1320) | (w1315 & w64487) | (w1320 & w64487);
assign w1327 = ~w1268 & w1274;
assign w1328 = ~w1287 & w1327;
assign w1329 = ~w1274 & w1281;
assign w1330 = ~w1268 & w1287;
assign w1331 = w1329 & w1330;
assign w1332 = ~w1328 & ~w1331;
assign w1333 = ~w1315 & ~w1332;
assign w1334 = ~w1268 & w1305;
assign w1335 = w1305 & w64488;
assign w1336 = w1306 & w1327;
assign w1337 = w1301 & w1329;
assign w1338 = ~w1335 & ~w1337;
assign w1339 = ~w1336 & w1338;
assign w1340 = ~w1333 & w1339;
assign w1341 = w1294 & ~w1340;
assign w1342 = ~w1274 & ~w1281;
assign w1343 = ~w1268 & w1288;
assign w1344 = w1288 & w1327;
assign w1345 = ~w1342 & ~w1344;
assign w1346 = w1287 & ~w1294;
assign w1347 = ~w1345 & w1346;
assign w1348 = w1268 & w1347;
assign w1349 = ~w1316 & ~w1348;
assign w1350 = ~w1326 & ~w1341;
assign w1351 = w1349 & w1350;
assign w1352 = ~pi0162 & ~w1351;
assign w1353 = pi0162 & w1351;
assign w1354 = ~w1352 & ~w1353;
assign w1355 = ~pi3114 & pi9040;
assign w1356 = ~pi3054 & ~pi9040;
assign w1357 = ~w1355 & ~w1356;
assign w1358 = pi0107 & ~w1357;
assign w1359 = ~pi0107 & w1357;
assign w1360 = ~w1358 & ~w1359;
assign w1361 = ~pi3057 & pi9040;
assign w1362 = ~pi3027 & ~pi9040;
assign w1363 = ~w1361 & ~w1362;
assign w1364 = pi0155 & ~w1363;
assign w1365 = ~pi0155 & w1363;
assign w1366 = ~w1364 & ~w1365;
assign w1367 = w1360 & w1366;
assign w1368 = ~pi3099 & pi9040;
assign w1369 = ~pi3165 & ~pi9040;
assign w1370 = ~w1368 & ~w1369;
assign w1371 = pi0142 & ~w1370;
assign w1372 = ~pi0142 & w1370;
assign w1373 = ~w1371 & ~w1372;
assign w1374 = ~pi3013 & pi9040;
assign w1375 = ~pi3035 & ~pi9040;
assign w1376 = ~w1374 & ~w1375;
assign w1377 = pi0143 & ~w1376;
assign w1378 = ~pi0143 & w1376;
assign w1379 = ~w1377 & ~w1378;
assign w1380 = ~w1373 & ~w1379;
assign w1381 = w1367 & w1380;
assign w1382 = ~pi3022 & pi9040;
assign w1383 = ~pi3048 & ~pi9040;
assign w1384 = ~w1382 & ~w1383;
assign w1385 = pi0127 & ~w1384;
assign w1386 = ~pi0127 & w1384;
assign w1387 = ~w1385 & ~w1386;
assign w1388 = w1360 & ~w1373;
assign w1389 = ~w1360 & ~w1373;
assign w1390 = ~w1360 & ~w1366;
assign w1391 = ~w1367 & ~w1390;
assign w1392 = ~w1379 & ~w1391;
assign w1393 = ~w1391 & w64489;
assign w1394 = ~pi3126 & pi9040;
assign w1395 = ~pi3114 & ~pi9040;
assign w1396 = ~w1394 & ~w1395;
assign w1397 = pi0149 & ~w1396;
assign w1398 = ~pi0149 & w1396;
assign w1399 = ~w1397 & ~w1398;
assign w1400 = ~w1393 & w1399;
assign w1401 = w1388 & w1400;
assign w1402 = w1360 & w1373;
assign w1403 = ~w1389 & ~w1402;
assign w1404 = ~w1366 & w1379;
assign w1405 = w1403 & w1404;
assign w1406 = ~w1401 & w1405;
assign w1407 = w1380 & w1390;
assign w1408 = w1366 & w1373;
assign w1409 = ~w1407 & ~w1408;
assign w1410 = w1399 & ~w1409;
assign w1411 = w1373 & w1379;
assign w1412 = ~w1360 & ~w1379;
assign w1413 = ~w1388 & ~w1412;
assign w1414 = w1391 & ~w1411;
assign w1415 = w1413 & w1414;
assign w1416 = ~w1381 & w1387;
assign w1417 = ~w1410 & w1416;
assign w1418 = ~w1415 & w1417;
assign w1419 = ~w1406 & w1418;
assign w1420 = ~w1373 & w1379;
assign w1421 = w1367 & w1420;
assign w1422 = w1373 & w1391;
assign w1423 = w1391 & w1411;
assign w1424 = ~w1421 & ~w1423;
assign w1425 = ~w1399 & ~w1424;
assign w1426 = w1373 & w1390;
assign w1427 = w1380 & w1391;
assign w1428 = ~w1421 & ~w1426;
assign w1429 = ~w1427 & w1428;
assign w1430 = w1412 & ~w1429;
assign w1431 = w1399 & ~w1404;
assign w1432 = ~w1403 & ~w1431;
assign w1433 = ~w1387 & ~w1421;
assign w1434 = ~w1432 & w1433;
assign w1435 = ~w1430 & w1434;
assign w1436 = w1435 & w64490;
assign w1437 = ~w1419 & ~w1436;
assign w1438 = ~pi0166 & w1437;
assign w1439 = pi0166 & ~w1437;
assign w1440 = ~w1438 & ~w1439;
assign w1441 = ~pi3037 & pi9040;
assign w1442 = ~pi3041 & ~pi9040;
assign w1443 = ~w1441 & ~w1442;
assign w1444 = pi0122 & ~w1443;
assign w1445 = ~pi0122 & w1443;
assign w1446 = ~w1444 & ~w1445;
assign w1447 = ~pi3098 & pi9040;
assign w1448 = ~pi3056 & ~pi9040;
assign w1449 = ~w1447 & ~w1448;
assign w1450 = pi0131 & ~w1449;
assign w1451 = ~pi0131 & w1449;
assign w1452 = ~w1450 & ~w1451;
assign w1453 = w1446 & ~w1452;
assign w1454 = ~pi3056 & pi9040;
assign w1455 = ~pi3102 & ~pi9040;
assign w1456 = ~w1454 & ~w1455;
assign w1457 = pi0157 & ~w1456;
assign w1458 = ~pi0157 & w1456;
assign w1459 = ~w1457 & ~w1458;
assign w1460 = ~pi3019 & pi9040;
assign w1461 = ~pi3024 & ~pi9040;
assign w1462 = ~w1460 & ~w1461;
assign w1463 = pi0140 & ~w1462;
assign w1464 = ~pi0140 & w1462;
assign w1465 = ~w1463 & ~w1464;
assign w1466 = ~w1459 & w1465;
assign w1467 = ~w1453 & w1466;
assign w1468 = ~pi3123 & pi9040;
assign w1469 = ~pi3032 & ~pi9040;
assign w1470 = ~w1468 & ~w1469;
assign w1471 = pi0145 & ~w1470;
assign w1472 = ~pi0145 & w1470;
assign w1473 = ~w1471 & ~w1472;
assign w1474 = w1452 & w1465;
assign w1475 = ~w1446 & ~w1459;
assign w1476 = w1474 & w1475;
assign w1477 = ~w1473 & ~w1476;
assign w1478 = w1467 & w1477;
assign w1479 = ~w1446 & w1465;
assign w1480 = w1446 & ~w1465;
assign w1481 = ~w1479 & ~w1480;
assign w1482 = ~w1459 & ~w1481;
assign w1483 = w1452 & w1473;
assign w1484 = ~w1446 & ~w1452;
assign w1485 = ~pi3041 & pi9040;
assign w1486 = ~pi3061 & ~pi9040;
assign w1487 = ~w1485 & ~w1486;
assign w1488 = pi0153 & ~w1487;
assign w1489 = ~pi0153 & w1487;
assign w1490 = ~w1488 & ~w1489;
assign w1491 = ~w1484 & ~w1490;
assign w1492 = ~w1483 & ~w1491;
assign w1493 = w1482 & ~w1492;
assign w1494 = w1446 & ~w1473;
assign w1495 = w1452 & ~w1465;
assign w1496 = ~w1459 & w1480;
assign w1497 = ~w1495 & ~w1496;
assign w1498 = w1494 & ~w1497;
assign w1499 = ~w1452 & w1498;
assign w1500 = w1446 & w1459;
assign w1501 = ~w1452 & ~w1500;
assign w1502 = ~w1473 & ~w1474;
assign w1503 = ~w1501 & w1502;
assign w1504 = w1475 & w1503;
assign w1505 = ~w1446 & w1473;
assign w1506 = ~w1494 & ~w1505;
assign w1507 = w1452 & ~w1506;
assign w1508 = w1452 & w1479;
assign w1509 = ~w1507 & ~w1508;
assign w1510 = w1459 & ~w1509;
assign w1511 = w1459 & w1465;
assign w1512 = w1453 & w1511;
assign w1513 = ~w1465 & ~w1473;
assign w1514 = ~w1511 & ~w1513;
assign w1515 = w1484 & w1514;
assign w1516 = w1490 & ~w1512;
assign w1517 = ~w1515 & w1516;
assign w1518 = ~w1504 & w1517;
assign w1519 = ~w1510 & w1518;
assign w1520 = ~w1467 & ~w1508;
assign w1521 = w1465 & w1473;
assign w1522 = w1520 & w1521;
assign w1523 = w1459 & w1481;
assign w1524 = w1452 & ~w1523;
assign w1525 = w1513 & ~w1524;
assign w1526 = ~w1490 & ~w1522;
assign w1527 = ~w1525 & w1526;
assign w1528 = ~w1519 & ~w1527;
assign w1529 = ~w1478 & ~w1493;
assign w1530 = ~w1499 & w1529;
assign w1531 = ~w1528 & w1530;
assign w1532 = pi0168 & ~w1531;
assign w1533 = ~pi0168 & w1531;
assign w1534 = ~w1532 & ~w1533;
assign w1535 = w1453 & w1466;
assign w1536 = w1473 & ~w1535;
assign w1537 = ~w1452 & ~w1465;
assign w1538 = ~w1475 & ~w1500;
assign w1539 = w1537 & ~w1538;
assign w1540 = w1536 & ~w1539;
assign w1541 = ~w1477 & ~w1540;
assign w1542 = ~w1481 & w64491;
assign w1543 = w1481 & w63521;
assign w1544 = w1475 & w1537;
assign w1545 = ~w1473 & ~w1544;
assign w1546 = ~w1543 & w1545;
assign w1547 = w1523 & w1546;
assign w1548 = w1546 & w64492;
assign w1549 = w1474 & ~w1538;
assign w1550 = ~w1474 & ~w1537;
assign w1551 = w1473 & w1481;
assign w1552 = w1550 & w1551;
assign w1553 = (w1490 & w1538) | (w1490 & w64493) | (w1538 & w64493);
assign w1554 = ~w1542 & w1553;
assign w1555 = ~w1552 & w1554;
assign w1556 = ~w1548 & w1555;
assign w1557 = w1505 & w1511;
assign w1558 = w1452 & w1496;
assign w1559 = w1484 & w1511;
assign w1560 = ~w1544 & ~w1559;
assign w1561 = ~w1550 & w1551;
assign w1562 = ~w1490 & ~w1557;
assign w1563 = ~w1503 & w1562;
assign w1564 = ~w1558 & w1560;
assign w1565 = w1563 & w1564;
assign w1566 = ~w1561 & w1565;
assign w1567 = ~w1556 & ~w1566;
assign w1568 = ~w1541 & ~w1567;
assign w1569 = pi0160 & w1568;
assign w1570 = ~pi0160 & ~w1568;
assign w1571 = ~w1569 & ~w1570;
assign w1572 = ~w1315 & w1330;
assign w1573 = w1342 & w1572;
assign w1574 = ~w1337 & ~w1343;
assign w1575 = ~w1287 & ~w1342;
assign w1576 = w1268 & ~w1575;
assign w1577 = ~w1328 & ~w1576;
assign w1578 = w1305 & w1577;
assign w1579 = ~w1294 & ~w1572;
assign w1580 = w1574 & w1579;
assign w1581 = ~w1578 & w1580;
assign w1582 = w1305 & w1327;
assign w1583 = w1315 & ~w1582;
assign w1584 = ~w1577 & ~w1583;
assign w1585 = w1294 & ~w1317;
assign w1586 = ~w1584 & w1585;
assign w1587 = ~w1581 & ~w1586;
assign w1588 = ~w1268 & ~w1297;
assign w1589 = w1323 & ~w1588;
assign w1590 = ~w1274 & ~w1287;
assign w1591 = w1321 & w1590;
assign w1592 = ~w1337 & ~w1591;
assign w1593 = ~w1344 & w1592;
assign w1594 = ~w1589 & w1593;
assign w1595 = w1315 & ~w1594;
assign w1596 = ~w1573 & ~w1595;
assign w1597 = ~w1587 & w1596;
assign w1598 = ~pi0190 & w1597;
assign w1599 = pi0190 & ~w1597;
assign w1600 = ~w1598 & ~w1599;
assign w1601 = w1275 & w1318;
assign w1602 = ~w1334 & ~w1601;
assign w1603 = w1325 & ~w1602;
assign w1604 = ~w1281 & w1327;
assign w1605 = ~w1322 & ~w1604;
assign w1606 = w1300 & ~w1605;
assign w1607 = w1329 & w1574;
assign w1608 = w1583 & ~w1606;
assign w1609 = w1608 & w64494;
assign w1610 = w1287 & w1298;
assign w1611 = ~w1343 & ~w1610;
assign w1612 = w1294 & ~w1611;
assign w1613 = ~w1287 & ~w1294;
assign w1614 = w1298 & w1613;
assign w1615 = ~w1315 & ~w1614;
assign w1616 = w1274 & ~w1294;
assign w1617 = ~w1301 & ~w1616;
assign w1618 = w1306 & ~w1617;
assign w1619 = ~w1331 & ~w1601;
assign w1620 = ~w1335 & w1619;
assign w1621 = w1615 & ~w1618;
assign w1622 = w1620 & w1621;
assign w1623 = ~w1612 & w1622;
assign w1624 = ~w1609 & ~w1623;
assign w1625 = ~w1603 & ~w1624;
assign w1626 = ~pi0191 & w1625;
assign w1627 = pi0191 & ~w1625;
assign w1628 = ~w1626 & ~w1627;
assign w1629 = ~pi3164 & pi9040;
assign w1630 = ~pi3026 & ~pi9040;
assign w1631 = ~w1629 & ~w1630;
assign w1632 = pi0120 & ~w1631;
assign w1633 = ~pi0120 & w1631;
assign w1634 = ~w1632 & ~w1633;
assign w1635 = ~pi3095 & pi9040;
assign w1636 = ~pi3012 & ~pi9040;
assign w1637 = ~w1635 & ~w1636;
assign w1638 = pi0144 & ~w1637;
assign w1639 = ~pi0144 & w1637;
assign w1640 = ~w1638 & ~w1639;
assign w1641 = ~w1634 & ~w1640;
assign w1642 = ~pi3012 & pi9040;
assign w1643 = ~pi3164 & ~pi9040;
assign w1644 = ~w1642 & ~w1643;
assign w1645 = pi0119 & ~w1644;
assign w1646 = ~pi0119 & w1644;
assign w1647 = ~w1645 & ~w1646;
assign w1648 = ~w1640 & w1647;
assign w1649 = ~w1641 & ~w1648;
assign w1650 = ~pi3061 & pi9040;
assign w1651 = ~pi3019 & ~pi9040;
assign w1652 = ~w1650 & ~w1651;
assign w1653 = pi0152 & ~w1652;
assign w1654 = ~pi0152 & w1652;
assign w1655 = ~w1653 & ~w1654;
assign w1656 = w1634 & ~w1655;
assign w1657 = ~pi3052 & pi9040;
assign w1658 = ~pi3020 & ~pi9040;
assign w1659 = ~w1657 & ~w1658;
assign w1660 = pi0151 & ~w1659;
assign w1661 = ~pi0151 & w1659;
assign w1662 = ~w1660 & ~w1661;
assign w1663 = ~w1634 & w1662;
assign w1664 = ~w1647 & ~w1663;
assign w1665 = (w1662 & w1663) | (w1662 & w63522) | (w1663 & w63522);
assign w1666 = w1656 & w1665;
assign w1667 = ~w1634 & w1647;
assign w1668 = ~w1634 & ~w1655;
assign w1669 = ~w1667 & ~w1668;
assign w1670 = w1647 & ~w1662;
assign w1671 = w1634 & w1655;
assign w1672 = ~w1668 & ~w1671;
assign w1673 = w1670 & ~w1672;
assign w1674 = ~pi3051 & pi9040;
assign w1675 = ~pi3059 & ~pi9040;
assign w1676 = ~w1674 & ~w1675;
assign w1677 = pi0148 & ~w1676;
assign w1678 = ~pi0148 & w1676;
assign w1679 = ~w1677 & ~w1678;
assign w1680 = (~w1679 & w1673) | (~w1679 & w63523) | (w1673 & w63523);
assign w1681 = ~w1647 & w1662;
assign w1682 = ~w1666 & ~w1681;
assign w1683 = ~w1680 & w1682;
assign w1684 = ~w1649 & ~w1683;
assign w1685 = ~w1655 & ~w1662;
assign w1686 = ~w1671 & ~w1685;
assign w1687 = ~w1640 & ~w1647;
assign w1688 = w1655 & w1662;
assign w1689 = ~w1647 & w1688;
assign w1690 = ~w1634 & w1689;
assign w1691 = ~w1647 & ~w1656;
assign w1692 = w1672 & ~w1681;
assign w1693 = w1640 & ~w1691;
assign w1694 = ~w1692 & w1693;
assign w1695 = (~w1640 & w1669) | (~w1640 & w64495) | (w1669 & w64495);
assign w1696 = w1670 & ~w1695;
assign w1697 = (w1679 & w1686) | (w1679 & w64496) | (w1686 & w64496);
assign w1698 = ~w1690 & w1697;
assign w1699 = ~w1694 & w1698;
assign w1700 = ~w1696 & w1699;
assign w1701 = w1668 & w1681;
assign w1702 = w1667 & w1688;
assign w1703 = ~w1679 & ~w1702;
assign w1704 = w1640 & ~w1647;
assign w1705 = ~w1686 & w1704;
assign w1706 = ~w1701 & w1703;
assign w1707 = ~w1705 & w1706;
assign w1708 = ~w1666 & w1707;
assign w1709 = ~w1700 & ~w1708;
assign w1710 = ~w1684 & ~w1709;
assign w1711 = pi0174 & w1710;
assign w1712 = ~pi0174 & ~w1710;
assign w1713 = ~w1711 & ~w1712;
assign w1714 = w1424 & w63348;
assign w1715 = w1366 & w1399;
assign w1716 = ~w1373 & w1715;
assign w1717 = (~w1420 & w1714) | (~w1420 & w63524) | (w1714 & w63524);
assign w1718 = ~w1389 & ~w1404;
assign w1719 = w1390 & w1420;
assign w1720 = ~w1718 & ~w1719;
assign w1721 = ~w1392 & ~w1399;
assign w1722 = ~w1720 & w1721;
assign w1723 = (~w1387 & w1717) | (~w1387 & w64497) | (w1717 & w64497);
assign w1724 = ~w1388 & w1399;
assign w1725 = w1380 & w1724;
assign w1726 = w1424 & w64498;
assign w1727 = w1720 & w1726;
assign w1728 = w1388 & w1404;
assign w1729 = w1366 & ~w1379;
assign w1730 = w1402 & w1729;
assign w1731 = (w1715 & w1730) | (w1715 & w63525) | (w1730 & w63525);
assign w1732 = ~w1366 & w1402;
assign w1733 = ~w1381 & ~w1732;
assign w1734 = ~w1399 & ~w1733;
assign w1735 = ~w1407 & ~w1728;
assign w1736 = ~w1731 & w1735;
assign w1737 = ~w1734 & w1736;
assign w1738 = w1373 & ~w1399;
assign w1739 = ~w1404 & w1738;
assign w1740 = ~w1729 & w1739;
assign w1741 = ~w1725 & ~w1740;
assign w1742 = (w1741 & w1737) | (w1741 & w64499) | (w1737 & w64499);
assign w1743 = ~w1727 & w1742;
assign w1744 = ~w1723 & w1743;
assign w1745 = pi0171 & ~w1744;
assign w1746 = ~pi0171 & w1744;
assign w1747 = ~w1745 & ~w1746;
assign w1748 = ~w1506 & w64500;
assign w1749 = w1446 & w1514;
assign w1750 = ~w1558 & w1749;
assign w1751 = w1560 & ~w1748;
assign w1752 = ~w1750 & w1751;
assign w1753 = ~w1548 & w1752;
assign w1754 = ~w1490 & ~w1753;
assign w1755 = w1453 & ~w1466;
assign w1756 = ~w1476 & ~w1755;
assign w1757 = ~w1473 & ~w1756;
assign w1758 = (w1490 & w1757) | (w1490 & w64501) | (w1757 & w64501);
assign w1759 = ~w1536 & ~w1546;
assign w1760 = ~w1484 & ~w1496;
assign w1761 = w1473 & w1490;
assign w1762 = ~w1537 & w1761;
assign w1763 = ~w1760 & w1762;
assign w1764 = ~w1557 & ~w1763;
assign w1765 = ~w1758 & w1764;
assign w1766 = ~w1759 & w1765;
assign w1767 = ~w1754 & w1766;
assign w1768 = pi0163 & ~w1767;
assign w1769 = ~pi0163 & w1767;
assign w1770 = ~w1768 & ~w1769;
assign w1771 = ~w1497 & w1761;
assign w1772 = ~w1473 & ~w1520;
assign w1773 = ~w1474 & w1523;
assign w1774 = w1490 & ~w1772;
assign w1775 = ~w1773 & w1774;
assign w1776 = ~w1490 & ~w1535;
assign w1777 = ~w1549 & w1776;
assign w1778 = ~w1498 & w1777;
assign w1779 = ~w1775 & ~w1778;
assign w1780 = ~w1452 & ~w1490;
assign w1781 = ~w1511 & w1780;
assign w1782 = ~w1538 & w1781;
assign w1783 = ~w1559 & ~w1782;
assign w1784 = ~w1543 & w1783;
assign w1785 = w1473 & ~w1784;
assign w1786 = ~w1547 & ~w1771;
assign w1787 = ~w1785 & w1786;
assign w1788 = ~w1779 & w1787;
assign w1789 = pi0167 & w1788;
assign w1790 = ~pi0167 & ~w1788;
assign w1791 = ~w1789 & ~w1790;
assign w1792 = w1634 & w1640;
assign w1793 = ~w1681 & w1792;
assign w1794 = ~w1647 & ~w1655;
assign w1795 = w1634 & ~w1662;
assign w1796 = w1794 & ~w1795;
assign w1797 = ~w1702 & ~w1796;
assign w1798 = ~w1640 & ~w1797;
assign w1799 = w1679 & ~w1793;
assign w1800 = ~w1673 & w1799;
assign w1801 = ~w1798 & w1800;
assign w1802 = ~w1667 & w1672;
assign w1803 = w1672 & w64502;
assign w1804 = ~w1649 & ~w1670;
assign w1805 = w1797 & w1804;
assign w1806 = (~w1679 & ~w1702) | (~w1679 & w64503) | (~w1702 & w64503);
assign w1807 = ~w1803 & w1806;
assign w1808 = ~w1805 & w1807;
assign w1809 = ~w1801 & ~w1808;
assign w1810 = w1655 & ~w1665;
assign w1811 = ~w1641 & ~w1662;
assign w1812 = w1810 & ~w1811;
assign w1813 = w1679 & ~w1695;
assign w1814 = w1812 & ~w1813;
assign w1815 = ~w1701 & ~w1795;
assign w1816 = w1634 & w1647;
assign w1817 = (~w1816 & w1673) | (~w1816 & w64504) | (w1673 & w64504);
assign w1818 = w1640 & ~w1817;
assign w1819 = ~w1815 & w1818;
assign w1820 = ~w1809 & ~w1814;
assign w1821 = ~w1819 & w1820;
assign w1822 = pi0179 & ~w1821;
assign w1823 = ~pi0179 & w1821;
assign w1824 = ~w1822 & ~w1823;
assign w1825 = ~pi3100 & pi9040;
assign w1826 = ~pi3124 & ~pi9040;
assign w1827 = ~w1825 & ~w1826;
assign w1828 = pi0114 & ~w1827;
assign w1829 = ~pi0114 & w1827;
assign w1830 = ~w1828 & ~w1829;
assign w1831 = ~pi3055 & pi9040;
assign w1832 = ~pi3039 & ~pi9040;
assign w1833 = ~w1831 & ~w1832;
assign w1834 = pi0147 & ~w1833;
assign w1835 = ~pi0147 & w1833;
assign w1836 = ~w1834 & ~w1835;
assign w1837 = ~w1830 & w1836;
assign w1838 = ~pi3124 & pi9040;
assign w1839 = ~pi3015 & ~pi9040;
assign w1840 = ~w1838 & ~w1839;
assign w1841 = pi0142 & ~w1840;
assign w1842 = ~pi0142 & w1840;
assign w1843 = ~w1841 & ~w1842;
assign w1844 = ~pi3015 & pi9040;
assign w1845 = ~pi3031 & ~pi9040;
assign w1846 = ~w1844 & ~w1845;
assign w1847 = pi0141 & ~w1846;
assign w1848 = ~pi0141 & w1846;
assign w1849 = ~w1847 & ~w1848;
assign w1850 = w1843 & w1849;
assign w1851 = w1837 & w1850;
assign w1852 = ~pi3017 & pi9040;
assign w1853 = ~pi3101 & ~pi9040;
assign w1854 = ~w1852 & ~w1853;
assign w1855 = pi0132 & ~w1854;
assign w1856 = ~pi0132 & w1854;
assign w1857 = ~w1855 & ~w1856;
assign w1858 = ~w1843 & w1857;
assign w1859 = ~w1836 & w1858;
assign w1860 = w1858 & w64505;
assign w1861 = ~w1830 & ~w1849;
assign w1862 = w1858 & w1861;
assign w1863 = ~pi3067 & pi9040;
assign w1864 = ~pi3017 & ~pi9040;
assign w1865 = ~w1863 & ~w1864;
assign w1866 = pi0155 & ~w1865;
assign w1867 = ~pi0155 & w1865;
assign w1868 = ~w1866 & ~w1867;
assign w1869 = w1830 & ~w1836;
assign w1870 = w1843 & w1857;
assign w1871 = w1869 & w1870;
assign w1872 = ~w1836 & ~w1857;
assign w1873 = w1843 & ~w1869;
assign w1874 = w1872 & w1873;
assign w1875 = ~w1843 & ~w1857;
assign w1876 = w1869 & w1875;
assign w1877 = w1843 & ~w1857;
assign w1878 = ~w1830 & ~w1857;
assign w1879 = ~w1877 & ~w1878;
assign w1880 = w1858 & w64506;
assign w1881 = (w1849 & w1879) | (w1849 & w64507) | (w1879 & w64507);
assign w1882 = ~w1880 & w1881;
assign w1883 = ~w1837 & w1875;
assign w1884 = w1830 & w1870;
assign w1885 = ~w1849 & ~w1883;
assign w1886 = ~w1884 & w1885;
assign w1887 = ~w1882 & ~w1886;
assign w1888 = ~w1862 & w1868;
assign w1889 = ~w1871 & ~w1876;
assign w1890 = w1888 & w1889;
assign w1891 = ~w1874 & w1890;
assign w1892 = ~w1887 & w1891;
assign w1893 = w1869 & w1877;
assign w1894 = w1836 & w1870;
assign w1895 = ~w1859 & ~w1894;
assign w1896 = (~w1876 & ~w1895) | (~w1876 & w63526) | (~w1895 & w63526);
assign w1897 = w1849 & ~w1896;
assign w1898 = ~w1858 & ~w1872;
assign w1899 = ~w1830 & w1898;
assign w1900 = ~w1849 & ~w1880;
assign w1901 = ~w1899 & w1900;
assign w1902 = ~w1868 & ~w1893;
assign w1903 = (w1902 & w1897) | (w1902 & w64508) | (w1897 & w64508);
assign w1904 = ~w1892 & ~w1903;
assign w1905 = ~w1851 & ~w1860;
assign w1906 = ~w1904 & w1905;
assign w1907 = pi0164 & ~w1906;
assign w1908 = ~pi0164 & w1906;
assign w1909 = ~w1907 & ~w1908;
assign w1910 = w1308 & ~w1339;
assign w1911 = w1321 & w1329;
assign w1912 = w1301 & w1616;
assign w1913 = w1303 & ~w1575;
assign w1914 = ~w1334 & ~w1610;
assign w1915 = ~w1294 & ~w1914;
assign w1916 = w1315 & ~w1317;
assign w1917 = ~w1331 & ~w1604;
assign w1918 = ~w1912 & w1917;
assign w1919 = w1916 & w1918;
assign w1920 = ~w1913 & ~w1915;
assign w1921 = w1919 & w1920;
assign w1922 = ~w1328 & ~w1346;
assign w1923 = w1297 & ~w1922;
assign w1924 = ~w1297 & ~w1327;
assign w1925 = w1300 & w1924;
assign w1926 = w1615 & ~w1923;
assign w1927 = ~w1925 & w1926;
assign w1928 = ~w1921 & ~w1927;
assign w1929 = ~w1348 & ~w1911;
assign w1930 = ~w1910 & w1929;
assign w1931 = ~w1928 & w1930;
assign w1932 = ~pi0195 & ~w1931;
assign w1933 = pi0195 & w1931;
assign w1934 = ~w1932 & ~w1933;
assign w1935 = ~w1360 & w1366;
assign w1936 = w1411 & w1935;
assign w1937 = ~w1399 & ~w1429;
assign w1938 = w1360 & w1379;
assign w1939 = ~w1379 & w1935;
assign w1940 = ~w1426 & ~w1938;
assign w1941 = w1724 & ~w1939;
assign w1942 = w1940 & w1941;
assign w1943 = ~w1936 & ~w1942;
assign w1944 = ~w1937 & w1943;
assign w1945 = ~w1399 & ~w1403;
assign w1946 = ~w1939 & w1945;
assign w1947 = w1424 & w64509;
assign w1948 = ~w1413 & w1715;
assign w1949 = ~w1405 & ~w1948;
assign w1950 = ~w1946 & w1949;
assign w1951 = ~w1947 & w1950;
assign w1952 = ~w1387 & ~w1951;
assign w1953 = (~w1399 & ~w1411) | (~w1399 & w64510) | (~w1411 & w64510);
assign w1954 = ~w1730 & w1953;
assign w1955 = w1399 & ~w1728;
assign w1956 = ~w1954 & ~w1955;
assign w1957 = (~w1956 & w1944) | (~w1956 & w64511) | (w1944 & w64511);
assign w1958 = ~w1952 & w1957;
assign w1959 = pi0197 & w1958;
assign w1960 = ~pi0197 & ~w1958;
assign w1961 = ~w1959 & ~w1960;
assign w1962 = w1387 & ~w1399;
assign w1963 = w1719 & ~w1962;
assign w1964 = ~w1380 & ~w1935;
assign w1965 = ~w1729 & ~w1964;
assign w1966 = ~w1422 & w1953;
assign w1967 = ~w1965 & w1966;
assign w1968 = ~w1400 & ~w1967;
assign w1969 = w1387 & w1424;
assign w1970 = ~w1968 & w1969;
assign w1971 = w1393 & ~w1399;
assign w1972 = ~w1387 & ~w1971;
assign w1973 = ~w1726 & w1972;
assign w1974 = ~w1425 & ~w1963;
assign w1975 = (w1974 & w1970) | (w1974 & w64512) | (w1970 & w64512);
assign w1976 = ~pi0200 & w1975;
assign w1977 = pi0200 & ~w1975;
assign w1978 = ~w1976 & ~w1977;
assign w1979 = ~pi3023 & pi9040;
assign w1980 = ~pi3036 & ~pi9040;
assign w1981 = ~w1979 & ~w1980;
assign w1982 = pi0133 & ~w1981;
assign w1983 = ~pi0133 & w1981;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = ~pi3102 & pi9040;
assign w1986 = ~pi3051 & ~pi9040;
assign w1987 = ~w1985 & ~w1986;
assign w1988 = pi0159 & ~w1987;
assign w1989 = ~pi0159 & w1987;
assign w1990 = ~w1988 & ~w1989;
assign w1991 = ~w1984 & w1990;
assign w1992 = ~pi3014 & pi9040;
assign w1993 = ~pi3023 & ~pi9040;
assign w1994 = ~w1992 & ~w1993;
assign w1995 = pi0150 & ~w1994;
assign w1996 = ~pi0150 & w1994;
assign w1997 = ~w1995 & ~w1996;
assign w1998 = ~pi3034 & pi9040;
assign w1999 = ~pi3098 & ~pi9040;
assign w2000 = ~w1998 & ~w1999;
assign w2001 = pi0120 & ~w2000;
assign w2002 = ~pi0120 & w2000;
assign w2003 = ~w2001 & ~w2002;
assign w2004 = w1997 & w2003;
assign w2005 = ~pi3032 & pi9040;
assign w2006 = ~pi3014 & ~pi9040;
assign w2007 = ~w2005 & ~w2006;
assign w2008 = pi0146 & ~w2007;
assign w2009 = ~pi0146 & w2007;
assign w2010 = ~w2008 & ~w2009;
assign w2011 = ~w2003 & ~w2010;
assign w2012 = w2003 & w2010;
assign w2013 = ~w2011 & ~w2012;
assign w2014 = ~w2004 & w2013;
assign w2015 = ~w1991 & w2014;
assign w2016 = w1984 & ~w1990;
assign w2017 = ~w1984 & ~w2003;
assign w2018 = w2010 & w2017;
assign w2019 = ~w2016 & ~w2018;
assign w2020 = w2010 & ~w2017;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = w2015 & w2021;
assign w2023 = ~w1984 & ~w2010;
assign w2024 = w1990 & w1997;
assign w2025 = w2023 & w2024;
assign w2026 = w2004 & w2016;
assign w2027 = w2010 & w2026;
assign w2028 = ~w2025 & ~w2027;
assign w2029 = w1984 & w2011;
assign w2030 = w1990 & ~w1997;
assign w2031 = w2029 & w2030;
assign w2032 = ~w1997 & ~w2003;
assign w2033 = ~w2004 & ~w2032;
assign w2034 = (w1984 & ~w2033) | (w1984 & w64513) | (~w2033 & w64513);
assign w2035 = ~w1984 & ~w2004;
assign w2036 = w1990 & ~w2035;
assign w2037 = ~w2034 & w2036;
assign w2038 = ~w1997 & ~w2010;
assign w2039 = ~w1990 & ~w2038;
assign w2040 = w2029 & w2039;
assign w2041 = w2004 & w2023;
assign w2042 = ~w2040 & ~w2041;
assign w2043 = ~pi3021 & pi9040;
assign w2044 = ~pi3096 & ~pi9040;
assign w2045 = ~w2043 & ~w2044;
assign w2046 = pi0119 & ~w2045;
assign w2047 = ~pi0119 & w2045;
assign w2048 = ~w2046 & ~w2047;
assign w2049 = w2003 & ~w2010;
assign w2050 = ~w1984 & ~w1990;
assign w2051 = ~w2018 & ~w2050;
assign w2052 = ~w1997 & ~w2049;
assign w2053 = ~w2051 & w2052;
assign w2054 = ~w2040 & w64514;
assign w2055 = ~w2053 & w2054;
assign w2056 = ~w2037 & w2055;
assign w2057 = ~w2011 & ~w2030;
assign w2058 = ~w1984 & ~w2032;
assign w2059 = ~w2057 & w2058;
assign w2060 = ~w2032 & ~w2049;
assign w2061 = ~w2017 & ~w2039;
assign w2062 = ~w2060 & w2061;
assign w2063 = ~w2059 & ~w2062;
assign w2064 = w1997 & w2010;
assign w2065 = ~w1990 & w2064;
assign w2066 = w2048 & ~w2065;
assign w2067 = w2063 & w2066;
assign w2068 = ~w2056 & ~w2067;
assign w2069 = w2028 & ~w2031;
assign w2070 = ~w2022 & w2069;
assign w2071 = ~w2068 & w2070;
assign w2072 = ~pi0172 & ~w2071;
assign w2073 = pi0172 & w2071;
assign w2074 = ~w2072 & ~w2073;
assign w2075 = w1850 & w1872;
assign w2076 = ~w1837 & ~w1861;
assign w2077 = w1858 & ~w2076;
assign w2078 = ~w2075 & ~w2077;
assign w2079 = w1836 & ~w1878;
assign w2080 = ~w1837 & w1857;
assign w2081 = w2079 & ~w2080;
assign w2082 = ~w1849 & ~w2081;
assign w2083 = w1857 & w1869;
assign w2084 = w1849 & ~w1878;
assign w2085 = ~w2083 & w2084;
assign w2086 = ~w2082 & ~w2085;
assign w2087 = ~w2077 & w64515;
assign w2088 = (~w1868 & w2086) | (~w1868 & w64516) | (w2086 & w64516);
assign w2089 = ~w1858 & w2079;
assign w2090 = (w1868 & w2089) | (w1868 & w64517) | (w2089 & w64517);
assign w2091 = w1837 & w1875;
assign w2092 = ~w1884 & ~w2091;
assign w2093 = ~w2090 & w2092;
assign w2094 = w1849 & ~w2093;
assign w2095 = ~w2078 & w2086;
assign w2096 = w1861 & w1875;
assign w2097 = ~w1836 & w2096;
assign w2098 = w1836 & ~w1877;
assign w2099 = w1899 & ~w2098;
assign w2100 = w1830 & ~w1898;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = ~w1849 & w1868;
assign w2103 = ~w2101 & w2102;
assign w2104 = (~w2097 & ~w2086) | (~w2097 & w64518) | (~w2086 & w64518);
assign w2105 = ~w2103 & w2104;
assign w2106 = ~w2088 & ~w2094;
assign w2107 = w2105 & w2106;
assign w2108 = pi0161 & ~w2107;
assign w2109 = ~pi0161 & w2107;
assign w2110 = ~w2108 & ~w2109;
assign w2111 = ~pi3018 & pi9040;
assign w2112 = ~pi3099 & ~pi9040;
assign w2113 = ~w2111 & ~w2112;
assign w2114 = pi0131 & ~w2113;
assign w2115 = ~pi0131 & w2113;
assign w2116 = ~w2114 & ~w2115;
assign w2117 = ~pi3027 & pi9040;
assign w2118 = ~pi3030 & ~pi9040;
assign w2119 = ~w2117 & ~w2118;
assign w2120 = pi0153 & ~w2119;
assign w2121 = ~pi0153 & w2119;
assign w2122 = ~w2120 & ~w2121;
assign w2123 = ~w2116 & w2122;
assign w2124 = ~pi3101 & pi9040;
assign w2125 = ~pi3018 & ~pi9040;
assign w2126 = ~w2124 & ~w2125;
assign w2127 = pi0147 & ~w2126;
assign w2128 = ~pi0147 & w2126;
assign w2129 = ~w2127 & ~w2128;
assign w2130 = w2123 & w2129;
assign w2131 = ~pi3039 & pi9040;
assign w2132 = ~pi3022 & ~pi9040;
assign w2133 = ~w2131 & ~w2132;
assign w2134 = pi0112 & ~w2133;
assign w2135 = ~pi0112 & w2133;
assign w2136 = ~w2134 & ~w2135;
assign w2137 = (~w2136 & ~w2123) | (~w2136 & w63527) | (~w2123 & w63527);
assign w2138 = ~w2116 & ~w2137;
assign w2139 = ~pi3048 & pi9040;
assign w2140 = ~pi3126 & ~pi9040;
assign w2141 = ~w2139 & ~w2140;
assign w2142 = pi0154 & ~w2141;
assign w2143 = ~pi0154 & w2141;
assign w2144 = ~w2142 & ~w2143;
assign w2145 = ~w2122 & w2144;
assign w2146 = ~w2129 & w2144;
assign w2147 = w2129 & ~w2144;
assign w2148 = ~w2146 & ~w2147;
assign w2149 = w2116 & ~w2148;
assign w2150 = ~w2145 & w2149;
assign w2151 = w2122 & ~w2129;
assign w2152 = w2116 & ~w2122;
assign w2153 = ~w2123 & ~w2152;
assign w2154 = (~w2151 & w2153) | (~w2151 & w63349) | (w2153 & w63349);
assign w2155 = ~w2129 & ~w2144;
assign w2156 = w2123 & w2155;
assign w2157 = w2136 & ~w2156;
assign w2158 = ~w2154 & w2157;
assign w2159 = ~w2144 & w2152;
assign w2160 = w2137 & ~w2159;
assign w2161 = ~w2158 & ~w2160;
assign w2162 = w2122 & ~w2136;
assign w2163 = (w2116 & w2161) | (w2116 & w64519) | (w2161 & w64519);
assign w2164 = ~w2116 & w2144;
assign w2165 = ~w2151 & w2164;
assign w2166 = ~pi3127 & pi9040;
assign w2167 = ~pi3057 & ~pi9040;
assign w2168 = ~w2166 & ~w2167;
assign w2169 = pi0132 & ~w2168;
assign w2170 = ~pi0132 & w2168;
assign w2171 = ~w2169 & ~w2170;
assign w2172 = ~w2165 & ~w2171;
assign w2173 = ~w2138 & w2172;
assign w2174 = ~w2163 & w2173;
assign w2175 = (w2136 & ~w2152) | (w2136 & w64520) | (~w2152 & w64520);
assign w2176 = w2146 & w2153;
assign w2177 = ~w2122 & w2147;
assign w2178 = ~w2176 & ~w2177;
assign w2179 = w2175 & ~w2178;
assign w2180 = w2162 & w2164;
assign w2181 = (w2171 & w2161) | (w2171 & w64521) | (w2161 & w64521);
assign w2182 = w2116 & w2122;
assign w2183 = w2147 & w2182;
assign w2184 = ~w2180 & ~w2183;
assign w2185 = ~w2179 & w2184;
assign w2186 = ~w2181 & w2185;
assign w2187 = ~w2174 & w2186;
assign w2188 = ~pi0169 & ~w2187;
assign w2189 = pi0169 & w2187;
assign w2190 = ~w2188 & ~w2189;
assign w2191 = ~w1849 & w1895;
assign w2192 = w1830 & ~w2191;
assign w2193 = ~w2096 & ~w2192;
assign w2194 = (w1849 & ~w1858) | (w1849 & w64507) | (~w1858 & w64507);
assign w2195 = ~w1836 & ~w1875;
assign w2196 = ~w2098 & ~w2195;
assign w2197 = w2194 & ~w2196;
assign w2198 = ~w2193 & ~w2197;
assign w2199 = ~w1861 & ~w1873;
assign w2200 = w1850 & w1878;
assign w2201 = w1861 & w1870;
assign w2202 = ~w2200 & ~w2201;
assign w2203 = ~w1860 & w2202;
assign w2204 = ~w2199 & w2203;
assign w2205 = w1868 & ~w2091;
assign w2206 = ~w2204 & w2205;
assign w2207 = ~w1871 & w2194;
assign w2208 = w1836 & w1875;
assign w2209 = ~w1849 & ~w1893;
assign w2210 = ~w2208 & w2209;
assign w2211 = ~w2207 & ~w2210;
assign w2212 = ~w1868 & w2203;
assign w2213 = ~w2211 & w2212;
assign w2214 = ~w2206 & ~w2213;
assign w2215 = ~w2198 & ~w2214;
assign w2216 = ~pi0165 & w2215;
assign w2217 = pi0165 & ~w2215;
assign w2218 = ~w2216 & ~w2217;
assign w2219 = w2010 & ~w2063;
assign w2220 = w2038 & w2050;
assign w2221 = ~w2023 & w2030;
assign w2222 = w1997 & ~w2019;
assign w2223 = w1984 & w2012;
assign w2224 = (w2048 & ~w2012) | (w2048 & w64522) | (~w2012 & w64522);
assign w2225 = w2003 & w2025;
assign w2226 = ~w2220 & ~w2221;
assign w2227 = w2224 & w2226;
assign w2228 = ~w2225 & w2227;
assign w2229 = ~w2222 & w2228;
assign w2230 = ~w2013 & w2024;
assign w2231 = ~w1990 & ~w2020;
assign w2232 = ~w2033 & w2231;
assign w2233 = w1984 & ~w2032;
assign w2234 = w2014 & w2233;
assign w2235 = ~w2048 & ~w2230;
assign w2236 = ~w2232 & w2235;
assign w2237 = ~w2234 & w2236;
assign w2238 = ~w2229 & ~w2237;
assign w2239 = ~w2219 & ~w2238;
assign w2240 = ~pi0173 & w2239;
assign w2241 = pi0173 & ~w2239;
assign w2242 = ~w2240 & ~w2241;
assign w2243 = ~w1685 & w1816;
assign w2244 = ~w1688 & w2243;
assign w2245 = (~w1816 & w1665) | (~w1816 & w64523) | (w1665 & w64523);
assign w2246 = (~w2244 & ~w1680) | (~w2244 & w64524) | (~w1680 & w64524);
assign w2247 = ~w1640 & ~w2246;
assign w2248 = ~w1634 & w1685;
assign w2249 = (w1640 & ~w1688) | (w1640 & w64525) | (~w1688 & w64525);
assign w2250 = ~w2248 & w2249;
assign w2251 = ~w1695 & ~w2250;
assign w2252 = w1794 & w1795;
assign w2253 = ~w2244 & ~w2252;
assign w2254 = ~w1812 & w2253;
assign w2255 = (w1679 & ~w2254) | (w1679 & w64526) | (~w2254 & w64526);
assign w2256 = ~w1810 & ~w1818;
assign w2257 = ~w1679 & w2254;
assign w2258 = ~w2256 & w2257;
assign w2259 = ~w2247 & ~w2255;
assign w2260 = ~w2258 & w2259;
assign w2261 = ~pi0192 & ~w2260;
assign w2262 = pi0192 & w2260;
assign w2263 = ~w2261 & ~w2262;
assign w2264 = ~w1836 & w2201;
assign w2265 = w1843 & ~w2084;
assign w2266 = w1837 & ~w2265;
assign w2267 = ~w2080 & ~w2208;
assign w2268 = w1849 & ~w2267;
assign w2269 = (w2195 & w2267) | (w2195 & w64527) | (w2267 & w64527);
assign w2270 = ~w2211 & w2269;
assign w2271 = (w1868 & ~w2196) | (w1868 & w64528) | (~w2196 & w64528);
assign w2272 = ~w2266 & w2271;
assign w2273 = ~w2270 & w2272;
assign w2274 = w1830 & w1894;
assign w2275 = ~w1849 & w2196;
assign w2276 = ~w1868 & ~w2274;
assign w2277 = ~w2268 & w2276;
assign w2278 = ~w2275 & w2277;
assign w2279 = ~w2273 & ~w2278;
assign w2280 = ~w2095 & ~w2264;
assign w2281 = ~w2279 & w64529;
assign w2282 = (pi0175 & w2279) | (pi0175 & w64530) | (w2279 & w64530);
assign w2283 = ~w2281 & ~w2282;
assign w2284 = w2123 & w2146;
assign w2285 = ~w2136 & w2284;
assign w2286 = w2153 & w2155;
assign w2287 = ~w2130 & ~w2286;
assign w2288 = w2129 & w2136;
assign w2289 = w2182 & ~w2288;
assign w2290 = w2148 & w2289;
assign w2291 = w2136 & ~w2290;
assign w2292 = ~w2287 & w2291;
assign w2293 = w2129 & w2152;
assign w2294 = ~w2129 & ~w2182;
assign w2295 = w2153 & w2294;
assign w2296 = ~w2293 & ~w2295;
assign w2297 = ~w2295 & w64531;
assign w2298 = ~w2136 & ~w2144;
assign w2299 = w2122 & w2298;
assign w2300 = ~w2292 & w64532;
assign w2301 = w2171 & ~w2300;
assign w2302 = w2129 & w2182;
assign w2303 = w2157 & ~w2302;
assign w2304 = w2137 & ~w2177;
assign w2305 = ~w2303 & ~w2304;
assign w2306 = ~w2136 & w2293;
assign w2307 = ~w2159 & ~w2176;
assign w2308 = ~w2306 & w2307;
assign w2309 = ~w2305 & w2308;
assign w2310 = ~w2171 & ~w2309;
assign w2311 = w2288 & w2297;
assign w2312 = (~w2285 & ~w2303) | (~w2285 & w64533) | (~w2303 & w64533);
assign w2313 = ~w2311 & w2312;
assign w2314 = ~w2310 & w2313;
assign w2315 = (pi0170 & ~w2314) | (pi0170 & w64534) | (~w2314 & w64534);
assign w2316 = w2314 & w64535;
assign w2317 = ~w2315 & ~w2316;
assign w2318 = ~pi3050 & pi9040;
assign w2319 = ~pi3123 & ~pi9040;
assign w2320 = ~w2318 & ~w2319;
assign w2321 = pi0148 & ~w2320;
assign w2322 = ~pi0148 & w2320;
assign w2323 = ~w2321 & ~w2322;
assign w2324 = ~pi3036 & pi9040;
assign w2325 = ~pi3034 & ~pi9040;
assign w2326 = ~w2324 & ~w2325;
assign w2327 = pi0140 & ~w2326;
assign w2328 = ~pi0140 & w2326;
assign w2329 = ~w2327 & ~w2328;
assign w2330 = ~w2323 & ~w2329;
assign w2331 = ~pi3020 & pi9040;
assign w2332 = ~pi3025 & ~pi9040;
assign w2333 = ~w2331 & ~w2332;
assign w2334 = pi0134 & ~w2333;
assign w2335 = ~pi0134 & w2333;
assign w2336 = ~w2334 & ~w2335;
assign w2337 = w2330 & w2336;
assign w2338 = ~w2323 & ~w2336;
assign w2339 = w2329 & w2338;
assign w2340 = ~w2337 & ~w2339;
assign w2341 = ~pi3049 & pi9040;
assign w2342 = ~pi3037 & ~pi9040;
assign w2343 = ~w2341 & ~w2342;
assign w2344 = pi0152 & ~w2343;
assign w2345 = ~pi0152 & w2343;
assign w2346 = ~w2344 & ~w2345;
assign w2347 = ~w2323 & ~w2346;
assign w2348 = ~w2336 & ~w2346;
assign w2349 = w2336 & w2346;
assign w2350 = ~w2348 & ~w2349;
assign w2351 = ~pi3024 & pi9040;
assign w2352 = ~pi3021 & ~pi9040;
assign w2353 = ~w2351 & ~w2352;
assign w2354 = pi0106 & ~w2353;
assign w2355 = ~pi0106 & w2353;
assign w2356 = ~w2354 & ~w2355;
assign w2357 = (w2356 & ~w2350) | (w2356 & w64536) | (~w2350 & w64536);
assign w2358 = w2340 & w2357;
assign w2359 = ~w2323 & w2329;
assign w2360 = w2323 & ~w2329;
assign w2361 = ~w2359 & ~w2360;
assign w2362 = ~w2348 & ~w2361;
assign w2363 = w2348 & w2361;
assign w2364 = (~w2356 & ~w2361) | (~w2356 & w64537) | (~w2361 & w64537);
assign w2365 = ~w2360 & ~w2364;
assign w2366 = ~w2362 & ~w2365;
assign w2367 = ~w2358 & ~w2366;
assign w2368 = ~pi3096 & pi9040;
assign w2369 = ~pi3050 & ~pi9040;
assign w2370 = ~w2368 & ~w2369;
assign w2371 = pi0122 & ~w2370;
assign w2372 = ~pi0122 & w2370;
assign w2373 = ~w2371 & ~w2372;
assign w2374 = ~w2367 & w2373;
assign w2375 = w2323 & w2336;
assign w2376 = ~w2329 & w2346;
assign w2377 = ~w2375 & ~w2376;
assign w2378 = w2356 & w2377;
assign w2379 = w2323 & ~w2336;
assign w2380 = ~w2329 & ~w2346;
assign w2381 = w2379 & w2380;
assign w2382 = w2346 & w2356;
assign w2383 = w2338 & w2382;
assign w2384 = ~w2381 & ~w2383;
assign w2385 = w2378 & ~w2384;
assign w2386 = ~w2347 & w2377;
assign w2387 = ~w2356 & ~w2386;
assign w2388 = ~w2329 & ~w2356;
assign w2389 = w2361 & w64538;
assign w2390 = w2387 & w2389;
assign w2391 = w2340 & w63529;
assign w2392 = w2364 & ~w2391;
assign w2393 = w2356 & w2379;
assign w2394 = ~w2373 & ~w2393;
assign w2395 = ~w2358 & w2394;
assign w2396 = ~w2392 & w2395;
assign w2397 = ~w2385 & ~w2390;
assign w2398 = ~w2396 & w2397;
assign w2399 = ~w2374 & w2398;
assign w2400 = pi0186 & ~w2399;
assign w2401 = ~pi0186 & w2399;
assign w2402 = ~w2400 & ~w2401;
assign w2403 = ~w2013 & ~w2064;
assign w2404 = ~w2013 & w64539;
assign w2405 = (w2010 & w2032) | (w2010 & w64540) | (w2032 & w64540);
assign w2406 = ~w2033 & ~w2405;
assign w2407 = w2034 & ~w2406;
assign w2408 = w2017 & w2064;
assign w2409 = ~w2404 & ~w2408;
assign w2410 = ~w2407 & w2409;
assign w2411 = w2048 & ~w2410;
assign w2412 = ~w1990 & w2403;
assign w2413 = ~w2023 & w2406;
assign w2414 = ~w2412 & ~w2413;
assign w2415 = ~w2065 & w2224;
assign w2416 = ~w2414 & ~w2415;
assign w2417 = w1990 & ~w2048;
assign w2418 = w2013 & w2417;
assign w2419 = ~w2408 & w2418;
assign w2420 = ~w2411 & ~w2419;
assign w2421 = ~w2416 & w2420;
assign w2422 = pi0189 & ~w2421;
assign w2423 = ~pi0189 & w2421;
assign w2424 = ~w2422 & ~w2423;
assign w2425 = ~w2136 & ~w2297;
assign w2426 = w2144 & w2295;
assign w2427 = w2291 & ~w2426;
assign w2428 = ~w2425 & ~w2427;
assign w2429 = w2123 & ~w2148;
assign w2430 = ~w2290 & ~w2429;
assign w2431 = w2296 & w2430;
assign w2432 = ~w2136 & ~w2431;
assign w2433 = ~w2147 & ~w2151;
assign w2434 = w2122 & w2433;
assign w2435 = w2175 & ~w2434;
assign w2436 = (~w2171 & ~w2435) | (~w2171 & w64541) | (~w2435 & w64541);
assign w2437 = ~w2432 & w2436;
assign w2438 = (w2298 & w2295) | (w2298 & w64542) | (w2295 & w64542);
assign w2439 = ~w2294 & w2435;
assign w2440 = w2430 & ~w2438;
assign w2441 = ~w2439 & w2440;
assign w2442 = w2171 & ~w2441;
assign w2443 = ~w2428 & ~w2437;
assign w2444 = (pi0178 & ~w2443) | (pi0178 & w64543) | (~w2443 & w64543);
assign w2445 = w2443 & w64544;
assign w2446 = ~w2444 & ~w2445;
assign w2447 = ~w2013 & w2221;
assign w2448 = w2048 & ~w2447;
assign w2449 = w2042 & w2448;
assign w2450 = ~w1984 & w2003;
assign w2451 = ~w2029 & ~w2450;
assign w2452 = ~w2057 & w2451;
assign w2453 = ~w2026 & ~w2048;
assign w2454 = ~w2065 & ~w2223;
assign w2455 = w2453 & w2454;
assign w2456 = ~w2452 & w2455;
assign w2457 = ~w2449 & ~w2456;
assign w2458 = w1991 & w2053;
assign w2459 = (~w2058 & ~w2228) | (~w2058 & w64545) | (~w2228 & w64545);
assign w2460 = w2015 & ~w2459;
assign w2461 = w2028 & ~w2458;
assign w2462 = ~w2457 & w2461;
assign w2463 = ~w2460 & w2462;
assign w2464 = pi0194 & ~w2463;
assign w2465 = ~pi0194 & w2463;
assign w2466 = ~w2464 & ~w2465;
assign w2467 = w2337 & w2346;
assign w2468 = w2356 & ~w2380;
assign w2469 = (w2468 & w2391) | (w2468 & w64546) | (w2391 & w64546);
assign w2470 = ~w2467 & ~w2469;
assign w2471 = w2373 & ~w2470;
assign w2472 = w2350 & w2361;
assign w2473 = w2336 & w2376;
assign w2474 = w2376 & w2375;
assign w2475 = ~w2472 & ~w2474;
assign w2476 = ~w2356 & w2359;
assign w2477 = ~w2350 & w2476;
assign w2478 = w2384 & ~w2477;
assign w2479 = w2475 & w2478;
assign w2480 = w2329 & ~w2346;
assign w2481 = w2336 & w2480;
assign w2482 = w2330 & w2348;
assign w2483 = ~w2481 & ~w2482;
assign w2484 = w2356 & ~w2483;
assign w2485 = (~w2380 & w2391) | (~w2380 & w64547) | (w2391 & w64547);
assign w2486 = ~w2356 & w2373;
assign w2487 = ~w2330 & w2486;
assign w2488 = ~w2485 & w2487;
assign w2489 = (~w2484 & w2479) | (~w2484 & w64548) | (w2479 & w64548);
assign w2490 = ~w2488 & w2489;
assign w2491 = ~w2471 & w2490;
assign w2492 = pi0199 & ~w2491;
assign w2493 = ~pi0199 & w2491;
assign w2494 = ~w2492 & ~w2493;
assign w2495 = ~w2346 & ~w2356;
assign w2496 = w2375 & w2495;
assign w2497 = w2357 & ~w2475;
assign w2498 = ~w2338 & ~w2375;
assign w2499 = w2388 & w2498;
assign w2500 = ~w2346 & ~w2361;
assign w2501 = ~w2389 & ~w2500;
assign w2502 = ~w2336 & ~w2501;
assign w2503 = w2349 & w2359;
assign w2504 = w2373 & ~w2503;
assign w2505 = ~w2499 & w2504;
assign w2506 = ~w2502 & w2505;
assign w2507 = (~w2347 & ~w2361) | (~w2347 & w63530) | (~w2361 & w63530);
assign w2508 = (~w2468 & w2507) | (~w2468 & w64549) | (w2507 & w64549);
assign w2509 = w2356 & ~w2507;
assign w2510 = ~w2508 & ~w2509;
assign w2511 = ~w2373 & ~w2482;
assign w2512 = ~w2510 & w2511;
assign w2513 = ~w2506 & ~w2512;
assign w2514 = ~w2496 & ~w2497;
assign w2515 = ~w2513 & w2514;
assign w2516 = pi0183 & ~w2515;
assign w2517 = ~pi0183 & w2515;
assign w2518 = ~w2516 & ~w2517;
assign w2519 = (w2373 & ~w2340) | (w2373 & w64550) | (~w2340 & w64550);
assign w2520 = w2375 & w2480;
assign w2521 = ~w2519 & ~w2520;
assign w2522 = w2356 & ~w2521;
assign w2523 = ~w2373 & ~w2388;
assign w2524 = ~w2473 & ~w2503;
assign w2525 = ~w2523 & ~w2524;
assign w2526 = ~w2379 & w2486;
assign w2527 = ~w2377 & w2526;
assign w2528 = ~w2323 & w2481;
assign w2529 = ~w2378 & ~w2473;
assign w2530 = ~w2387 & w2529;
assign w2531 = ~w2363 & ~w2528;
assign w2532 = ~w2530 & w2531;
assign w2533 = ~w2373 & ~w2532;
assign w2534 = ~w2525 & ~w2527;
assign w2535 = ~w2522 & w2534;
assign w2536 = ~w2533 & w2535;
assign w2537 = pi0187 & ~w2536;
assign w2538 = ~pi0187 & w2536;
assign w2539 = ~w2537 & ~w2538;
assign w2540 = w1671 & w1687;
assign w2541 = ~w1688 & ~w2252;
assign w2542 = w2250 & ~w2541;
assign w2543 = w1648 & ~w1656;
assign w2544 = w2243 & ~w2543;
assign w2545 = ~w1792 & ~w1795;
assign w2546 = w1664 & w2545;
assign w2547 = w1703 & ~w2248;
assign w2548 = ~w2544 & ~w2546;
assign w2549 = w2547 & w2548;
assign w2550 = w1640 & w1802;
assign w2551 = ~w1688 & w2543;
assign w2552 = w1679 & ~w1701;
assign w2553 = ~w2551 & w2552;
assign w2554 = ~w2550 & w2553;
assign w2555 = ~w2549 & ~w2554;
assign w2556 = ~w2540 & ~w2542;
assign w2557 = ~w2555 & w2556;
assign w2558 = pi0210 & ~w2557;
assign w2559 = ~pi0210 & w2557;
assign w2560 = ~w2558 & ~w2559;
assign w2561 = ~w2137 & ~w2298;
assign w2562 = ~w2286 & ~w2561;
assign w2563 = ~w2157 & ~w2562;
assign w2564 = w2137 & ~w2433;
assign w2565 = w2136 & ~w2177;
assign w2566 = ~w2289 & w2565;
assign w2567 = ~w2564 & ~w2566;
assign w2568 = w2172 & ~w2567;
assign w2569 = w2116 & ~w2129;
assign w2570 = ~w2147 & ~w2569;
assign w2571 = w2566 & ~w2570;
assign w2572 = w2171 & ~w2183;
assign w2573 = ~w2284 & w2572;
assign w2574 = ~w2306 & w2573;
assign w2575 = ~w2571 & w2574;
assign w2576 = ~w2568 & ~w2575;
assign w2577 = ~w2311 & ~w2563;
assign w2578 = ~w2576 & w2577;
assign w2579 = pi0188 & w2578;
assign w2580 = ~pi0188 & ~w2578;
assign w2581 = ~w2579 & ~w2580;
assign w2582 = ~pi3115 & pi9040;
assign w2583 = ~pi3153 & ~pi9040;
assign w2584 = ~w2582 & ~w2583;
assign w2585 = pi0211 & ~w2584;
assign w2586 = ~pi0211 & w2584;
assign w2587 = ~w2585 & ~w2586;
assign w2588 = ~pi3172 & pi9040;
assign w2589 = ~pi3228 & ~pi9040;
assign w2590 = ~w2588 & ~w2589;
assign w2591 = pi0201 & ~w2590;
assign w2592 = ~pi0201 & w2590;
assign w2593 = ~w2591 & ~w2592;
assign w2594 = ~pi3116 & pi9040;
assign w2595 = ~pi3172 & ~pi9040;
assign w2596 = ~w2594 & ~w2595;
assign w2597 = pi0177 & ~w2596;
assign w2598 = ~pi0177 & w2596;
assign w2599 = ~w2597 & ~w2598;
assign w2600 = w2593 & w2599;
assign w2601 = ~w2593 & ~w2599;
assign w2602 = ~pi3188 & pi9040;
assign w2603 = ~pi3110 & ~pi9040;
assign w2604 = ~w2602 & ~w2603;
assign w2605 = pi0209 & ~w2604;
assign w2606 = ~pi0209 & w2604;
assign w2607 = ~w2605 & ~w2606;
assign w2608 = ~pi3104 & pi9040;
assign w2609 = ~pi3115 & ~pi9040;
assign w2610 = ~w2608 & ~w2609;
assign w2611 = pi0216 & ~w2610;
assign w2612 = ~pi0216 & w2610;
assign w2613 = ~w2611 & ~w2612;
assign w2614 = ~w2607 & w2613;
assign w2615 = ~w2600 & w2614;
assign w2616 = ~w2601 & w2615;
assign w2617 = ~pi3089 & pi9040;
assign w2618 = ~pi3169 & ~pi9040;
assign w2619 = ~w2617 & ~w2618;
assign w2620 = pi0196 & ~w2619;
assign w2621 = ~pi0196 & w2619;
assign w2622 = ~w2620 & ~w2621;
assign w2623 = ~w2599 & ~w2622;
assign w2624 = ~w2593 & ~w2622;
assign w2625 = ~w2613 & w2622;
assign w2626 = w2613 & ~w2622;
assign w2627 = ~w2625 & ~w2626;
assign w2628 = (~w2624 & w2627) | (~w2624 & w63531) | (w2627 & w63531);
assign w2629 = w2599 & w2627;
assign w2630 = ~w2593 & w2613;
assign w2631 = w2623 & ~w2630;
assign w2632 = ~w2629 & ~w2631;
assign w2633 = ~w2628 & w2632;
assign w2634 = w2632 & w63532;
assign w2635 = w2593 & ~w2613;
assign w2636 = ~w2601 & ~w2635;
assign w2637 = w2607 & ~w2636;
assign w2638 = w2593 & ~w2599;
assign w2639 = ~w2636 & w64551;
assign w2640 = w2600 & w2625;
assign w2641 = w2599 & ~w2607;
assign w2642 = w2624 & w2641;
assign w2643 = ~w2640 & ~w2642;
assign w2644 = ~w2616 & w2643;
assign w2645 = ~w2639 & w2644;
assign w2646 = ~w2634 & w2645;
assign w2647 = ~w2587 & ~w2646;
assign w2648 = w2623 & w2635;
assign w2649 = w2601 & w2625;
assign w2650 = ~w2648 & ~w2649;
assign w2651 = w2643 & w2650;
assign w2652 = w2633 & ~w2651;
assign w2653 = (~w2607 & ~w2627) | (~w2607 & w64552) | (~w2627 & w64552);
assign w2654 = w2600 & w2622;
assign w2655 = ~w2653 & ~w2654;
assign w2656 = w2627 & ~w2655;
assign w2657 = (~w2628 & w2652) | (~w2628 & w64553) | (w2652 & w64553);
assign w2658 = ~w2599 & w2626;
assign w2659 = ~w2593 & w2658;
assign w2660 = ~w2654 & ~w2659;
assign w2661 = w2607 & ~w2660;
assign w2662 = w2599 & w2622;
assign w2663 = ~w2599 & w2613;
assign w2664 = ~w2662 & ~w2663;
assign w2665 = ~w2593 & ~w2664;
assign w2666 = (w2622 & ~w2627) | (w2622 & w63533) | (~w2627 & w63533);
assign w2667 = w2665 & w2666;
assign w2668 = (~w2607 & ~w2664) | (~w2607 & w2692) | (~w2664 & w2692);
assign w2669 = ~w2667 & w2668;
assign w2670 = ~w2627 & w64554;
assign w2671 = w2587 & ~w2637;
assign w2672 = ~w2670 & w2671;
assign w2673 = ~w2669 & w2672;
assign w2674 = ~w2661 & ~w2673;
assign w2675 = ~w2647 & w2674;
assign w2676 = (pi0233 & ~w2675) | (pi0233 & w64555) | (~w2675 & w64555);
assign w2677 = w2675 & w64556;
assign w2678 = ~w2676 & ~w2677;
assign w2679 = w2600 & w2626;
assign w2680 = ~w2631 & w2663;
assign w2681 = w2607 & ~w2679;
assign w2682 = ~w2680 & w2681;
assign w2683 = ~w2607 & ~w2631;
assign w2684 = ~w2654 & w2683;
assign w2685 = ~w2682 & ~w2684;
assign w2686 = (w2587 & w2685) | (w2587 & w64557) | (w2685 & w64557);
assign w2687 = ~w2665 & ~w2679;
assign w2688 = ~w2607 & ~w2687;
assign w2689 = w2625 & w2638;
assign w2690 = ~w2688 & ~w2689;
assign w2691 = ~w2587 & ~w2690;
assign w2692 = ~w2593 & ~w2607;
assign w2693 = w2622 & ~w2692;
assign w2694 = w2630 & w2693;
assign w2695 = w2599 & ~w2613;
assign w2696 = w2624 & w2695;
assign w2697 = ~w2587 & w2607;
assign w2698 = ~w2648 & w2697;
assign w2699 = ~w2632 & w2698;
assign w2700 = ~w2694 & ~w2696;
assign w2701 = ~w2699 & w2700;
assign w2702 = ~w2686 & w2701;
assign w2703 = ~w2691 & w2702;
assign w2704 = pi0234 & ~w2703;
assign w2705 = ~pi0234 & w2703;
assign w2706 = ~w2704 & ~w2705;
assign w2707 = w2636 & w2693;
assign w2708 = w2599 & ~w2630;
assign w2709 = w2707 & ~w2708;
assign w2710 = ~w2613 & w2641;
assign w2711 = w2650 & ~w2710;
assign w2712 = ~w2709 & w2711;
assign w2713 = ~w2633 & w2712;
assign w2714 = (~w2587 & w2652) | (~w2587 & w64558) | (w2652 & w64558);
assign w2715 = ~w2658 & ~w2708;
assign w2716 = w2662 & w2692;
assign w2717 = ~w2697 & ~w2716;
assign w2718 = ~w2715 & ~w2717;
assign w2719 = (~w2718 & w2713) | (~w2718 & w64559) | (w2713 & w64559);
assign w2720 = ~w2714 & w2719;
assign w2721 = ~pi0241 & w2720;
assign w2722 = pi0241 & ~w2720;
assign w2723 = ~w2721 & ~w2722;
assign w2724 = ~pi3088 & pi9040;
assign w2725 = ~pi3108 & ~pi9040;
assign w2726 = ~w2724 & ~w2725;
assign w2727 = pi0184 & ~w2726;
assign w2728 = ~pi0184 & w2726;
assign w2729 = ~w2727 & ~w2728;
assign w2730 = ~pi3228 & pi9040;
assign w2731 = ~pi3077 & ~pi9040;
assign w2732 = ~w2730 & ~w2731;
assign w2733 = pi0211 & ~w2732;
assign w2734 = ~pi0211 & w2732;
assign w2735 = ~w2733 & ~w2734;
assign w2736 = ~w2729 & ~w2735;
assign w2737 = w2729 & w2735;
assign w2738 = ~w2736 & ~w2737;
assign w2739 = ~pi3160 & pi9040;
assign w2740 = ~pi3113 & ~pi9040;
assign w2741 = ~w2739 & ~w2740;
assign w2742 = pi0196 & ~w2741;
assign w2743 = ~pi0196 & w2741;
assign w2744 = ~w2742 & ~w2743;
assign w2745 = ~w2738 & w2744;
assign w2746 = ~pi3078 & pi9040;
assign w2747 = ~pi3160 & ~pi9040;
assign w2748 = ~w2746 & ~w2747;
assign w2749 = pi0218 & ~w2748;
assign w2750 = ~pi0218 & w2748;
assign w2751 = ~w2749 & ~w2750;
assign w2752 = ~w2745 & ~w2751;
assign w2753 = ~pi3137 & pi9040;
assign w2754 = ~pi3180 & ~pi9040;
assign w2755 = ~w2753 & ~w2754;
assign w2756 = pi0182 & ~w2755;
assign w2757 = ~pi0182 & w2755;
assign w2758 = ~w2756 & ~w2757;
assign w2759 = ~w2735 & ~w2758;
assign w2760 = w2729 & ~w2744;
assign w2761 = w2759 & w2760;
assign w2762 = ~w2744 & ~w2758;
assign w2763 = w2729 & w2744;
assign w2764 = w2759 & w2763;
assign w2765 = ~w2762 & ~w2764;
assign w2766 = ~w2761 & ~w2765;
assign w2767 = ~w2735 & w2758;
assign w2768 = w2760 & w2767;
assign w2769 = w2751 & ~w2768;
assign w2770 = ~w2766 & w2769;
assign w2771 = ~w2752 & ~w2770;
assign w2772 = w2744 & ~w2758;
assign w2773 = ~w2761 & ~w2772;
assign w2774 = w2735 & w2758;
assign w2775 = w2760 & w2774;
assign w2776 = ~w2735 & w2772;
assign w2777 = ~w2775 & ~w2776;
assign w2778 = ~w2751 & w2777;
assign w2779 = ~w2773 & w2778;
assign w2780 = ~w2744 & w2751;
assign w2781 = w2758 & ~w2780;
assign w2782 = ~w2738 & w2781;
assign w2783 = ~w2751 & w2758;
assign w2784 = ~w2729 & ~w2744;
assign w2785 = w2735 & w2784;
assign w2786 = ~w2783 & w2785;
assign w2787 = ~pi3074 & pi9040;
assign w2788 = ~pi3084 & ~pi9040;
assign w2789 = ~w2787 & ~w2788;
assign w2790 = pi0207 & ~w2789;
assign w2791 = ~pi0207 & w2789;
assign w2792 = ~w2790 & ~w2791;
assign w2793 = ~w2782 & ~w2792;
assign w2794 = ~w2786 & w2793;
assign w2795 = ~w2779 & w2794;
assign w2796 = ~w2759 & ~w2774;
assign w2797 = w2744 & w2796;
assign w2798 = ~w2785 & ~w2797;
assign w2799 = w2783 & ~w2798;
assign w2800 = w2736 & w2762;
assign w2801 = w2735 & w2751;
assign w2802 = w2744 & w2758;
assign w2803 = ~w2729 & w2802;
assign w2804 = ~w2760 & ~w2803;
assign w2805 = w2801 & ~w2804;
assign w2806 = ~w2768 & w2792;
assign w2807 = ~w2800 & w2806;
assign w2808 = ~w2805 & w2807;
assign w2809 = ~w2799 & w2808;
assign w2810 = ~w2795 & ~w2809;
assign w2811 = ~w2771 & ~w2810;
assign w2812 = ~pi0225 & w2811;
assign w2813 = pi0225 & ~w2811;
assign w2814 = ~w2812 & ~w2813;
assign w2815 = ~w2601 & ~w2626;
assign w2816 = ~w2623 & ~w2815;
assign w2817 = ~w2640 & ~w2816;
assign w2818 = w2697 & ~w2817;
assign w2819 = w2587 & ~w2815;
assign w2820 = ~w2623 & ~w2819;
assign w2821 = w2692 & ~w2820;
assign w2822 = w2593 & ~w2682;
assign w2823 = ~w2648 & ~w2822;
assign w2824 = ~w2653 & ~w2823;
assign w2825 = w2587 & ~w2659;
assign w2826 = ~w2707 & w2825;
assign w2827 = ~w2658 & ~w2689;
assign w2828 = ~w2607 & ~w2827;
assign w2829 = ~w2587 & ~w2696;
assign w2830 = ~w2716 & w2829;
assign w2831 = ~w2828 & w2830;
assign w2832 = ~w2826 & ~w2831;
assign w2833 = ~w2818 & ~w2821;
assign w2834 = ~w2832 & w2833;
assign w2835 = ~w2824 & w2834;
assign w2836 = ~pi0236 & ~w2835;
assign w2837 = pi0236 & w2835;
assign w2838 = ~w2836 & ~w2837;
assign w2839 = ~pi3069 & pi9040;
assign w2840 = ~pi3107 & ~pi9040;
assign w2841 = ~w2839 & ~w2840;
assign w2842 = pi0202 & ~w2841;
assign w2843 = ~pi0202 & w2841;
assign w2844 = ~w2842 & ~w2843;
assign w2845 = ~pi3108 & pi9040;
assign w2846 = ~pi3137 & ~pi9040;
assign w2847 = ~w2845 & ~w2846;
assign w2848 = pi0193 & ~w2847;
assign w2849 = ~pi0193 & w2847;
assign w2850 = ~w2848 & ~w2849;
assign w2851 = ~pi3113 & pi9040;
assign w2852 = ~pi3076 & ~pi9040;
assign w2853 = ~w2851 & ~w2852;
assign w2854 = pi0182 & ~w2853;
assign w2855 = ~pi0182 & w2853;
assign w2856 = ~w2854 & ~w2855;
assign w2857 = ~w2850 & w2856;
assign w2858 = ~pi3070 & pi9040;
assign w2859 = ~pi3080 & ~pi9040;
assign w2860 = ~w2858 & ~w2859;
assign w2861 = pi0212 & ~w2860;
assign w2862 = ~pi0212 & w2860;
assign w2863 = ~w2861 & ~w2862;
assign w2864 = ~pi3180 & pi9040;
assign w2865 = ~pi3088 & ~pi9040;
assign w2866 = ~w2864 & ~w2865;
assign w2867 = pi0207 & ~w2866;
assign w2868 = ~pi0207 & w2866;
assign w2869 = ~w2867 & ~w2868;
assign w2870 = ~w2863 & w2869;
assign w2871 = w2857 & w2870;
assign w2872 = ~w2844 & ~w2871;
assign w2873 = ~w2857 & ~w2870;
assign w2874 = w2856 & ~w2863;
assign w2875 = w2856 & ~w2869;
assign w2876 = ~w2850 & ~w2875;
assign w2877 = ~w2874 & ~w2876;
assign w2878 = ~w2873 & w2877;
assign w2879 = ~w2856 & ~w2869;
assign w2880 = ~w2850 & ~w2863;
assign w2881 = w2850 & w2863;
assign w2882 = ~w2856 & w2881;
assign w2883 = (w2879 & w2882) | (w2879 & w64560) | (w2882 & w64560);
assign w2884 = (w2844 & ~w2877) | (w2844 & w63534) | (~w2877 & w63534);
assign w2885 = (~w2872 & ~w2884) | (~w2872 & w64561) | (~w2884 & w64561);
assign w2886 = ~pi3107 & pi9040;
assign w2887 = ~pi3070 & ~pi9040;
assign w2888 = ~w2886 & ~w2887;
assign w2889 = pi0223 & ~w2888;
assign w2890 = ~pi0223 & w2888;
assign w2891 = ~w2889 & ~w2890;
assign w2892 = w2863 & ~w2869;
assign w2893 = ~w2870 & ~w2892;
assign w2894 = (~w2844 & w2893) | (~w2844 & w63351) | (w2893 & w63351);
assign w2895 = w2844 & ~w2869;
assign w2896 = (w2844 & ~w2880) | (w2844 & w63535) | (~w2880 & w63535);
assign w2897 = ~w2895 & ~w2896;
assign w2898 = ~w2873 & ~w2897;
assign w2899 = w2875 & w2881;
assign w2900 = (~w2899 & ~w2894) | (~w2899 & w63536) | (~w2894 & w63536);
assign w2901 = ~w2898 & w2900;
assign w2902 = w2891 & ~w2901;
assign w2903 = ~w2885 & ~w2902;
assign w2904 = ~w2881 & ~w2893;
assign w2905 = w2897 & w2904;
assign w2906 = w2850 & w2879;
assign w2907 = ~w2850 & ~w2856;
assign w2908 = w2863 & w2907;
assign w2909 = w2907 & w64562;
assign w2910 = ~w2906 & ~w2909;
assign w2911 = w2844 & ~w2910;
assign w2912 = ~w2844 & w2850;
assign w2913 = ~w2875 & w2881;
assign w2914 = ~w2912 & ~w2913;
assign w2915 = w2856 & ~w2914;
assign w2916 = ~w2905 & ~w2915;
assign w2917 = ~w2911 & w2916;
assign w2918 = ~w2891 & ~w2917;
assign w2919 = w2903 & ~w2918;
assign w2920 = ~pi0227 & w2919;
assign w2921 = pi0227 & ~w2919;
assign w2922 = ~w2920 & ~w2921;
assign w2923 = w2736 & w2758;
assign w2924 = (w2744 & w2923) | (w2744 & w64563) | (w2923 & w64563);
assign w2925 = w2737 & ~w2758;
assign w2926 = w2751 & ~w2925;
assign w2927 = w2760 & w2796;
assign w2928 = ~w2926 & w2927;
assign w2929 = ~w2762 & ~w2802;
assign w2930 = ~w2737 & w2929;
assign w2931 = ~w2751 & ~w2930;
assign w2932 = w2784 & ~w2796;
assign w2933 = ~w2931 & w2932;
assign w2934 = ~w2764 & ~w2924;
assign w2935 = ~w2928 & w2934;
assign w2936 = ~w2933 & w2935;
assign w2937 = w2792 & ~w2936;
assign w2938 = w2738 & w2762;
assign w2939 = ~w2931 & ~w2938;
assign w2940 = ~w2738 & ~w2777;
assign w2941 = ~w2763 & ~w2780;
assign w2942 = w2767 & ~w2941;
assign w2943 = ~w2940 & ~w2942;
assign w2944 = w2939 & w2943;
assign w2945 = ~w2792 & ~w2944;
assign w2946 = ~w2937 & ~w2945;
assign w2947 = pi0224 & ~w2946;
assign w2948 = ~pi0224 & w2946;
assign w2949 = ~w2947 & ~w2948;
assign w2950 = ~pi3109 & pi9040;
assign w2951 = ~pi3157 & ~pi9040;
assign w2952 = ~w2950 & ~w2951;
assign w2953 = pi0198 & ~w2952;
assign w2954 = ~pi0198 & w2952;
assign w2955 = ~w2953 & ~w2954;
assign w2956 = ~pi3111 & pi9040;
assign w2957 = ~pi3109 & ~pi9040;
assign w2958 = ~w2956 & ~w2957;
assign w2959 = pi0214 & ~w2958;
assign w2960 = ~pi0214 & w2958;
assign w2961 = ~w2959 & ~w2960;
assign w2962 = ~w2955 & w2961;
assign w2963 = ~pi3163 & pi9040;
assign w2964 = ~pi3085 & ~pi9040;
assign w2965 = ~w2963 & ~w2964;
assign w2966 = pi0180 & ~w2965;
assign w2967 = ~pi0180 & w2965;
assign w2968 = ~w2966 & ~w2967;
assign w2969 = ~pi3083 & pi9040;
assign w2970 = ~pi3118 & ~pi9040;
assign w2971 = ~w2969 & ~w2970;
assign w2972 = pi0219 & ~w2971;
assign w2973 = ~pi0219 & w2971;
assign w2974 = ~w2972 & ~w2973;
assign w2975 = ~w2968 & w2974;
assign w2976 = w2962 & w2975;
assign w2977 = ~pi3085 & pi9040;
assign w2978 = ~pi3081 & ~pi9040;
assign w2979 = ~w2977 & ~w2978;
assign w2980 = pi0205 & ~w2979;
assign w2981 = ~pi0205 & w2979;
assign w2982 = ~w2980 & ~w2981;
assign w2983 = w2962 & w2968;
assign w2984 = ~w2955 & ~w2961;
assign w2985 = ~w2974 & w2984;
assign w2986 = ~w2983 & ~w2985;
assign w2987 = ~pi3075 & pi9040;
assign w2988 = ~pi3091 & ~pi9040;
assign w2989 = ~w2987 & ~w2988;
assign w2990 = pi0220 & ~w2989;
assign w2991 = ~pi0220 & w2989;
assign w2992 = ~w2990 & ~w2991;
assign w2993 = w2986 & ~w2992;
assign w2994 = ~w2955 & ~w2968;
assign w2995 = w2955 & w2968;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = w2968 & ~w2974;
assign w2998 = ~w2961 & ~w2997;
assign w2999 = w2996 & w2998;
assign w3000 = w2992 & ~w2999;
assign w3001 = ~w2993 & ~w3000;
assign w3002 = w2955 & w2961;
assign w3003 = ~w2968 & w3002;
assign w3004 = ~w2992 & ~w3003;
assign w3005 = w2955 & ~w2974;
assign w3006 = ~w3004 & w3005;
assign w3007 = w2968 & w2992;
assign w3008 = w3002 & w3007;
assign w3009 = ~w2976 & w2982;
assign w3010 = ~w3008 & w3009;
assign w3011 = ~w3006 & w3010;
assign w3012 = ~w3001 & w3011;
assign w3013 = w3002 & w2975;
assign w3014 = ~w2982 & ~w3013;
assign w3015 = ~w2986 & w2992;
assign w3016 = ~w2961 & w2974;
assign w3017 = ~w2996 & w3016;
assign w3018 = w3014 & ~w3017;
assign w3019 = ~w3015 & w3018;
assign w3020 = ~w3012 & ~w3019;
assign w3021 = ~w2961 & ~w2974;
assign w3022 = w2996 & ~w3021;
assign w3023 = ~w2982 & ~w2984;
assign w3024 = ~w3022 & w3023;
assign w3025 = ~w2976 & ~w3017;
assign w3026 = ~w3024 & w3025;
assign w3027 = ~w2992 & ~w3026;
assign w3028 = ~w3020 & ~w3027;
assign w3029 = ~pi0231 & w3028;
assign w3030 = pi0231 & ~w3028;
assign w3031 = ~w3029 & ~w3030;
assign w3032 = ~pi3157 & pi9040;
assign w3033 = ~pi3112 & ~pi9040;
assign w3034 = ~w3032 & ~w3033;
assign w3035 = pi0213 & ~w3034;
assign w3036 = ~pi0213 & w3034;
assign w3037 = ~w3035 & ~w3036;
assign w3038 = ~pi3093 & pi9040;
assign w3039 = ~pi3225 & ~pi9040;
assign w3040 = ~w3038 & ~w3039;
assign w3041 = pi0180 & ~w3040;
assign w3042 = ~pi0180 & w3040;
assign w3043 = ~w3041 & ~w3042;
assign w3044 = ~pi3112 & pi9040;
assign w3045 = ~pi3111 & ~pi9040;
assign w3046 = ~w3044 & ~w3045;
assign w3047 = pi0193 & ~w3046;
assign w3048 = ~pi0193 & w3046;
assign w3049 = ~w3047 & ~w3048;
assign w3050 = w3043 & ~w3049;
assign w3051 = ~pi3072 & pi9040;
assign w3052 = ~pi3168 & ~pi9040;
assign w3053 = ~w3051 & ~w3052;
assign w3054 = pi0208 & ~w3053;
assign w3055 = ~pi0208 & w3053;
assign w3056 = ~w3054 & ~w3055;
assign w3057 = ~w3050 & ~w3056;
assign w3058 = ~w3043 & w3049;
assign w3059 = ~w3050 & ~w3058;
assign w3060 = ~pi3081 & pi9040;
assign w3061 = ~pi3073 & ~pi9040;
assign w3062 = ~w3060 & ~w3061;
assign w3063 = pi0223 & ~w3062;
assign w3064 = ~pi0223 & w3062;
assign w3065 = ~w3063 & ~w3064;
assign w3066 = w3049 & w3065;
assign w3067 = ~w3037 & ~w3066;
assign w3068 = w3043 & w3065;
assign w3069 = ~w3056 & w3068;
assign w3070 = ~w3067 & ~w3069;
assign w3071 = w3059 & ~w3070;
assign w3072 = (w3057 & w3070) | (w3057 & w64564) | (w3070 & w64564);
assign w3073 = ~w3043 & ~w3065;
assign w3074 = ~w3068 & ~w3073;
assign w3075 = ~w3059 & w3074;
assign w3076 = w3056 & w3075;
assign w3077 = ~pi3086 & pi9040;
assign w3078 = ~pi3121 & ~pi9040;
assign w3079 = ~w3077 & ~w3078;
assign w3080 = pi0198 & ~w3079;
assign w3081 = ~pi0198 & w3079;
assign w3082 = ~w3080 & ~w3081;
assign w3083 = (~w3065 & w3076) | (~w3065 & w63537) | (w3076 & w63537);
assign w3084 = (~w3037 & w3083) | (~w3037 & w64565) | (w3083 & w64565);
assign w3085 = ~w3049 & ~w3056;
assign w3086 = ~w3065 & ~w3085;
assign w3087 = w3068 & w3085;
assign w3088 = ~w3086 & ~w3087;
assign w3089 = w3037 & ~w3088;
assign w3090 = ~w3088 & w64566;
assign w3091 = ~w3043 & w3090;
assign w3092 = w3037 & w3065;
assign w3093 = w3085 & w3092;
assign w3094 = ~w3037 & w3066;
assign w3095 = w3043 & w3056;
assign w3096 = w3094 & w3095;
assign w3097 = ~w3093 & ~w3096;
assign w3098 = ~w3049 & ~w3065;
assign w3099 = ~w3037 & ~w3098;
assign w3100 = ~w3057 & ~w3099;
assign w3101 = w3049 & w3074;
assign w3102 = w3100 & w3101;
assign w3103 = ~w3049 & ~w3074;
assign w3104 = (w3056 & ~w3074) | (w3056 & w63538) | (~w3074 & w63538);
assign w3105 = ~w3103 & w3104;
assign w3106 = w3071 & w3105;
assign w3107 = ~w3102 & ~w3106;
assign w3108 = w3037 & w3049;
assign w3109 = w3059 & ~w3108;
assign w3110 = ~w3074 & ~w3109;
assign w3111 = ~w3109 & w63539;
assign w3112 = ~w3082 & ~w3111;
assign w3113 = w3107 & w3112;
assign w3114 = ~w3050 & ~w3073;
assign w3115 = w3100 & ~w3114;
assign w3116 = ~w3037 & ~w3065;
assign w3117 = ~w3056 & ~w3066;
assign w3118 = ~w3116 & w3117;
assign w3119 = w3074 & w3118;
assign w3120 = ~w3115 & ~w3119;
assign w3121 = w3082 & ~w3094;
assign w3122 = w3120 & w3121;
assign w3123 = ~w3113 & ~w3122;
assign w3124 = ~w3091 & w3097;
assign w3125 = ~w3084 & w3124;
assign w3126 = (pi0228 & w3123) | (pi0228 & w64567) | (w3123 & w64567);
assign w3127 = ~w3123 & w64568;
assign w3128 = ~w3126 & ~w3127;
assign w3129 = w3108 & ~w3120;
assign w3130 = (~w3037 & w3111) | (~w3037 & w64569) | (w3111 & w64569);
assign w3131 = w3059 & w3092;
assign w3132 = ~w3076 & ~w3131;
assign w3133 = ~w3130 & w3132;
assign w3134 = ~w3082 & ~w3133;
assign w3135 = w3049 & w3095;
assign w3136 = ~w3056 & w3065;
assign w3137 = w3058 & w3136;
assign w3138 = ~w3037 & ~w3136;
assign w3139 = ~w3086 & w3138;
assign w3140 = ~w3135 & ~w3137;
assign w3141 = ~w3139 & w3140;
assign w3142 = ~w3089 & w3141;
assign w3143 = w3082 & ~w3142;
assign w3144 = ~w3129 & ~w3143;
assign w3145 = ~w3134 & w3144;
assign w3146 = ~pi0229 & w3145;
assign w3147 = pi0229 & ~w3145;
assign w3148 = ~w3146 & ~w3147;
assign w3149 = ~pi3087 & pi9040;
assign w3150 = ~pi3075 & ~pi9040;
assign w3151 = ~w3149 & ~w3150;
assign w3152 = pi0221 & ~w3151;
assign w3153 = ~pi0221 & w3151;
assign w3154 = ~w3152 & ~w3153;
assign w3155 = ~pi3122 & pi9040;
assign w3156 = ~pi3079 & ~pi9040;
assign w3157 = ~w3155 & ~w3156;
assign w3158 = pi0203 & ~w3157;
assign w3159 = ~pi0203 & w3157;
assign w3160 = ~w3158 & ~w3159;
assign w3161 = ~pi3073 & pi9040;
assign w3162 = ~pi3163 & ~pi9040;
assign w3163 = ~w3161 & ~w3162;
assign w3164 = pi0217 & ~w3163;
assign w3165 = ~pi0217 & w3163;
assign w3166 = ~w3164 & ~w3165;
assign w3167 = ~w3160 & ~w3166;
assign w3168 = ~pi3071 & pi9040;
assign w3169 = ~pi3082 & ~pi9040;
assign w3170 = ~w3168 & ~w3169;
assign w3171 = pi0204 & ~w3170;
assign w3172 = ~pi0204 & w3170;
assign w3173 = ~w3171 & ~w3172;
assign w3174 = ~pi3184 & pi9040;
assign w3175 = ~pi3087 & ~pi9040;
assign w3176 = ~w3174 & ~w3175;
assign w3177 = pi0215 & ~w3176;
assign w3178 = ~pi0215 & w3176;
assign w3179 = ~w3177 & ~w3178;
assign w3180 = ~w3173 & w3179;
assign w3181 = w3167 & w3180;
assign w3182 = ~w3160 & w3166;
assign w3183 = ~pi3091 & pi9040;
assign w3184 = ~pi3184 & ~pi9040;
assign w3185 = ~w3183 & ~w3184;
assign w3186 = pi0206 & ~w3185;
assign w3187 = ~pi0206 & w3185;
assign w3188 = ~w3186 & ~w3187;
assign w3189 = ~w3173 & w3188;
assign w3190 = w3182 & w3189;
assign w3191 = ~w3173 & ~w3188;
assign w3192 = w3167 & w3191;
assign w3193 = ~w3190 & ~w3192;
assign w3194 = w3166 & w3179;
assign w3195 = w3160 & ~w3188;
assign w3196 = ~w3160 & w3188;
assign w3197 = ~w3195 & ~w3196;
assign w3198 = w3173 & ~w3188;
assign w3199 = w3194 & ~w3198;
assign w3200 = ~w3197 & w3199;
assign w3201 = w3166 & ~w3188;
assign w3202 = ~w3173 & ~w3179;
assign w3203 = w3160 & ~w3201;
assign w3204 = w3202 & w3203;
assign w3205 = ~w3200 & ~w3204;
assign w3206 = w3167 & w3202;
assign w3207 = w3188 & w3206;
assign w3208 = ~w3167 & ~w3180;
assign w3209 = w3160 & w3166;
assign w3210 = ~w3166 & ~w3179;
assign w3211 = w3173 & ~w3210;
assign w3212 = ~w3209 & ~w3211;
assign w3213 = ~w3208 & ~w3212;
assign w3214 = w3166 & w3173;
assign w3215 = w3197 & w3214;
assign w3216 = ~w3167 & ~w3209;
assign w3217 = ~w3179 & ~w3188;
assign w3218 = w3216 & w3217;
assign w3219 = ~w3207 & ~w3215;
assign w3220 = ~w3218 & w3219;
assign w3221 = w3220 & w63540;
assign w3222 = ~w3166 & w3195;
assign w3223 = ~w3194 & ~w3222;
assign w3224 = (w3160 & w3222) | (w3160 & w63541) | (w3222 & w63541);
assign w3225 = (w3173 & w3224) | (w3173 & w64570) | (w3224 & w64570);
assign w3226 = ~w3181 & w3193;
assign w3227 = ~w3225 & w3226;
assign w3228 = (~w3154 & w3221) | (~w3154 & w64571) | (w3221 & w64571);
assign w3229 = ~w3179 & w3198;
assign w3230 = ~w3180 & ~w3229;
assign w3231 = ~w3160 & w3198;
assign w3232 = w3160 & ~w3198;
assign w3233 = ~w3231 & ~w3232;
assign w3234 = w3166 & ~w3189;
assign w3235 = ~w3233 & w3234;
assign w3236 = ~w3230 & w3235;
assign w3237 = (w3154 & ~w3220) | (w3154 & w64572) | (~w3220 & w64572);
assign w3238 = w3179 & ~w3209;
assign w3239 = ~w3173 & w3197;
assign w3240 = w3238 & w3239;
assign w3241 = w3160 & ~w3179;
assign w3242 = ~w3189 & ~w3214;
assign w3243 = w3241 & w3242;
assign w3244 = ~w3240 & ~w3243;
assign w3245 = ~w3233 & w3238;
assign w3246 = w3193 & ~w3206;
assign w3247 = ~w3245 & w3246;
assign w3248 = ~w3244 & ~w3247;
assign w3249 = ~w3236 & ~w3248;
assign w3250 = ~w3237 & w3249;
assign w3251 = (pi0226 & ~w3250) | (pi0226 & w64573) | (~w3250 & w64573);
assign w3252 = w3250 & w64574;
assign w3253 = ~w3251 & ~w3252;
assign w3254 = ~w2984 & ~w3013;
assign w3255 = w2993 & ~w3254;
assign w3256 = ~w2968 & w3021;
assign w3257 = w3021 & w63542;
assign w3258 = ~w2968 & ~w2992;
assign w3259 = w2984 & w3258;
assign w3260 = w2974 & w2992;
assign w3261 = ~w2955 & ~w3260;
assign w3262 = ~w2955 & w2974;
assign w3263 = ~w3258 & ~w3262;
assign w3264 = w2961 & ~w2975;
assign w3265 = ~w3263 & w3264;
assign w3266 = w3261 & w3265;
assign w3267 = w2997 & w3002;
assign w3268 = w2982 & ~w3267;
assign w3269 = w3007 & ~w3262;
assign w3270 = ~w3259 & ~w3269;
assign w3271 = ~w3257 & w3270;
assign w3272 = w3268 & w3271;
assign w3273 = ~w3266 & w3272;
assign w3274 = ~w3255 & w3273;
assign w3275 = ~w2961 & w2968;
assign w3276 = ~w3005 & w3275;
assign w3277 = ~w3267 & ~w3276;
assign w3278 = ~w3257 & w3277;
assign w3279 = ~w2962 & w2992;
assign w3280 = w3277 & w63543;
assign w3281 = (~w2982 & ~w3263) | (~w2982 & w64575) | (~w3263 & w64575);
assign w3282 = ~w3280 & w3281;
assign w3283 = (~w3014 & w3280) | (~w3014 & w64576) | (w3280 & w64576);
assign w3284 = w2961 & w2994;
assign w3285 = ~w3275 & ~w3284;
assign w3286 = (~w2974 & w3284) | (~w2974 & w64577) | (w3284 & w64577);
assign w3287 = w2986 & w63544;
assign w3288 = w3254 & w3287;
assign w3289 = ~w3265 & ~w3286;
assign w3290 = ~w3288 & w3289;
assign w3291 = ~w3283 & w3290;
assign w3292 = ~w3274 & ~w3291;
assign w3293 = w2961 & w3262;
assign w3294 = w2992 & ~w3293;
assign w3295 = ~w2975 & ~w2997;
assign w3296 = ~w2996 & ~w3295;
assign w3297 = w3294 & w3296;
assign w3298 = ~w3292 & w64578;
assign w3299 = (~pi0235 & w3292) | (~pi0235 & w64579) | (w3292 & w64579);
assign w3300 = ~w3298 & ~w3299;
assign w3301 = ~w3201 & ~w3229;
assign w3302 = w3160 & ~w3301;
assign w3303 = (~w3154 & ~w3247) | (~w3154 & w64580) | (~w3247 & w64580);
assign w3304 = w3182 & ~w3230;
assign w3305 = w3211 & w3222;
assign w3306 = w3173 & w3188;
assign w3307 = ~w3216 & w3306;
assign w3308 = ~w3204 & ~w3305;
assign w3309 = ~w3307 & w3308;
assign w3310 = (w3154 & ~w3309) | (w3154 & w64581) | (~w3309 & w64581);
assign w3311 = ~w3192 & ~w3307;
assign w3312 = ~w3179 & ~w3311;
assign w3313 = ~w3200 & ~w3312;
assign w3314 = ~w3303 & w3313;
assign w3315 = ~w3310 & w3314;
assign w3316 = pi0230 & ~w3315;
assign w3317 = ~pi0230 & w3315;
assign w3318 = ~w3316 & ~w3317;
assign w3319 = ~w3256 & w3294;
assign w3320 = ~w2961 & w2975;
assign w3321 = w3004 & ~w3320;
assign w3322 = ~w3319 & ~w3321;
assign w3323 = w2995 & w3016;
assign w3324 = w3268 & ~w3323;
assign w3325 = w2984 & w2997;
assign w3326 = ~w3265 & ~w3325;
assign w3327 = w3324 & w3326;
assign w3328 = ~w3322 & w3327;
assign w3329 = ~w3282 & ~w3328;
assign w3330 = ~w2976 & w3278;
assign w3331 = ~w2992 & ~w3324;
assign w3332 = ~w3330 & w3331;
assign w3333 = ~w3329 & ~w3332;
assign w3334 = ~pi0248 & w3333;
assign w3335 = pi0248 & ~w3333;
assign w3336 = ~w3334 & ~w3335;
assign w3337 = ~w3074 & w63538;
assign w3338 = ~w3071 & ~w3337;
assign w3339 = ~w3071 & w63545;
assign w3340 = ~w3090 & ~w3339;
assign w3341 = w3107 & w3340;
assign w3342 = w3082 & ~w3341;
assign w3343 = ~w3094 & ~w3135;
assign w3344 = ~w3043 & w3085;
assign w3345 = w3073 & w3108;
assign w3346 = ~w3095 & ~w3345;
assign w3347 = ~w3092 & ~w3116;
assign w3348 = ~w3346 & w3347;
assign w3349 = w3343 & ~w3344;
assign w3350 = ~w3348 & w3349;
assign w3351 = ~w3037 & w3075;
assign w3352 = ~w3345 & ~w3351;
assign w3353 = ~w3056 & ~w3352;
assign w3354 = (w3097 & w3350) | (w3097 & w64582) | (w3350 & w64582);
assign w3355 = ~w3353 & w3354;
assign w3356 = ~w3342 & w64583;
assign w3357 = (pi0238 & w3342) | (pi0238 & w64584) | (w3342 & w64584);
assign w3358 = ~w3356 & ~w3357;
assign w3359 = ~pi3120 & pi9040;
assign w3360 = ~pi3188 & ~pi9040;
assign w3361 = ~w3359 & ~w3360;
assign w3362 = pi0204 & ~w3361;
assign w3363 = ~pi0204 & w3361;
assign w3364 = ~w3362 & ~w3363;
assign w3365 = ~pi3119 & pi9040;
assign w3366 = ~pi3120 & ~pi9040;
assign w3367 = ~w3365 & ~w3366;
assign w3368 = pi0222 & ~w3367;
assign w3369 = ~pi0222 & w3367;
assign w3370 = ~w3368 & ~w3369;
assign w3371 = w3364 & w3370;
assign w3372 = ~pi3084 & pi9040;
assign w3373 = ~pi3089 & ~pi9040;
assign w3374 = ~w3372 & ~w3373;
assign w3375 = pi0216 & ~w3374;
assign w3376 = ~pi0216 & w3374;
assign w3377 = ~w3375 & ~w3376;
assign w3378 = w3364 & w3377;
assign w3379 = ~w3371 & ~w3378;
assign w3380 = ~pi3169 & pi9040;
assign w3381 = ~pi3074 & ~pi9040;
assign w3382 = ~w3380 & ~w3381;
assign w3383 = pi0221 & ~w3382;
assign w3384 = ~pi0221 & w3382;
assign w3385 = ~w3383 & ~w3384;
assign w3386 = ~w3377 & w3385;
assign w3387 = ~w3370 & w3377;
assign w3388 = ~w3386 & ~w3387;
assign w3389 = ~w3379 & ~w3388;
assign w3390 = ~w3370 & ~w3385;
assign w3391 = w3364 & w3390;
assign w3392 = w3377 & ~w3385;
assign w3393 = ~w3364 & ~w3392;
assign w3394 = ~w3392 & w64585;
assign w3395 = ~pi3077 & pi9040;
assign w3396 = ~pi3116 & ~pi9040;
assign w3397 = ~w3395 & ~w3396;
assign w3398 = pi0185 & ~w3397;
assign w3399 = ~pi0185 & w3397;
assign w3400 = ~w3398 & ~w3399;
assign w3401 = ~w3394 & ~w3400;
assign w3402 = ~w3391 & w3401;
assign w3403 = ~w3370 & w3385;
assign w3404 = w3364 & w3385;
assign w3405 = ~w3377 & ~w3404;
assign w3406 = w3403 & w3405;
assign w3407 = (w3400 & ~w3405) | (w3400 & w63546) | (~w3405 & w63546);
assign w3408 = w3377 & w3404;
assign w3409 = w3407 & ~w3408;
assign w3410 = w3371 & ~w3385;
assign w3411 = w3371 & w64586;
assign w3412 = ~w3364 & ~w3385;
assign w3413 = ~w3411 & ~w3412;
assign w3414 = w3409 & w3413;
assign w3415 = (~w3389 & w3414) | (~w3389 & w64587) | (w3414 & w64587);
assign w3416 = ~pi3117 & pi9040;
assign w3417 = ~pi3104 & ~pi9040;
assign w3418 = ~w3416 & ~w3417;
assign w3419 = pi0177 & ~w3418;
assign w3420 = ~pi0177 & w3418;
assign w3421 = ~w3419 & ~w3420;
assign w3422 = ~w3415 & w3421;
assign w3423 = ~w3377 & w3400;
assign w3424 = w3410 & ~w3423;
assign w3425 = ~w3364 & ~w3400;
assign w3426 = ~w3386 & ~w3390;
assign w3427 = w3425 & ~w3426;
assign w3428 = ~w3424 & ~w3427;
assign w3429 = ~w3421 & ~w3428;
assign w3430 = w3387 & w3404;
assign w3431 = w3370 & w3385;
assign w3432 = w3425 & w3431;
assign w3433 = ~w3404 & ~w3412;
assign w3434 = ~w3377 & ~w3433;
assign w3435 = w3370 & w3434;
assign w3436 = w3364 & w3421;
assign w3437 = ~w3370 & ~w3378;
assign w3438 = ~w3436 & w3437;
assign w3439 = ~w3393 & w3438;
assign w3440 = ~w3435 & ~w3439;
assign w3441 = w3400 & ~w3440;
assign w3442 = ~w3430 & ~w3432;
assign w3443 = ~w3429 & w3442;
assign w3444 = ~w3441 & w3443;
assign w3445 = ~w3422 & w3444;
assign w3446 = pi0242 & ~w3445;
assign w3447 = ~pi0242 & w3445;
assign w3448 = ~w3446 & ~w3447;
assign w3449 = ~w3232 & w3234;
assign w3450 = ~w3223 & ~w3449;
assign w3451 = w3173 & ~w3196;
assign w3452 = w3210 & ~w3451;
assign w3453 = ~w3154 & ~w3452;
assign w3454 = ~w3450 & w3453;
assign w3455 = w3241 & w3306;
assign w3456 = ~w3160 & ~w3214;
assign w3457 = ~w3301 & w3456;
assign w3458 = ~w3189 & ~w3196;
assign w3459 = ~w3212 & ~w3458;
assign w3460 = w3154 & ~w3181;
assign w3461 = ~w3455 & w3460;
assign w3462 = ~w3457 & w3461;
assign w3463 = ~w3459 & w3462;
assign w3464 = ~w3454 & ~w3463;
assign w3465 = w3173 & ~w3209;
assign w3466 = ~w3218 & ~w3229;
assign w3467 = ~w3465 & ~w3466;
assign w3468 = w3182 & w3198;
assign w3469 = ~w3310 & w3468;
assign w3470 = ~w3305 & ~w3467;
assign w3471 = ~w3464 & w3470;
assign w3472 = w3471 & w64588;
assign w3473 = (~pi0239 & ~w3471) | (~pi0239 & w64589) | (~w3471 & w64589);
assign w3474 = ~w3472 & ~w3473;
assign w3475 = w2759 & w2780;
assign w3476 = w2763 & w2796;
assign w3477 = ~w3476 & w63547;
assign w3478 = ~w2939 & ~w3477;
assign w3479 = ~w2729 & ~w2796;
assign w3480 = ~w3476 & w64590;
assign w3481 = ~w3479 & w3480;
assign w3482 = ~w2796 & w64591;
assign w3483 = ~w2751 & w3482;
assign w3484 = ~w2761 & ~w3483;
assign w3485 = ~w3481 & w3484;
assign w3486 = ~w2792 & ~w3485;
assign w3487 = (~w2751 & ~w2763) | (~w2751 & w64592) | (~w2763 & w64592);
assign w3488 = ~w2738 & ~w2744;
assign w3489 = ~w2797 & w3487;
assign w3490 = w3480 & ~w3482;
assign w3491 = (w2792 & ~w3489) | (w2792 & w64593) | (~w3489 & w64593);
assign w3492 = ~w3490 & w3491;
assign w3493 = ~w3478 & ~w3492;
assign w3494 = ~w3486 & w3493;
assign w3495 = pi0240 & ~w3494;
assign w3496 = ~pi0240 & w3494;
assign w3497 = ~w3495 & ~w3496;
assign w3498 = ~w2869 & ~w2880;
assign w3499 = w2856 & ~w3498;
assign w3500 = ~w2906 & ~w3499;
assign w3501 = ~w2856 & ~w2863;
assign w3502 = w2850 & w3501;
assign w3503 = w2891 & ~w3502;
assign w3504 = ~w3500 & ~w3503;
assign w3505 = ~w2899 & ~w3504;
assign w3506 = w2844 & ~w3505;
assign w3507 = w2894 & w3500;
assign w3508 = w2882 & ~w2895;
assign w3509 = ~w2893 & w63548;
assign w3510 = w2895 & w2907;
assign w3511 = ~w3508 & ~w3510;
assign w3512 = ~w3509 & w3511;
assign w3513 = w2891 & ~w3512;
assign w3514 = ~w2856 & w2869;
assign w3515 = w2844 & ~w2880;
assign w3516 = ~w2891 & w3514;
assign w3517 = ~w3515 & w3516;
assign w3518 = ~w3507 & ~w3517;
assign w3519 = ~w3513 & w3518;
assign w3520 = ~w3506 & w3519;
assign w3521 = ~pi0247 & w3520;
assign w3522 = pi0247 & ~w3520;
assign w3523 = ~w3521 & ~w3522;
assign w3524 = (~w3154 & ~w3244) | (~w3154 & w64594) | (~w3244 & w64594);
assign w3525 = ~w3190 & ~w3307;
assign w3526 = w3179 & ~w3525;
assign w3527 = ~w3154 & ~w3202;
assign w3528 = ~w3216 & ~w3458;
assign w3529 = ~w3527 & w3528;
assign w3530 = ~w3179 & ~w3449;
assign w3531 = ~w3194 & w3460;
assign w3532 = ~w3530 & w3531;
assign w3533 = ~w3248 & w3532;
assign w3534 = ~w3526 & ~w3529;
assign w3535 = ~w3524 & w3534;
assign w3536 = ~w3533 & w3535;
assign w3537 = pi0237 & w3536;
assign w3538 = ~pi0237 & ~w3536;
assign w3539 = ~w3537 & ~w3538;
assign w3540 = w2895 & w3501;
assign w3541 = ~w2891 & ~w3540;
assign w3542 = ~w2875 & w64595;
assign w3543 = ~w2844 & ~w2850;
assign w3544 = w2893 & ~w3543;
assign w3545 = w2893 & w63549;
assign w3546 = (~w3514 & w3545) | (~w3514 & w64596) | (w3545 & w64596);
assign w3547 = ~w2856 & w2863;
assign w3548 = w3515 & ~w3547;
assign w3549 = ~w3509 & w3548;
assign w3550 = ~w2844 & w2869;
assign w3551 = (w3550 & w2882) | (w3550 & w64597) | (w2882 & w64597);
assign w3552 = ~w3549 & ~w3551;
assign w3553 = (~w3541 & ~w3552) | (~w3541 & w64598) | (~w3552 & w64598);
assign w3554 = w2893 & w2907;
assign w3555 = ~w2875 & ~w2912;
assign w3556 = ~w3544 & ~w3555;
assign w3557 = w2844 & w2869;
assign w3558 = ~w2857 & ~w3547;
assign w3559 = w3557 & ~w3558;
assign w3560 = ~w3554 & ~w3559;
assign w3561 = ~w3556 & w3560;
assign w3562 = ~w2891 & ~w3561;
assign w3563 = w2850 & w3509;
assign w3564 = ~w2902 & w64599;
assign w3565 = ~w3553 & ~w3562;
assign w3566 = ~w3564 & w3565;
assign w3567 = ~pi0249 & w3566;
assign w3568 = pi0249 & ~w3566;
assign w3569 = ~w3567 & ~w3568;
assign w3570 = ~w3377 & w3432;
assign w3571 = ~w3364 & w3370;
assign w3572 = w3392 & ~w3571;
assign w3573 = w3401 & ~w3572;
assign w3574 = ~w3409 & ~w3573;
assign w3575 = ~w3391 & ~w3435;
assign w3576 = ~w3574 & w3575;
assign w3577 = ~w3421 & ~w3576;
assign w3578 = w3392 & w3571;
assign w3579 = ~w3411 & ~w3578;
assign w3580 = ~w3389 & w3579;
assign w3581 = w3409 & ~w3580;
assign w3582 = ~w3400 & w3403;
assign w3583 = ~w3390 & w3423;
assign w3584 = w3393 & ~w3583;
assign w3585 = w3407 & w3584;
assign w3586 = w3579 & ~w3582;
assign w3587 = ~w3585 & w3586;
assign w3588 = w3421 & ~w3587;
assign w3589 = ~w3570 & ~w3581;
assign w3590 = ~w3588 & w3589;
assign w3591 = ~w3577 & w3590;
assign w3592 = pi0243 & ~w3591;
assign w3593 = ~pi0243 & w3591;
assign w3594 = ~w3592 & ~w3593;
assign w3595 = w2872 & ~w2878;
assign w3596 = w2844 & ~w2908;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = ~w2877 & w2896;
assign w3599 = w2913 & ~w3557;
assign w3600 = w2875 & w3543;
assign w3601 = ~w2891 & ~w3600;
assign w3602 = ~w3599 & w3601;
assign w3603 = ~w3598 & w3602;
assign w3604 = w2857 & w2869;
assign w3605 = ~w2869 & w3558;
assign w3606 = ~w3604 & ~w3605;
assign w3607 = ~w2844 & ~w3606;
assign w3608 = w2844 & ~w3604;
assign w3609 = w3499 & w3608;
assign w3610 = ~w2899 & ~w2909;
assign w3611 = w3503 & w3610;
assign w3612 = ~w3609 & w3611;
assign w3613 = ~w3607 & w3612;
assign w3614 = ~w3603 & ~w3613;
assign w3615 = ~w3597 & ~w3614;
assign w3616 = ~pi0252 & w3615;
assign w3617 = pi0252 & ~w3615;
assign w3618 = ~w3616 & ~w3617;
assign w3619 = w2784 & w2796;
assign w3620 = w2778 & ~w3619;
assign w3621 = ~w2803 & w2926;
assign w3622 = ~w3620 & ~w3621;
assign w3623 = ~w2744 & ~w2801;
assign w3624 = w2738 & ~w2758;
assign w3625 = ~w3623 & w3624;
assign w3626 = w2778 & w64600;
assign w3627 = w2774 & ~w2941;
assign w3628 = ~w2768 & ~w3627;
assign w3629 = ~w3625 & w3628;
assign w3630 = ~w3626 & w3629;
assign w3631 = ~w2792 & ~w3630;
assign w3632 = w2735 & w2803;
assign w3633 = w3487 & ~w3632;
assign w3634 = ~w2769 & ~w3633;
assign w3635 = (~w3622 & w64601) | (~w3622 & w64602) | (w64601 & w64602);
assign w3636 = ~w3631 & w3635;
assign w3637 = ~pi0244 & w3636;
assign w3638 = pi0244 & ~w3636;
assign w3639 = ~w3637 & ~w3638;
assign w3640 = ~pi3118 & pi9040;
assign w3641 = ~pi3086 & ~pi9040;
assign w3642 = ~w3640 & ~w3641;
assign w3643 = pi0217 & ~w3642;
assign w3644 = ~pi0217 & w3642;
assign w3645 = ~w3643 & ~w3644;
assign w3646 = ~pi3094 & pi9040;
assign w3647 = ~pi3093 & ~pi9040;
assign w3648 = ~w3646 & ~w3647;
assign w3649 = pi0181 & ~w3648;
assign w3650 = ~pi0181 & w3648;
assign w3651 = ~w3649 & ~w3650;
assign w3652 = w3645 & w3651;
assign w3653 = ~pi3082 & pi9040;
assign w3654 = ~pi3122 & ~pi9040;
assign w3655 = ~w3653 & ~w3654;
assign w3656 = pi0205 & ~w3655;
assign w3657 = ~pi0205 & w3655;
assign w3658 = ~w3656 & ~w3657;
assign w3659 = ~w3645 & ~w3658;
assign w3660 = ~w3651 & w3659;
assign w3661 = ~w3652 & ~w3660;
assign w3662 = ~pi3090 & pi9040;
assign w3663 = ~pi3094 & ~pi9040;
assign w3664 = ~w3662 & ~w3663;
assign w3665 = pi0214 & ~w3664;
assign w3666 = ~pi0214 & w3664;
assign w3667 = ~w3665 & ~w3666;
assign w3668 = ~w3661 & ~w3667;
assign w3669 = w3645 & ~w3667;
assign w3670 = w3652 & ~w3658;
assign w3671 = ~w3645 & w3667;
assign w3672 = w3658 & w3671;
assign w3673 = ~w3670 & ~w3672;
assign w3674 = ~w3669 & w3673;
assign w3675 = ~pi3225 & pi9040;
assign w3676 = ~pi3090 & ~pi9040;
assign w3677 = ~w3675 & ~w3676;
assign w3678 = pi0203 & ~w3677;
assign w3679 = ~pi0203 & w3677;
assign w3680 = ~w3678 & ~w3679;
assign w3681 = (w3680 & ~w3673) | (w3680 & w64603) | (~w3673 & w64603);
assign w3682 = ~w3668 & ~w3681;
assign w3683 = ~pi3168 & pi9040;
assign w3684 = ~pi3092 & ~pi9040;
assign w3685 = ~w3683 & ~w3684;
assign w3686 = pi0176 & ~w3685;
assign w3687 = ~pi0176 & w3685;
assign w3688 = ~w3686 & ~w3687;
assign w3689 = ~w3682 & w3688;
assign w3690 = w3645 & w3658;
assign w3691 = ~w3659 & ~w3690;
assign w3692 = ~w3658 & w3688;
assign w3693 = w3691 & ~w3692;
assign w3694 = ~w3651 & w3667;
assign w3695 = ~w3693 & w3694;
assign w3696 = w3652 & w64604;
assign w3697 = w3667 & ~w3690;
assign w3698 = ~w3667 & w3690;
assign w3699 = ~w3697 & ~w3698;
assign w3700 = ~w3659 & ~w3699;
assign w3701 = (~w3651 & w3699) | (~w3651 & w3660) | (w3699 & w3660);
assign w3702 = (w3693 & w3701) | (w3693 & w63551) | (w3701 & w63551);
assign w3703 = ~w3667 & ~w3691;
assign w3704 = (w3651 & w3703) | (w3651 & w64605) | (w3703 & w64605);
assign w3705 = ~w3695 & ~w3704;
assign w3706 = ~w3702 & w3705;
assign w3707 = ~w3680 & ~w3706;
assign w3708 = w3680 & ~w3688;
assign w3709 = ~w3659 & w3708;
assign w3710 = w3674 & w3709;
assign w3711 = ~w3658 & w3671;
assign w3712 = w3651 & w3680;
assign w3713 = w3711 & w3712;
assign w3714 = ~w3710 & ~w3713;
assign w3715 = ~w3689 & w3714;
assign w3716 = ~w3707 & w3715;
assign w3717 = pi0259 & ~w3716;
assign w3718 = ~pi0259 & w3716;
assign w3719 = ~w3717 & ~w3718;
assign w3720 = w3072 & ~w3110;
assign w3721 = ~w3105 & ~w3720;
assign w3722 = w3082 & ~w3721;
assign w3723 = w3082 & w3343;
assign w3724 = w3037 & ~w3059;
assign w3725 = ~w3137 & w3724;
assign w3726 = w3338 & ~w3725;
assign w3727 = ~w3723 & ~w3726;
assign w3728 = ~w3722 & ~w3727;
assign w3729 = ~pi0232 & w3728;
assign w3730 = pi0232 & ~w3728;
assign w3731 = ~w3729 & ~w3730;
assign w3732 = w3651 & w3658;
assign w3733 = ~w3671 & ~w3732;
assign w3734 = w3688 & ~w3733;
assign w3735 = (w3659 & w3733) | (w3659 & w64606) | (w3733 & w64606);
assign w3736 = w3701 & ~w3735;
assign w3737 = (~w3688 & ~w3659) | (~w3688 & w63552) | (~w3659 & w63552);
assign w3738 = ~w3645 & w3737;
assign w3739 = w3737 & w64607;
assign w3740 = ~w3696 & ~w3739;
assign w3741 = (w3680 & w3736) | (w3680 & w64608) | (w3736 & w64608);
assign w3742 = ~w3667 & w3732;
assign w3743 = ~w3680 & ~w3738;
assign w3744 = ~w3699 & w3737;
assign w3745 = w3743 & ~w3744;
assign w3746 = ~w3742 & ~w3745;
assign w3747 = ~w3691 & w63553;
assign w3748 = (~w3680 & w3700) | (~w3680 & w64609) | (w3700 & w64609);
assign w3749 = w3688 & ~w3748;
assign w3750 = ~w3746 & ~w3749;
assign w3751 = ~w3645 & w3688;
assign w3752 = w3704 & w3751;
assign w3753 = ~w3741 & ~w3752;
assign w3754 = ~w3750 & w3753;
assign w3755 = ~pi0253 & w3754;
assign w3756 = pi0253 & ~w3754;
assign w3757 = ~w3755 & ~w3756;
assign w3758 = w2983 & ~w2992;
assign w3759 = w2961 & w2974;
assign w3760 = ~w3325 & ~w3759;
assign w3761 = w3319 & ~w3760;
assign w3762 = w2955 & ~w2992;
assign w3763 = ~w3262 & ~w3762;
assign w3764 = ~w3275 & ~w3759;
assign w3765 = ~w3763 & w3764;
assign w3766 = w2992 & ~w3285;
assign w3767 = w2982 & ~w3765;
assign w3768 = ~w3766 & w3767;
assign w3769 = ~w3021 & ~w3261;
assign w3770 = w3295 & ~w3769;
assign w3771 = ~w3008 & ~w3323;
assign w3772 = w3014 & w3771;
assign w3773 = ~w3770 & w3772;
assign w3774 = ~w3768 & ~w3773;
assign w3775 = ~w3758 & ~w3761;
assign w3776 = ~w3774 & w3775;
assign w3777 = ~pi0267 & ~w3776;
assign w3778 = pi0267 & w3776;
assign w3779 = ~w3777 & ~w3778;
assign w3780 = ~w3688 & ~w3691;
assign w3781 = w3694 & ~w3780;
assign w3782 = ~w3660 & w64610;
assign w3783 = w3673 & ~w3747;
assign w3784 = ~w3688 & ~w3783;
assign w3785 = ~w3711 & ~w3742;
assign w3786 = ~w3780 & ~w3785;
assign w3787 = ~w3782 & ~w3786;
assign w3788 = ~w3784 & w3787;
assign w3789 = w3680 & ~w3781;
assign w3790 = ~w3680 & ~w3788;
assign w3791 = w3651 & w3688;
assign w3792 = ~w3692 & ~w3732;
assign w3793 = w3645 & w3667;
assign w3794 = ~w3791 & w3793;
assign w3795 = ~w3792 & w3794;
assign w3796 = w3688 & w3702;
assign w3797 = (~w3795 & ~w3788) | (~w3795 & w64611) | (~w3788 & w64611);
assign w3798 = ~w3790 & ~w3796;
assign w3799 = (pi0260 & ~w3798) | (pi0260 & w64612) | (~w3798 & w64612);
assign w3800 = w3798 & w64613;
assign w3801 = ~w3799 & ~w3800;
assign w3802 = w3645 & w3786;
assign w3803 = w3651 & w3697;
assign w3804 = ~w3743 & w3803;
assign w3805 = ~w3711 & ~w3732;
assign w3806 = w3708 & ~w3805;
assign w3807 = w3680 & ~w3782;
assign w3808 = (w3807 & ~w3702) | (w3807 & w64614) | (~w3702 & w64614);
assign w3809 = w3734 & ~w3803;
assign w3810 = ~w3667 & ~w3783;
assign w3811 = ~w3658 & ~w3667;
assign w3812 = ~w3688 & ~w3811;
assign w3813 = w3733 & w3812;
assign w3814 = ~w3680 & ~w3813;
assign w3815 = ~w3809 & w3814;
assign w3816 = ~w3810 & w3815;
assign w3817 = ~w3808 & ~w3816;
assign w3818 = ~w3802 & ~w3806;
assign w3819 = ~w3804 & w3818;
assign w3820 = ~w3817 & w3819;
assign w3821 = pi0268 & ~w3820;
assign w3822 = ~pi0268 & w3820;
assign w3823 = ~w3821 & ~w3822;
assign w3824 = ~w3400 & ~w3579;
assign w3825 = w3378 & ~w3400;
assign w3826 = w3431 & w3825;
assign w3827 = w3377 & ~w3403;
assign w3828 = ~w3412 & ~w3827;
assign w3829 = (~w3392 & w3827) | (~w3392 & w64615) | (w3827 & w64615);
assign w3830 = ~w3391 & w3400;
assign w3831 = ~w3829 & w3830;
assign w3832 = ~w3405 & w3831;
assign w3833 = w3386 & w3571;
assign w3834 = ~w3403 & ~w3833;
assign w3835 = ~w3406 & ~w3430;
assign w3836 = ~w3834 & w3835;
assign w3837 = ~w3377 & w3425;
assign w3838 = ~w3825 & ~w3837;
assign w3839 = w3390 & ~w3838;
assign w3840 = ~w3826 & ~w3839;
assign w3841 = ~w3836 & w3840;
assign w3842 = (w3421 & ~w3841) | (w3421 & w64616) | (~w3841 & w64616);
assign w3843 = ~w3582 & w3838;
assign w3844 = w3835 & ~w3843;
assign w3845 = ~w3421 & ~w3831;
assign w3846 = ~w3844 & w3845;
assign w3847 = ~w3371 & ~w3433;
assign w3848 = w3583 & w3847;
assign w3849 = ~w3824 & ~w3848;
assign w3850 = ~w3846 & w3849;
assign w3851 = ~w3842 & w3850;
assign w3852 = pi0246 & ~w3851;
assign w3853 = ~pi0246 & w3851;
assign w3854 = ~w3852 & ~w3853;
assign w3855 = w3407 & ~w3578;
assign w3856 = ~w3370 & w3434;
assign w3857 = ~w3401 & ~w3582;
assign w3858 = ~w3856 & ~w3857;
assign w3859 = ~w3855 & ~w3858;
assign w3860 = ~w3386 & w3571;
assign w3861 = ~w3405 & ~w3426;
assign w3862 = w3400 & ~w3861;
assign w3863 = ~w3388 & w3401;
assign w3864 = ~w3862 & ~w3863;
assign w3865 = ~w3421 & ~w3860;
assign w3866 = ~w3864 & w3865;
assign w3867 = ~w3386 & w3400;
assign w3868 = w3828 & w3867;
assign w3869 = ~w3385 & w3825;
assign w3870 = w3421 & ~w3430;
assign w3871 = ~w3833 & w3870;
assign w3872 = ~w3869 & w3871;
assign w3873 = ~w3868 & w3872;
assign w3874 = ~w3866 & ~w3873;
assign w3875 = ~w3859 & ~w3874;
assign w3876 = ~pi0258 & w3875;
assign w3877 = pi0258 & ~w3875;
assign w3878 = ~w3876 & ~w3877;
assign w3879 = ~pi3171 & pi9040;
assign w3880 = ~pi3181 & ~pi9040;
assign w3881 = ~w3879 & ~w3880;
assign w3882 = pi0279 & ~w3881;
assign w3883 = ~pi0279 & w3881;
assign w3884 = ~w3882 & ~w3883;
assign w3885 = ~pi3158 & pi9040;
assign w3886 = ~pi3128 & ~pi9040;
assign w3887 = ~w3885 & ~w3886;
assign w3888 = pi0272 & ~w3887;
assign w3889 = ~pi0272 & w3887;
assign w3890 = ~w3888 & ~w3889;
assign w3891 = w3884 & w3890;
assign w3892 = ~pi3151 & pi9040;
assign w3893 = ~pi3235 & ~pi9040;
assign w3894 = ~w3892 & ~w3893;
assign w3895 = pi0256 & ~w3894;
assign w3896 = ~pi0256 & w3894;
assign w3897 = ~w3895 & ~w3896;
assign w3898 = w3891 & ~w3897;
assign w3899 = ~w3890 & ~w3897;
assign w3900 = ~w3884 & w3899;
assign w3901 = ~w3898 & ~w3900;
assign w3902 = ~pi3182 & pi9040;
assign w3903 = ~pi3152 & ~pi9040;
assign w3904 = ~w3902 & ~w3903;
assign w3905 = pi0264 & ~w3904;
assign w3906 = ~pi0264 & w3904;
assign w3907 = ~w3905 & ~w3906;
assign w3908 = w3901 & w3907;
assign w3909 = ~pi3196 & pi9040;
assign w3910 = ~pi3171 & ~pi9040;
assign w3911 = ~w3909 & ~w3910;
assign w3912 = pi0245 & ~w3911;
assign w3913 = ~pi0245 & w3911;
assign w3914 = ~w3912 & ~w3913;
assign w3915 = ~w3897 & ~w3914;
assign w3916 = w3897 & w3914;
assign w3917 = ~w3915 & ~w3916;
assign w3918 = ~w3890 & w3897;
assign w3919 = ~w3917 & ~w3918;
assign w3920 = w3908 & w3919;
assign w3921 = ~pi3136 & pi9040;
assign w3922 = ~pi3183 & ~pi9040;
assign w3923 = ~w3921 & ~w3922;
assign w3924 = pi0285 & ~w3923;
assign w3925 = ~pi0285 & w3923;
assign w3926 = ~w3924 & ~w3925;
assign w3927 = ~w3907 & ~w3926;
assign w3928 = w3884 & w3927;
assign w3929 = w3917 & w3928;
assign w3930 = ~w3907 & ~w3914;
assign w3931 = ~w3884 & w3897;
assign w3932 = w3890 & w3897;
assign w3933 = ~w3931 & ~w3932;
assign w3934 = w3930 & w3933;
assign w3935 = ~w3884 & w3914;
assign w3936 = w3899 & w3935;
assign w3937 = w3884 & ~w3914;
assign w3938 = w3899 & ~w3937;
assign w3939 = w3890 & w3916;
assign w3940 = ~w3938 & ~w3939;
assign w3941 = ~w3907 & ~w3940;
assign w3942 = w3918 & w3930;
assign w3943 = w3932 & w3935;
assign w3944 = ~w3942 & ~w3943;
assign w3945 = ~w3936 & w3944;
assign w3946 = ~w3941 & w3945;
assign w3947 = w3934 & ~w3946;
assign w3948 = w3884 & w3918;
assign w3949 = w3890 & w3931;
assign w3950 = ~w3948 & ~w3949;
assign w3951 = ~w3915 & ~w3935;
assign w3952 = w3950 & w3951;
assign w3953 = (w3907 & ~w3950) | (w3907 & w64617) | (~w3950 & w64617);
assign w3954 = w3930 & ~w3949;
assign w3955 = ~w3907 & w3914;
assign w3956 = ~w3884 & ~w3897;
assign w3957 = ~w3918 & w3955;
assign w3958 = ~w3956 & w3957;
assign w3959 = ~w3954 & ~w3958;
assign w3960 = w3891 & w3915;
assign w3961 = ~w3959 & ~w3960;
assign w3962 = (w3926 & w3961) | (w3926 & w64618) | (w3961 & w64618);
assign w3963 = w3907 & w3935;
assign w3964 = ~w3890 & w3937;
assign w3965 = ~w3963 & ~w3964;
assign w3966 = w3897 & ~w3965;
assign w3967 = w3890 & w3914;
assign w3968 = w3956 & w3967;
assign w3969 = ~w3915 & ~w3968;
assign w3970 = w3907 & ~w3969;
assign w3971 = ~w3926 & w3944;
assign w3972 = ~w3966 & w3971;
assign w3973 = ~w3970 & w3972;
assign w3974 = ~w3962 & ~w3973;
assign w3975 = ~w3920 & ~w3929;
assign w3976 = ~w3947 & w3975;
assign w3977 = ~w3974 & w3976;
assign w3978 = pi0291 & ~w3977;
assign w3979 = ~pi0291 & w3977;
assign w3980 = ~w3978 & ~w3979;
assign w3981 = ~pi3147 & pi9040;
assign w3982 = ~pi3308 & ~pi9040;
assign w3983 = ~w3981 & ~w3982;
assign w3984 = pi0276 & ~w3983;
assign w3985 = ~pi0276 & w3983;
assign w3986 = ~w3984 & ~w3985;
assign w3987 = ~pi3175 & pi9040;
assign w3988 = ~pi3154 & ~pi9040;
assign w3989 = ~w3987 & ~w3988;
assign w3990 = pi0278 & ~w3989;
assign w3991 = ~pi0278 & w3989;
assign w3992 = ~w3990 & ~w3991;
assign w3993 = w3986 & w3992;
assign w3994 = ~pi3198 & pi9040;
assign w3995 = ~pi3159 & ~pi9040;
assign w3996 = ~w3994 & ~w3995;
assign w3997 = pi0255 & ~w3996;
assign w3998 = ~pi0255 & w3996;
assign w3999 = ~w3997 & ~w3998;
assign w4000 = w3992 & w3999;
assign w4001 = ~w3993 & ~w4000;
assign w4002 = ~pi3224 & pi9040;
assign w4003 = ~pi3167 & ~pi9040;
assign w4004 = ~w4002 & ~w4003;
assign w4005 = pi0251 & ~w4004;
assign w4006 = ~pi0251 & w4004;
assign w4007 = ~w4005 & ~w4006;
assign w4008 = ~w3999 & ~w4007;
assign w4009 = ~pi3156 & pi9040;
assign w4010 = ~pi3224 & ~pi9040;
assign w4011 = ~w4009 & ~w4010;
assign w4012 = pi0277 & ~w4011;
assign w4013 = ~pi0277 & w4011;
assign w4014 = ~w4012 & ~w4013;
assign w4015 = w4008 & ~w4014;
assign w4016 = ~w3999 & w4014;
assign w4017 = w4007 & w4016;
assign w4018 = ~w4015 & ~w4017;
assign w4019 = w3999 & ~w4007;
assign w4020 = w4014 & ~w4019;
assign w4021 = w3993 & w4020;
assign w4022 = w3999 & w4007;
assign w4023 = w3999 & ~w4014;
assign w4024 = ~w3986 & ~w3992;
assign w4025 = ~w4022 & ~w4023;
assign w4026 = w4024 & w4025;
assign w4027 = ~w4021 & ~w4026;
assign w4028 = w3992 & ~w4018;
assign w4029 = w4027 & w4028;
assign w4030 = w4001 & w4029;
assign w4031 = ~w3999 & w4007;
assign w4032 = w3993 & w4031;
assign w4033 = ~w4014 & w4032;
assign w4034 = w3986 & ~w4007;
assign w4035 = w4023 & w4034;
assign w4036 = ~w3992 & w4035;
assign w4037 = w3992 & w4014;
assign w4038 = w4034 & w4037;
assign w4039 = w4016 & w4034;
assign w4040 = ~pi3155 & pi9040;
assign w4041 = ~pi3198 & ~pi9040;
assign w4042 = ~w4040 & ~w4041;
assign w4043 = pi0286 & ~w4042;
assign w4044 = ~pi0286 & w4042;
assign w4045 = ~w4043 & ~w4044;
assign w4046 = ~w4039 & ~w4045;
assign w4047 = ~w3986 & w3999;
assign w4048 = ~w4017 & ~w4047;
assign w4049 = ~w3992 & ~w4048;
assign w4050 = ~w3992 & w4014;
assign w4051 = ~w3986 & w4008;
assign w4052 = ~w4050 & w4051;
assign w4053 = ~w3986 & w4007;
assign w4054 = ~w4014 & w4053;
assign w4055 = ~w3993 & ~w4054;
assign w4056 = w4022 & ~w4055;
assign w4057 = ~w4038 & w4046;
assign w4058 = ~w4052 & w4057;
assign w4059 = ~w4049 & ~w4056;
assign w4060 = w4058 & w4059;
assign w4061 = ~w4034 & ~w4053;
assign w4062 = ~w3992 & ~w4014;
assign w4063 = ~w4061 & w4062;
assign w4064 = ~w4022 & ~w4034;
assign w4065 = ~w4001 & w4064;
assign w4066 = w4050 & w4051;
assign w4067 = w4014 & ~w4022;
assign w4068 = ~w4014 & ~w4019;
assign w4069 = ~w4067 & ~w4068;
assign w4070 = w3986 & w4069;
assign w4071 = w4045 & ~w4063;
assign w4072 = ~w4065 & ~w4066;
assign w4073 = w4071 & w4072;
assign w4074 = ~w4070 & w4073;
assign w4075 = ~w4060 & ~w4074;
assign w4076 = ~w4033 & ~w4036;
assign w4077 = ~w4030 & w4076;
assign w4078 = ~w4075 & w4077;
assign w4079 = pi0293 & w4078;
assign w4080 = ~pi0293 & ~w4078;
assign w4081 = ~w4079 & ~w4080;
assign w4082 = ~pi3296 & pi9040;
assign w4083 = ~pi3176 & ~pi9040;
assign w4084 = ~w4082 & ~w4083;
assign w4085 = pi0262 & ~w4084;
assign w4086 = ~pi0262 & w4084;
assign w4087 = ~w4085 & ~w4086;
assign w4088 = ~pi3132 & pi9040;
assign w4089 = ~pi3129 & ~pi9040;
assign w4090 = ~w4088 & ~w4089;
assign w4091 = pi0266 & ~w4090;
assign w4092 = ~pi0266 & w4090;
assign w4093 = ~w4091 & ~w4092;
assign w4094 = w4087 & w4093;
assign w4095 = ~pi3148 & pi9040;
assign w4096 = ~pi3240 & ~pi9040;
assign w4097 = ~w4095 & ~w4096;
assign w4098 = pi0271 & ~w4097;
assign w4099 = ~pi0271 & w4097;
assign w4100 = ~w4098 & ~w4099;
assign w4101 = ~pi3183 & pi9040;
assign w4102 = ~pi3194 & ~pi9040;
assign w4103 = ~w4101 & ~w4102;
assign w4104 = pi0287 & ~w4103;
assign w4105 = ~pi0287 & w4103;
assign w4106 = ~w4104 & ~w4105;
assign w4107 = ~w4100 & ~w4106;
assign w4108 = ~pi3145 & pi9040;
assign w4109 = ~pi3134 & ~pi9040;
assign w4110 = ~w4108 & ~w4109;
assign w4111 = pi0254 & ~w4110;
assign w4112 = ~pi0254 & w4110;
assign w4113 = ~w4111 & ~w4112;
assign w4114 = w4107 & ~w4113;
assign w4115 = w4094 & w4114;
assign w4116 = ~w4087 & ~w4093;
assign w4117 = ~w4106 & w4116;
assign w4118 = ~w4093 & w4106;
assign w4119 = w4087 & w4118;
assign w4120 = ~w4117 & ~w4119;
assign w4121 = ~w4100 & ~w4120;
assign w4122 = w4093 & ~w4100;
assign w4123 = ~w4087 & w4106;
assign w4124 = w4122 & w4123;
assign w4125 = w4100 & w4116;
assign w4126 = ~w4124 & ~w4125;
assign w4127 = ~pi3181 & pi9040;
assign w4128 = ~pi3132 & ~pi9040;
assign w4129 = ~w4127 & ~w4128;
assign w4130 = pi0273 & ~w4129;
assign w4131 = ~pi0273 & w4129;
assign w4132 = ~w4130 & ~w4131;
assign w4133 = ~w4126 & ~w4132;
assign w4134 = ~w4087 & w4100;
assign w4135 = w4093 & w4123;
assign w4136 = ~w4117 & ~w4135;
assign w4137 = w4134 & w4136;
assign w4138 = ~w4121 & ~w4133;
assign w4139 = (w4113 & ~w4138) | (w4113 & w64619) | (~w4138 & w64619);
assign w4140 = w4093 & ~w4106;
assign w4141 = w4087 & w4107;
assign w4142 = w4113 & ~w4141;
assign w4143 = w4140 & ~w4142;
assign w4144 = ~w4113 & w4118;
assign w4145 = ~w4100 & w4144;
assign w4146 = w4087 & w4100;
assign w4147 = w4094 & w4106;
assign w4148 = w4113 & ~w4147;
assign w4149 = w4146 & ~w4148;
assign w4150 = ~w4132 & ~w4145;
assign w4151 = ~w4143 & w4150;
assign w4152 = ~w4149 & w4151;
assign w4153 = w4118 & w4146;
assign w4154 = ~w4113 & ~w4136;
assign w4155 = w4087 & ~w4100;
assign w4156 = ~w4140 & ~w4155;
assign w4157 = w4113 & ~w4122;
assign w4158 = ~w4142 & ~w4157;
assign w4159 = ~w4156 & ~w4158;
assign w4160 = w4132 & ~w4153;
assign w4161 = ~w4154 & w4160;
assign w4162 = ~w4159 & w4161;
assign w4163 = ~w4152 & ~w4162;
assign w4164 = ~w4115 & ~w4139;
assign w4165 = ~w4163 & w4164;
assign w4166 = ~pi0288 & w4165;
assign w4167 = pi0288 & ~w4165;
assign w4168 = ~w4166 & ~w4167;
assign w4169 = ~w4037 & w4051;
assign w4170 = w4022 & w4062;
assign w4171 = w3992 & ~w4023;
assign w4172 = w4053 & w4171;
assign w4173 = ~w4000 & ~w4007;
assign w4174 = ~w4014 & ~w4053;
assign w4175 = ~w4173 & w4174;
assign w4176 = w4046 & ~w4170;
assign w4177 = ~w4169 & ~w4172;
assign w4178 = ~w4175 & w4177;
assign w4179 = w4176 & w4178;
assign w4180 = ~w4024 & ~w4050;
assign w4181 = w4031 & ~w4180;
assign w4182 = ~w4008 & ~w4054;
assign w4183 = ~w4001 & ~w4182;
assign w4184 = w3999 & w4014;
assign w4185 = w4061 & w4184;
assign w4186 = ~w4036 & w4045;
assign w4187 = ~w4181 & ~w4185;
assign w4188 = w4186 & w4187;
assign w4189 = ~w4183 & w4188;
assign w4190 = ~w4179 & ~w4189;
assign w4191 = ~w4015 & ~w4185;
assign w4192 = ~w4180 & ~w4191;
assign w4193 = ~w4033 & ~w4038;
assign w4194 = ~w4192 & w4193;
assign w4195 = ~w4190 & w4194;
assign w4196 = pi0300 & ~w4195;
assign w4197 = ~pi0300 & w4195;
assign w4198 = ~w4196 & ~w4197;
assign w4199 = w3899 & w3937;
assign w4200 = w3914 & w3948;
assign w4201 = ~w3898 & ~w4199;
assign w4202 = ~w4200 & w4201;
assign w4203 = w3907 & ~w4202;
assign w4204 = w3890 & w3915;
assign w4205 = w3915 & w64620;
assign w4206 = w3926 & ~w4205;
assign w4207 = w3946 & w4206;
assign w4208 = ~w4203 & w4207;
assign w4209 = ~w3933 & ~w3949;
assign w4210 = ~w3938 & ~w4209;
assign w4211 = w3907 & ~w3936;
assign w4212 = ~w4210 & w4211;
assign w4213 = ~w3926 & ~w3968;
assign w4214 = ~w4212 & w4213;
assign w4215 = ~w4208 & ~w4214;
assign w4216 = w3890 & ~w3930;
assign w4217 = w3937 & w4216;
assign w4218 = ~w3884 & w3952;
assign w4219 = ~w3932 & w4202;
assign w4220 = w3927 & ~w3967;
assign w4221 = ~w4219 & w4220;
assign w4222 = ~w4217 & ~w4218;
assign w4223 = ~w4221 & w4222;
assign w4224 = (pi0290 & w4215) | (pi0290 & w64621) | (w4215 & w64621);
assign w4225 = ~w4215 & w64622;
assign w4226 = ~w4224 & ~w4225;
assign w4227 = w4069 & ~w4180;
assign w4228 = w3986 & ~w4018;
assign w4229 = w3986 & ~w3999;
assign w4230 = ~w4024 & ~w4229;
assign w4231 = ~w4007 & ~w4023;
assign w4232 = w4230 & w4231;
assign w4233 = ~w4227 & ~w4232;
assign w4234 = (w4045 & ~w4233) | (w4045 & w64623) | (~w4233 & w64623);
assign w4235 = w3986 & ~w3992;
assign w4236 = ~w4031 & w4235;
assign w4237 = ~w4181 & ~w4236;
assign w4238 = w4068 & ~w4237;
assign w4239 = ~w4000 & w4045;
assign w4240 = ~w4027 & ~w4045;
assign w4241 = ~w4032 & ~w4035;
assign w4242 = ~w4054 & w4241;
assign w4243 = ~w4240 & w4242;
assign w4244 = ~w4239 & ~w4243;
assign w4245 = ~w4234 & ~w4238;
assign w4246 = ~w4244 & w4245;
assign w4247 = pi0310 & w4246;
assign w4248 = ~pi0310 & ~w4246;
assign w4249 = ~w4247 & ~w4248;
assign w4250 = w3930 & ~w3950;
assign w4251 = w3884 & w3939;
assign w4252 = w3897 & w3937;
assign w4253 = ~w3956 & ~w4252;
assign w4254 = w3908 & w4253;
assign w4255 = ~w3901 & ~w3907;
assign w4256 = ~w3926 & ~w4251;
assign w4257 = ~w4255 & w4256;
assign w4258 = ~w4254 & w4257;
assign w4259 = ~w3901 & w3914;
assign w4260 = ~w3907 & w3931;
assign w4261 = w3908 & ~w4253;
assign w4262 = ~w3964 & ~w4260;
assign w4263 = w4206 & w4262;
assign w4264 = ~w4259 & w4263;
assign w4265 = ~w4261 & w4264;
assign w4266 = ~w4258 & ~w4265;
assign w4267 = w3907 & w4205;
assign w4268 = ~w4250 & ~w4267;
assign w4269 = ~w4266 & w4268;
assign w4270 = pi0296 & ~w4269;
assign w4271 = ~pi0296 & w4269;
assign w4272 = ~w4270 & ~w4271;
assign w4273 = ~w4047 & ~w4054;
assign w4274 = w4045 & ~w4273;
assign w4275 = ~w4039 & ~w4185;
assign w4276 = ~w4274 & w4275;
assign w4277 = w3992 & ~w4276;
assign w4278 = w4045 & w4067;
assign w4279 = ~w3992 & w4016;
assign w4280 = ~w4278 & ~w4279;
assign w4281 = w4061 & ~w4280;
assign w4282 = ~w4020 & w4045;
assign w4283 = w4236 & w4282;
assign w4284 = w4007 & ~w4016;
assign w4285 = ~w4230 & w4284;
assign w4286 = ~w4070 & ~w4285;
assign w4287 = ~w4029 & w4286;
assign w4288 = ~w4045 & ~w4287;
assign w4289 = ~w4281 & ~w4283;
assign w4290 = ~w4277 & w4289;
assign w4291 = ~w4288 & w4290;
assign w4292 = pi0306 & ~w4291;
assign w4293 = ~pi0306 & w4291;
assign w4294 = ~w4292 & ~w4293;
assign w4295 = ~pi3176 & pi9040;
assign w4296 = ~pi3158 & ~pi9040;
assign w4297 = ~w4295 & ~w4296;
assign w4298 = pi0282 & ~w4297;
assign w4299 = ~pi0282 & w4297;
assign w4300 = ~w4298 & ~w4299;
assign w4301 = ~pi3128 & pi9040;
assign w4302 = ~pi3142 & ~pi9040;
assign w4303 = ~w4301 & ~w4302;
assign w4304 = pi0270 & ~w4303;
assign w4305 = ~pi0270 & w4303;
assign w4306 = ~w4304 & ~w4305;
assign w4307 = ~pi3150 & pi9040;
assign w4308 = ~pi3251 & ~pi9040;
assign w4309 = ~w4307 & ~w4308;
assign w4310 = pi0279 & ~w4309;
assign w4311 = ~pi0279 & w4309;
assign w4312 = ~w4310 & ~w4311;
assign w4313 = w4306 & ~w4312;
assign w4314 = ~pi3174 & pi9040;
assign w4315 = ~pi3139 & ~pi9040;
assign w4316 = ~w4314 & ~w4315;
assign w4317 = pi0255 & ~w4316;
assign w4318 = ~pi0255 & w4316;
assign w4319 = ~w4317 & ~w4318;
assign w4320 = ~pi3139 & pi9040;
assign w4321 = ~pi3151 & ~pi9040;
assign w4322 = ~w4320 & ~w4321;
assign w4323 = pi0286 & ~w4322;
assign w4324 = ~pi0286 & w4322;
assign w4325 = ~w4323 & ~w4324;
assign w4326 = ~w4319 & w4325;
assign w4327 = w4319 & ~w4325;
assign w4328 = ~w4326 & ~w4327;
assign w4329 = w4313 & w4328;
assign w4330 = w4312 & w4325;
assign w4331 = ~w4312 & ~w4325;
assign w4332 = ~w4330 & ~w4331;
assign w4333 = ~w4312 & ~w4319;
assign w4334 = w4306 & ~w4333;
assign w4335 = w4300 & w4330;
assign w4336 = w4334 & ~w4335;
assign w4337 = ~w4332 & w4336;
assign w4338 = ~pi3235 & pi9040;
assign w4339 = ~pi3145 & ~pi9040;
assign w4340 = ~w4338 & ~w4339;
assign w4341 = pi0256 & ~w4340;
assign w4342 = ~pi0256 & w4340;
assign w4343 = ~w4341 & ~w4342;
assign w4344 = w4327 & ~w4343;
assign w4345 = (w4344 & ~w4336) | (w4344 & w64624) | (~w4336 & w64624);
assign w4346 = ~w4329 & ~w4345;
assign w4347 = w4300 & ~w4346;
assign w4348 = ~w4306 & ~w4319;
assign w4349 = ~w4300 & w4319;
assign w4350 = w4313 & w4349;
assign w4351 = ~w4348 & ~w4350;
assign w4352 = w4300 & ~w4325;
assign w4353 = ~w4330 & ~w4352;
assign w4354 = ~w4343 & w4353;
assign w4355 = ~w4351 & w4354;
assign w4356 = ~w4312 & w4325;
assign w4357 = ~w4300 & w4312;
assign w4358 = ~w4356 & ~w4357;
assign w4359 = w4300 & ~w4319;
assign w4360 = ~w4349 & ~w4359;
assign w4361 = w4356 & ~w4360;
assign w4362 = w4319 & ~w4358;
assign w4363 = ~w4361 & w4362;
assign w4364 = ~w4319 & w4330;
assign w4365 = ~w4325 & w4349;
assign w4366 = ~w4364 & ~w4365;
assign w4367 = ~w4306 & ~w4366;
assign w4368 = w4300 & ~w4312;
assign w4369 = ~w4319 & ~w4368;
assign w4370 = w4332 & ~w4369;
assign w4371 = w4306 & w4366;
assign w4372 = ~w4370 & w4371;
assign w4373 = ~w4363 & ~w4367;
assign w4374 = ~w4372 & w4373;
assign w4375 = w4343 & ~w4374;
assign w4376 = ~w4306 & w4325;
assign w4377 = w4359 & w4376;
assign w4378 = ~w4319 & ~w4325;
assign w4379 = w4334 & w4378;
assign w4380 = w4334 & w64625;
assign w4381 = w4330 & w4349;
assign w4382 = ~w4377 & ~w4381;
assign w4383 = ~w4380 & w4382;
assign w4384 = ~w4355 & w4383;
assign w4385 = ~w4347 & w4384;
assign w4386 = ~w4375 & w4385;
assign w4387 = ~pi0309 & w4386;
assign w4388 = pi0309 & ~w4386;
assign w4389 = ~w4387 & ~w4388;
assign w4390 = w3955 & w4209;
assign w4391 = ~w3943 & ~w3948;
assign w4392 = (~w3926 & ~w4391) | (~w3926 & w64626) | (~w4391 & w64626);
assign w4393 = ~w4200 & ~w4259;
assign w4394 = (w3907 & ~w4393) | (w3907 & w64627) | (~w4393 & w64627);
assign w4395 = w3927 & w3968;
assign w4396 = ~w3928 & ~w3930;
assign w4397 = w3899 & ~w4396;
assign w4398 = w3930 & w3932;
assign w4399 = ~w3926 & ~w4398;
assign w4400 = ~w4218 & w4399;
assign w4401 = w3951 & w4216;
assign w4402 = w3926 & ~w4199;
assign w4403 = ~w3934 & w4402;
assign w4404 = ~w4401 & w4403;
assign w4405 = ~w4400 & ~w4404;
assign w4406 = ~w4390 & ~w4395;
assign w4407 = ~w4397 & w4406;
assign w4408 = ~w4394 & w4407;
assign w4409 = ~w4405 & w4408;
assign w4410 = pi0295 & ~w4409;
assign w4411 = ~pi0295 & w4409;
assign w4412 = ~w4410 & ~w4411;
assign w4413 = ~pi3251 & pi9040;
assign w4414 = ~pi3136 & ~pi9040;
assign w4415 = ~w4413 & ~w4414;
assign w4416 = pi0285 & ~w4415;
assign w4417 = ~pi0285 & w4415;
assign w4418 = ~w4416 & ~w4417;
assign w4419 = ~pi3179 & pi9040;
assign w4420 = ~pi3182 & ~pi9040;
assign w4421 = ~w4419 & ~w4420;
assign w4422 = pi0281 & ~w4421;
assign w4423 = ~pi0281 & w4421;
assign w4424 = ~w4422 & ~w4423;
assign w4425 = w4418 & w4424;
assign w4426 = ~pi3134 & pi9040;
assign w4427 = ~pi3296 & ~pi9040;
assign w4428 = ~w4426 & ~w4427;
assign w4429 = pi0262 & ~w4428;
assign w4430 = ~pi0262 & w4428;
assign w4431 = ~w4429 & ~w4430;
assign w4432 = ~pi3240 & pi9040;
assign w4433 = ~pi3130 & ~pi9040;
assign w4434 = ~w4432 & ~w4433;
assign w4435 = pi0272 & ~w4434;
assign w4436 = ~pi0272 & w4434;
assign w4437 = ~w4435 & ~w4436;
assign w4438 = ~w4431 & ~w4437;
assign w4439 = ~pi3194 & pi9040;
assign w4440 = ~pi3179 & ~pi9040;
assign w4441 = ~w4439 & ~w4440;
assign w4442 = pi0265 & ~w4441;
assign w4443 = ~pi0265 & w4441;
assign w4444 = ~w4442 & ~w4443;
assign w4445 = ~w4418 & w4444;
assign w4446 = w4418 & ~w4431;
assign w4447 = ~w4445 & ~w4446;
assign w4448 = w4437 & w4444;
assign w4449 = w4447 & ~w4448;
assign w4450 = (~w4438 & ~w4447) | (~w4438 & w63554) | (~w4447 & w63554);
assign w4451 = ~w4437 & ~w4444;
assign w4452 = ~w4450 & ~w4451;
assign w4453 = ~w4450 & w64628;
assign w4454 = ~w4418 & w4431;
assign w4455 = ~w4446 & ~w4454;
assign w4456 = w4448 & ~w4455;
assign w4457 = w4450 & ~w4456;
assign w4458 = w4454 & w4457;
assign w4459 = w4438 & w4447;
assign w4460 = ~pi3152 & pi9040;
assign w4461 = ~pi3196 & ~pi9040;
assign w4462 = ~w4460 & ~w4461;
assign w4463 = pi0266 & ~w4462;
assign w4464 = ~pi0266 & w4462;
assign w4465 = ~w4463 & ~w4464;
assign w4466 = ~w4459 & w4465;
assign w4467 = ~w4453 & w4466;
assign w4468 = ~w4458 & w4467;
assign w4469 = w4438 & w4445;
assign w4470 = ~w4438 & ~w4445;
assign w4471 = ~w4469 & ~w4470;
assign w4472 = ~w4424 & ~w4471;
assign w4473 = w4418 & w4451;
assign w4474 = (w4473 & w4471) | (w4473 & w64629) | (w4471 & w64629);
assign w4475 = ~w4438 & ~w4444;
assign w4476 = w4455 & w4475;
assign w4477 = w4472 & ~w4476;
assign w4478 = w4431 & w4437;
assign w4479 = w4418 & ~w4444;
assign w4480 = ~w4445 & ~w4479;
assign w4481 = w4478 & w4480;
assign w4482 = ~w4465 & ~w4481;
assign w4483 = ~w4474 & w4482;
assign w4484 = ~w4477 & w4483;
assign w4485 = ~w4468 & ~w4484;
assign w4486 = w4424 & ~w4478;
assign w4487 = w4471 & w4486;
assign w4488 = w4454 & w4465;
assign w4489 = ~w4480 & ~w4488;
assign w4490 = w4437 & ~w4489;
assign w4491 = w4431 & w4473;
assign w4492 = w4465 & w4491;
assign w4493 = ~w4490 & ~w4492;
assign w4494 = ~w4424 & ~w4493;
assign w4495 = ~w4487 & ~w4494;
assign w4496 = ~w4485 & w4495;
assign w4497 = pi0292 & ~w4496;
assign w4498 = ~pi0292 & w4496;
assign w4499 = ~w4497 & ~w4498;
assign w4500 = ~pi3166 & pi9040;
assign w4501 = ~pi3177 & ~pi9040;
assign w4502 = ~w4500 & ~w4501;
assign w4503 = pi0271 & ~w4502;
assign w4504 = ~pi0271 & w4502;
assign w4505 = ~w4503 & ~w4504;
assign w4506 = ~pi3167 & pi9040;
assign w4507 = ~pi3227 & ~pi9040;
assign w4508 = ~w4506 & ~w4507;
assign w4509 = pi0250 & ~w4508;
assign w4510 = ~pi0250 & w4508;
assign w4511 = ~w4509 & ~w4510;
assign w4512 = ~w4505 & w4511;
assign w4513 = w4505 & ~w4511;
assign w4514 = ~w4512 & ~w4513;
assign w4515 = ~pi3308 & pi9040;
assign w4516 = ~pi3155 & ~pi9040;
assign w4517 = ~w4515 & ~w4516;
assign w4518 = pi0283 & ~w4517;
assign w4519 = ~pi0283 & w4517;
assign w4520 = ~w4518 & ~w4519;
assign w4521 = w4514 & w4520;
assign w4522 = ~pi3178 & pi9040;
assign w4523 = ~pi3140 & ~pi9040;
assign w4524 = ~w4522 & ~w4523;
assign w4525 = pi0273 & ~w4524;
assign w4526 = ~pi0273 & w4524;
assign w4527 = ~w4525 & ~w4526;
assign w4528 = ~w4511 & ~w4527;
assign w4529 = ~pi3133 & pi9040;
assign w4530 = ~pi3141 & ~pi9040;
assign w4531 = ~w4529 & ~w4530;
assign w4532 = pi0263 & ~w4531;
assign w4533 = ~pi0263 & w4531;
assign w4534 = ~w4532 & ~w4533;
assign w4535 = w4528 & w4534;
assign w4536 = w4521 & w4535;
assign w4537 = w4511 & w4534;
assign w4538 = w4505 & w4527;
assign w4539 = ~w4520 & w4538;
assign w4540 = w4537 & w4539;
assign w4541 = ~w4505 & ~w4534;
assign w4542 = w4520 & w4527;
assign w4543 = w4541 & w4542;
assign w4544 = ~w4540 & ~w4543;
assign w4545 = w4505 & w4534;
assign w4546 = ~w4541 & ~w4545;
assign w4547 = w4511 & w4527;
assign w4548 = ~w4528 & ~w4547;
assign w4549 = ~w4534 & w4548;
assign w4550 = ~w4514 & ~w4520;
assign w4551 = w4549 & w4550;
assign w4552 = ~w4527 & w4550;
assign w4553 = ~w4551 & ~w4552;
assign w4554 = w4546 & ~w4553;
assign w4555 = ~pi3143 & pi9040;
assign w4556 = ~pi3195 & ~pi9040;
assign w4557 = ~w4555 & ~w4556;
assign w4558 = pi0275 & ~w4557;
assign w4559 = ~pi0275 & w4557;
assign w4560 = ~w4558 & ~w4559;
assign w4561 = ~w4520 & ~w4527;
assign w4562 = ~w4538 & ~w4561;
assign w4563 = ~w4505 & ~w4527;
assign w4564 = ~w4520 & ~w4563;
assign w4565 = ~w4512 & ~w4535;
assign w4566 = ~w4564 & ~w4565;
assign w4567 = (~w4539 & ~w4549) | (~w4539 & w64630) | (~w4549 & w64630);
assign w4568 = ~w4566 & w4567;
assign w4569 = w4560 & w4568;
assign w4570 = ~w4514 & w4527;
assign w4571 = ~w4539 & ~w4546;
assign w4572 = w4570 & w4571;
assign w4573 = w4514 & w4562;
assign w4574 = w4527 & ~w4534;
assign w4575 = w4513 & w4574;
assign w4576 = w4511 & w4545;
assign w4577 = ~w4527 & ~w4541;
assign w4578 = ~w4520 & ~w4574;
assign w4579 = ~w4577 & w4578;
assign w4580 = ~w4575 & ~w4576;
assign w4581 = ~w4579 & w4580;
assign w4582 = w4573 & ~w4581;
assign w4583 = w4511 & ~w4534;
assign w4584 = w4542 & w4583;
assign w4585 = ~w4527 & ~w4534;
assign w4586 = ~w4512 & w4585;
assign w4587 = ~w4521 & w4586;
assign w4588 = ~w4560 & ~w4584;
assign w4589 = ~w4572 & w4588;
assign w4590 = ~w4587 & w4589;
assign w4591 = ~w4582 & w4590;
assign w4592 = ~w4569 & ~w4591;
assign w4593 = ~w4536 & w4544;
assign w4594 = ~w4554 & w4593;
assign w4595 = (pi0299 & w4592) | (pi0299 & w64631) | (w4592 & w64631);
assign w4596 = ~w4592 & w64632;
assign w4597 = ~w4595 & ~w4596;
assign w4598 = w4445 & w64633;
assign w4599 = w4438 & ~w4479;
assign w4600 = w4424 & w4444;
assign w4601 = ~w4486 & ~w4600;
assign w4602 = ~w4599 & ~w4601;
assign w4603 = (~w4448 & w4601) | (~w4448 & w63352) | (w4601 & w63352);
assign w4604 = w4454 & ~w4603;
assign w4605 = w4418 & ~w4600;
assign w4606 = ~w4475 & w4605;
assign w4607 = w4424 & ~w4469;
assign w4608 = ~w4438 & ~w4478;
assign w4609 = ~w4607 & ~w4608;
assign w4610 = ~w4451 & ~w4478;
assign w4611 = w4447 & w4610;
assign w4612 = ~w4606 & ~w4611;
assign w4613 = ~w4609 & w4612;
assign w4614 = ~w4604 & w4613;
assign w4615 = ~w4477 & w4614;
assign w4616 = w4452 & ~w4455;
assign w4617 = ~w4491 & ~w4598;
assign w4618 = (w4465 & w4615) | (w4465 & w63555) | (w4615 & w63555);
assign w4619 = ~w4465 & ~w4614;
assign w4620 = (pi0289 & w4618) | (pi0289 & w64634) | (w4618 & w64634);
assign w4621 = ~w4618 & w64635;
assign w4622 = ~w4620 & ~w4621;
assign w4623 = ~w4577 & ~w4584;
assign w4624 = w4562 & ~w4623;
assign w4625 = w4581 & ~w4624;
assign w4626 = w4560 & ~w4625;
assign w4627 = w4513 & w4520;
assign w4628 = ~w4586 & ~w4627;
assign w4629 = ~w4568 & ~w4628;
assign w4630 = ~w4520 & ~w4545;
assign w4631 = ~w4548 & ~w4630;
assign w4632 = w4514 & ~w4528;
assign w4633 = ~w4549 & ~w4631;
assign w4634 = ~w4632 & w4633;
assign w4635 = w4514 & w4542;
assign w4636 = ~w4634 & ~w4635;
assign w4637 = ~w4560 & ~w4636;
assign w4638 = ~w4626 & ~w4629;
assign w4639 = ~w4637 & w4638;
assign w4640 = ~pi0301 & w4639;
assign w4641 = pi0301 & ~w4639;
assign w4642 = ~w4640 & ~w4641;
assign w4643 = ~w4306 & w4312;
assign w4644 = w4328 & ~w4353;
assign w4645 = w4643 & ~w4644;
assign w4646 = w4328 & w4368;
assign w4647 = w4371 & w64636;
assign w4648 = ~w4365 & ~w4646;
assign w4649 = ~w4645 & w4648;
assign w4650 = ~w4647 & w4649;
assign w4651 = ~w4343 & ~w4650;
assign w4652 = ~w4300 & w4325;
assign w4653 = w4343 & w4652;
assign w4654 = w4326 & w4368;
assign w4655 = ~w4653 & ~w4654;
assign w4656 = ~w4306 & ~w4655;
assign w4657 = ~w4368 & ~w4378;
assign w4658 = ~w4333 & ~w4657;
assign w4659 = w4358 & w4658;
assign w4660 = w4306 & ~w4332;
assign w4661 = w4369 & w4660;
assign w4662 = ~w4659 & ~w4661;
assign w4663 = w4336 & w4383;
assign w4664 = ~w4374 & w4663;
assign w4665 = (~w4656 & w4662) | (~w4656 & w64637) | (w4662 & w64637);
assign w4666 = ~w4664 & w4665;
assign w4667 = (pi0297 & ~w4666) | (pi0297 & w64638) | (~w4666 & w64638);
assign w4668 = w4666 & w64639;
assign w4669 = ~w4667 & ~w4668;
assign w4670 = w4329 & ~w4360;
assign w4671 = w4327 & w4643;
assign w4672 = ~w4319 & w4331;
assign w4673 = ~w4671 & ~w4672;
assign w4674 = ~w4300 & ~w4673;
assign w4675 = ~w4659 & ~w4674;
assign w4676 = ~w4306 & ~w4675;
assign w4677 = ~w4357 & ~w4643;
assign w4678 = w4325 & w4360;
assign w4679 = ~w4677 & w4678;
assign w4680 = ~w4335 & ~w4365;
assign w4681 = ~w4331 & w4334;
assign w4682 = w4680 & w4681;
assign w4683 = (w4343 & w4360) | (w4343 & w64640) | (w4360 & w64640);
assign w4684 = ~w4679 & w4683;
assign w4685 = ~w4682 & w4684;
assign w4686 = ~w4676 & w4685;
assign w4687 = ~w4672 & w4680;
assign w4688 = w4680 & w64641;
assign w4689 = w4333 & w4652;
assign w4690 = ~w4306 & ~w4381;
assign w4691 = ~w4689 & w4690;
assign w4692 = ~w4658 & w4691;
assign w4693 = ~w4688 & ~w4692;
assign w4694 = w4358 & ~w4366;
assign w4695 = ~w4343 & ~w4694;
assign w4696 = ~w4693 & w4695;
assign w4697 = ~w4686 & ~w4696;
assign w4698 = ~w4697 & w64642;
assign w4699 = (pi0307 & w4697) | (pi0307 & w64643) | (w4697 & w64643);
assign w4700 = ~w4698 & ~w4699;
assign w4701 = ~pi3177 & pi9040;
assign w4702 = ~pi3161 & ~pi9040;
assign w4703 = ~w4701 & ~w4702;
assign w4704 = pi0269 & ~w4703;
assign w4705 = ~pi0269 & w4703;
assign w4706 = ~w4704 & ~w4705;
assign w4707 = ~pi3138 & pi9040;
assign w4708 = ~pi3146 & ~pi9040;
assign w4709 = ~w4707 & ~w4708;
assign w4710 = pi0284 & ~w4709;
assign w4711 = ~pi0284 & w4709;
assign w4712 = ~w4710 & ~w4711;
assign w4713 = ~pi3149 & pi9040;
assign w4714 = ~pi3156 & ~pi9040;
assign w4715 = ~w4713 & ~w4714;
assign w4716 = pi0274 & ~w4715;
assign w4717 = ~pi0274 & w4715;
assign w4718 = ~w4716 & ~w4717;
assign w4719 = ~w4712 & ~w4718;
assign w4720 = ~pi3140 & pi9040;
assign w4721 = ~pi3175 & ~pi9040;
assign w4722 = ~w4720 & ~w4721;
assign w4723 = pi0275 & ~w4722;
assign w4724 = ~pi0275 & w4722;
assign w4725 = ~w4723 & ~w4724;
assign w4726 = ~pi3141 & pi9040;
assign w4727 = ~pi3166 & ~pi9040;
assign w4728 = ~w4726 & ~w4727;
assign w4729 = pi0250 & ~w4728;
assign w4730 = ~pi0250 & w4728;
assign w4731 = ~w4729 & ~w4730;
assign w4732 = ~w4725 & w4731;
assign w4733 = w4719 & w4732;
assign w4734 = w4706 & ~w4733;
assign w4735 = w4725 & ~w4731;
assign w4736 = ~w4732 & ~w4735;
assign w4737 = ~w4718 & ~w4736;
assign w4738 = w4734 & w4737;
assign w4739 = w4718 & w4732;
assign w4740 = w4719 & ~w4725;
assign w4741 = ~w4739 & ~w4740;
assign w4742 = ~w4706 & ~w4741;
assign w4743 = w4718 & ~w4731;
assign w4744 = w4712 & ~w4725;
assign w4745 = w4743 & w4744;
assign w4746 = ~pi3135 & pi9040;
assign w4747 = ~pi3149 & ~pi9040;
assign w4748 = ~w4746 & ~w4747;
assign w4749 = pi0280 & ~w4748;
assign w4750 = ~pi0280 & w4748;
assign w4751 = ~w4749 & ~w4750;
assign w4752 = w4718 & w4725;
assign w4753 = ~w4731 & w4752;
assign w4754 = (~w4706 & ~w4752) | (~w4706 & w64644) | (~w4752 & w64644);
assign w4755 = ~w4712 & w4725;
assign w4756 = ~w4754 & w4755;
assign w4757 = w4706 & w4731;
assign w4758 = w4752 & w4757;
assign w4759 = ~w4745 & w4751;
assign w4760 = ~w4758 & w4759;
assign w4761 = ~w4738 & w4760;
assign w4762 = ~w4742 & ~w4756;
assign w4763 = w4761 & w4762;
assign w4764 = w4712 & w4725;
assign w4765 = ~w4718 & w4731;
assign w4766 = w4764 & w4765;
assign w4767 = w4712 & ~w4731;
assign w4768 = w4752 & w4767;
assign w4769 = ~w4751 & ~w4766;
assign w4770 = ~w4768 & w4769;
assign w4771 = w4706 & ~w4741;
assign w4772 = ~w4718 & ~w4725;
assign w4773 = w4767 & w4772;
assign w4774 = w4770 & ~w4773;
assign w4775 = ~w4771 & w4774;
assign w4776 = ~w4763 & ~w4775;
assign w4777 = w4725 & ~w4765;
assign w4778 = w4712 & ~w4777;
assign w4779 = ~w4718 & w4767;
assign w4780 = ~w4751 & ~w4779;
assign w4781 = ~w4753 & ~w4772;
assign w4782 = w4780 & w4781;
assign w4783 = ~w4778 & ~w4782;
assign w4784 = ~w4706 & ~w4732;
assign w4785 = ~w4783 & w4784;
assign w4786 = ~w4776 & ~w4785;
assign w4787 = ~pi0294 & w4786;
assign w4788 = pi0294 & ~w4786;
assign w4789 = ~w4787 & ~w4788;
assign w4790 = ~w4712 & w4731;
assign w4791 = w4772 & ~w4790;
assign w4792 = ~w4768 & ~w4791;
assign w4793 = ~w4706 & ~w4792;
assign w4794 = ~w4743 & ~w4764;
assign w4795 = w4777 & w4794;
assign w4796 = ~w4767 & ~w4790;
assign w4797 = w4706 & ~w4712;
assign w4798 = w4718 & ~w4764;
assign w4799 = ~w4797 & w4798;
assign w4800 = w4796 & w4799;
assign w4801 = ~w4725 & ~w4757;
assign w4802 = w4800 & w4801;
assign w4803 = ~w4744 & w4757;
assign w4804 = w4751 & ~w4803;
assign w4805 = ~w4795 & w4804;
assign w4806 = ~w4793 & w4805;
assign w4807 = ~w4802 & w4806;
assign w4808 = w4754 & ~w4794;
assign w4809 = w4718 & ~w4725;
assign w4810 = ~w4790 & ~w4797;
assign w4811 = ~w4765 & ~w4809;
assign w4812 = ~w4755 & ~w4811;
assign w4813 = w4706 & ~w4795;
assign w4814 = ~w4812 & w4813;
assign w4815 = (~w4751 & w4810) | (~w4751 & w64645) | (w4810 & w64645);
assign w4816 = ~w4814 & w4815;
assign w4817 = (~w4770 & w4814) | (~w4770 & w63556) | (w4814 & w63556);
assign w4818 = ~w4739 & ~w4811;
assign w4819 = ~w4712 & w4818;
assign w4820 = ~w4800 & ~w4808;
assign w4821 = ~w4819 & w4820;
assign w4822 = ~w4817 & w4821;
assign w4823 = (w4706 & ~w4798) | (w4706 & w64646) | (~w4798 & w64646);
assign w4824 = w4736 & ~w4796;
assign w4825 = w4823 & w4824;
assign w4826 = (~w4825 & w4822) | (~w4825 & w64647) | (w4822 & w64647);
assign w4827 = ~pi0316 & w4826;
assign w4828 = pi0316 & ~w4826;
assign w4829 = ~w4827 & ~w4828;
assign w4830 = w4573 & ~w4625;
assign w4831 = ~w4552 & ~w4572;
assign w4832 = (w4560 & w4830) | (w4560 & w64648) | (w4830 & w64648);
assign w4833 = w4534 & w4560;
assign w4834 = ~w4537 & ~w4627;
assign w4835 = ~w4542 & ~w4561;
assign w4836 = ~w4833 & w4835;
assign w4837 = ~w4834 & w4836;
assign w4838 = w4514 & ~w4546;
assign w4839 = ~w4539 & ~w4838;
assign w4840 = ~w4560 & ~w4839;
assign w4841 = w4544 & ~w4551;
assign w4842 = ~w4837 & w4841;
assign w4843 = ~w4840 & w4842;
assign w4844 = ~w4832 & w4843;
assign w4845 = pi0311 & w4844;
assign w4846 = ~pi0311 & ~w4844;
assign w4847 = ~w4845 & ~w4846;
assign w4848 = ~pi3131 & pi9040;
assign w4849 = ~pi3143 & ~pi9040;
assign w4850 = ~w4848 & ~w4849;
assign w4851 = pi0257 & ~w4850;
assign w4852 = ~pi0257 & w4850;
assign w4853 = ~w4851 & ~w4852;
assign w4854 = ~pi3161 & pi9040;
assign w4855 = ~pi3131 & ~pi9040;
assign w4856 = ~w4854 & ~w4855;
assign w4857 = pi0280 & ~w4856;
assign w4858 = ~pi0280 & w4856;
assign w4859 = ~w4857 & ~w4858;
assign w4860 = w4853 & ~w4859;
assign w4861 = ~pi3144 & pi9040;
assign w4862 = ~pi3170 & ~pi9040;
assign w4863 = ~w4861 & ~w4862;
assign w4864 = pi0276 & ~w4863;
assign w4865 = ~pi0276 & w4863;
assign w4866 = ~w4864 & ~w4865;
assign w4867 = ~pi3159 & pi9040;
assign w4868 = ~pi3144 & ~pi9040;
assign w4869 = ~w4867 & ~w4868;
assign w4870 = pi0274 & ~w4869;
assign w4871 = ~pi0274 & w4869;
assign w4872 = ~w4870 & ~w4871;
assign w4873 = w4866 & ~w4872;
assign w4874 = ~w4860 & ~w4873;
assign w4875 = w4859 & ~w4866;
assign w4876 = ~w4859 & w4866;
assign w4877 = ~w4875 & ~w4876;
assign w4878 = ~pi3146 & pi9040;
assign w4879 = ~pi3135 & ~pi9040;
assign w4880 = ~w4878 & ~w4879;
assign w4881 = pi0261 & ~w4880;
assign w4882 = ~pi0261 & w4880;
assign w4883 = ~w4881 & ~w4882;
assign w4884 = w4877 & ~w4883;
assign w4885 = w4874 & w4884;
assign w4886 = w4853 & w4885;
assign w4887 = ~w4875 & ~w4883;
assign w4888 = ~w4859 & w4872;
assign w4889 = ~w4866 & w4888;
assign w4890 = ~w4853 & w4876;
assign w4891 = w4860 & ~w4866;
assign w4892 = ~w4890 & ~w4891;
assign w4893 = w4853 & w4859;
assign w4894 = ~w4872 & w4893;
assign w4895 = ~w4889 & ~w4894;
assign w4896 = w4892 & w4895;
assign w4897 = ~w4887 & ~w4896;
assign w4898 = ~w4859 & ~w4866;
assign w4899 = ~w4866 & w4872;
assign w4900 = w4874 & ~w4899;
assign w4901 = w4874 & w63557;
assign w4902 = ~w4853 & ~w4872;
assign w4903 = w4898 & ~w4902;
assign w4904 = ~w4901 & ~w4903;
assign w4905 = w4896 & w4904;
assign w4906 = ~w4883 & w4905;
assign w4907 = ~pi3217 & pi9040;
assign w4908 = ~pi3138 & ~pi9040;
assign w4909 = ~w4907 & ~w4908;
assign w4910 = pi0251 & ~w4909;
assign w4911 = ~pi0251 & w4909;
assign w4912 = ~w4910 & ~w4911;
assign w4913 = (~w4912 & w4906) | (~w4912 & w64649) | (w4906 & w64649);
assign w4914 = w4875 & w4902;
assign w4915 = w4853 & w4883;
assign w4916 = ~w4914 & ~w4915;
assign w4917 = w4896 & ~w4916;
assign w4918 = (~w4902 & ~w4877) | (~w4902 & w64650) | (~w4877 & w64650);
assign w4919 = w4876 & ~w4883;
assign w4920 = ~w4876 & w4883;
assign w4921 = w4902 & ~w4919;
assign w4922 = ~w4920 & w4921;
assign w4923 = ~w4918 & ~w4922;
assign w4924 = ~w4917 & ~w4923;
assign w4925 = w4912 & ~w4924;
assign w4926 = (w4883 & ~w4892) | (w4883 & w64651) | (~w4892 & w64651);
assign w4927 = w4853 & w4872;
assign w4928 = ~w4902 & ~w4927;
assign w4929 = ~w4875 & ~w4919;
assign w4930 = ~w4853 & w4883;
assign w4931 = w4888 & w4930;
assign w4932 = (~w4931 & w4929) | (~w4931 & w64652) | (w4929 & w64652);
assign w4933 = w4926 & ~w4932;
assign w4934 = ~w4886 & ~w4933;
assign w4935 = ~w4925 & w4934;
assign w4936 = (pi0298 & ~w4935) | (pi0298 & w64653) | (~w4935 & w64653);
assign w4937 = w4935 & w64654;
assign w4938 = ~w4936 & ~w4937;
assign w4939 = w4853 & ~w4883;
assign w4940 = w4899 & w4939;
assign w4941 = ~w4893 & ~w4899;
assign w4942 = ~w4859 & ~w4872;
assign w4943 = ~w4883 & ~w4942;
assign w4944 = w4941 & w4943;
assign w4945 = ~w4872 & w4905;
assign w4946 = w4893 & w4899;
assign w4947 = w4883 & ~w4946;
assign w4948 = ~w4891 & ~w4941;
assign w4949 = w4947 & w4948;
assign w4950 = ~w4944 & ~w4949;
assign w4951 = (~w4912 & w4945) | (~w4912 & w64655) | (w4945 & w64655);
assign w4952 = ~w4900 & w4927;
assign w4953 = ~w4926 & ~w4952;
assign w4954 = w4912 & ~w4953;
assign w4955 = ~w4883 & w4912;
assign w4956 = ~w4889 & ~w4893;
assign w4957 = w4955 & ~w4956;
assign w4958 = w4873 & w4915;
assign w4959 = w4859 & w4958;
assign w4960 = ~w4940 & ~w4959;
assign w4961 = ~w4957 & w4960;
assign w4962 = ~w4954 & w4961;
assign w4963 = ~w4951 & w4962;
assign w4964 = pi0319 & ~w4963;
assign w4965 = ~pi0319 & w4963;
assign w4966 = ~w4964 & ~w4965;
assign w4967 = w4379 & w4383;
assign w4968 = w4349 & w4356;
assign w4969 = w4369 & ~w4687;
assign w4970 = ~w4968 & ~w4969;
assign w4971 = ~w4306 & ~w4970;
assign w4972 = w4306 & w4689;
assign w4973 = ~w4381 & ~w4654;
assign w4974 = ~w4671 & w4973;
assign w4975 = ~w4337 & w4974;
assign w4976 = w4343 & ~w4975;
assign w4977 = w4354 & w4681;
assign w4978 = w4306 & ~w4359;
assign w4979 = ~w4358 & ~w4364;
assign w4980 = ~w4343 & ~w4978;
assign w4981 = ~w4979 & w4980;
assign w4982 = ~w4972 & ~w4977;
assign w4983 = ~w4981 & w4982;
assign w4984 = ~w4967 & w4983;
assign w4985 = ~w4976 & w4984;
assign w4986 = (~pi0320 & ~w4985) | (~pi0320 & w64656) | (~w4985 & w64656);
assign w4987 = w4985 & w64657;
assign w4988 = ~w4986 & ~w4987;
assign w4989 = ~w4535 & ~w4547;
assign w4990 = w4546 & ~w4989;
assign w4991 = ~w4521 & ~w4575;
assign w4992 = ~w4539 & ~w4550;
assign w4993 = w4991 & w4992;
assign w4994 = ~w4990 & ~w4993;
assign w4995 = ~w4539 & w4560;
assign w4996 = ~w4576 & w4995;
assign w4997 = ~w4994 & ~w4996;
assign w4998 = ~w4534 & w4560;
assign w4999 = ~w4547 & w4998;
assign w5000 = ~w4991 & w4999;
assign w5001 = w4514 & ~w4527;
assign w5002 = ~w4570 & w4833;
assign w5003 = ~w5001 & w5002;
assign w5004 = ~w5000 & ~w5003;
assign w5005 = ~w4997 & w5004;
assign w5006 = pi0321 & ~w5005;
assign w5007 = ~pi0321 & w5005;
assign w5008 = ~w5006 & ~w5007;
assign w5009 = ~w4106 & w4134;
assign w5010 = ~w4093 & w4146;
assign w5011 = ~w4147 & ~w5009;
assign w5012 = ~w5010 & w5011;
assign w5013 = w4113 & ~w5012;
assign w5014 = ~w4120 & w5013;
assign w5015 = w4094 & ~w4106;
assign w5016 = ~w4094 & ~w4141;
assign w5017 = (w4113 & ~w5016) | (w4113 & w64658) | (~w5016 & w64658);
assign w5018 = w4106 & w4134;
assign w5019 = ~w5017 & w5018;
assign w5020 = w4113 & w4116;
assign w5021 = ~w4119 & ~w5020;
assign w5022 = ~w4100 & ~w5021;
assign w5023 = w4132 & ~w5015;
assign w5024 = ~w5022 & w5023;
assign w5025 = ~w5019 & w5024;
assign w5026 = ~w4087 & w4093;
assign w5027 = w4107 & w5026;
assign w5028 = ~w4132 & ~w5027;
assign w5029 = ~w5017 & w5028;
assign w5030 = ~w5025 & ~w5029;
assign w5031 = ~w4106 & w5010;
assign w5032 = ~w4123 & w4132;
assign w5033 = w5026 & ~w5032;
assign w5034 = ~w5031 & ~w5033;
assign w5035 = ~w4121 & w5034;
assign w5036 = ~w4113 & ~w5035;
assign w5037 = ~w5014 & ~w5036;
assign w5038 = ~w5030 & w5037;
assign w5039 = pi0305 & ~w5038;
assign w5040 = ~pi0305 & w5038;
assign w5041 = ~w5039 & ~w5040;
assign w5042 = ~w4106 & w5020;
assign w5043 = ~w4132 & ~w5042;
assign w5044 = w4093 & ~w4113;
assign w5045 = ~w4107 & ~w5018;
assign w5046 = w5044 & ~w5045;
assign w5047 = ~w4116 & ~w4147;
assign w5048 = w4100 & w4106;
assign w5049 = ~w4114 & ~w5048;
assign w5050 = ~w5047 & w5049;
assign w5051 = ~w5046 & ~w5050;
assign w5052 = ~w5013 & w5051;
assign w5053 = ~w5043 & ~w5052;
assign w5054 = w4100 & ~w4106;
assign w5055 = w5044 & w5054;
assign w5056 = w4087 & w5055;
assign w5057 = w4132 & ~w5056;
assign w5058 = ~w4144 & ~w5015;
assign w5059 = w4100 & ~w5058;
assign w5060 = ~w4093 & ~w4113;
assign w5061 = w4155 & w5060;
assign w5062 = ~w5055 & ~w5061;
assign w5063 = ~w4100 & ~w4136;
assign w5064 = w4094 & ~w4100;
assign w5065 = ~w4135 & ~w5064;
assign w5066 = w4113 & ~w5065;
assign w5067 = ~w4119 & w5062;
assign w5068 = ~w5059 & w5067;
assign w5069 = ~w5063 & ~w5066;
assign w5070 = w5068 & w5069;
assign w5071 = ~w5057 & ~w5070;
assign w5072 = ~w5053 & ~w5071;
assign w5073 = ~pi0308 & w5072;
assign w5074 = pi0308 & ~w5072;
assign w5075 = ~w5073 & ~w5074;
assign w5076 = w4752 & w4790;
assign w5077 = ~w4766 & ~w5076;
assign w5078 = ~w4737 & ~w4745;
assign w5079 = w4780 & ~w5078;
assign w5080 = w5077 & ~w5079;
assign w5081 = ~w4706 & ~w5080;
assign w5082 = w4719 & ~w4731;
assign w5083 = w4823 & ~w5082;
assign w5084 = w4754 & ~w4779;
assign w5085 = ~w5083 & ~w5084;
assign w5086 = ~w4733 & w4751;
assign w5087 = w5077 & w5086;
assign w5088 = ~w4800 & w5087;
assign w5089 = ~w5085 & w5088;
assign w5090 = ~w4816 & ~w5089;
assign w5091 = ~w5081 & ~w5090;
assign w5092 = pi0303 & w5091;
assign w5093 = ~pi0303 & ~w5091;
assign w5094 = ~w5092 & ~w5093;
assign w5095 = ~w4116 & ~w5044;
assign w5096 = w5048 & ~w5095;
assign w5097 = ~w5061 & ~w5096;
assign w5098 = ~w4132 & ~w5097;
assign w5099 = w5016 & ~w5062;
assign w5100 = ~w4134 & ~w5048;
assign w5101 = ~w4119 & w5100;
assign w5102 = ~w5032 & w5101;
assign w5103 = w4142 & w5102;
assign w5104 = ~w4117 & ~w5010;
assign w5105 = ~w5064 & w5104;
assign w5106 = ~w4113 & ~w5105;
assign w5107 = w4157 & ~w5016;
assign w5108 = ~w4124 & ~w4153;
assign w5109 = ~w5009 & w5108;
assign w5110 = ~w5107 & w5109;
assign w5111 = ~w5106 & w5110;
assign w5112 = w4132 & ~w5111;
assign w5113 = ~w4115 & ~w5099;
assign w5114 = ~w5098 & w5113;
assign w5115 = ~w5103 & w5114;
assign w5116 = ~w5112 & w5115;
assign w5117 = pi0317 & ~w5116;
assign w5118 = ~pi0317 & w5116;
assign w5119 = ~w5117 & ~w5118;
assign w5120 = w4877 & w4928;
assign w5121 = w4932 & ~w5120;
assign w5122 = ~w4912 & ~w5121;
assign w5123 = w4889 & w4954;
assign w5124 = w4901 & w4955;
assign w5125 = w4898 & w4902;
assign w5126 = ~w4912 & ~w5125;
assign w5127 = w4883 & ~w5126;
assign w5128 = w4904 & w5127;
assign w5129 = ~w4958 & ~w5124;
assign w5130 = ~w5128 & w5129;
assign w5131 = ~w5122 & w5130;
assign w5132 = ~w5123 & w5131;
assign w5133 = ~pi0313 & ~w5132;
assign w5134 = pi0313 & w5132;
assign w5135 = ~w5133 & ~w5134;
assign w5136 = w4431 & w4611;
assign w5137 = ~w4456 & ~w5136;
assign w5138 = w4424 & ~w4476;
assign w5139 = (~w4424 & ~w4445) | (~w4424 & w64659) | (~w4445 & w64659);
assign w5140 = ~w4418 & ~w4610;
assign w5141 = w4446 & ~w4451;
assign w5142 = w5139 & ~w5141;
assign w5143 = ~w5140 & w5142;
assign w5144 = ~w5138 & ~w5143;
assign w5145 = w5137 & ~w5144;
assign w5146 = w4465 & ~w5145;
assign w5147 = w4449 & ~w4454;
assign w5148 = ~w4456 & ~w4465;
assign w5149 = ~w5147 & w5148;
assign w5150 = w4607 & ~w5149;
assign w5151 = ~w4469 & ~w4476;
assign w5152 = ~w4465 & ~w5151;
assign w5153 = ~w5136 & w64660;
assign w5154 = ~w5152 & w5153;
assign w5155 = ~w5150 & ~w5154;
assign w5156 = ~w5146 & ~w5155;
assign w5157 = ~pi0314 & w5156;
assign w5158 = pi0314 & ~w5156;
assign w5159 = ~w5157 & ~w5158;
assign w5160 = ~w4883 & ~w4894;
assign w5161 = ~w4866 & ~w4872;
assign w5162 = w4860 & w5161;
assign w5163 = w4947 & ~w5162;
assign w5164 = ~w5160 & ~w5163;
assign w5165 = w4883 & w4899;
assign w5166 = ~w5165 & w64661;
assign w5167 = (w4859 & w5165) | (w4859 & w64662) | (w5165 & w64662);
assign w5168 = ~w5166 & ~w5167;
assign w5169 = w4883 & ~w5161;
assign w5170 = ~w5168 & w5169;
assign w5171 = ~w4872 & w4919;
assign w5172 = w5126 & ~w5171;
assign w5173 = ~w4885 & w5172;
assign w5174 = ~w5170 & w5173;
assign w5175 = ~w4927 & ~w4939;
assign w5176 = w5166 & ~w5175;
assign w5177 = ~w4853 & w5168;
assign w5178 = w4912 & ~w5176;
assign w5179 = ~w5177 & w5178;
assign w5180 = ~w5174 & ~w5179;
assign w5181 = ~w5164 & ~w5180;
assign w5182 = ~pi0304 & w5181;
assign w5183 = pi0304 & ~w5181;
assign w5184 = ~w5182 & ~w5183;
assign w5185 = w4718 & w4764;
assign w5186 = w4734 & ~w5185;
assign w5187 = w4751 & w4777;
assign w5188 = ~w5185 & w5187;
assign w5189 = ~w4706 & ~w4739;
assign w5190 = ~w5188 & w5189;
assign w5191 = ~w5186 & ~w5190;
assign w5192 = ~w4719 & ~w4801;
assign w5193 = w4796 & ~w5192;
assign w5194 = ~w4758 & w4770;
assign w5195 = ~w5193 & w5194;
assign w5196 = w4706 & w4818;
assign w5197 = w4751 & ~w4773;
assign w5198 = ~w5196 & w5197;
assign w5199 = ~w5195 & ~w5198;
assign w5200 = ~w5191 & ~w5199;
assign w5201 = ~pi0340 & w5200;
assign w5202 = pi0340 & ~w5200;
assign w5203 = ~w5201 & ~w5202;
assign w5204 = w4446 & w4448;
assign w5205 = w4478 & w4479;
assign w5206 = w5139 & ~w5205;
assign w5207 = (w4424 & ~w4457) | (w4424 & w64663) | (~w4457 & w64663);
assign w5208 = ~w5206 & ~w5207;
assign w5209 = w4451 & ~w4455;
assign w5210 = ~w4424 & ~w4598;
assign w5211 = ~w4611 & ~w5209;
assign w5212 = w5210 & w5211;
assign w5213 = w4465 & ~w5204;
assign w5214 = (w5213 & w5212) | (w5213 & w64664) | (w5212 & w64664);
assign w5215 = ~w5208 & w5214;
assign w5216 = w4425 & ~w4448;
assign w5217 = w4602 & w5216;
assign w5218 = ~w4608 & w5212;
assign w5219 = ~w4457 & ~w4465;
assign w5220 = ~w5217 & w5219;
assign w5221 = ~w5218 & w5220;
assign w5222 = ~w5215 & ~w5221;
assign w5223 = ~pi0318 & w5222;
assign w5224 = pi0318 & ~w5222;
assign w5225 = ~w5223 & ~w5224;
assign w5226 = ~pi3295 & pi9040;
assign w5227 = ~pi3232 & ~pi9040;
assign w5228 = ~w5226 & ~w5227;
assign w5229 = pi0336 & ~w5228;
assign w5230 = ~pi0336 & w5228;
assign w5231 = ~w5229 & ~w5230;
assign w5232 = ~pi3230 & pi9040;
assign w5233 = ~pi3250 & ~pi9040;
assign w5234 = ~w5232 & ~w5233;
assign w5235 = pi0312 & ~w5234;
assign w5236 = ~pi0312 & w5234;
assign w5237 = ~w5235 & ~w5236;
assign w5238 = ~w5231 & ~w5237;
assign w5239 = ~pi3208 & pi9040;
assign w5240 = ~pi3201 & ~pi9040;
assign w5241 = ~w5239 & ~w5240;
assign w5242 = pi0334 & ~w5241;
assign w5243 = ~pi0334 & w5241;
assign w5244 = ~w5242 & ~w5243;
assign w5245 = ~w5238 & ~w5244;
assign w5246 = ~pi3199 & pi9040;
assign w5247 = ~pi3255 & ~pi9040;
assign w5248 = ~w5246 & ~w5247;
assign w5249 = pi0341 & ~w5248;
assign w5250 = ~pi0341 & w5248;
assign w5251 = ~w5249 & ~w5250;
assign w5252 = ~w5237 & w5251;
assign w5253 = w5231 & w5252;
assign w5254 = w5244 & ~w5251;
assign w5255 = w5238 & w5254;
assign w5256 = ~w5253 & ~w5255;
assign w5257 = (w5244 & ~w5256) | (w5244 & w64665) | (~w5256 & w64665);
assign w5258 = ~w5245 & ~w5257;
assign w5259 = ~w5231 & w5244;
assign w5260 = w5237 & ~w5251;
assign w5261 = w5259 & w5260;
assign w5262 = ~pi3211 & pi9040;
assign w5263 = ~pi3333 & ~pi9040;
assign w5264 = ~w5262 & ~w5263;
assign w5265 = pi0345 & ~w5264;
assign w5266 = ~pi0345 & w5264;
assign w5267 = ~w5265 & ~w5266;
assign w5268 = ~w5261 & w5267;
assign w5269 = ~w5258 & w5268;
assign w5270 = ~w5244 & w5251;
assign w5271 = ~w5254 & ~w5270;
assign w5272 = w5231 & w5271;
assign w5273 = ~w5267 & ~w5272;
assign w5274 = ~w5269 & ~w5273;
assign w5275 = w5251 & w5267;
assign w5276 = w5231 & w5237;
assign w5277 = ~w5244 & w5276;
assign w5278 = ~w5259 & ~w5277;
assign w5279 = w5275 & ~w5278;
assign w5280 = ~w5231 & ~w5244;
assign w5281 = w5237 & w5251;
assign w5282 = w5280 & w5281;
assign w5283 = ~w5251 & w5276;
assign w5284 = ~w5282 & ~w5283;
assign w5285 = ~w5267 & ~w5284;
assign w5286 = w5238 & ~w5251;
assign w5287 = ~w5244 & w5286;
assign w5288 = ~pi3232 & pi9040;
assign w5289 = ~pi3322 & ~pi9040;
assign w5290 = ~w5288 & ~w5289;
assign w5291 = pi0335 & ~w5290;
assign w5292 = ~pi0335 & w5290;
assign w5293 = ~w5291 & ~w5292;
assign w5294 = ~w5261 & w5293;
assign w5295 = ~w5287 & w5294;
assign w5296 = ~w5279 & ~w5285;
assign w5297 = w5295 & w5296;
assign w5298 = ~w5231 & w5267;
assign w5299 = w5237 & ~w5298;
assign w5300 = w5271 & w5299;
assign w5301 = ~w5256 & ~w5267;
assign w5302 = ~w5238 & ~w5298;
assign w5303 = w5270 & ~w5302;
assign w5304 = ~w5293 & ~w5300;
assign w5305 = ~w5303 & w5304;
assign w5306 = ~w5301 & w5305;
assign w5307 = ~w5297 & ~w5306;
assign w5308 = ~w5274 & ~w5307;
assign w5309 = ~pi0359 & w5308;
assign w5310 = pi0359 & ~w5308;
assign w5311 = ~w5309 & ~w5310;
assign w5312 = ~pi3255 & pi9040;
assign w5313 = ~pi3345 & ~pi9040;
assign w5314 = ~w5312 & ~w5313;
assign w5315 = pi0350 & ~w5314;
assign w5316 = ~pi0350 & w5314;
assign w5317 = ~w5315 & ~w5316;
assign w5318 = ~pi3258 & pi9040;
assign w5319 = ~pi3219 & ~pi9040;
assign w5320 = ~w5318 & ~w5319;
assign w5321 = pi0347 & ~w5320;
assign w5322 = ~pi0347 & w5320;
assign w5323 = ~w5321 & ~w5322;
assign w5324 = ~pi3215 & pi9040;
assign w5325 = ~pi3214 & ~pi9040;
assign w5326 = ~w5324 & ~w5325;
assign w5327 = pi0335 & ~w5326;
assign w5328 = ~pi0335 & w5326;
assign w5329 = ~w5327 & ~w5328;
assign w5330 = w5323 & w5329;
assign w5331 = ~pi3345 & pi9040;
assign w5332 = ~pi3252 & ~pi9040;
assign w5333 = ~w5331 & ~w5332;
assign w5334 = pi0312 & ~w5333;
assign w5335 = ~pi0312 & w5333;
assign w5336 = ~w5334 & ~w5335;
assign w5337 = w5330 & ~w5336;
assign w5338 = ~pi3218 & pi9040;
assign w5339 = ~pi3282 & ~pi9040;
assign w5340 = ~w5338 & ~w5339;
assign w5341 = pi0342 & ~w5340;
assign w5342 = ~pi0342 & w5340;
assign w5343 = ~w5341 & ~w5342;
assign w5344 = w5337 & ~w5343;
assign w5345 = ~w5329 & ~w5336;
assign w5346 = w5343 & w5345;
assign w5347 = ~w5344 & ~w5346;
assign w5348 = ~pi3213 & pi9040;
assign w5349 = ~pi3295 & ~pi9040;
assign w5350 = ~w5348 & ~w5349;
assign w5351 = pi0325 & ~w5350;
assign w5352 = ~pi0325 & w5350;
assign w5353 = ~w5351 & ~w5352;
assign w5354 = ~w5347 & w5353;
assign w5355 = w5336 & ~w5343;
assign w5356 = ~w5323 & w5329;
assign w5357 = w5355 & w5356;
assign w5358 = w5353 & ~w5357;
assign w5359 = w5323 & ~w5329;
assign w5360 = ~w5356 & ~w5359;
assign w5361 = w5323 & w5343;
assign w5362 = ~w5360 & ~w5361;
assign w5363 = ~w5358 & w5362;
assign w5364 = w5336 & w5343;
assign w5365 = ~w5330 & w5353;
assign w5366 = w5364 & ~w5365;
assign w5367 = ~w5317 & ~w5366;
assign w5368 = ~w5363 & w5367;
assign w5369 = ~w5354 & w5368;
assign w5370 = ~w5336 & ~w5353;
assign w5371 = w5360 & w5370;
assign w5372 = ~w5355 & ~w5356;
assign w5373 = w5358 & ~w5372;
assign w5374 = w5359 & w5364;
assign w5375 = w5317 & ~w5374;
assign w5376 = ~w5371 & w5375;
assign w5377 = ~w5373 & w5376;
assign w5378 = ~w5369 & ~w5377;
assign w5379 = ~w5353 & ~w5357;
assign w5380 = w5336 & w5359;
assign w5381 = ~w5323 & w5345;
assign w5382 = ~w5380 & ~w5381;
assign w5383 = ~w5343 & ~w5382;
assign w5384 = ~w5336 & w5343;
assign w5385 = ~w5360 & w5384;
assign w5386 = w5353 & ~w5385;
assign w5387 = ~w5383 & w5386;
assign w5388 = ~w5379 & ~w5387;
assign w5389 = ~w5378 & ~w5388;
assign w5390 = pi0352 & w5389;
assign w5391 = ~pi0352 & ~w5389;
assign w5392 = ~w5390 & ~w5391;
assign w5393 = ~w5277 & ~w5286;
assign w5394 = (w5293 & w5393) | (w5293 & w5959) | (w5393 & w5959);
assign w5395 = ~w5295 & ~w5394;
assign w5396 = ~w5261 & ~w5275;
assign w5397 = ~w5298 & ~w5396;
assign w5398 = ~w5244 & w5284;
assign w5399 = ~w5257 & ~w5398;
assign w5400 = ~w5395 & ~w5397;
assign w5401 = ~w5399 & w5400;
assign w5402 = ~w5238 & ~w5276;
assign w5403 = ~w5267 & ~w5402;
assign w5404 = w5259 & w5281;
assign w5405 = w5244 & w5251;
assign w5406 = ~w5267 & w5405;
assign w5407 = ~w5231 & ~w5271;
assign w5408 = ~w5252 & ~w5254;
assign w5409 = ~w5280 & w5408;
assign w5410 = ~w5407 & ~w5409;
assign w5411 = ~w5237 & ~w5410;
assign w5412 = w5231 & w5244;
assign w5413 = ~w5298 & ~w5412;
assign w5414 = w5260 & ~w5413;
assign w5415 = ~w5293 & ~w5404;
assign w5416 = ~w5406 & w5415;
assign w5417 = ~w5403 & ~w5414;
assign w5418 = w5416 & w5417;
assign w5419 = ~w5411 & w5418;
assign w5420 = ~w5401 & ~w5419;
assign w5421 = ~pi0355 & w5420;
assign w5422 = pi0355 & ~w5420;
assign w5423 = ~w5421 & ~w5422;
assign w5424 = ~pi3298 & pi9040;
assign w5425 = ~pi3239 & ~pi9040;
assign w5426 = ~w5424 & ~w5425;
assign w5427 = pi0348 & ~w5426;
assign w5428 = ~pi0348 & w5426;
assign w5429 = ~w5427 & ~w5428;
assign w5430 = ~pi3222 & pi9040;
assign w5431 = ~pi3207 & ~pi9040;
assign w5432 = ~w5430 & ~w5431;
assign w5433 = pi0342 & ~w5432;
assign w5434 = ~pi0342 & w5432;
assign w5435 = ~w5433 & ~w5434;
assign w5436 = w5429 & ~w5435;
assign w5437 = ~pi3226 & pi9040;
assign w5438 = ~pi3257 & ~pi9040;
assign w5439 = ~w5437 & ~w5438;
assign w5440 = pi0302 & ~w5439;
assign w5441 = ~pi0302 & w5439;
assign w5442 = ~w5440 & ~w5441;
assign w5443 = ~pi3307 & pi9040;
assign w5444 = ~pi3234 & ~pi9040;
assign w5445 = ~w5443 & ~w5444;
assign w5446 = pi0350 & ~w5445;
assign w5447 = ~pi0350 & w5445;
assign w5448 = ~w5446 & ~w5447;
assign w5449 = ~w5442 & ~w5448;
assign w5450 = ~pi3212 & pi9040;
assign w5451 = ~pi3298 & ~pi9040;
assign w5452 = ~w5450 & ~w5451;
assign w5453 = pi0343 & ~w5452;
assign w5454 = ~pi0343 & w5452;
assign w5455 = ~w5453 & ~w5454;
assign w5456 = w5449 & w5455;
assign w5457 = w5436 & w5456;
assign w5458 = w5435 & w5455;
assign w5459 = ~w5435 & ~w5455;
assign w5460 = ~w5458 & ~w5459;
assign w5461 = w5442 & w5448;
assign w5462 = ~w5435 & w5442;
assign w5463 = w5435 & ~w5442;
assign w5464 = ~w5462 & ~w5463;
assign w5465 = ~w5461 & w5464;
assign w5466 = ~w5429 & ~w5465;
assign w5467 = w5460 & ~w5461;
assign w5468 = w5466 & w5467;
assign w5469 = ~w5429 & w5448;
assign w5470 = w5442 & w5458;
assign w5471 = w5469 & w5470;
assign w5472 = w5448 & ~w5455;
assign w5473 = w5436 & w5472;
assign w5474 = ~w5471 & ~w5473;
assign w5475 = ~pi3229 & pi9040;
assign w5476 = ~pi3307 & ~pi9040;
assign w5477 = ~w5475 & ~w5476;
assign w5478 = pi0329 & ~w5477;
assign w5479 = ~pi0329 & w5477;
assign w5480 = ~w5478 & ~w5479;
assign w5481 = w5435 & w5469;
assign w5482 = w5480 & ~w5481;
assign w5483 = w5429 & w5442;
assign w5484 = w5448 & w5464;
assign w5485 = (~w5483 & ~w5464) | (~w5483 & w64666) | (~w5464 & w64666);
assign w5486 = ~w5455 & ~w5461;
assign w5487 = ~w5485 & w5486;
assign w5488 = ~w5456 & ~w5462;
assign w5489 = ~w5429 & w5435;
assign w5490 = ~w5469 & ~w5489;
assign w5491 = ~w5488 & w5490;
assign w5492 = ~w5487 & ~w5491;
assign w5493 = w5482 & w5492;
assign w5494 = w5429 & w5435;
assign w5495 = ~w5448 & ~w5464;
assign w5496 = ~w5484 & ~w5495;
assign w5497 = w5455 & w5496;
assign w5498 = w5496 & w64667;
assign w5499 = w5488 & w5495;
assign w5500 = w5442 & w5472;
assign w5501 = ~w5429 & ~w5472;
assign w5502 = ~w5458 & w5501;
assign w5503 = w5488 & w5502;
assign w5504 = (~w5480 & ~w5500) | (~w5480 & w64668) | (~w5500 & w64668);
assign w5505 = ~w5499 & w5504;
assign w5506 = ~w5503 & w5505;
assign w5507 = ~w5498 & w5506;
assign w5508 = ~w5457 & w5474;
assign w5509 = ~w5468 & w5508;
assign w5510 = (w5509 & w5507) | (w5509 & w64669) | (w5507 & w64669);
assign w5511 = pi0373 & ~w5510;
assign w5512 = ~pi0373 & w5510;
assign w5513 = ~w5511 & ~w5512;
assign w5514 = ~w5492 & w5494;
assign w5515 = w5429 & w5484;
assign w5516 = ~w5449 & ~w5461;
assign w5517 = ~w5464 & w5516;
assign w5518 = w5455 & w5517;
assign w5519 = w5435 & ~w5486;
assign w5520 = ~w5429 & ~w5516;
assign w5521 = ~w5519 & w5520;
assign w5522 = ~w5480 & ~w5515;
assign w5523 = ~w5518 & ~w5521;
assign w5524 = w5522 & w5523;
assign w5525 = w5463 & w5472;
assign w5526 = ~w5448 & ~w5459;
assign w5527 = w5462 & w5472;
assign w5528 = ~w5526 & ~w5527;
assign w5529 = w5429 & ~w5528;
assign w5530 = w5501 & ~w5526;
assign w5531 = ~w5470 & w5480;
assign w5532 = ~w5525 & w5531;
assign w5533 = ~w5530 & w5532;
assign w5534 = ~w5529 & w5533;
assign w5535 = ~w5524 & ~w5534;
assign w5536 = ~w5514 & ~w5535;
assign w5537 = ~pi0374 & w5536;
assign w5538 = pi0374 & ~w5536;
assign w5539 = ~w5537 & ~w5538;
assign w5540 = ~pi3294 & pi9040;
assign w5541 = ~pi3229 & ~pi9040;
assign w5542 = ~w5540 & ~w5541;
assign w5543 = pi0323 & ~w5542;
assign w5544 = ~pi0323 & w5542;
assign w5545 = ~w5543 & ~w5544;
assign w5546 = ~pi3234 & pi9040;
assign w5547 = ~pi3263 & ~pi9040;
assign w5548 = ~w5546 & ~w5547;
assign w5549 = pi0331 & ~w5548;
assign w5550 = ~pi0331 & w5548;
assign w5551 = ~w5549 & ~w5550;
assign w5552 = w5545 & w5551;
assign w5553 = ~w5545 & ~w5551;
assign w5554 = ~w5552 & ~w5553;
assign w5555 = ~pi3207 & pi9040;
assign w5556 = ~pi3206 & ~pi9040;
assign w5557 = ~w5555 & ~w5556;
assign w5558 = pi0328 & ~w5557;
assign w5559 = ~pi0328 & w5557;
assign w5560 = ~w5558 & ~w5559;
assign w5561 = ~w5554 & ~w5560;
assign w5562 = ~pi3200 & pi9040;
assign w5563 = ~pi3292 & ~pi9040;
assign w5564 = ~w5562 & ~w5563;
assign w5565 = pi0344 & ~w5564;
assign w5566 = ~pi0344 & w5564;
assign w5567 = ~w5565 & ~w5566;
assign w5568 = ~pi3292 & pi9040;
assign w5569 = ~pi3226 & ~pi9040;
assign w5570 = ~w5568 & ~w5569;
assign w5571 = pi0332 & ~w5570;
assign w5572 = ~pi0332 & w5570;
assign w5573 = ~w5571 & ~w5572;
assign w5574 = ~w5567 & w5573;
assign w5575 = w5561 & w5574;
assign w5576 = ~pi3202 & pi9040;
assign w5577 = ~pi3210 & ~pi9040;
assign w5578 = ~w5576 & ~w5577;
assign w5579 = pi0346 & ~w5578;
assign w5580 = ~pi0346 & w5578;
assign w5581 = ~w5579 & ~w5580;
assign w5582 = ~w5552 & ~w5560;
assign w5583 = w5560 & w5567;
assign w5584 = ~w5573 & ~w5583;
assign w5585 = ~w5582 & w5584;
assign w5586 = w5567 & w5573;
assign w5587 = w5545 & w5567;
assign w5588 = ~w5545 & ~w5567;
assign w5589 = ~w5587 & ~w5588;
assign w5590 = ~w5551 & w5589;
assign w5591 = ~w5545 & w5560;
assign w5592 = w5545 & ~w5560;
assign w5593 = ~w5591 & ~w5592;
assign w5594 = w5573 & ~w5589;
assign w5595 = ~w5593 & w5594;
assign w5596 = ~w5590 & ~w5595;
assign w5597 = ~w5595 & w64670;
assign w5598 = ~w5551 & ~w5567;
assign w5599 = ~w5567 & ~w5573;
assign w5600 = ~w5545 & w5551;
assign w5601 = ~w5599 & w5600;
assign w5602 = ~w5598 & ~w5601;
assign w5603 = w5593 & ~w5602;
assign w5604 = ~w5585 & ~w5603;
assign w5605 = ~w5597 & w5604;
assign w5606 = ~w5581 & ~w5605;
assign w5607 = ~w5554 & w5583;
assign w5608 = ~w5560 & ~w5573;
assign w5609 = w5551 & ~w5589;
assign w5610 = ~w5589 & w64671;
assign w5611 = ~w5567 & w5610;
assign w5612 = ~w5607 & ~w5611;
assign w5613 = w5581 & ~w5612;
assign w5614 = ~w5551 & w5567;
assign w5615 = ~w5593 & w5614;
assign w5616 = (~w5581 & w5593) | (~w5581 & w64672) | (w5593 & w64672);
assign w5617 = w5573 & w5589;
assign w5618 = ~w5616 & ~w5617;
assign w5619 = (~w5575 & w5596) | (~w5575 & w64673) | (w5596 & w64673);
assign w5620 = ~w5613 & w5619;
assign w5621 = ~w5606 & w5620;
assign w5622 = ~pi0361 & ~w5621;
assign w5623 = pi0361 & w5621;
assign w5624 = ~w5622 & ~w5623;
assign w5625 = ~w5545 & ~w5560;
assign w5626 = w5553 & w5585;
assign w5627 = w5561 & w5567;
assign w5628 = w5560 & w5601;
assign w5629 = w5560 & ~w5573;
assign w5630 = w5552 & w5629;
assign w5631 = w5574 & w5625;
assign w5632 = ~w5630 & ~w5631;
assign w5633 = ~w5628 & w5632;
assign w5634 = ~w5626 & w5633;
assign w5635 = ~w5627 & w5634;
assign w5636 = w5634 & w63320;
assign w5637 = ~w5551 & w5560;
assign w5638 = w5545 & w5574;
assign w5639 = ~w5637 & w5638;
assign w5640 = ~w5551 & ~w5591;
assign w5641 = w5589 & ~w5629;
assign w5642 = w5640 & ~w5641;
assign w5643 = w5560 & w5573;
assign w5644 = w5553 & w5643;
assign w5645 = ~w5639 & ~w5644;
assign w5646 = ~w5642 & w5645;
assign w5647 = (~w5581 & w5636) | (~w5581 & w63558) | (w5636 & w63558);
assign w5648 = w5561 & ~w5581;
assign w5649 = (w5561 & w64674) | (w5561 & w64675) | (w64674 & w64675);
assign w5650 = w5586 & ~w5649;
assign w5651 = w5637 & w5638;
assign w5652 = ~w5589 & w63560;
assign w5653 = w5545 & ~w5614;
assign w5654 = w5608 & w5653;
assign w5655 = ~w5651 & ~w5654;
assign w5656 = ~w5652 & w5655;
assign w5657 = (w5581 & ~w5656) | (w5581 & w63561) | (~w5656 & w63561);
assign w5658 = w5551 & ~w5560;
assign w5659 = (~w5652 & ~w5634) | (~w5652 & w63353) | (~w5634 & w63353);
assign w5660 = ~w5573 & ~w5658;
assign w5661 = ~w5659 & w5660;
assign w5662 = ~w5650 & ~w5657;
assign w5663 = ~w5647 & w5662;
assign w5664 = w5663 & w64676;
assign w5665 = (~pi0367 & ~w5663) | (~pi0367 & w64677) | (~w5663 & w64677);
assign w5666 = ~w5664 & ~w5665;
assign w5667 = ~pi3197 & pi9040;
assign w5668 = ~pi3213 & ~pi9040;
assign w5669 = ~w5667 & ~w5668;
assign w5670 = pi0322 & ~w5669;
assign w5671 = ~pi0322 & w5669;
assign w5672 = ~w5670 & ~w5671;
assign w5673 = ~pi3282 & pi9040;
assign w5674 = ~pi3209 & ~pi9040;
assign w5675 = ~w5673 & ~w5674;
assign w5676 = pi0337 & ~w5675;
assign w5677 = ~pi0337 & w5675;
assign w5678 = ~w5676 & ~w5677;
assign w5679 = ~w5672 & ~w5678;
assign w5680 = ~pi3254 & pi9040;
assign w5681 = ~pi3205 & ~pi9040;
assign w5682 = ~w5680 & ~w5681;
assign w5683 = pi0336 & ~w5682;
assign w5684 = ~pi0336 & w5682;
assign w5685 = ~w5683 & ~w5684;
assign w5686 = ~pi3209 & pi9040;
assign w5687 = ~pi3256 & ~pi9040;
assign w5688 = ~w5686 & ~w5687;
assign w5689 = pi0326 & ~w5688;
assign w5690 = ~pi0326 & w5688;
assign w5691 = ~w5689 & ~w5690;
assign w5692 = ~w5685 & ~w5691;
assign w5693 = ~pi3385 & pi9040;
assign w5694 = ~pi3230 & ~pi9040;
assign w5695 = ~w5693 & ~w5694;
assign w5696 = pi0333 & ~w5695;
assign w5697 = ~pi0333 & w5695;
assign w5698 = ~w5696 & ~w5697;
assign w5699 = w5692 & ~w5698;
assign w5700 = w5679 & w5699;
assign w5701 = ~w5679 & ~w5685;
assign w5702 = ~w5685 & w5691;
assign w5703 = w5691 & ~w5698;
assign w5704 = w5672 & w5703;
assign w5705 = ~w5702 & ~w5704;
assign w5706 = ~w5701 & ~w5705;
assign w5707 = ~w5691 & ~w5698;
assign w5708 = w5685 & ~w5707;
assign w5709 = ~w5672 & w5698;
assign w5710 = w5678 & w5685;
assign w5711 = ~w5709 & ~w5710;
assign w5712 = ~w5708 & ~w5711;
assign w5713 = ~w5672 & ~w5691;
assign w5714 = w5678 & ~w5713;
assign w5715 = ~w5704 & w5714;
assign w5716 = ~w5712 & w5715;
assign w5717 = w5672 & w5698;
assign w5718 = ~w5691 & w5717;
assign w5719 = w5691 & w5709;
assign w5720 = ~w5718 & ~w5719;
assign w5721 = ~w5678 & ~w5720;
assign w5722 = (w5678 & ~w5717) | (w5678 & w63354) | (~w5717 & w63354);
assign w5723 = ~w5698 & w5702;
assign w5724 = w5702 & w63562;
assign w5725 = w5691 & w5698;
assign w5726 = w5685 & w5725;
assign w5727 = w5722 & ~w5726;
assign w5728 = ~w5724 & w5727;
assign w5729 = ~w5721 & ~w5728;
assign w5730 = (~w5706 & w5729) | (~w5706 & w63563) | (w5729 & w63563);
assign w5731 = ~pi3205 & pi9040;
assign w5732 = ~pi3215 & ~pi9040;
assign w5733 = ~w5731 & ~w5732;
assign w5734 = pi0341 & ~w5733;
assign w5735 = ~pi0341 & w5733;
assign w5736 = ~w5734 & ~w5735;
assign w5737 = ~w5730 & ~w5736;
assign w5738 = ~w5723 & ~w5726;
assign w5739 = w5672 & ~w5698;
assign w5740 = w5692 & ~w5709;
assign w5741 = ~w5739 & w5740;
assign w5742 = w5738 & ~w5741;
assign w5743 = w5672 & w5685;
assign w5744 = w5707 & ~w5743;
assign w5745 = w5742 & w5744;
assign w5746 = ~w5706 & ~w5745;
assign w5747 = (w5712 & w5745) | (w5712 & w63564) | (w5745 & w63564);
assign w5748 = w5692 & w5709;
assign w5749 = w5691 & w5743;
assign w5750 = ~w5748 & ~w5749;
assign w5751 = w5678 & ~w5750;
assign w5752 = (~w5751 & ~w5729) | (~w5751 & w64678) | (~w5729 & w64678);
assign w5753 = ~w5672 & w5708;
assign w5754 = w5685 & w5691;
assign w5755 = w5672 & ~w5754;
assign w5756 = ~w5678 & ~w5755;
assign w5757 = ~w5753 & w5756;
assign w5758 = ~w5752 & ~w5757;
assign w5759 = ~w5700 & ~w5747;
assign w5760 = ~w5737 & w5759;
assign w5761 = (pi0360 & ~w5760) | (pi0360 & w64679) | (~w5760 & w64679);
assign w5762 = w5760 & w64680;
assign w5763 = ~w5761 & ~w5762;
assign w5764 = ~w5678 & ~w5736;
assign w5765 = w5702 & w5717;
assign w5766 = ~w5748 & ~w5765;
assign w5767 = ~w5753 & w5766;
assign w5768 = w5764 & ~w5767;
assign w5769 = ~w5678 & ~w5740;
assign w5770 = ~w5749 & w5769;
assign w5771 = w5685 & ~w5691;
assign w5772 = w5698 & w5771;
assign w5773 = w5678 & ~w5772;
assign w5774 = w5766 & w5773;
assign w5775 = ~w5770 & ~w5774;
assign w5776 = (w5736 & ~w5746) | (w5736 & w64681) | (~w5746 & w64681);
assign w5777 = w5709 & w5710;
assign w5778 = w5678 & ~w5736;
assign w5779 = ~w5742 & w5778;
assign w5780 = ~w5736 & w5743;
assign w5781 = w5707 & w5780;
assign w5782 = ~w5724 & ~w5777;
assign w5783 = ~w5781 & w5782;
assign w5784 = ~w5768 & w5783;
assign w5785 = ~w5779 & w5784;
assign w5786 = ~w5776 & w5785;
assign w5787 = pi0354 & ~w5786;
assign w5788 = ~pi0354 & w5786;
assign w5789 = ~w5787 & ~w5788;
assign w5790 = ~pi3290 & pi9040;
assign w5791 = ~pi3202 & ~pi9040;
assign w5792 = ~w5790 & ~w5791;
assign w5793 = pi0302 & ~w5792;
assign w5794 = ~pi0302 & w5792;
assign w5795 = ~w5793 & ~w5794;
assign w5796 = ~pi3221 & pi9040;
assign w5797 = ~pi3203 & ~pi9040;
assign w5798 = ~w5796 & ~w5797;
assign w5799 = pi0349 & ~w5798;
assign w5800 = ~pi0349 & w5798;
assign w5801 = ~w5799 & ~w5800;
assign w5802 = ~w5795 & w5801;
assign w5803 = w5795 & ~w5801;
assign w5804 = ~w5802 & ~w5803;
assign w5805 = ~pi3238 & pi9040;
assign w5806 = ~pi3294 & ~pi9040;
assign w5807 = ~w5805 & ~w5806;
assign w5808 = pi0329 & ~w5807;
assign w5809 = ~pi0329 & w5807;
assign w5810 = ~w5808 & ~w5809;
assign w5811 = w5801 & w5810;
assign w5812 = ~w5804 & ~w5811;
assign w5813 = ~pi3206 & pi9040;
assign w5814 = ~pi3290 & ~pi9040;
assign w5815 = ~w5813 & ~w5814;
assign w5816 = pi0338 & ~w5815;
assign w5817 = ~pi0338 & w5815;
assign w5818 = ~w5816 & ~w5817;
assign w5819 = w5812 & ~w5818;
assign w5820 = w5810 & w5818;
assign w5821 = ~w5802 & w5820;
assign w5822 = w5801 & ~w5810;
assign w5823 = ~w5795 & w5822;
assign w5824 = ~w5821 & ~w5823;
assign w5825 = ~pi3204 & pi9040;
assign w5826 = ~pi3223 & ~pi9040;
assign w5827 = ~w5825 & ~w5826;
assign w5828 = pi0339 & ~w5827;
assign w5829 = ~pi0339 & w5827;
assign w5830 = ~w5828 & ~w5829;
assign w5831 = ~w5824 & ~w5830;
assign w5832 = ~w5795 & w5818;
assign w5833 = w5795 & ~w5818;
assign w5834 = ~w5818 & w5830;
assign w5835 = ~w5833 & ~w5834;
assign w5836 = w5801 & ~w5832;
assign w5837 = w5835 & w5836;
assign w5838 = ~w5820 & w5837;
assign w5839 = ~w5831 & ~w5838;
assign w5840 = ~pi3216 & pi9040;
assign w5841 = ~pi3204 & ~pi9040;
assign w5842 = ~w5840 & ~w5841;
assign w5843 = pi0330 & ~w5842;
assign w5844 = ~pi0330 & w5842;
assign w5845 = ~w5843 & ~w5844;
assign w5846 = w5811 & w5832;
assign w5847 = ~w5845 & ~w5846;
assign w5848 = ~w5822 & w5830;
assign w5849 = w5810 & ~w5818;
assign w5850 = ~w5804 & w5849;
assign w5851 = ~w5803 & ~w5849;
assign w5852 = ~w5850 & ~w5851;
assign w5853 = (w5848 & w5850) | (w5848 & w63565) | (w5850 & w63565);
assign w5854 = (~w5845 & w5835) | (~w5845 & w64682) | (w5835 & w64682);
assign w5855 = ~w5853 & w5854;
assign w5856 = (~w5847 & w5853) | (~w5847 & w64683) | (w5853 & w64683);
assign w5857 = ~w5819 & w5839;
assign w5858 = ~w5856 & w5857;
assign w5859 = w5818 & ~w5830;
assign w5860 = w5839 & w5859;
assign w5861 = ~w5810 & w5818;
assign w5862 = w5830 & ~w5861;
assign w5863 = w5795 & w5862;
assign w5864 = w5811 & w5833;
assign w5865 = w5845 & ~w5864;
assign w5866 = ~w5795 & ~w5801;
assign w5867 = ~w5810 & w5830;
assign w5868 = ~w5820 & w5866;
assign w5869 = ~w5867 & w5868;
assign w5870 = ~w5863 & w5865;
assign w5871 = ~w5869 & w5870;
assign w5872 = ~w5860 & w5871;
assign w5873 = ~w5858 & ~w5872;
assign w5874 = ~w5810 & ~w5830;
assign w5875 = w5837 & w5874;
assign w5876 = ~w5801 & w5818;
assign w5877 = ~w5849 & ~w5876;
assign w5878 = w5830 & ~w5877;
assign w5879 = w5861 & w5866;
assign w5880 = ~w5833 & ~w5879;
assign w5881 = w5878 & ~w5880;
assign w5882 = ~w5875 & ~w5881;
assign w5883 = (pi0364 & w5873) | (pi0364 & w64684) | (w5873 & w64684);
assign w5884 = ~w5873 & w64685;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = w5429 & w5464;
assign w5887 = ~w5527 & ~w5886;
assign w5888 = ~w5461 & w5501;
assign w5889 = ~w5496 & w5888;
assign w5890 = (w5480 & w5887) | (w5480 & w63566) | (w5887 & w63566);
assign w5891 = ~w5889 & w5890;
assign w5892 = ~w5498 & w5891;
assign w5893 = ~w5460 & w5464;
assign w5894 = w5461 & w5501;
assign w5895 = ~w5458 & ~w5495;
assign w5896 = w5529 & ~w5895;
assign w5897 = ~w5480 & ~w5481;
assign w5898 = ~w5893 & w5897;
assign w5899 = ~w5894 & w5898;
assign w5900 = ~w5896 & w5899;
assign w5901 = ~w5892 & ~w5900;
assign w5902 = ~w5429 & ~w5455;
assign w5903 = ~w5517 & w5902;
assign w5904 = w5474 & ~w5902;
assign w5905 = ~w5499 & w5904;
assign w5906 = ~w5903 & ~w5905;
assign w5907 = (pi0381 & w5901) | (pi0381 & w64686) | (w5901 & w64686);
assign w5908 = ~w5901 & w64687;
assign w5909 = ~w5907 & ~w5908;
assign w5910 = w5567 & ~w5573;
assign w5911 = ~w5592 & w5910;
assign w5912 = ~w5654 & ~w5911;
assign w5913 = w5640 & ~w5912;
assign w5914 = w5581 & ~w5635;
assign w5915 = w5560 & ~w5600;
assign w5916 = w5599 & ~w5915;
assign w5917 = w5551 & w5586;
assign w5918 = ~w5591 & w5917;
assign w5919 = ~w5916 & ~w5918;
assign w5920 = ~w5581 & ~w5919;
assign w5921 = ~w5615 & ~w5653;
assign w5922 = w5581 & ~w5643;
assign w5923 = ~w5921 & ~w5922;
assign w5924 = ~w5596 & w5923;
assign w5925 = ~w5913 & ~w5920;
assign w5926 = ~w5924 & w5925;
assign w5927 = ~w5914 & w5926;
assign w5928 = pi0357 & ~w5927;
assign w5929 = ~pi0357 & w5927;
assign w5930 = ~w5928 & ~w5929;
assign w5931 = w5803 & w5820;
assign w5932 = ~w5879 & ~w5931;
assign w5933 = ~w5802 & ~w5832;
assign w5934 = w5810 & w5933;
assign w5935 = ~w5823 & ~w5934;
assign w5936 = ~w5845 & ~w5935;
assign w5937 = w5822 & w5832;
assign w5938 = w5932 & ~w5937;
assign w5939 = ~w5936 & w5938;
assign w5940 = ~w5830 & ~w5939;
assign w5941 = ~w5802 & ~w5876;
assign w5942 = w5874 & w5941;
assign w5943 = w5878 & w5932;
assign w5944 = w5795 & ~w5830;
assign w5945 = w5811 & ~w5944;
assign w5946 = ~w5832 & w5945;
assign w5947 = w5845 & ~w5937;
assign w5948 = ~w5942 & w5947;
assign w5949 = ~w5946 & w5948;
assign w5950 = ~w5943 & w5949;
assign w5951 = w5867 & w5941;
assign w5952 = w5847 & w5932;
assign w5953 = ~w5951 & w5952;
assign w5954 = ~w5950 & ~w5953;
assign w5955 = ~w5940 & ~w5954;
assign w5956 = ~pi0358 & w5955;
assign w5957 = pi0358 & ~w5955;
assign w5958 = ~w5956 & ~w5957;
assign w5959 = ~w5267 & w5293;
assign w5960 = ~w5283 & w5959;
assign w5961 = ~w5410 & w5960;
assign w5962 = ~w5252 & ~w5260;
assign w5963 = w5245 & w5962;
assign w5964 = ~w5255 & ~w5959;
assign w5965 = ~w5963 & w5964;
assign w5966 = ~w5961 & ~w5965;
assign w5967 = w5267 & ~w5293;
assign w5968 = w5412 & ~w5962;
assign w5969 = ~w5404 & ~w5967;
assign w5970 = ~w5968 & w5969;
assign w5971 = ~w5966 & w5970;
assign w5972 = w5281 & w5412;
assign w5973 = ~w5254 & w5962;
assign w5974 = ~w5968 & ~w5973;
assign w5975 = w5967 & ~w5972;
assign w5976 = ~w5974 & w5975;
assign w5977 = ~w5971 & ~w5976;
assign w5978 = ~pi0385 & w5977;
assign w5979 = pi0385 & ~w5977;
assign w5980 = ~w5978 & ~w5979;
assign w5981 = w5725 & w5780;
assign w5982 = ~w5679 & ~w5713;
assign w5983 = ~w5710 & ~w5754;
assign w5984 = ~w5982 & ~w5983;
assign w5985 = w5703 & w5984;
assign w5986 = ~w5699 & ~w5772;
assign w5987 = w5764 & ~w5986;
assign w5988 = ~w5707 & ~w5771;
assign w5989 = w5778 & w5988;
assign w5990 = ~w5719 & w5989;
assign w5991 = ~w5736 & ~w5747;
assign w5992 = ~w5722 & ~w5771;
assign w5993 = ~w5720 & ~w5992;
assign w5994 = ~w5678 & w5703;
assign w5995 = ~w5712 & ~w5994;
assign w5996 = ~w5745 & w64688;
assign w5997 = ~w5981 & ~w5985;
assign w5998 = ~w5987 & ~w5990;
assign w5999 = w5997 & w5998;
assign w6000 = (w5999 & w5991) | (w5999 & w64689) | (w5991 & w64689);
assign w6001 = pi0366 & ~w6000;
assign w6002 = ~pi0366 & w6000;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = ~w5581 & ~w5610;
assign w6005 = ~w5589 & w64690;
assign w6006 = (w5574 & w5554) | (w5574 & w64691) | (w5554 & w64691);
assign w6007 = ~w6005 & ~w6006;
assign w6008 = (w5659 & w64692) | (w5659 & w64693) | (w64692 & w64693);
assign w6009 = ~w5574 & ~w5581;
assign w6010 = ~w5658 & w6009;
assign w6011 = ~w5921 & w6010;
assign w6012 = (w5659 & w64694) | (w5659 & w64695) | (w64694 & w64695);
assign w6013 = ~w6008 & w6012;
assign w6014 = pi0375 & w6013;
assign w6015 = ~pi0375 & ~w6013;
assign w6016 = ~w6014 & ~w6015;
assign w6017 = ~pi3214 & pi9040;
assign w6018 = ~pi3199 & ~pi9040;
assign w6019 = ~w6017 & ~w6018;
assign w6020 = pi0351 & ~w6019;
assign w6021 = ~pi0351 & w6019;
assign w6022 = ~w6020 & ~w6021;
assign w6023 = ~pi3201 & pi9040;
assign w6024 = ~pi3302 & ~pi9040;
assign w6025 = ~w6023 & ~w6024;
assign w6026 = pi0328 & ~w6025;
assign w6027 = ~pi0328 & w6025;
assign w6028 = ~w6026 & ~w6027;
assign w6029 = ~w6022 & w6028;
assign w6030 = ~pi3252 & pi9040;
assign w6031 = ~pi3385 & ~pi9040;
assign w6032 = ~w6030 & ~w6031;
assign w6033 = pi0333 & ~w6032;
assign w6034 = ~pi0333 & w6032;
assign w6035 = ~w6033 & ~w6034;
assign w6036 = ~pi3333 & pi9040;
assign w6037 = ~pi3253 & ~pi9040;
assign w6038 = ~w6036 & ~w6037;
assign w6039 = pi0346 & ~w6038;
assign w6040 = ~pi0346 & w6038;
assign w6041 = ~w6039 & ~w6040;
assign w6042 = w6035 & w6041;
assign w6043 = w6029 & w6042;
assign w6044 = ~pi3322 & pi9040;
assign w6045 = ~pi3218 & ~pi9040;
assign w6046 = ~w6044 & ~w6045;
assign w6047 = pi0326 & ~w6046;
assign w6048 = ~pi0326 & w6046;
assign w6049 = ~w6047 & ~w6048;
assign w6050 = ~w6022 & w6035;
assign w6051 = w6028 & w6035;
assign w6052 = ~w6041 & w6051;
assign w6053 = ~pi3302 & pi9040;
assign w6054 = ~pi3258 & ~pi9040;
assign w6055 = ~w6053 & ~w6054;
assign w6056 = pi0324 & ~w6055;
assign w6057 = ~pi0324 & w6055;
assign w6058 = ~w6056 & ~w6057;
assign w6059 = w6029 & w6058;
assign w6060 = ~w6052 & ~w6059;
assign w6061 = ~w6050 & ~w6060;
assign w6062 = w6029 & ~w6041;
assign w6063 = ~w6028 & w6042;
assign w6064 = ~w6062 & ~w6063;
assign w6065 = ~w6058 & w6064;
assign w6066 = w6028 & w6041;
assign w6067 = ~w6035 & w6041;
assign w6068 = w6022 & ~w6028;
assign w6069 = ~w6067 & w6068;
assign w6070 = ~w6066 & ~w6069;
assign w6071 = w6065 & w6070;
assign w6072 = (~w6049 & w6071) | (~w6049 & w64696) | (w6071 & w64696);
assign w6073 = ~w6022 & ~w6028;
assign w6074 = ~w6035 & w6066;
assign w6075 = w6066 & w64697;
assign w6076 = ~w6050 & ~w6075;
assign w6077 = ~w6073 & ~w6076;
assign w6078 = ~w6028 & ~w6041;
assign w6079 = w6067 & w6073;
assign w6080 = (w6058 & ~w6051) | (w6058 & w63569) | (~w6051 & w63569);
assign w6081 = ~w6079 & w6080;
assign w6082 = ~w6078 & w6081;
assign w6083 = w6022 & ~w6041;
assign w6084 = ~w6051 & w6083;
assign w6085 = w6081 & w64698;
assign w6086 = ~w6065 & ~w6085;
assign w6087 = ~w6077 & ~w6086;
assign w6088 = w6049 & ~w6087;
assign w6089 = ~w6035 & w6078;
assign w6090 = w6078 & w64697;
assign w6091 = ~w6075 & ~w6090;
assign w6092 = ~w6041 & w6050;
assign w6093 = w6091 & ~w6092;
assign w6094 = w6022 & w6042;
assign w6095 = (w6058 & ~w6029) | (w6058 & w63355) | (~w6029 & w63355);
assign w6096 = ~w6094 & w6095;
assign w6097 = ~w6093 & w6096;
assign w6098 = w6041 & ~w6058;
assign w6099 = w6068 & w6098;
assign w6100 = ~w6043 & ~w6099;
assign w6101 = ~w6097 & w6100;
assign w6102 = ~w6072 & w6101;
assign w6103 = ~w6088 & w6102;
assign w6104 = ~pi0356 & w6103;
assign w6105 = pi0356 & ~w6103;
assign w6106 = ~w6104 & ~w6105;
assign w6107 = w5231 & ~w5271;
assign w6108 = ~w5252 & w6107;
assign w6109 = ~w5267 & ~w6108;
assign w6110 = ~w5268 & ~w6109;
assign w6111 = w5244 & w5252;
assign w6112 = ~w5413 & w6111;
assign w6113 = w5280 & ~w5962;
assign w6114 = ~w5280 & w5402;
assign w6115 = w5962 & w6114;
assign w6116 = (~w5267 & w6115) | (~w5267 & w64699) | (w6115 & w64699);
assign w6117 = w5394 & ~w6112;
assign w6118 = ~w6116 & w6117;
assign w6119 = w5403 & ~w6113;
assign w6120 = w5275 & ~w6111;
assign w6121 = ~w6107 & ~w6120;
assign w6122 = ~w5276 & ~w6121;
assign w6123 = ~w5261 & ~w5293;
assign w6124 = ~w5972 & w6123;
assign w6125 = ~w6119 & w6124;
assign w6126 = ~w6122 & w6125;
assign w6127 = ~w6118 & ~w6126;
assign w6128 = ~w6110 & ~w6127;
assign w6129 = ~pi0390 & w6128;
assign w6130 = pi0390 & ~w6128;
assign w6131 = ~w6129 & ~w6130;
assign w6132 = ~w5470 & w5482;
assign w6133 = ~w5525 & ~w5886;
assign w6134 = ~w5466 & w6133;
assign w6135 = w5460 & ~w5486;
assign w6136 = ~w5516 & w6135;
assign w6137 = ~w6134 & ~w6136;
assign w6138 = ~w6132 & ~w6137;
assign w6139 = ~w5455 & w6133;
assign w6140 = w5480 & ~w5500;
assign w6141 = ~w5497 & w6140;
assign w6142 = ~w6139 & w6141;
assign w6143 = ~w6138 & ~w6142;
assign w6144 = ~pi0370 & w6143;
assign w6145 = pi0370 & ~w6143;
assign w6146 = ~w6144 & ~w6145;
assign w6147 = ~w5724 & ~w5984;
assign w6148 = (~w5736 & w5984) | (~w5736 & w63570) | (w5984 & w63570);
assign w6149 = (w5715 & ~w5746) | (w5715 & w64700) | (~w5746 & w64700);
assign w6150 = w5698 & w5764;
assign w6151 = (w5692 & w6150) | (w5692 & w64701) | (w6150 & w64701);
assign w6152 = w5672 & ~w5738;
assign w6153 = (~w5678 & w6152) | (~w5678 & w63571) | (w6152 & w63571);
assign w6154 = ~w5701 & ~w5739;
assign w6155 = (~w5748 & ~w6147) | (~w5748 & w63572) | (~w6147 & w63572);
assign w6156 = w5736 & ~w6155;
assign w6157 = w5742 & w5989;
assign w6158 = w6155 & w6157;
assign w6159 = ~w6148 & ~w6151;
assign w6160 = ~w6153 & w6159;
assign w6161 = ~w6156 & w6160;
assign w6162 = ~w6158 & w6161;
assign w6163 = (pi0362 & ~w6162) | (pi0362 & w64702) | (~w6162 & w64702);
assign w6164 = w6162 & w64703;
assign w6165 = ~w6163 & ~w6164;
assign w6166 = ~w5810 & w5833;
assign w6167 = ~w5830 & ~w5933;
assign w6168 = ~w6166 & ~w6167;
assign w6169 = ~w5822 & ~w6168;
assign w6170 = w5865 & ~w5931;
assign w6171 = ~w5861 & ~w5866;
assign w6172 = w5830 & ~w5876;
assign w6173 = ~w6171 & w6172;
assign w6174 = ~w5838 & ~w6173;
assign w6175 = w6170 & w6174;
assign w6176 = (~w5855 & ~w6175) | (~w5855 & w64704) | (~w6175 & w64704);
assign w6177 = ~w5852 & ~w5937;
assign w6178 = ~w5830 & ~w6170;
assign w6179 = ~w6177 & w6178;
assign w6180 = ~w6176 & ~w6179;
assign w6181 = ~pi0380 & w6180;
assign w6182 = pi0380 & ~w6180;
assign w6183 = ~w6181 & ~w6182;
assign w6184 = w6084 & ~w6089;
assign w6185 = ~w6058 & w6184;
assign w6186 = ~w6050 & ~w6067;
assign w6187 = ~w6064 & w6186;
assign w6188 = ~w6089 & w6096;
assign w6189 = w6035 & w6078;
assign w6190 = ~w6079 & ~w6189;
assign w6191 = w6028 & ~w6035;
assign w6192 = w6022 & w6191;
assign w6193 = ~w6043 & ~w6058;
assign w6194 = ~w6192 & w6193;
assign w6195 = w6190 & w6194;
assign w6196 = (~w6187 & w6195) | (~w6187 & w63356) | (w6195 & w63356);
assign w6197 = w6078 & w64705;
assign w6198 = ~w6063 & ~w6197;
assign w6199 = ~w6062 & w6198;
assign w6200 = w6196 & ~w6199;
assign w6201 = ~w6035 & ~w6066;
assign w6202 = w6096 & ~w6201;
assign w6203 = w6029 & w6067;
assign w6204 = (~w6058 & ~w6042) | (~w6058 & w64706) | (~w6042 & w64706);
assign w6205 = w6094 & w6204;
assign w6206 = w6067 & w6068;
assign w6207 = ~w6203 & ~w6206;
assign w6208 = ~w6205 & w6207;
assign w6209 = (w6049 & w6200) | (w6049 & w63573) | (w6200 & w63573);
assign w6210 = ~w6090 & ~w6203;
assign w6211 = w6058 & ~w6210;
assign w6212 = ~w6185 & ~w6211;
assign w6213 = (w6212 & w6196) | (w6212 & w64707) | (w6196 & w64707);
assign w6214 = ~w6209 & w64708;
assign w6215 = (pi0365 & w6209) | (pi0365 & w64709) | (w6209 & w64709);
assign w6216 = ~w6214 & ~w6215;
assign w6217 = ~w5336 & ~w5343;
assign w6218 = (w5353 & ~w6217) | (w5353 & w64710) | (~w6217 & w64710);
assign w6219 = w5336 & w5362;
assign w6220 = ~w5323 & ~w5343;
assign w6221 = w5323 & w5384;
assign w6222 = ~w6220 & ~w6221;
assign w6223 = w6218 & w6222;
assign w6224 = ~w6219 & w6223;
assign w6225 = ~w5343 & w5345;
assign w6226 = w5353 & w6225;
assign w6227 = (w5336 & w6220) | (w5336 & w64711) | (w6220 & w64711);
assign w6228 = ~w5346 & ~w6227;
assign w6229 = w5353 & ~w6228;
assign w6230 = w6221 & ~w6229;
assign w6231 = w5317 & ~w6226;
assign w6232 = ~w6219 & w6231;
assign w6233 = ~w6230 & w6232;
assign w6234 = w5356 & w6217;
assign w6235 = ~w5317 & ~w6234;
assign w6236 = ~w6229 & w6235;
assign w6237 = ~w6233 & ~w6236;
assign w6238 = ~w5360 & ~w5383;
assign w6239 = ~w5353 & w6228;
assign w6240 = ~w6238 & w6239;
assign w6241 = w5329 & ~w5353;
assign w6242 = ~w5317 & ~w5336;
assign w6243 = w6241 & w6242;
assign w6244 = (~w6243 & ~w6224) | (~w6243 & w64712) | (~w6224 & w64712);
assign w6245 = ~w6240 & w6244;
assign w6246 = ~w6237 & w6245;
assign w6247 = pi0379 & ~w6246;
assign w6248 = ~pi0379 & w6246;
assign w6249 = ~w6247 & ~w6248;
assign w6250 = w5353 & w5381;
assign w6251 = ~w5317 & ~w6250;
assign w6252 = w5329 & w5355;
assign w6253 = ~w5381 & ~w6252;
assign w6254 = ~w6225 & w6253;
assign w6255 = ~w6220 & ~w6254;
assign w6256 = (w6241 & w6221) | (w6241 & w64713) | (w6221 & w64713);
assign w6257 = ~w6226 & ~w6256;
assign w6258 = ~w6224 & w6257;
assign w6259 = (~w6251 & ~w6258) | (~w6251 & w64714) | (~w6258 & w64714);
assign w6260 = w5356 & w5364;
assign w6261 = ~w5353 & w6260;
assign w6262 = w5317 & ~w6261;
assign w6263 = ~w5344 & ~w5374;
assign w6264 = ~w5329 & ~w5353;
assign w6265 = w5355 & w6264;
assign w6266 = w5343 & ~w5360;
assign w6267 = ~w5353 & ~w6266;
assign w6268 = w5353 & ~w6252;
assign w6269 = ~w5337 & w6268;
assign w6270 = ~w6267 & ~w6269;
assign w6271 = ~w6260 & ~w6265;
assign w6272 = ~w5383 & w6271;
assign w6273 = w6263 & w6272;
assign w6274 = (~w6262 & ~w6273) | (~w6262 & w64715) | (~w6273 & w64715);
assign w6275 = ~w6259 & ~w6274;
assign w6276 = pi0368 & ~w6275;
assign w6277 = ~pi0368 & w6275;
assign w6278 = ~w6276 & ~w6277;
assign w6279 = ~w6022 & w6098;
assign w6280 = (w6058 & ~w6066) | (w6058 & w64716) | (~w6066 & w64716);
assign w6281 = ~w6092 & w6280;
assign w6282 = ~w6198 & w6281;
assign w6283 = w6049 & ~w6279;
assign w6284 = ~w6184 & w6283;
assign w6285 = ~w6282 & w6284;
assign w6286 = w6051 & w64717;
assign w6287 = ~w6092 & w6204;
assign w6288 = ~w6081 & ~w6287;
assign w6289 = (~w6049 & ~w6029) | (~w6049 & w64718) | (~w6029 & w64718);
assign w6290 = ~w6286 & w6289;
assign w6291 = w6091 & w6290;
assign w6292 = ~w6288 & w6291;
assign w6293 = ~w6285 & ~w6292;
assign w6294 = w6082 & ~w6087;
assign w6295 = ~w6186 & w6204;
assign w6296 = ~w6202 & ~w6295;
assign w6297 = w6068 & ~w6296;
assign w6298 = ~w6293 & ~w6297;
assign w6299 = ~w6294 & w6298;
assign w6300 = pi0353 & ~w6299;
assign w6301 = ~pi0353 & w6299;
assign w6302 = ~w6300 & ~w6301;
assign w6303 = ~w5323 & w5384;
assign w6304 = ~w5380 & ~w6303;
assign w6305 = ~w5372 & ~w6304;
assign w6306 = w5379 & ~w6305;
assign w6307 = ~w6218 & ~w6306;
assign w6308 = w5364 & w6264;
assign w6309 = ~w5353 & ~w6253;
assign w6310 = w6227 & w6268;
assign w6311 = w5317 & ~w6303;
assign w6312 = ~w6308 & w6311;
assign w6313 = w6263 & w6312;
assign w6314 = ~w6309 & ~w6310;
assign w6315 = w6313 & w6314;
assign w6316 = (w5353 & ~w6220) | (w5353 & w64719) | (~w6220 & w64719);
assign w6317 = (~w5361 & ~w6304) | (~w5361 & w64720) | (~w6304 & w64720);
assign w6318 = ~w5345 & w5361;
assign w6319 = ~w6241 & w6318;
assign w6320 = ~w6317 & ~w6319;
assign w6321 = ~w5317 & ~w6265;
assign w6322 = ~w6320 & w6321;
assign w6323 = ~w6315 & ~w6322;
assign w6324 = ~w6307 & ~w6323;
assign w6325 = pi0377 & w6324;
assign w6326 = ~pi0377 & ~w6324;
assign w6327 = ~w6325 & ~w6326;
assign w6328 = w5822 & w5944;
assign w6329 = ~w5795 & ~w5818;
assign w6330 = ~w5945 & ~w6329;
assign w6331 = ~w5850 & ~w6330;
assign w6332 = w5861 & w5944;
assign w6333 = ~w5931 & ~w6332;
assign w6334 = ~w6331 & w6333;
assign w6335 = ~w5845 & ~w6334;
assign w6336 = w5848 & ~w6329;
assign w6337 = w5877 & w6336;
assign w6338 = ~w5862 & ~w5877;
assign w6339 = ~w5812 & ~w6338;
assign w6340 = w5812 & ~w5830;
assign w6341 = w5845 & ~w6339;
assign w6342 = ~w6340 & w6341;
assign w6343 = ~w6328 & ~w6337;
assign w6344 = ~w6335 & w6343;
assign w6345 = ~w6342 & w6344;
assign w6346 = pi0398 & ~w6345;
assign w6347 = ~pi0398 & w6345;
assign w6348 = ~w6346 & ~w6347;
assign w6349 = ~w6050 & ~w6191;
assign w6350 = w6281 & ~w6349;
assign w6351 = ~w6043 & ~w6206;
assign w6352 = ~w6286 & w6351;
assign w6353 = ~w6350 & w6352;
assign w6354 = w6049 & ~w6353;
assign w6355 = ~w6281 & ~w6295;
assign w6356 = ~w6069 & ~w6355;
assign w6357 = ~w6049 & ~w6356;
assign w6358 = ~w6190 & w6281;
assign w6359 = ~w6074 & w6198;
assign w6360 = ~w6058 & w6076;
assign w6361 = ~w6359 & w6360;
assign w6362 = ~w6358 & ~w6361;
assign w6363 = ~w6354 & w6362;
assign w6364 = ~w6357 & w6363;
assign w6365 = pi0378 & ~w6364;
assign w6366 = ~pi0378 & w6364;
assign w6367 = ~w6365 & ~w6366;
assign w6368 = ~pi3220 & pi9040;
assign w6369 = ~pi3216 & ~pi9040;
assign w6370 = ~w6368 & ~w6369;
assign w6371 = pi0344 & ~w6370;
assign w6372 = ~pi0344 & w6370;
assign w6373 = ~w6371 & ~w6372;
assign w6374 = ~pi3223 & pi9040;
assign w6375 = ~pi3259 & ~pi9040;
assign w6376 = ~w6374 & ~w6375;
assign w6377 = pi0349 & ~w6376;
assign w6378 = ~pi0349 & w6376;
assign w6379 = ~w6377 & ~w6378;
assign w6380 = ~w6373 & w6379;
assign w6381 = ~pi3203 & pi9040;
assign w6382 = ~pi3220 & ~pi9040;
assign w6383 = ~w6381 & ~w6382;
assign w6384 = pi0330 & ~w6383;
assign w6385 = ~pi0330 & w6383;
assign w6386 = ~w6384 & ~w6385;
assign w6387 = ~pi3263 & pi9040;
assign w6388 = ~pi3233 & ~pi9040;
assign w6389 = ~w6387 & ~w6388;
assign w6390 = pi0327 & ~w6389;
assign w6391 = ~pi0327 & w6389;
assign w6392 = ~w6390 & ~w6391;
assign w6393 = w6386 & w6392;
assign w6394 = ~w6380 & w6393;
assign w6395 = w6380 & ~w6392;
assign w6396 = ~w6394 & ~w6395;
assign w6397 = ~w6373 & ~w6386;
assign w6398 = w6373 & w6386;
assign w6399 = ~w6397 & ~w6398;
assign w6400 = ~w6379 & ~w6392;
assign w6401 = ~w6399 & ~w6400;
assign w6402 = ~w6373 & ~w6379;
assign w6403 = ~w6386 & ~w6392;
assign w6404 = ~w6402 & ~w6403;
assign w6405 = ~w6397 & ~w6404;
assign w6406 = ~w6401 & ~w6405;
assign w6407 = ~pi3210 & pi9040;
assign w6408 = ~pi3212 & ~pi9040;
assign w6409 = ~w6407 & ~w6408;
assign w6410 = pi0323 & ~w6409;
assign w6411 = ~pi0323 & w6409;
assign w6412 = ~w6410 & ~w6411;
assign w6413 = ~w6398 & w6412;
assign w6414 = w6396 & w6413;
assign w6415 = ~w6406 & w6414;
assign w6416 = w6379 & w6397;
assign w6417 = w6415 & w6416;
assign w6418 = ~pi3259 & pi9040;
assign w6419 = ~pi3222 & ~pi9040;
assign w6420 = ~w6418 & ~w6419;
assign w6421 = pi0315 & ~w6420;
assign w6422 = ~pi0315 & w6420;
assign w6423 = ~w6421 & ~w6422;
assign w6424 = w6373 & ~w6379;
assign w6425 = w6392 & w6424;
assign w6426 = w6399 & w6404;
assign w6427 = ~w6424 & ~w6426;
assign w6428 = (w6412 & w6426) | (w6412 & w64721) | (w6426 & w64721);
assign w6429 = w6402 & w6403;
assign w6430 = ~w6425 & ~w6429;
assign w6431 = ~w6428 & w6430;
assign w6432 = w6423 & ~w6431;
assign w6433 = w6379 & ~w6392;
assign w6434 = ~w6386 & w6423;
assign w6435 = (w6433 & ~w6399) | (w6433 & w64722) | (~w6399 & w64722);
assign w6436 = w6399 & w64723;
assign w6437 = ~w6435 & ~w6436;
assign w6438 = ~w6379 & ~w6386;
assign w6439 = ~w6380 & ~w6438;
assign w6440 = w6426 & w6439;
assign w6441 = ~w6423 & w6440;
assign w6442 = ~w6373 & w6386;
assign w6443 = w6379 & ~w6442;
assign w6444 = ~w6379 & w6399;
assign w6445 = w6392 & ~w6443;
assign w6446 = ~w6444 & w6445;
assign w6447 = w6437 & ~w6446;
assign w6448 = ~w6441 & w6447;
assign w6449 = ~w6412 & ~w6448;
assign w6450 = w6412 & ~w6423;
assign w6451 = ~w6397 & w6450;
assign w6452 = w6427 & w6451;
assign w6453 = ~w6417 & ~w6452;
assign w6454 = ~w6432 & w6453;
assign w6455 = (~pi0369 & ~w6454) | (~pi0369 & w64724) | (~w6454 & w64724);
assign w6456 = w6454 & w64725;
assign w6457 = ~w6455 & ~w6456;
assign w6458 = w6379 & w6392;
assign w6459 = w6379 & w6398;
assign w6460 = ~w6373 & ~w6403;
assign w6461 = ~w6439 & ~w6460;
assign w6462 = (~w6423 & w6461) | (~w6423 & w63574) | (w6461 & w63574);
assign w6463 = w6458 & w6462;
assign w6464 = ~w6379 & w6393;
assign w6465 = w6423 & ~w6464;
assign w6466 = (w6465 & w6406) | (w6465 & w63357) | (w6406 & w63357);
assign w6467 = ~w6406 & ~w6423;
assign w6468 = ~w6466 & ~w6467;
assign w6469 = w6392 & ~w6466;
assign w6470 = w6412 & ~w6433;
assign w6471 = ~w6468 & w6470;
assign w6472 = ~w6469 & w6471;
assign w6473 = ~w6373 & w6464;
assign w6474 = ~w6468 & ~w6473;
assign w6475 = w6401 & w6450;
assign w6476 = ~w6397 & w6423;
assign w6477 = ~w6459 & w6476;
assign w6478 = ~w6437 & w6477;
assign w6479 = ~w6463 & ~w6475;
assign w6480 = ~w6478 & w6479;
assign w6481 = ~w6472 & w6480;
assign w6482 = (~pi0371 & ~w6481) | (~pi0371 & w63575) | (~w6481 & w63575);
assign w6483 = w6481 & w63576;
assign w6484 = ~w6482 & ~w6483;
assign w6485 = w6446 & w6465;
assign w6486 = ~w6423 & w6464;
assign w6487 = ~w6393 & ~w6423;
assign w6488 = w6460 & w6487;
assign w6489 = ~w6373 & ~w6423;
assign w6490 = w6379 & ~w6489;
assign w6491 = ~w6399 & w6490;
assign w6492 = ~w6444 & ~w6491;
assign w6493 = ~w6392 & ~w6492;
assign w6494 = w6412 & ~w6488;
assign w6495 = ~w6440 & w6494;
assign w6496 = ~w6493 & w6495;
assign w6497 = w6476 & w6492;
assign w6498 = ~w6412 & ~w6429;
assign w6499 = ~w6462 & w6498;
assign w6500 = ~w6497 & w6499;
assign w6501 = ~w6496 & ~w6500;
assign w6502 = ~w6485 & ~w6486;
assign w6503 = ~w6501 & w6502;
assign w6504 = ~pi0363 & w6503;
assign w6505 = pi0363 & ~w6503;
assign w6506 = ~w6504 & ~w6505;
assign w6507 = w6412 & ~w6424;
assign w6508 = ~w6396 & ~w6507;
assign w6509 = (w6423 & w6415) | (w6423 & w64726) | (w6415 & w64726);
assign w6510 = ~w6379 & w6406;
assign w6511 = w6439 & w6487;
assign w6512 = ~w6510 & ~w6511;
assign w6513 = ~w6412 & ~w6512;
assign w6514 = ~w6393 & ~w6416;
assign w6515 = w6450 & ~w6514;
assign w6516 = ~w6413 & ~w6489;
assign w6517 = w6458 & ~w6516;
assign w6518 = ~w6515 & ~w6517;
assign w6519 = ~w6509 & w6518;
assign w6520 = ~w6513 & w6519;
assign w6521 = pi0372 & ~w6520;
assign w6522 = ~pi0372 & w6520;
assign w6523 = ~w6521 & ~w6522;
assign w6524 = ~pi3289 & pi9040;
assign w6525 = ~pi3280 & ~pi9040;
assign w6526 = ~w6524 & ~w6525;
assign w6527 = pi0401 & ~w6526;
assign w6528 = ~pi0401 & w6526;
assign w6529 = ~w6527 & ~w6528;
assign w6530 = ~pi3283 & pi9040;
assign w6531 = ~pi3335 & ~pi9040;
assign w6532 = ~w6530 & ~w6531;
assign w6533 = pi0405 & ~w6532;
assign w6534 = ~pi0405 & w6532;
assign w6535 = ~w6533 & ~w6534;
assign w6536 = ~w6529 & ~w6535;
assign w6537 = w6529 & w6535;
assign w6538 = ~w6536 & ~w6537;
assign w6539 = ~pi3334 & pi9040;
assign w6540 = ~pi3352 & ~pi9040;
assign w6541 = ~w6539 & ~w6540;
assign w6542 = pi0389 & ~w6541;
assign w6543 = ~pi0389 & w6541;
assign w6544 = ~w6542 & ~w6543;
assign w6545 = ~pi3287 & pi9040;
assign w6546 = ~pi3315 & ~pi9040;
assign w6547 = ~w6545 & ~w6546;
assign w6548 = pi0382 & ~w6547;
assign w6549 = ~pi0382 & w6547;
assign w6550 = ~w6548 & ~w6549;
assign w6551 = ~w6544 & ~w6550;
assign w6552 = ~w6538 & w6551;
assign w6553 = w6544 & w6550;
assign w6554 = w6535 & ~w6544;
assign w6555 = ~w6553 & ~w6554;
assign w6556 = w6529 & ~w6550;
assign w6557 = ~w6536 & ~w6556;
assign w6558 = w6555 & w6557;
assign w6559 = ~w6552 & ~w6558;
assign w6560 = ~pi3321 & pi9040;
assign w6561 = ~pi3402 & ~pi9040;
assign w6562 = ~w6560 & ~w6561;
assign w6563 = pi0402 & ~w6562;
assign w6564 = ~pi0402 & w6562;
assign w6565 = ~w6563 & ~w6564;
assign w6566 = ~w6559 & w6565;
assign w6567 = ~w6529 & w6544;
assign w6568 = ~w6535 & w6550;
assign w6569 = w6567 & ~w6568;
assign w6570 = w6565 & ~w6569;
assign w6571 = w6544 & ~w6550;
assign w6572 = w6538 & w6571;
assign w6573 = ~w6550 & w6554;
assign w6574 = ~w6572 & ~w6573;
assign w6575 = w6570 & ~w6574;
assign w6576 = (w6565 & w6538) | (w6565 & w63358) | (w6538 & w63358);
assign w6577 = w6535 & w6550;
assign w6578 = w6529 & ~w6544;
assign w6579 = ~w6567 & ~w6578;
assign w6580 = ~w6537 & ~w6579;
assign w6581 = (~w6577 & w6579) | (~w6577 & w63359) | (w6579 & w63359);
assign w6582 = ~w6576 & ~w6581;
assign w6583 = ~pi3285 & pi9040;
assign w6584 = ~pi3421 & ~pi9040;
assign w6585 = ~w6583 & ~w6584;
assign w6586 = pi0415 & ~w6585;
assign w6587 = ~pi0415 & w6585;
assign w6588 = ~w6586 & ~w6587;
assign w6589 = (~w6588 & w6575) | (~w6588 & w64727) | (w6575 & w64727);
assign w6590 = w6544 & ~w6577;
assign w6591 = ~w6538 & ~w6565;
assign w6592 = w6590 & w6591;
assign w6593 = w6550 & w6592;
assign w6594 = w6567 & w6577;
assign w6595 = w6529 & w6550;
assign w6596 = w6535 & ~w6565;
assign w6597 = ~w6595 & ~w6596;
assign w6598 = ~w6579 & ~w6597;
assign w6599 = ~w6544 & w6568;
assign w6600 = ~w6565 & w6599;
assign w6601 = ~w6594 & ~w6598;
assign w6602 = ~w6600 & w6601;
assign w6603 = ~w6567 & w6568;
assign w6604 = w6570 & ~w6603;
assign w6605 = w6602 & w6604;
assign w6606 = w6550 & ~w6578;
assign w6607 = ~w6577 & ~w6579;
assign w6608 = ~w6606 & ~w6607;
assign w6609 = ~w6565 & ~w6608;
assign w6610 = w6588 & ~w6609;
assign w6611 = ~w6605 & w6610;
assign w6612 = ~w6566 & ~w6593;
assign w6613 = ~w6589 & w6612;
assign w6614 = ~w6611 & w6613;
assign w6615 = pi0421 & ~w6614;
assign w6616 = ~pi0421 & w6614;
assign w6617 = ~w6615 & ~w6616;
assign w6618 = ~pi3286 & pi9040;
assign w6619 = ~pi3287 & ~pi9040;
assign w6620 = ~w6618 & ~w6619;
assign w6621 = pi0400 & ~w6620;
assign w6622 = ~pi0400 & w6620;
assign w6623 = ~w6621 & ~w6622;
assign w6624 = ~pi3284 & pi9040;
assign w6625 = ~pi3401 & ~pi9040;
assign w6626 = ~w6624 & ~w6625;
assign w6627 = pi0391 & ~w6626;
assign w6628 = ~pi0391 & w6626;
assign w6629 = ~w6627 & ~w6628;
assign w6630 = ~pi3417 & pi9040;
assign w6631 = ~pi3313 & ~pi9040;
assign w6632 = ~w6630 & ~w6631;
assign w6633 = pi0397 & ~w6632;
assign w6634 = ~pi0397 & w6632;
assign w6635 = ~w6633 & ~w6634;
assign w6636 = ~w6629 & ~w6635;
assign w6637 = ~pi3339 & pi9040;
assign w6638 = ~pi3285 & ~pi9040;
assign w6639 = ~w6637 & ~w6638;
assign w6640 = pi0383 & ~w6639;
assign w6641 = ~pi0383 & w6639;
assign w6642 = ~w6640 & ~w6641;
assign w6643 = w6636 & w6642;
assign w6644 = ~pi3315 & pi9040;
assign w6645 = ~pi3283 & ~pi9040;
assign w6646 = ~w6644 & ~w6645;
assign w6647 = pi0387 & ~w6646;
assign w6648 = ~pi0387 & w6646;
assign w6649 = ~w6647 & ~w6648;
assign w6650 = w6643 & w6649;
assign w6651 = ~w6635 & ~w6642;
assign w6652 = w6629 & ~w6642;
assign w6653 = ~w6629 & ~w6649;
assign w6654 = w6635 & ~w6653;
assign w6655 = ~pi3402 & pi9040;
assign w6656 = ~pi3277 & ~pi9040;
assign w6657 = ~w6655 & ~w6656;
assign w6658 = pi0411 & ~w6657;
assign w6659 = ~pi0411 & w6657;
assign w6660 = ~w6658 & ~w6659;
assign w6661 = (w6660 & ~w6654) | (w6660 & w63360) | (~w6654 & w63360);
assign w6662 = ~w6651 & w6661;
assign w6663 = ~w6653 & w6660;
assign w6664 = w6629 & w6649;
assign w6665 = w6635 & ~w6642;
assign w6666 = w6664 & w6665;
assign w6667 = w6635 & w6642;
assign w6668 = ~w6651 & ~w6667;
assign w6669 = ~w6629 & ~w6668;
assign w6670 = (w6663 & w6669) | (w6663 & w63577) | (w6669 & w63577);
assign w6671 = ~w6636 & ~w6652;
assign w6672 = ~w6649 & w6671;
assign w6673 = ~w6660 & ~w6666;
assign w6674 = ~w6672 & w6673;
assign w6675 = ~w6662 & ~w6674;
assign w6676 = ~w6623 & ~w6650;
assign w6677 = (w6676 & ~w6675) | (w6676 & w64728) | (~w6675 & w64728);
assign w6678 = w6642 & w6664;
assign w6679 = w6635 & ~w6649;
assign w6680 = ~w6629 & ~w6642;
assign w6681 = ~w6679 & w6680;
assign w6682 = ~w6678 & ~w6681;
assign w6683 = (~w6682 & ~w6675) | (~w6682 & w63578) | (~w6675 & w63578);
assign w6684 = w6629 & w6660;
assign w6685 = ~w6649 & ~w6684;
assign w6686 = w6652 & w6685;
assign w6687 = w6642 & ~w6649;
assign w6688 = w6636 & w6687;
assign w6689 = ~w6686 & ~w6688;
assign w6690 = w6623 & w6689;
assign w6691 = ~w6683 & w6690;
assign w6692 = ~w6677 & ~w6691;
assign w6693 = w6629 & ~w6649;
assign w6694 = w6651 & w6693;
assign w6695 = w6623 & ~w6693;
assign w6696 = w6682 & w6695;
assign w6697 = ~w6687 & ~w6696;
assign w6698 = w6635 & w6660;
assign w6699 = ~w6697 & w6698;
assign w6700 = ~w6694 & ~w6699;
assign w6701 = (pi0422 & w6692) | (pi0422 & w64729) | (w6692 & w64729);
assign w6702 = ~w6692 & w64730;
assign w6703 = ~w6701 & ~w6702;
assign w6704 = (~w6660 & ~w6654) | (~w6660 & w64731) | (~w6654 & w64731);
assign w6705 = ~w6689 & ~w6704;
assign w6706 = ~w6635 & w6649;
assign w6707 = w6684 & w6706;
assign w6708 = ~w6643 & w6663;
assign w6709 = ~w6704 & ~w6708;
assign w6710 = w6649 & ~w6671;
assign w6711 = w6642 & ~w6706;
assign w6712 = ~w6651 & ~w6711;
assign w6713 = ~w6711 & w64732;
assign w6714 = ~w6710 & w6713;
assign w6715 = ~w6686 & ~w6707;
assign w6716 = ~w6709 & w6715;
assign w6717 = ~w6714 & w6716;
assign w6718 = ~w6623 & ~w6717;
assign w6719 = w6629 & ~w6660;
assign w6720 = w6687 & w6719;
assign w6721 = ~w6635 & w6720;
assign w6722 = w6642 & w6653;
assign w6723 = w6653 & w6667;
assign w6724 = (~w6660 & w6671) | (~w6660 & w64733) | (w6671 & w64733);
assign w6725 = ~w6721 & ~w6723;
assign w6726 = w6661 & ~w6694;
assign w6727 = (w6623 & ~w6725) | (w6623 & w64734) | (~w6725 & w64734);
assign w6728 = ~w6726 & w6727;
assign w6729 = ~w6629 & ~w6660;
assign w6730 = ~w6665 & ~w6729;
assign w6731 = w6685 & ~w6730;
assign w6732 = w6681 & w6731;
assign w6733 = (w6660 & w6668) | (w6660 & w6684) | (w6668 & w6684);
assign w6734 = ~w6678 & ~w6731;
assign w6735 = w6733 & ~w6734;
assign w6736 = ~w6705 & ~w6732;
assign w6737 = ~w6735 & w6736;
assign w6738 = ~w6728 & w6737;
assign w6739 = w6738 & w64735;
assign w6740 = (~pi0420 & ~w6738) | (~pi0420 & w64736) | (~w6738 & w64736);
assign w6741 = ~w6739 & ~w6740;
assign w6742 = ~pi3401 & pi9040;
assign w6743 = ~pi3339 & ~pi9040;
assign w6744 = ~w6742 & ~w6743;
assign w6745 = pi0384 & ~w6744;
assign w6746 = ~pi0384 & w6744;
assign w6747 = ~w6745 & ~w6746;
assign w6748 = ~pi3303 & pi9040;
assign w6749 = ~pi3340 & ~pi9040;
assign w6750 = ~w6748 & ~w6749;
assign w6751 = pi0400 & ~w6750;
assign w6752 = ~pi0400 & w6750;
assign w6753 = ~w6751 & ~w6752;
assign w6754 = ~w6747 & w6753;
assign w6755 = w6747 & ~w6753;
assign w6756 = ~w6754 & ~w6755;
assign w6757 = ~pi3313 & pi9040;
assign w6758 = ~pi3284 & ~pi9040;
assign w6759 = ~w6757 & ~w6758;
assign w6760 = pi0383 & ~w6759;
assign w6761 = ~pi0383 & w6759;
assign w6762 = ~w6760 & ~w6761;
assign w6763 = ~pi3288 & pi9040;
assign w6764 = ~pi3291 & ~pi9040;
assign w6765 = ~w6763 & ~w6764;
assign w6766 = pi0406 & ~w6765;
assign w6767 = ~pi0406 & w6765;
assign w6768 = ~w6766 & ~w6767;
assign w6769 = w6762 & ~w6768;
assign w6770 = w6756 & w6769;
assign w6771 = ~pi3293 & pi9040;
assign w6772 = ~pi3342 & ~pi9040;
assign w6773 = ~w6771 & ~w6772;
assign w6774 = pi0389 & ~w6773;
assign w6775 = ~pi0389 & w6773;
assign w6776 = ~w6774 & ~w6775;
assign w6777 = ~w6768 & w6776;
assign w6778 = ~pi3340 & pi9040;
assign w6779 = ~pi3293 & ~pi9040;
assign w6780 = ~w6778 & ~w6779;
assign w6781 = pi0382 & ~w6780;
assign w6782 = ~pi0382 & w6780;
assign w6783 = ~w6781 & ~w6782;
assign w6784 = w6762 & w6783;
assign w6785 = ~w6754 & ~w6784;
assign w6786 = ~w6747 & ~w6783;
assign w6787 = w6753 & w6762;
assign w6788 = ~w6786 & ~w6787;
assign w6789 = w6777 & ~w6785;
assign w6790 = w6788 & w6789;
assign w6791 = ~w6762 & ~w6783;
assign w6792 = ~w6755 & ~w6791;
assign w6793 = w6755 & w6791;
assign w6794 = ~w6792 & ~w6793;
assign w6795 = w6768 & ~w6784;
assign w6796 = w6794 & w6795;
assign w6797 = ~w6768 & ~w6794;
assign w6798 = w6753 & ~w6783;
assign w6799 = ~w6753 & w6783;
assign w6800 = ~w6798 & ~w6799;
assign w6801 = ~w6747 & w6800;
assign w6802 = ~w6791 & w6801;
assign w6803 = w6797 & ~w6802;
assign w6804 = w6756 & w6784;
assign w6805 = ~w6747 & ~w6762;
assign w6806 = w6753 & w6768;
assign w6807 = ~w6798 & ~w6806;
assign w6808 = w6805 & ~w6807;
assign w6809 = ~w6776 & ~w6804;
assign w6810 = ~w6808 & w6809;
assign w6811 = ~w6803 & w6810;
assign w6812 = w6747 & w6762;
assign w6813 = ~w6805 & ~w6812;
assign w6814 = ~w6786 & w6806;
assign w6815 = w6813 & w6814;
assign w6816 = ~w6753 & ~w6762;
assign w6817 = w6794 & w6816;
assign w6818 = w6776 & ~w6815;
assign w6819 = ~w6817 & w6818;
assign w6820 = ~w6811 & ~w6819;
assign w6821 = ~w6770 & ~w6790;
assign w6822 = ~w6796 & w6821;
assign w6823 = ~w6820 & w6822;
assign w6824 = pi0435 & ~w6823;
assign w6825 = ~pi0435 & w6823;
assign w6826 = ~w6824 & ~w6825;
assign w6827 = ~w6762 & w6783;
assign w6828 = w6768 & ~w6827;
assign w6829 = w6747 & w6753;
assign w6830 = w6762 & ~w6783;
assign w6831 = ~w6827 & ~w6830;
assign w6832 = ~w6829 & ~w6831;
assign w6833 = ~w6753 & w6830;
assign w6834 = ~w6800 & w6805;
assign w6835 = ~w6833 & ~w6834;
assign w6836 = (w6786 & w6834) | (w6786 & w64737) | (w6834 & w64737);
assign w6837 = (w6799 & w6795) | (w6799 & w64738) | (w6795 & w64738);
assign w6838 = (~w6793 & w6832) | (~w6793 & w63579) | (w6832 & w63579);
assign w6839 = ~w6837 & w6838;
assign w6840 = ~w6836 & w6839;
assign w6841 = (~w6776 & ~w6839) | (~w6776 & w64739) | (~w6839 & w64739);
assign w6842 = w6776 & ~w6797;
assign w6843 = w6840 & w6842;
assign w6844 = w6747 & w6783;
assign w6845 = w6776 & ~w6844;
assign w6846 = w6788 & ~w6816;
assign w6847 = w6845 & w6846;
assign w6848 = ~w6841 & ~w6847;
assign w6849 = ~w6843 & w6848;
assign w6850 = pi0430 & w6849;
assign w6851 = ~pi0430 & ~w6849;
assign w6852 = ~w6850 & ~w6851;
assign w6853 = w6629 & w6679;
assign w6854 = ~w6643 & ~w6853;
assign w6855 = w6733 & w6854;
assign w6856 = ~w6678 & ~w6729;
assign w6857 = ~w6668 & ~w6856;
assign w6858 = ~w6855 & ~w6857;
assign w6859 = ~w6623 & ~w6858;
assign w6860 = ~w6642 & w6679;
assign w6861 = w6649 & w6669;
assign w6862 = w6660 & ~w6854;
assign w6863 = ~w6635 & w6719;
assign w6864 = ~w6688 & ~w6860;
assign w6865 = ~w6863 & w6864;
assign w6866 = ~w6861 & w6865;
assign w6867 = ~w6862 & w6866;
assign w6868 = w6623 & ~w6867;
assign w6869 = ~w6705 & ~w6721;
assign w6870 = ~w6859 & w6869;
assign w6871 = ~w6868 & w6870;
assign w6872 = pi0433 & ~w6871;
assign w6873 = ~pi0433 & w6871;
assign w6874 = ~w6872 & ~w6873;
assign w6875 = ~pi3276 & pi9040;
assign w6876 = ~pi3380 & ~pi9040;
assign w6877 = ~w6875 & ~w6876;
assign w6878 = pi0405 & ~w6877;
assign w6879 = ~pi0405 & w6877;
assign w6880 = ~w6878 & ~w6879;
assign w6881 = ~pi3319 & pi9040;
assign w6882 = ~pi3317 & ~pi9040;
assign w6883 = ~w6881 & ~w6882;
assign w6884 = pi0407 & ~w6883;
assign w6885 = ~pi0407 & w6883;
assign w6886 = ~w6884 & ~w6885;
assign w6887 = w6880 & ~w6886;
assign w6888 = ~pi3364 & pi9040;
assign w6889 = ~pi3278 & ~pi9040;
assign w6890 = ~w6888 & ~w6889;
assign w6891 = pi0415 & ~w6890;
assign w6892 = ~pi0415 & w6890;
assign w6893 = ~w6891 & ~w6892;
assign w6894 = w6887 & w6893;
assign w6895 = ~pi3320 & pi9040;
assign w6896 = ~pi3341 & ~pi9040;
assign w6897 = ~w6895 & ~w6896;
assign w6898 = pi0404 & ~w6897;
assign w6899 = ~pi0404 & w6897;
assign w6900 = ~w6898 & ~w6899;
assign w6901 = ~w6894 & w6900;
assign w6902 = ~pi3317 & pi9040;
assign w6903 = ~pi3364 & ~pi9040;
assign w6904 = ~w6902 & ~w6903;
assign w6905 = pi0376 & ~w6904;
assign w6906 = ~pi0376 & w6904;
assign w6907 = ~w6905 & ~w6906;
assign w6908 = w6880 & ~w6907;
assign w6909 = w6893 & w6907;
assign w6910 = ~w6908 & ~w6909;
assign w6911 = ~w6886 & ~w6910;
assign w6912 = ~w6880 & w6907;
assign w6913 = ~w6893 & ~w6907;
assign w6914 = ~pi3318 & pi9040;
assign w6915 = ~pi3414 & ~pi9040;
assign w6916 = ~w6914 & ~w6915;
assign w6917 = pi0392 & ~w6916;
assign w6918 = ~pi0392 & w6916;
assign w6919 = ~w6917 & ~w6918;
assign w6920 = w6913 & w6919;
assign w6921 = ~w6912 & ~w6920;
assign w6922 = ~w6911 & ~w6921;
assign w6923 = ~w6880 & ~w6907;
assign w6924 = w6886 & ~w6893;
assign w6925 = ~w6923 & ~w6924;
assign w6926 = ~w6913 & ~w6919;
assign w6927 = ~w6925 & w6926;
assign w6928 = ~w6922 & ~w6927;
assign w6929 = w6901 & w6928;
assign w6930 = w6880 & w6886;
assign w6931 = w6910 & w6930;
assign w6932 = ~w6886 & ~w6912;
assign w6933 = ~w6908 & ~w6932;
assign w6934 = ~w6913 & w6919;
assign w6935 = ~w6887 & w6934;
assign w6936 = ~w6933 & w6935;
assign w6937 = ~w6931 & ~w6936;
assign w6938 = (w6919 & w6936) | (w6919 & w64740) | (w6936 & w64740);
assign w6939 = ~w6893 & ~w6919;
assign w6940 = (w6939 & w6932) | (w6939 & w64741) | (w6932 & w64741);
assign w6941 = ~w6919 & ~w6932;
assign w6942 = w6909 & w6941;
assign w6943 = ~w6900 & ~w6940;
assign w6944 = ~w6942 & w6943;
assign w6945 = ~w6938 & w6944;
assign w6946 = ~w6929 & ~w6945;
assign w6947 = ~w6886 & ~w6919;
assign w6948 = w6908 & w6947;
assign w6949 = ~w6880 & w6886;
assign w6950 = ~w6939 & w6949;
assign w6951 = ~w6934 & w6950;
assign w6952 = ~w6908 & ~w6912;
assign w6953 = ~w6893 & ~w6952;
assign w6954 = w6893 & w6952;
assign w6955 = ~w6953 & ~w6954;
assign w6956 = ~w6886 & w6907;
assign w6957 = ~w6955 & w64742;
assign w6958 = ~w6948 & ~w6951;
assign w6959 = ~w6957 & w6958;
assign w6960 = ~w6946 & w6959;
assign w6961 = ~pi0418 & w6960;
assign w6962 = pi0418 & ~w6960;
assign w6963 = ~w6961 & ~w6962;
assign w6964 = ~pi3301 & pi9040;
assign w6965 = ~pi3354 & ~pi9040;
assign w6966 = ~w6964 & ~w6965;
assign w6967 = pi0409 & ~w6966;
assign w6968 = ~pi0409 & w6966;
assign w6969 = ~w6967 & ~w6968;
assign w6970 = ~pi3354 & pi9040;
assign w6971 = ~pi3305 & ~pi9040;
assign w6972 = ~w6970 & ~w6971;
assign w6973 = pi0395 & ~w6972;
assign w6974 = ~pi0395 & w6972;
assign w6975 = ~w6973 & ~w6974;
assign w6976 = ~w6969 & ~w6975;
assign w6977 = ~pi3338 & pi9040;
assign w6978 = ~pi3318 & ~pi9040;
assign w6979 = ~w6977 & ~w6978;
assign w6980 = pi0403 & ~w6979;
assign w6981 = ~pi0403 & w6979;
assign w6982 = ~w6980 & ~w6981;
assign w6983 = ~w6975 & ~w6982;
assign w6984 = w6969 & w6982;
assign w6985 = ~w6983 & ~w6984;
assign w6986 = w6969 & w6983;
assign w6987 = ~w6969 & w6975;
assign w6988 = ~pi3300 & pi9040;
assign w6989 = ~pi3299 & ~pi9040;
assign w6990 = ~w6988 & ~w6989;
assign w6991 = pi0394 & ~w6990;
assign w6992 = ~pi0394 & w6990;
assign w6993 = ~w6991 & ~w6992;
assign w6994 = w6987 & ~w6993;
assign w6995 = w6987 & w63361;
assign w6996 = ~pi3414 & pi9040;
assign w6997 = ~pi3320 & ~pi9040;
assign w6998 = ~w6996 & ~w6997;
assign w6999 = pi0410 & ~w6998;
assign w7000 = ~pi0410 & w6998;
assign w7001 = ~w6999 & ~w7000;
assign w7002 = ~w6995 & w7001;
assign w7003 = ~w6986 & w7002;
assign w7004 = ~w6982 & ~w6993;
assign w7005 = w6985 & ~w7004;
assign w7006 = ~w7003 & w7005;
assign w7007 = w6983 & w63580;
assign w7008 = w6976 & w7004;
assign w7009 = ~w7007 & ~w7008;
assign w7010 = w6969 & w6975;
assign w7011 = ~w6976 & ~w7010;
assign w7012 = ~w6993 & w7011;
assign w7013 = ~w6985 & w7001;
assign w7014 = ~w7012 & w7013;
assign w7015 = w7009 & ~w7014;
assign w7016 = ~w7006 & w7015;
assign w7017 = ~w6975 & ~w6993;
assign w7018 = w6975 & w6993;
assign w7019 = ~w7017 & ~w7018;
assign w7020 = w6984 & ~w7019;
assign w7021 = w7011 & w64743;
assign w7022 = ~w7020 & ~w7021;
assign w7023 = ~pi3274 & pi9040;
assign w7024 = ~pi3400 & ~pi9040;
assign w7025 = ~w7023 & ~w7024;
assign w7026 = pi0408 & ~w7025;
assign w7027 = ~pi0408 & w7025;
assign w7028 = ~w7026 & ~w7027;
assign w7029 = (w7016 & w64744) | (w7016 & w64745) | (w64744 & w64745);
assign w7030 = ~w6969 & w7001;
assign w7031 = ~w6982 & w7030;
assign w7032 = ~w7019 & w7031;
assign w7033 = ~w7016 & ~w7028;
assign w7034 = w6969 & w7001;
assign w7035 = w6975 & ~w6982;
assign w7036 = ~w6975 & w6982;
assign w7037 = w6993 & ~w7036;
assign w7038 = ~w7035 & ~w7037;
assign w7039 = (w7034 & w7037) | (w7034 & w64746) | (w7037 & w64746);
assign w7040 = w6969 & ~w6993;
assign w7041 = w6975 & w6982;
assign w7042 = w6993 & ~w7011;
assign w7043 = ~w6982 & ~w7001;
assign w7044 = ~w7028 & ~w7043;
assign w7045 = ~w7041 & ~w7044;
assign w7046 = w7042 & w7045;
assign w7047 = (w7039 & w7046) | (w7039 & w64747) | (w7046 & w64747);
assign w7048 = w7021 & w7036;
assign w7049 = ~w7032 & ~w7048;
assign w7050 = ~w7047 & w7049;
assign w7051 = ~w7033 & w7050;
assign w7052 = w7051 & w64748;
assign w7053 = (pi0429 & ~w7051) | (pi0429 & w64749) | (~w7051 & w64749);
assign w7054 = ~w7052 & ~w7053;
assign w7055 = ~w6969 & ~w7001;
assign w7056 = w6983 & w7055;
assign w7057 = ~w7001 & w7041;
assign w7058 = w6982 & w7001;
assign w7059 = ~w7010 & ~w7057;
assign w7060 = (~w6993 & ~w7059) | (~w6993 & w63582) | (~w7059 & w63582);
assign w7061 = w6987 & w7002;
assign w7062 = w7009 & ~w7056;
assign w7063 = ~w7060 & w7062;
assign w7064 = (~w7028 & ~w7063) | (~w7028 & w64750) | (~w7063 & w64750);
assign w7065 = w6982 & w7042;
assign w7066 = (~w7008 & ~w7042) | (~w7008 & w64751) | (~w7042 & w64751);
assign w7067 = ~w7001 & ~w7066;
assign w7068 = w7034 & ~w7041;
assign w7069 = w7019 & w7068;
assign w7070 = w7035 & ~w7040;
assign w7071 = ~w7001 & ~w7070;
assign w7072 = ~w7003 & ~w7071;
assign w7073 = ~w7048 & ~w7065;
assign w7074 = ~w7072 & w7073;
assign w7075 = w7028 & ~w7074;
assign w7076 = ~w7067 & ~w7069;
assign w7077 = ~w7064 & w7076;
assign w7078 = ~w7075 & w7077;
assign w7079 = pi0436 & ~w7078;
assign w7080 = ~pi0436 & w7078;
assign w7081 = ~w7079 & ~w7080;
assign w7082 = ~w6928 & w6930;
assign w7083 = w6886 & ~w6900;
assign w7084 = w6954 & w7083;
assign w7085 = ~w6909 & w6934;
assign w7086 = ~w6952 & w7085;
assign w7087 = w6880 & w6919;
assign w7088 = w6913 & ~w7087;
assign w7089 = ~w6880 & w6909;
assign w7090 = ~w7088 & ~w7089;
assign w7091 = ~w6886 & ~w7090;
assign w7092 = ~w6900 & ~w7086;
assign w7093 = ~w7091 & w7092;
assign w7094 = ~w6880 & ~w6919;
assign w7095 = ~w6893 & ~w7094;
assign w7096 = w6893 & ~w6919;
assign w7097 = w6912 & w7096;
assign w7098 = ~w7095 & ~w7097;
assign w7099 = w6886 & ~w7098;
assign w7100 = w6907 & w7087;
assign w7101 = w6908 & w7096;
assign w7102 = ~w6886 & ~w7096;
assign w7103 = ~w7095 & w7102;
assign w7104 = ~w7100 & ~w7101;
assign w7105 = ~w7103 & w7104;
assign w7106 = w6900 & ~w7099;
assign w7107 = w7105 & w7106;
assign w7108 = ~w7093 & ~w7107;
assign w7109 = ~w7082 & ~w7084;
assign w7110 = ~w7108 & w7109;
assign w7111 = pi0419 & ~w7110;
assign w7112 = ~pi0419 & w7110;
assign w7113 = ~w7111 & ~w7112;
assign w7114 = ~w6713 & ~w6722;
assign w7115 = w6660 & ~w7114;
assign w7116 = w6712 & w6729;
assign w7117 = ~w6694 & ~w6720;
assign w7118 = ~w7116 & w7117;
assign w7119 = ~w7115 & w7118;
assign w7120 = ~w6623 & ~w7119;
assign w7121 = ~w6685 & w6711;
assign w7122 = ~w6731 & ~w7121;
assign w7123 = w6623 & ~w7122;
assign w7124 = ~w6653 & ~w6664;
assign w7125 = ~w6660 & ~w7124;
assign w7126 = w7114 & w7125;
assign w7127 = ~w6670 & ~w7123;
assign w7128 = ~w7126 & w7127;
assign w7129 = ~w7120 & w7128;
assign w7130 = ~pi0424 & w7129;
assign w7131 = pi0424 & ~w7129;
assign w7132 = ~w7130 & ~w7131;
assign w7133 = ~pi3335 & pi9040;
assign w7134 = ~pi3289 & ~pi9040;
assign w7135 = ~w7133 & ~w7134;
assign w7136 = pi0408 & ~w7135;
assign w7137 = ~pi0408 & w7135;
assign w7138 = ~w7136 & ~w7137;
assign w7139 = ~pi3352 & pi9040;
assign w7140 = ~pi3321 & ~pi9040;
assign w7141 = ~w7139 & ~w7140;
assign w7142 = pi0397 & ~w7141;
assign w7143 = ~pi0397 & w7141;
assign w7144 = ~w7142 & ~w7143;
assign w7145 = w7138 & ~w7144;
assign w7146 = ~pi3355 & pi9040;
assign w7147 = ~pi3286 & ~pi9040;
assign w7148 = ~w7146 & ~w7147;
assign w7149 = pi0403 & ~w7148;
assign w7150 = ~pi0403 & w7148;
assign w7151 = ~w7149 & ~w7150;
assign w7152 = w7145 & w7151;
assign w7153 = ~w7138 & ~w7151;
assign w7154 = w7144 & w7153;
assign w7155 = ~w7138 & w7151;
assign w7156 = ~w7144 & w7155;
assign w7157 = ~w7154 & ~w7156;
assign w7158 = ~pi3291 & pi9040;
assign w7159 = ~pi3334 & ~pi9040;
assign w7160 = ~w7158 & ~w7159;
assign w7161 = pi0396 & ~w7160;
assign w7162 = ~pi0396 & w7160;
assign w7163 = ~w7161 & ~w7162;
assign w7164 = (w7163 & ~w7157) | (w7163 & w64752) | (~w7157 & w64752);
assign w7165 = ~w7151 & ~w7163;
assign w7166 = w7145 & w7165;
assign w7167 = ~w7164 & ~w7166;
assign w7168 = ~pi3280 & pi9040;
assign w7169 = ~pi3417 & ~pi9040;
assign w7170 = ~w7168 & ~w7169;
assign w7171 = pi0414 & ~w7170;
assign w7172 = ~pi0414 & w7170;
assign w7173 = ~w7171 & ~w7172;
assign w7174 = ~w7167 & w7173;
assign w7175 = w7138 & w7144;
assign w7176 = ~w7151 & w7175;
assign w7177 = ~w7144 & w7153;
assign w7178 = ~w7152 & ~w7177;
assign w7179 = (~w7176 & w7178) | (~w7176 & w64753) | (w7178 & w64753);
assign w7180 = w7144 & ~w7173;
assign w7181 = ~w7138 & w7180;
assign w7182 = ~w7152 & w7163;
assign w7183 = ~w7181 & w7182;
assign w7184 = ~w7179 & w7183;
assign w7185 = ~w7157 & w7173;
assign w7186 = ~w7163 & ~w7173;
assign w7187 = w7138 & w7186;
assign w7188 = ~pi3337 & pi9040;
assign w7189 = ~pi3288 & ~pi9040;
assign w7190 = ~w7188 & ~w7189;
assign w7191 = pi0391 & ~w7190;
assign w7192 = ~pi0391 & w7190;
assign w7193 = ~w7191 & ~w7192;
assign w7194 = ~w7187 & w7193;
assign w7195 = ~w7185 & w7194;
assign w7196 = ~w7184 & w7195;
assign w7197 = w7151 & ~w7173;
assign w7198 = w7163 & ~w7197;
assign w7199 = w7138 & w7173;
assign w7200 = w7198 & ~w7199;
assign w7201 = w7198 & w64754;
assign w7202 = w7173 & ~w7178;
assign w7203 = ~w7138 & w7197;
assign w7204 = ~w7176 & ~w7203;
assign w7205 = ~w7181 & w7204;
assign w7206 = ~w7198 & ~w7205;
assign w7207 = w7144 & ~w7163;
assign w7208 = w7155 & w7207;
assign w7209 = ~w7193 & ~w7208;
assign w7210 = ~w7201 & w7209;
assign w7211 = ~w7202 & w7210;
assign w7212 = ~w7206 & w7211;
assign w7213 = ~w7196 & ~w7212;
assign w7214 = w7175 & ~w7193;
assign w7215 = ~w7181 & ~w7214;
assign w7216 = w7151 & w7163;
assign w7217 = ~w7215 & w7216;
assign w7218 = ~w7174 & ~w7217;
assign w7219 = ~w7213 & w7218;
assign w7220 = pi0427 & ~w7219;
assign w7221 = ~pi0427 & w7219;
assign w7222 = ~w7220 & ~w7221;
assign w7223 = ~w7163 & w7185;
assign w7224 = ~w7151 & w7173;
assign w7225 = ~w7197 & ~w7224;
assign w7226 = w7163 & w7173;
assign w7227 = w7175 & ~w7226;
assign w7228 = w7225 & ~w7227;
assign w7229 = ~w7145 & ~w7225;
assign w7230 = ~w7228 & ~w7229;
assign w7231 = (w7157 & w7230) | (w7157 & w63583) | (w7230 & w63583);
assign w7232 = w7186 & w7231;
assign w7233 = ~w7144 & ~w7152;
assign w7234 = w7173 & w7175;
assign w7235 = (w7163 & ~w7153) | (w7163 & w63584) | (~w7153 & w63584);
assign w7236 = ~w7203 & ~w7234;
assign w7237 = w7235 & w7236;
assign w7238 = ~w7233 & w7237;
assign w7239 = ~w7230 & ~w7238;
assign w7240 = ~w7232 & w7239;
assign w7241 = w7193 & ~w7240;
assign w7242 = (~w7193 & ~w7236) | (~w7193 & w63585) | (~w7236 & w63585);
assign w7243 = ~w7178 & ~w7225;
assign w7244 = ~w7242 & ~w7243;
assign w7245 = w7163 & ~w7244;
assign w7246 = ~w7231 & w7242;
assign w7247 = ~w7223 & ~w7245;
assign w7248 = ~w7246 & w7247;
assign w7249 = ~w7241 & w7248;
assign w7250 = pi0437 & ~w7249;
assign w7251 = ~pi0437 & w7249;
assign w7252 = ~w7250 & ~w7251;
assign w7253 = w6550 & w6580;
assign w7254 = w6544 & w6596;
assign w7255 = ~w6573 & ~w7254;
assign w7256 = ~w6529 & w6551;
assign w7257 = (~w7256 & ~w7255) | (~w7256 & w63362) | (~w7255 & w63362);
assign w7258 = ~w6565 & ~w7257;
assign w7259 = ~w6554 & w6606;
assign w7260 = w6544 & w6568;
assign w7261 = w6565 & ~w7260;
assign w7262 = w7259 & w7261;
assign w7263 = ~w7258 & ~w7262;
assign w7264 = ~w6575 & w63363;
assign w7265 = w7263 & w7264;
assign w7266 = (w6588 & w7265) | (w6588 & w63586) | (w7265 & w63586);
assign w7267 = ~w6607 & w64755;
assign w7268 = ~w6573 & ~w7259;
assign w7269 = (~w6588 & w7259) | (~w6588 & w64756) | (w7259 & w64756);
assign w7270 = ~w7267 & ~w7269;
assign w7271 = w6565 & ~w7270;
assign w7272 = ~w6537 & w6588;
assign w7273 = ~w6536 & w6565;
assign w7274 = ~w6588 & w7273;
assign w7275 = w6571 & ~w7272;
assign w7276 = ~w7274 & w7275;
assign w7277 = ~w6579 & ~w6599;
assign w7278 = ~w6565 & ~w7277;
assign w7279 = w7268 & w7278;
assign w7280 = ~w7276 & ~w7279;
assign w7281 = ~w7271 & w7280;
assign w7282 = (pi0445 & w7266) | (pi0445 & w64757) | (w7266 & w64757);
assign w7283 = ~w7266 & w64758;
assign w7284 = ~w7282 & ~w7283;
assign w7285 = ~w6594 & ~w7256;
assign w7286 = w7263 & ~w7285;
assign w7287 = ~w6551 & ~w7260;
assign w7288 = w6538 & ~w7287;
assign w7289 = w6557 & w6565;
assign w7290 = ~w7253 & w7289;
assign w7291 = (w6588 & ~w6591) | (w6588 & w64759) | (~w6591 & w64759);
assign w7292 = ~w7288 & w7291;
assign w7293 = ~w7290 & w7292;
assign w7294 = w6570 & w6590;
assign w7295 = ~w6535 & ~w6550;
assign w7296 = w6579 & w7295;
assign w7297 = ~w6588 & ~w7296;
assign w7298 = ~w7294 & w7297;
assign w7299 = w6602 & w7298;
assign w7300 = ~w7293 & ~w7299;
assign w7301 = ~w7286 & ~w7300;
assign w7302 = ~pi0447 & w7301;
assign w7303 = pi0447 & ~w7301;
assign w7304 = ~w7302 & ~w7303;
assign w7305 = ~w7030 & w7035;
assign w7306 = (~w7055 & w7305) | (~w7055 & w63587) | (w7305 & w63587);
assign w7307 = (w6993 & w7306) | (w6993 & w64760) | (w7306 & w64760);
assign w7308 = w7006 & w7017;
assign w7309 = ~w7030 & ~w7040;
assign w7310 = w6983 & ~w7309;
assign w7311 = ~w7307 & ~w7310;
assign w7312 = (w7028 & w7308) | (w7028 & w64761) | (w7308 & w64761);
assign w7313 = w7040 & w7057;
assign w7314 = ~w7043 & ~w7058;
assign w7315 = w7012 & ~w7314;
assign w7316 = (w6982 & w7011) | (w6982 & w63361) | (w7011 & w63361);
assign w7317 = w7055 & ~w7316;
assign w7318 = w7011 & w64762;
assign w7319 = ~w7039 & ~w7318;
assign w7320 = ~w7317 & w7319;
assign w7321 = ~w7028 & ~w7320;
assign w7322 = ~w7313 & ~w7315;
assign w7323 = ~w7321 & w7322;
assign w7324 = ~w7312 & w7323;
assign w7325 = ~pi0432 & w7324;
assign w7326 = pi0432 & ~w7324;
assign w7327 = ~w7325 & ~w7326;
assign w7328 = ~pi3304 & pi9040;
assign w7329 = ~pi3306 & ~pi9040;
assign w7330 = ~w7328 & ~w7329;
assign w7331 = pi0376 & ~w7330;
assign w7332 = ~pi0376 & w7330;
assign w7333 = ~w7331 & ~w7332;
assign w7334 = ~pi3297 & pi9040;
assign w7335 = ~pi3386 & ~pi9040;
assign w7336 = ~w7334 & ~w7335;
assign w7337 = pi0404 & ~w7336;
assign w7338 = ~pi0404 & w7336;
assign w7339 = ~w7337 & ~w7338;
assign w7340 = w7333 & ~w7339;
assign w7341 = ~pi3281 & pi9040;
assign w7342 = ~pi3275 & ~pi9040;
assign w7343 = ~w7341 & ~w7342;
assign w7344 = pi0412 & ~w7343;
assign w7345 = ~pi0412 & w7343;
assign w7346 = ~w7344 & ~w7345;
assign w7347 = ~w7340 & ~w7346;
assign w7348 = ~pi3341 & pi9040;
assign w7349 = ~pi3312 & ~pi9040;
assign w7350 = ~w7348 & ~w7349;
assign w7351 = pi0413 & ~w7350;
assign w7352 = ~pi0413 & w7350;
assign w7353 = ~w7351 & ~w7352;
assign w7354 = ~w7339 & ~w7353;
assign w7355 = ~w7333 & w7339;
assign w7356 = ~w7333 & ~w7353;
assign w7357 = ~pi3275 & pi9040;
assign w7358 = ~pi3319 & ~pi9040;
assign w7359 = ~w7357 & ~w7358;
assign w7360 = pi0399 & ~w7359;
assign w7361 = ~pi0399 & w7359;
assign w7362 = ~w7360 & ~w7361;
assign w7363 = w7356 & ~w7362;
assign w7364 = ~pi3316 & pi9040;
assign w7365 = ~pi3338 & ~pi9040;
assign w7366 = ~w7364 & ~w7365;
assign w7367 = pi0386 & ~w7366;
assign w7368 = ~pi0386 & w7366;
assign w7369 = ~w7367 & ~w7368;
assign w7370 = (~w7369 & w7363) | (~w7369 & w64763) | (w7363 & w64763);
assign w7371 = ~w7354 & w7370;
assign w7372 = w7339 & w7353;
assign w7373 = ~w7355 & w7362;
assign w7374 = ~w7372 & w7373;
assign w7375 = ~w7371 & ~w7374;
assign w7376 = w7347 & ~w7375;
assign w7377 = w7339 & ~w7362;
assign w7378 = w7353 & w7355;
assign w7379 = ~w7346 & ~w7378;
assign w7380 = w7377 & ~w7379;
assign w7381 = ~w7339 & w7362;
assign w7382 = w7353 & w7381;
assign w7383 = w7381 & w7384;
assign w7384 = ~w7333 & w7353;
assign w7385 = ~w7353 & w7362;
assign w7386 = ~w7339 & ~w7384;
assign w7387 = ~w7385 & w7386;
assign w7388 = ~w7346 & w7387;
assign w7389 = w7333 & w7346;
assign w7390 = w7372 & w7389;
assign w7391 = ~w7340 & ~w7355;
assign w7392 = ~w7353 & ~w7391;
assign w7393 = w7333 & ~w7362;
assign w7394 = w7354 & w7393;
assign w7395 = w7346 & ~w7394;
assign w7396 = w7392 & w7395;
assign w7397 = w7369 & ~w7390;
assign w7398 = ~w7383 & w7397;
assign w7399 = ~w7380 & w7398;
assign w7400 = ~w7388 & ~w7396;
assign w7401 = w7399 & w7400;
assign w7402 = w7339 & w7362;
assign w7403 = w7333 & ~w7353;
assign w7404 = ~w7384 & ~w7403;
assign w7405 = w7402 & ~w7404;
assign w7406 = w7346 & w7387;
assign w7407 = w7356 & w7381;
assign w7408 = ~w7369 & ~w7407;
assign w7409 = ~w7405 & w7408;
assign w7410 = ~w7406 & w7409;
assign w7411 = ~w7401 & ~w7410;
assign w7412 = ~w7376 & ~w7411;
assign w7413 = ~pi0416 & w7412;
assign w7414 = pi0416 & ~w7412;
assign w7415 = ~w7413 & ~w7414;
assign w7416 = ~w7163 & ~w7204;
assign w7417 = (~w7230 & w63588) | (~w7230 & w63589) | (w63588 & w63589);
assign w7418 = w7144 & ~w7153;
assign w7419 = w7200 & ~w7418;
assign w7420 = ~w7416 & ~w7419;
assign w7421 = ~w7417 & w7420;
assign w7422 = w7193 & ~w7421;
assign w7423 = ~w7178 & w7226;
assign w7424 = ~w7166 & ~w7227;
assign w7425 = ~w7225 & ~w7424;
assign w7426 = ~w7154 & w7193;
assign w7427 = ~w7173 & ~w7426;
assign w7428 = w7164 & w7427;
assign w7429 = ~w7193 & w7228;
assign w7430 = w7421 & w7429;
assign w7431 = ~w7423 & ~w7425;
assign w7432 = ~w7428 & w7431;
assign w7433 = ~w7422 & w7432;
assign w7434 = (pi0431 & ~w7433) | (pi0431 & w64764) | (~w7433 & w64764);
assign w7435 = w7433 & w64765;
assign w7436 = ~w7434 & ~w7435;
assign w7437 = ~w7087 & ~w7094;
assign w7438 = ~w6959 & ~w7437;
assign w7439 = w6930 & w7088;
assign w7440 = ~w6948 & ~w6953;
assign w7441 = ~w7105 & ~w7440;
assign w7442 = w6952 & ~w7437;
assign w7443 = w6911 & w7098;
assign w7444 = w6919 & w6924;
assign w7445 = ~w7088 & w7444;
assign w7446 = ~w6900 & ~w7442;
assign w7447 = ~w7445 & w7446;
assign w7448 = ~w7443 & w7447;
assign w7449 = ~w6952 & w64766;
assign w7450 = w6923 & w7444;
assign w7451 = w6900 & ~w7097;
assign w7452 = ~w7450 & w7451;
assign w7453 = ~w7449 & w7452;
assign w7454 = w6937 & w7453;
assign w7455 = ~w7448 & ~w7454;
assign w7456 = ~w7439 & ~w7441;
assign w7457 = ~w7455 & w7456;
assign w7458 = w7457 & w64767;
assign w7459 = (pi0426 & ~w7457) | (pi0426 & w64768) | (~w7457 & w64768);
assign w7460 = ~w7458 & ~w7459;
assign w7461 = ~pi3380 & pi9040;
assign w7462 = ~pi3301 & ~pi9040;
assign w7463 = ~w7461 & ~w7462;
assign w7464 = pi0395 & ~w7463;
assign w7465 = ~pi0395 & w7463;
assign w7466 = ~w7464 & ~w7465;
assign w7467 = ~pi3299 & pi9040;
assign w7468 = ~pi3276 & ~pi9040;
assign w7469 = ~w7467 & ~w7468;
assign w7470 = pi0409 & ~w7469;
assign w7471 = ~pi0409 & w7469;
assign w7472 = ~w7470 & ~w7471;
assign w7473 = ~pi3312 & pi9040;
assign w7474 = ~pi3304 & ~pi9040;
assign w7475 = ~w7473 & ~w7474;
assign w7476 = pi0413 & ~w7475;
assign w7477 = ~pi0413 & w7475;
assign w7478 = ~w7476 & ~w7477;
assign w7479 = w7472 & ~w7478;
assign w7480 = ~pi3278 & pi9040;
assign w7481 = ~pi3279 & ~pi9040;
assign w7482 = ~w7480 & ~w7481;
assign w7483 = pi0386 & ~w7482;
assign w7484 = ~pi0386 & w7482;
assign w7485 = ~w7483 & ~w7484;
assign w7486 = ~w7472 & ~w7485;
assign w7487 = ~pi3386 & pi9040;
assign w7488 = ~pi3316 & ~pi9040;
assign w7489 = ~w7487 & ~w7488;
assign w7490 = pi0393 & ~w7489;
assign w7491 = ~pi0393 & w7489;
assign w7492 = ~w7490 & ~w7491;
assign w7493 = ~w7485 & ~w7492;
assign w7494 = ~w7486 & ~w7493;
assign w7495 = ~w7472 & w7478;
assign w7496 = w7485 & ~w7495;
assign w7497 = w7494 & ~w7496;
assign w7498 = ~pi3279 & pi9040;
assign w7499 = ~pi3274 & ~pi9040;
assign w7500 = ~w7498 & ~w7499;
assign w7501 = pi0388 & ~w7500;
assign w7502 = ~pi0388 & w7500;
assign w7503 = ~w7501 & ~w7502;
assign w7504 = (w7503 & w7497) | (w7503 & w63590) | (w7497 & w63590);
assign w7505 = w7478 & w7486;
assign w7506 = w7492 & w7505;
assign w7507 = ~w7486 & ~w7503;
assign w7508 = ~w7497 & w64769;
assign w7509 = ~w7504 & ~w7506;
assign w7510 = (w7466 & ~w7509) | (w7466 & w64770) | (~w7509 & w64770);
assign w7511 = w7479 & w7492;
assign w7512 = ~w7478 & ~w7492;
assign w7513 = w7486 & w7512;
assign w7514 = ~w7511 & ~w7513;
assign w7515 = w7503 & ~w7514;
assign w7516 = w7472 & w7485;
assign w7517 = ~w7486 & ~w7516;
assign w7518 = ~w7485 & w7503;
assign w7519 = w7517 & w63591;
assign w7520 = w7478 & ~w7492;
assign w7521 = (w7520 & ~w7517) | (w7520 & w64771) | (~w7517 & w64771);
assign w7522 = ~w7519 & ~w7521;
assign w7523 = w7478 & w7492;
assign w7524 = ~w7516 & w7523;
assign w7525 = w7472 & w7524;
assign w7526 = ~w7503 & w7525;
assign w7527 = ~w7472 & ~w7492;
assign w7528 = ~w7479 & ~w7527;
assign w7529 = ~w7485 & ~w7528;
assign w7530 = w7478 & w7516;
assign w7531 = ~w7478 & ~w7516;
assign w7532 = ~w7530 & ~w7531;
assign w7533 = ~w7486 & ~w7532;
assign w7534 = ~w7478 & ~w7485;
assign w7535 = w7485 & w7492;
assign w7536 = ~w7534 & ~w7535;
assign w7537 = ~w7529 & ~w7536;
assign w7538 = ~w7533 & w7537;
assign w7539 = w7522 & ~w7526;
assign w7540 = ~w7538 & w7539;
assign w7541 = ~w7466 & ~w7540;
assign w7542 = ~w7510 & ~w7515;
assign w7543 = ~w7541 & w7542;
assign w7544 = pi0444 & w7543;
assign w7545 = ~pi0444 & ~w7543;
assign w7546 = ~w7544 & ~w7545;
assign w7547 = w6768 & ~w6776;
assign w7548 = w6827 & w6829;
assign w7549 = ~w6800 & w6812;
assign w7550 = ~w7548 & ~w7549;
assign w7551 = ~w6801 & w7550;
assign w7552 = w7547 & ~w7551;
assign w7553 = ~w6753 & ~w6813;
assign w7554 = ~w6762 & ~w6829;
assign w7555 = ~w6800 & ~w7554;
assign w7556 = w6777 & ~w7553;
assign w7557 = ~w7555 & w7556;
assign w7558 = ~w6777 & ~w7547;
assign w7559 = ~w6793 & w7558;
assign w7560 = ~w6802 & w7559;
assign w7561 = ~w7557 & ~w7560;
assign w7562 = w7550 & ~w7561;
assign w7563 = ~w7552 & ~w7562;
assign w7564 = ~pi0452 & w7563;
assign w7565 = pi0452 & ~w7563;
assign w7566 = ~w7564 & ~w7565;
assign w7567 = ~w7494 & ~w7527;
assign w7568 = ~w7519 & ~w7567;
assign w7569 = w7503 & ~w7568;
assign w7570 = ~w7522 & w7569;
assign w7571 = ~w7478 & w7535;
assign w7572 = ~w7472 & w7571;
assign w7573 = w7512 & ~w7517;
assign w7574 = ~w7497 & ~w7573;
assign w7575 = ~w7503 & w7574;
assign w7576 = w7503 & ~w7505;
assign w7577 = ~w7567 & ~w7571;
assign w7578 = w7576 & w7577;
assign w7579 = ~w7575 & ~w7578;
assign w7580 = ~w7572 & ~w7579;
assign w7581 = (~w7466 & w7579) | (~w7466 & w63592) | (w7579 & w63592);
assign w7582 = (~w7503 & w7529) | (~w7503 & w64772) | (w7529 & w64772);
assign w7583 = w7520 & ~w7582;
assign w7584 = w7466 & ~w7583;
assign w7585 = w7580 & w7584;
assign w7586 = w7523 & w7582;
assign w7587 = ~w7570 & ~w7586;
assign w7588 = ~w7581 & w7587;
assign w7589 = ~w7585 & w7588;
assign w7590 = pi0434 & ~w7589;
assign w7591 = ~pi0434 & w7589;
assign w7592 = ~w7590 & ~w7591;
assign w7593 = w6969 & w7028;
assign w7594 = w7038 & w7593;
assign w7595 = ~w7001 & ~w7594;
assign w7596 = ~w7031 & ~w7034;
assign w7597 = (w7028 & w7596) | (w7028 & w64773) | (w7596 & w64773);
assign w7598 = (~w7007 & ~w7042) | (~w7007 & w64774) | (~w7042 & w64774);
assign w7599 = ~w7597 & w7598;
assign w7600 = ~w7595 & ~w7599;
assign w7601 = w7041 & w7055;
assign w7602 = (~w7305 & w7596) | (~w7305 & w64775) | (w7596 & w64775);
assign w7603 = w7004 & ~w7602;
assign w7604 = w7018 & w7031;
assign w7605 = ~w7020 & ~w7601;
assign w7606 = ~w7604 & w7605;
assign w7607 = ~w7603 & w7606;
assign w7608 = ~w7028 & ~w7607;
assign w7609 = ~w7046 & ~w7600;
assign w7610 = ~w7608 & w7609;
assign w7611 = pi0441 & ~w7610;
assign w7612 = ~pi0441 & w7610;
assign w7613 = ~w7611 & ~w7612;
assign w7614 = ~w7384 & ~w7402;
assign w7615 = w7379 & ~w7614;
assign w7616 = ~w7355 & ~w7404;
assign w7617 = ~w7362 & w7616;
assign w7618 = ~w7333 & w7362;
assign w7619 = w7372 & w7618;
assign w7620 = w7346 & w7619;
assign w7621 = ~w7615 & ~w7620;
assign w7622 = ~w7617 & w7621;
assign w7623 = ~w7369 & ~w7622;
assign w7624 = ~w7381 & w7389;
assign w7625 = w7377 & w7404;
assign w7626 = ~w7354 & ~w7619;
assign w7627 = ~w7346 & ~w7393;
assign w7628 = ~w7626 & w7627;
assign w7629 = ~w7624 & ~w7625;
assign w7630 = ~w7628 & w7629;
assign w7631 = w7369 & ~w7630;
assign w7632 = ~w7339 & ~w7389;
assign w7633 = w7369 & ~w7632;
assign w7634 = w7381 & w64776;
assign w7635 = ~w7346 & ~w7362;
assign w7636 = w7384 & w7635;
assign w7637 = ~w7634 & ~w7636;
assign w7638 = ~w7633 & ~w7637;
assign w7639 = w7346 & ~w7363;
assign w7640 = ~w7340 & w7614;
assign w7641 = w7639 & w7640;
assign w7642 = ~w7638 & ~w7641;
assign w7643 = ~w7631 & w7642;
assign w7644 = ~w7623 & w7643;
assign w7645 = pi0423 & ~w7644;
assign w7646 = ~pi0423 & w7644;
assign w7647 = ~w7645 & ~w7646;
assign w7648 = w7353 & w7377;
assign w7649 = (w7333 & w7405) | (w7333 & w64777) | (w7405 & w64777);
assign w7650 = ~w7383 & ~w7392;
assign w7651 = w7370 & ~w7650;
assign w7652 = (~w7346 & w7651) | (~w7346 & w64778) | (w7651 & w64778);
assign w7653 = ~w7377 & w7403;
assign w7654 = ~w7347 & ~w7369;
assign w7655 = ~w7382 & ~w7653;
assign w7656 = w7654 & w7655;
assign w7657 = ~w7625 & w7656;
assign w7658 = ~w7382 & w7639;
assign w7659 = w7356 & w7362;
assign w7660 = w7379 & ~w7659;
assign w7661 = ~w7658 & ~w7660;
assign w7662 = ~w7394 & w7637;
assign w7663 = ~w7649 & w7662;
assign w7664 = ~w7661 & w7663;
assign w7665 = w7369 & ~w7664;
assign w7666 = ~w7652 & ~w7657;
assign w7667 = ~w7665 & w7666;
assign w7668 = pi0425 & w7667;
assign w7669 = ~pi0425 & ~w7667;
assign w7670 = ~w7668 & ~w7669;
assign w7671 = w6565 & w7295;
assign w7672 = w6529 & w7671;
assign w7673 = ~w6572 & ~w7267;
assign w7674 = (w6588 & ~w7263) | (w6588 & w64779) | (~w7263 & w64779);
assign w7675 = w6595 & ~w7260;
assign w7676 = ~w6536 & w64780;
assign w7677 = ~w7671 & ~w7676;
assign w7678 = ~w7675 & ~w7677;
assign w7679 = w6529 & ~w7255;
assign w7680 = ~w6600 & ~w7679;
assign w7681 = (~w6588 & ~w7680) | (~w6588 & w64781) | (~w7680 & w64781);
assign w7682 = w6558 & ~w6565;
assign w7683 = ~w7672 & ~w7682;
assign w7684 = ~w6593 & w7683;
assign w7685 = ~w7681 & w7684;
assign w7686 = ~w7674 & w7685;
assign w7687 = pi0449 & ~w7686;
assign w7688 = ~pi0449 & w7686;
assign w7689 = ~w7687 & ~w7688;
assign w7690 = ~w7495 & w7535;
assign w7691 = w7503 & ~w7690;
assign w7692 = w7538 & w7691;
assign w7693 = ~w7503 & w7571;
assign w7694 = w7495 & w7518;
assign w7695 = (~w7694 & w7532) | (~w7694 & w64782) | (w7532 & w64782);
assign w7696 = ~w7492 & ~w7695;
assign w7697 = ~w7472 & ~w7503;
assign w7698 = ~w7493 & ~w7535;
assign w7699 = w7697 & w7698;
assign w7700 = w7466 & ~w7525;
assign w7701 = ~w7699 & w7700;
assign w7702 = ~w7696 & w7701;
assign w7703 = w7532 & w7576;
assign w7704 = ~w7466 & ~w7513;
assign w7705 = ~w7703 & w7704;
assign w7706 = ~w7582 & w7705;
assign w7707 = ~w7702 & ~w7706;
assign w7708 = ~w7692 & ~w7693;
assign w7709 = ~w7707 & w7708;
assign w7710 = pi0428 & ~w7709;
assign w7711 = ~pi0428 & w7709;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = w7523 & w7697;
assign w7714 = ~w7466 & ~w7713;
assign w7715 = (~w7524 & w7568) | (~w7524 & w64783) | (w7568 & w64783);
assign w7716 = ~w7714 & ~w7715;
assign w7717 = ~w7466 & ~w7478;
assign w7718 = ~w7574 & w7717;
assign w7719 = w7466 & ~w7511;
assign w7720 = (~w7503 & ~w7536) | (~w7503 & w64784) | (~w7536 & w64784);
assign w7721 = w7478 & w7527;
assign w7722 = w7691 & ~w7721;
assign w7723 = ~w7719 & ~w7720;
assign w7724 = ~w7722 & w7723;
assign w7725 = ~w7534 & w7720;
assign w7726 = w7584 & w7725;
assign w7727 = ~w7718 & ~w7724;
assign w7728 = ~w7716 & w7727;
assign w7729 = ~w7726 & w7728;
assign w7730 = pi0438 & ~w7729;
assign w7731 = ~pi0438 & w7729;
assign w7732 = ~w7730 & ~w7731;
assign w7733 = w7154 & w7226;
assign w7734 = w7138 & w7180;
assign w7735 = ~w7163 & ~w7734;
assign w7736 = ~w7179 & w7735;
assign w7737 = ~w7145 & ~w7180;
assign w7738 = ~w7163 & ~w7176;
assign w7739 = ~w7737 & w7738;
assign w7740 = ~w7145 & w7224;
assign w7741 = w7183 & ~w7740;
assign w7742 = ~w7193 & ~w7739;
assign w7743 = ~w7741 & w7742;
assign w7744 = ~w7156 & ~w7734;
assign w7745 = w7163 & ~w7744;
assign w7746 = w7138 & ~w7225;
assign w7747 = w7179 & w7746;
assign w7748 = ~w7208 & ~w7745;
assign w7749 = ~w7747 & w7748;
assign w7750 = w7193 & ~w7749;
assign w7751 = ~w7201 & ~w7733;
assign w7752 = ~w7736 & w7751;
assign w7753 = ~w7743 & w7752;
assign w7754 = ~w7750 & w7753;
assign w7755 = pi0439 & ~w7754;
assign w7756 = ~pi0439 & w7754;
assign w7757 = ~w7755 & ~w7756;
assign w7758 = w6901 & ~w7100;
assign w7759 = ~w6909 & ~w6920;
assign w7760 = w7437 & ~w7759;
assign w7761 = w6910 & w6932;
assign w7762 = ~w6952 & w7083;
assign w7763 = ~w7101 & w7762;
assign w7764 = ~w7760 & ~w7761;
assign w7765 = ~w7763 & w7764;
assign w7766 = ~w7758 & ~w7765;
assign w7767 = ~w6923 & ~w6931;
assign w7768 = w6941 & ~w7767;
assign w7769 = (~w7101 & w6955) | (~w7101 & w64785) | (w6955 & w64785);
assign w7770 = ~w7768 & w7769;
assign w7771 = w6900 & ~w7770;
assign w7772 = ~w7766 & ~w7771;
assign w7773 = ~pi0417 & w7772;
assign w7774 = pi0417 & ~w7772;
assign w7775 = ~w7773 & ~w7774;
assign w7776 = w6794 & w64786;
assign w7777 = ~w6747 & w6798;
assign w7778 = w6828 & ~w7777;
assign w7779 = w6806 & ~w7778;
assign w7780 = w6844 & w7550;
assign w7781 = ~w6768 & w6831;
assign w7782 = ~w7777 & w7781;
assign w7783 = ~w7779 & ~w7782;
assign w7784 = ~w7780 & w7783;
assign w7785 = ~w6776 & ~w7784;
assign w7786 = w6835 & ~w7548;
assign w7787 = w6777 & ~w7786;
assign w7788 = w6769 & ~w6786;
assign w7789 = ~w6776 & w6830;
assign w7790 = ~w7788 & ~w7789;
assign w7791 = ~w6756 & ~w7790;
assign w7792 = ~w6812 & ~w7778;
assign w7793 = ~w6833 & w6845;
assign w7794 = ~w7792 & w7793;
assign w7795 = ~w7776 & ~w7791;
assign w7796 = ~w7794 & w7795;
assign w7797 = ~w7787 & w7796;
assign w7798 = ~w7785 & w7797;
assign w7799 = pi0458 & ~w7798;
assign w7800 = ~pi0458 & w7798;
assign w7801 = ~w7799 & ~w7800;
assign w7802 = w7346 & w7394;
assign w7803 = w7346 & w7616;
assign w7804 = ~w7392 & ~w7648;
assign w7805 = w7347 & ~w7804;
assign w7806 = ~w7407 & ~w7803;
assign w7807 = ~w7805 & w7806;
assign w7808 = w7369 & ~w7807;
assign w7809 = ~w7356 & ~w7632;
assign w7810 = ~w7393 & ~w7618;
assign w7811 = ~w7809 & w7810;
assign w7812 = ~w7390 & ~w7405;
assign w7813 = ~w7811 & w7812;
assign w7814 = ~w7369 & ~w7813;
assign w7815 = w7346 & ~w7402;
assign w7816 = ~w7347 & w7353;
assign w7817 = ~w7815 & w7816;
assign w7818 = ~w7802 & ~w7817;
assign w7819 = ~w7814 & w7818;
assign w7820 = ~w7808 & w7819;
assign w7821 = pi0454 & w7820;
assign w7822 = ~pi0454 & ~w7820;
assign w7823 = ~w7821 & ~w7822;
assign w7824 = ~pi3418 & pi9040;
assign w7825 = ~pi3411 & ~pi9040;
assign w7826 = ~w7824 & ~w7825;
assign w7827 = pi0443 & ~w7826;
assign w7828 = ~pi0443 & w7826;
assign w7829 = ~w7827 & ~w7828;
assign w7830 = ~pi3412 & pi9040;
assign w7831 = ~pi3373 & ~pi9040;
assign w7832 = ~w7830 & ~w7831;
assign w7833 = pi0469 & ~w7832;
assign w7834 = ~pi0469 & w7832;
assign w7835 = ~w7833 & ~w7834;
assign w7836 = w7829 & ~w7835;
assign w7837 = ~w7829 & w7835;
assign w7838 = ~w7836 & ~w7837;
assign w7839 = ~pi3372 & pi9040;
assign w7840 = ~pi3395 & ~pi9040;
assign w7841 = ~w7839 & ~w7840;
assign w7842 = pi0450 & ~w7841;
assign w7843 = ~pi0450 & w7841;
assign w7844 = ~w7842 & ~w7843;
assign w7845 = ~pi3396 & pi9040;
assign w7846 = ~pi3464 & ~pi9040;
assign w7847 = ~w7845 & ~w7846;
assign w7848 = pi0473 & ~w7847;
assign w7849 = ~pi0473 & w7847;
assign w7850 = ~w7848 & ~w7849;
assign w7851 = ~w7844 & w7850;
assign w7852 = ~w7838 & w7851;
assign w7853 = w7844 & ~w7850;
assign w7854 = w7837 & w7853;
assign w7855 = ~w7829 & ~w7844;
assign w7856 = ~w7835 & ~w7850;
assign w7857 = w7855 & w7856;
assign w7858 = ~w7854 & ~w7857;
assign w7859 = ~w7852 & w7858;
assign w7860 = ~w7835 & w7851;
assign w7861 = w7835 & ~w7850;
assign w7862 = w7829 & ~w7844;
assign w7863 = w7861 & w7862;
assign w7864 = ~w7860 & ~w7863;
assign w7865 = ~pi3383 & pi9040;
assign w7866 = pi3361 & ~pi9040;
assign w7867 = ~w7865 & ~w7866;
assign w7868 = pi0479 & ~w7867;
assign w7869 = ~pi0479 & w7867;
assign w7870 = ~w7868 & ~w7869;
assign w7871 = ~w7864 & ~w7870;
assign w7872 = w7859 & ~w7871;
assign w7873 = ~pi3480 & pi9040;
assign w7874 = ~pi3415 & ~pi9040;
assign w7875 = ~w7873 & ~w7874;
assign w7876 = pi0440 & ~w7875;
assign w7877 = ~pi0440 & w7875;
assign w7878 = ~w7876 & ~w7877;
assign w7879 = ~w7872 & w7878;
assign w7880 = ~w7829 & ~w7878;
assign w7881 = w7861 & w7880;
assign w7882 = w7829 & w7853;
assign w7883 = ~w7835 & w7855;
assign w7884 = ~w7882 & ~w7883;
assign w7885 = w7878 & w7884;
assign w7886 = (w7836 & ~w7884) | (w7836 & w64787) | (~w7884 & w64787);
assign w7887 = w7844 & w7850;
assign w7888 = w7829 & w7835;
assign w7889 = w7878 & ~w7888;
assign w7890 = w7887 & ~w7889;
assign w7891 = ~w7881 & ~w7890;
assign w7892 = ~w7886 & w7891;
assign w7893 = ~w7870 & w7892;
assign w7894 = ~w7844 & ~w7878;
assign w7895 = w7838 & w7894;
assign w7896 = w7853 & w7878;
assign w7897 = ~w7836 & ~w7896;
assign w7898 = ~w7886 & ~w7897;
assign w7899 = w7837 & w7887;
assign w7900 = w7870 & ~w7899;
assign w7901 = ~w7895 & w7900;
assign w7902 = ~w7898 & w7901;
assign w7903 = ~w7893 & ~w7902;
assign w7904 = w7829 & ~w7878;
assign w7905 = w7851 & w7888;
assign w7906 = (w7904 & w7905) | (w7904 & w64788) | (w7905 & w64788);
assign w7907 = w7853 & w7906;
assign w7908 = ~w7879 & ~w7907;
assign w7909 = ~w7903 & w7908;
assign w7910 = ~pi0480 & ~w7909;
assign w7911 = pi0480 & w7909;
assign w7912 = ~w7910 & ~w7911;
assign w7913 = ~pi3409 & pi9040;
assign w7914 = ~pi3412 & ~pi9040;
assign w7915 = ~w7913 & ~w7914;
assign w7916 = pi0453 & ~w7915;
assign w7917 = ~pi0453 & w7915;
assign w7918 = ~w7916 & ~w7917;
assign w7919 = ~pi3368 & pi9040;
assign w7920 = ~pi3409 & ~pi9040;
assign w7921 = ~w7919 & ~w7920;
assign w7922 = pi0476 & ~w7921;
assign w7923 = ~pi0476 & w7921;
assign w7924 = ~w7922 & ~w7923;
assign w7925 = w7918 & w7924;
assign w7926 = ~pi3411 & pi9040;
assign w7927 = ~pi3392 & ~pi9040;
assign w7928 = ~w7926 & ~w7927;
assign w7929 = pi0462 & ~w7928;
assign w7930 = ~pi0462 & w7928;
assign w7931 = ~w7929 & ~w7930;
assign w7932 = ~pi3393 & pi9040;
assign w7933 = ~pi3413 & ~pi9040;
assign w7934 = ~w7932 & ~w7933;
assign w7935 = pi0457 & ~w7934;
assign w7936 = ~pi0457 & w7934;
assign w7937 = ~w7935 & ~w7936;
assign w7938 = ~w7931 & w7937;
assign w7939 = w7925 & w7938;
assign w7940 = ~pi3419 & pi9040;
assign w7941 = ~pi3458 & ~pi9040;
assign w7942 = ~w7940 & ~w7941;
assign w7943 = pi0461 & ~w7942;
assign w7944 = ~pi0461 & w7942;
assign w7945 = ~w7943 & ~w7944;
assign w7946 = ~pi3371 & pi9040;
assign w7947 = ~pi3398 & ~pi9040;
assign w7948 = ~w7946 & ~w7947;
assign w7949 = pi0463 & ~w7948;
assign w7950 = ~pi0463 & w7948;
assign w7951 = ~w7949 & ~w7950;
assign w7952 = ~w7937 & ~w7951;
assign w7953 = w7924 & ~w7951;
assign w7954 = ~w7952 & ~w7953;
assign w7955 = w7954 & w63593;
assign w7956 = ~w7924 & w7951;
assign w7957 = ~w7937 & w7956;
assign w7958 = w7924 & w7937;
assign w7959 = w7951 & w7958;
assign w7960 = ~w7957 & ~w7959;
assign w7961 = ~w7924 & w7931;
assign w7962 = w7924 & ~w7931;
assign w7963 = w7952 & ~w7962;
assign w7964 = ~w7961 & w7963;
assign w7965 = w7960 & ~w7964;
assign w7966 = w7918 & ~w7961;
assign w7967 = w7937 & w7951;
assign w7968 = w7931 & w7967;
assign w7969 = ~w7963 & ~w7968;
assign w7970 = ~w7966 & ~w7969;
assign w7971 = ~w7918 & ~w7931;
assign w7972 = ~w7967 & w7971;
assign w7973 = ~w7931 & ~w7951;
assign w7974 = ~w7972 & ~w7973;
assign w7975 = w7954 & ~w7974;
assign w7976 = ~w7970 & ~w7975;
assign w7977 = w7931 & w7953;
assign w7978 = ~w7918 & ~w7977;
assign w7979 = ~w7961 & w7978;
assign w7980 = w7976 & w7979;
assign w7981 = (~w7955 & w7965) | (~w7955 & w64789) | (w7965 & w64789);
assign w7982 = (~w7945 & w7980) | (~w7945 & w64790) | (w7980 & w64790);
assign w7983 = w7951 & w7962;
assign w7984 = w7925 & ~w7983;
assign w7985 = w7969 & w7984;
assign w7986 = (w7945 & ~w7976) | (w7945 & w64791) | (~w7976 & w64791);
assign w7987 = w7956 & w63594;
assign w7988 = ~w7939 & ~w7987;
assign w7989 = ~w7986 & w7988;
assign w7990 = ~w7982 & w7989;
assign w7991 = pi0491 & ~w7990;
assign w7992 = ~pi0491 & w7990;
assign w7993 = ~w7991 & ~w7992;
assign w7994 = ~pi3464 & pi9040;
assign w7995 = ~pi3372 & ~pi9040;
assign w7996 = ~w7994 & ~w7995;
assign w7997 = pi0459 & ~w7996;
assign w7998 = ~pi0459 & w7996;
assign w7999 = ~w7997 & ~w7998;
assign w8000 = ~pi3415 & pi9040;
assign w8001 = ~pi3418 & ~pi9040;
assign w8002 = ~w8000 & ~w8001;
assign w8003 = pi0468 & ~w8002;
assign w8004 = ~pi0468 & w8002;
assign w8005 = ~w8003 & ~w8004;
assign w8006 = ~pi3399 & pi9040;
assign w8007 = ~pi3480 & ~pi9040;
assign w8008 = ~w8006 & ~w8007;
assign w8009 = pi0471 & ~w8008;
assign w8010 = ~pi0471 & w8008;
assign w8011 = ~w8009 & ~w8010;
assign w8012 = w8005 & ~w8011;
assign w8013 = ~pi3375 & pi9040;
assign w8014 = ~pi3383 & ~pi9040;
assign w8015 = ~w8013 & ~w8014;
assign w8016 = pi0442 & ~w8015;
assign w8017 = ~pi0442 & w8015;
assign w8018 = ~w8016 & ~w8017;
assign w8019 = ~pi3373 & pi9040;
assign w8020 = ~pi3396 & ~pi9040;
assign w8021 = ~w8019 & ~w8020;
assign w8022 = pi0476 & ~w8021;
assign w8023 = ~pi0476 & w8021;
assign w8024 = ~w8022 & ~w8023;
assign w8025 = ~w8018 & w8024;
assign w8026 = w8018 & ~w8024;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = w8012 & w8027;
assign w8029 = w8018 & w8024;
assign w8030 = w8005 & w8011;
assign w8031 = w8029 & w8030;
assign w8032 = ~w8028 & ~w8031;
assign w8033 = ~w8005 & ~w8018;
assign w8034 = ~w8005 & w8011;
assign w8035 = ~w8027 & w8034;
assign w8036 = (~w8033 & w8027) | (~w8033 & w64792) | (w8027 & w64792);
assign w8037 = (w7999 & ~w8032) | (w7999 & w64793) | (~w8032 & w64793);
assign w8038 = ~w8005 & ~w8011;
assign w8039 = w8018 & w8038;
assign w8040 = w8005 & w8025;
assign w8041 = ~w8039 & ~w8040;
assign w8042 = ~w7999 & ~w8041;
assign w8043 = w8018 & ~w8034;
assign w8044 = ~w8011 & ~w8024;
assign w8045 = w8011 & w8024;
assign w8046 = ~w8044 & ~w8045;
assign w8047 = w8043 & w8046;
assign w8048 = ~w8042 & ~w8047;
assign w8049 = ~w8037 & w8048;
assign w8050 = ~pi3395 & pi9040;
assign w8051 = ~pi3375 & ~pi9040;
assign w8052 = ~w8050 & ~w8051;
assign w8053 = pi0463 & ~w8052;
assign w8054 = ~pi0463 & w8052;
assign w8055 = ~w8053 & ~w8054;
assign w8056 = ~w8049 & w8055;
assign w8057 = w8025 & w8038;
assign w8058 = ~w8018 & ~w8024;
assign w8059 = w8034 & w8058;
assign w8060 = w8026 & w8030;
assign w8061 = ~w8059 & ~w8060;
assign w8062 = ~w8057 & w8061;
assign w8063 = w7999 & ~w8062;
assign w8064 = w8012 & w8029;
assign w8065 = w8029 & w8034;
assign w8066 = ~w8025 & ~w8033;
assign w8067 = ~w7999 & ~w8043;
assign w8068 = w8066 & w8067;
assign w8069 = w7999 & ~w8058;
assign w8070 = w8044 & w8069;
assign w8071 = ~w7999 & ~w8018;
assign w8072 = w8038 & w8071;
assign w8073 = ~w8065 & ~w8072;
assign w8074 = ~w8070 & w8073;
assign w8075 = ~w8068 & w8074;
assign w8076 = ~w8055 & ~w8075;
assign w8077 = w8030 & w8071;
assign w8078 = ~w8064 & ~w8077;
assign w8079 = ~w8063 & w8078;
assign w8080 = ~w8076 & w8079;
assign w8081 = ~w8056 & w8080;
assign w8082 = pi0498 & w8081;
assign w8083 = ~pi0498 & ~w8081;
assign w8084 = ~w8082 & ~w8083;
assign w8085 = ~pi3410 & pi9040;
assign w8086 = ~pi3388 & ~pi9040;
assign w8087 = ~w8085 & ~w8086;
assign w8088 = pi0472 & ~w8087;
assign w8089 = ~pi0472 & w8087;
assign w8090 = ~w8088 & ~w8089;
assign w8091 = ~pi3376 & pi9040;
assign w8092 = ~pi3381 & ~pi9040;
assign w8093 = ~w8091 & ~w8092;
assign w8094 = pi0442 & ~w8093;
assign w8095 = ~pi0442 & w8093;
assign w8096 = ~w8094 & ~w8095;
assign w8097 = ~w8090 & w8096;
assign w8098 = ~pi3370 & pi9040;
assign w8099 = ~pi3397 & ~pi9040;
assign w8100 = ~w8098 & ~w8099;
assign w8101 = pi0465 & ~w8100;
assign w8102 = ~pi0465 & w8100;
assign w8103 = ~w8101 & ~w8102;
assign w8104 = ~w8097 & ~w8103;
assign w8105 = ~pi3381 & pi9040;
assign w8106 = ~pi3455 & ~pi9040;
assign w8107 = ~w8105 & ~w8106;
assign w8108 = pi0467 & ~w8107;
assign w8109 = ~pi0467 & w8107;
assign w8110 = ~w8108 & ~w8109;
assign w8111 = ~w8103 & w8110;
assign w8112 = ~pi3452 & pi9040;
assign w8113 = ~pi3377 & ~pi9040;
assign w8114 = ~w8112 & ~w8113;
assign w8115 = pi0475 & ~w8114;
assign w8116 = ~pi0475 & w8114;
assign w8117 = ~w8115 & ~w8116;
assign w8118 = ~w8111 & ~w8117;
assign w8119 = w8090 & ~w8096;
assign w8120 = w8118 & w8119;
assign w8121 = w8090 & w8096;
assign w8122 = w8103 & ~w8121;
assign w8123 = w8090 & ~w8110;
assign w8124 = ~w8119 & ~w8123;
assign w8125 = ~w8122 & ~w8124;
assign w8126 = ~w8117 & ~w8125;
assign w8127 = ~w8125 & w64794;
assign w8128 = ~w8120 & ~w8127;
assign w8129 = w8104 & ~w8128;
assign w8130 = ~w8117 & ~w8121;
assign w8131 = w8103 & ~w8110;
assign w8132 = ~w8096 & ~w8110;
assign w8133 = ~w8131 & ~w8132;
assign w8134 = w8130 & ~w8133;
assign w8135 = ~pi3367 & pi9040;
assign w8136 = ~pi3454 & ~pi9040;
assign w8137 = ~w8135 & ~w8136;
assign w8138 = pi0468 & ~w8137;
assign w8139 = ~pi0468 & w8137;
assign w8140 = ~w8138 & ~w8139;
assign w8141 = ~w8090 & ~w8096;
assign w8142 = ~w8090 & w8110;
assign w8143 = ~w8123 & ~w8142;
assign w8144 = ~w8103 & ~w8143;
assign w8145 = ~w8141 & w8144;
assign w8146 = w8110 & w8117;
assign w8147 = ~w8097 & w8103;
assign w8148 = w8146 & w8147;
assign w8149 = w8119 & w8146;
assign w8150 = ~w8140 & ~w8149;
assign w8151 = ~w8134 & w8150;
assign w8152 = ~w8148 & w8151;
assign w8153 = ~w8145 & w8152;
assign w8154 = w8117 & ~w8133;
assign w8155 = (~w8111 & w8133) | (~w8111 & w8118) | (w8133 & w8118);
assign w8156 = w8141 & w8155;
assign w8157 = ~w8121 & w64795;
assign w8158 = w8096 & w8117;
assign w8159 = (w8158 & w8144) | (w8158 & w63595) | (w8144 & w63595);
assign w8160 = ~w8141 & ~w8157;
assign w8161 = ~w8159 & w8160;
assign w8162 = ~w8156 & ~w8161;
assign w8163 = ~w8104 & ~w8122;
assign w8164 = w8118 & w8163;
assign w8165 = w8140 & ~w8164;
assign w8166 = ~w8162 & w8165;
assign w8167 = (~w8129 & w8166) | (~w8129 & w64796) | (w8166 & w64796);
assign w8168 = pi0489 & w8167;
assign w8169 = ~pi0489 & ~w8167;
assign w8170 = ~w8168 & ~w8169;
assign w8171 = w8005 & ~w8024;
assign w8172 = w7999 & ~w8171;
assign w8173 = ~w8005 & ~w8024;
assign w8174 = ~w8045 & ~w8173;
assign w8175 = ~w8039 & w8174;
assign w8176 = ~w8034 & ~w8175;
assign w8177 = ~w8175 & w63596;
assign w8178 = (~w8040 & w8175) | (~w8040 & w64797) | (w8175 & w64797);
assign w8179 = w8172 & ~w8178;
assign w8180 = ~w7999 & w8012;
assign w8181 = ~w8035 & ~w8180;
assign w8182 = ~w8179 & w8181;
assign w8183 = w8055 & ~w8182;
assign w8184 = w8069 & ~w8173;
assign w8185 = w8024 & ~w8038;
assign w8186 = w8184 & ~w8185;
assign w8187 = (~w8077 & ~w8184) | (~w8077 & w64798) | (~w8184 & w64798);
assign w8188 = w8027 & ~w8187;
assign w8189 = ~w8035 & ~w8060;
assign w8190 = w7999 & ~w8059;
assign w8191 = ~w8176 & w8190;
assign w8192 = ~w8189 & w8191;
assign w8193 = (w7999 & w8028) | (w7999 & w64799) | (w8028 & w64799);
assign w8194 = w8025 & ~w8034;
assign w8195 = ~w7999 & w8194;
assign w8196 = ~w7999 & ~w8005;
assign w8197 = w8029 & w8196;
assign w8198 = ~w8039 & ~w8197;
assign w8199 = w8061 & w8198;
assign w8200 = ~w8195 & w8199;
assign w8201 = (~w8055 & ~w8200) | (~w8055 & w64800) | (~w8200 & w64800);
assign w8202 = ~w8188 & ~w8192;
assign w8203 = ~w8201 & w8202;
assign w8204 = (~pi0490 & ~w8203) | (~pi0490 & w64801) | (~w8203 & w64801);
assign w8205 = w8203 & w64802;
assign w8206 = ~w8204 & ~w8205;
assign w8207 = ~pi3361 & pi9040;
assign w8208 = pi3407 & ~pi9040;
assign w8209 = ~w8207 & ~w8208;
assign w8210 = pi0443 & ~w8209;
assign w8211 = ~pi0443 & w8209;
assign w8212 = ~w8210 & ~w8211;
assign w8213 = ~pi3379 & pi9040;
assign w8214 = ~pi3363 & ~pi9040;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = pi0457 & ~w8215;
assign w8217 = ~pi0457 & w8215;
assign w8218 = ~w8216 & ~w8217;
assign w8219 = ~pi3407 & pi9040;
assign w8220 = ~pi3406 & ~pi9040;
assign w8221 = ~w8219 & ~w8220;
assign w8222 = pi0456 & ~w8221;
assign w8223 = ~pi0456 & w8221;
assign w8224 = ~w8222 & ~w8223;
assign w8225 = ~w8218 & ~w8224;
assign w8226 = ~pi3413 & pi9040;
assign w8227 = ~pi3371 & ~pi9040;
assign w8228 = ~w8226 & ~w8227;
assign w8229 = pi0450 & ~w8228;
assign w8230 = ~pi0450 & w8228;
assign w8231 = ~w8229 & ~w8230;
assign w8232 = ~pi3406 & pi9040;
assign w8233 = ~pi3379 & ~pi9040;
assign w8234 = ~w8232 & ~w8233;
assign w8235 = pi0461 & ~w8234;
assign w8236 = ~pi0461 & w8234;
assign w8237 = ~w8235 & ~w8236;
assign w8238 = ~w8231 & ~w8237;
assign w8239 = w8225 & w8238;
assign w8240 = ~pi3392 & pi9040;
assign w8241 = ~pi3419 & ~pi9040;
assign w8242 = ~w8240 & ~w8241;
assign w8243 = pi0477 & ~w8242;
assign w8244 = ~pi0477 & w8242;
assign w8245 = ~w8243 & ~w8244;
assign w8246 = w8231 & w8237;
assign w8247 = w8225 & w8246;
assign w8248 = w8231 & ~w8237;
assign w8249 = w8218 & w8248;
assign w8250 = ~w8247 & ~w8249;
assign w8251 = ~w8245 & ~w8250;
assign w8252 = w8237 & w8245;
assign w8253 = ~w8218 & w8224;
assign w8254 = ~w8224 & w8237;
assign w8255 = w8218 & w8231;
assign w8256 = w8254 & w8255;
assign w8257 = ~w8253 & ~w8256;
assign w8258 = w8252 & ~w8257;
assign w8259 = w8248 & w8253;
assign w8260 = ~w8239 & ~w8259;
assign w8261 = ~w8251 & w8260;
assign w8262 = (~w8212 & ~w8261) | (~w8212 & w64803) | (~w8261 & w64803);
assign w8263 = ~w8218 & ~w8231;
assign w8264 = ~w8224 & ~w8263;
assign w8265 = ~w8231 & w8237;
assign w8266 = w8224 & w8237;
assign w8267 = ~w8265 & ~w8266;
assign w8268 = ~w8263 & ~w8267;
assign w8269 = w8224 & ~w8237;
assign w8270 = w8263 & w8269;
assign w8271 = ~w8268 & ~w8270;
assign w8272 = w8245 & ~w8255;
assign w8273 = ~w8264 & w8272;
assign w8274 = w8271 & w8273;
assign w8275 = w8218 & w8269;
assign w8276 = ~w8245 & ~w8275;
assign w8277 = w8218 & ~w8254;
assign w8278 = w8276 & w8277;
assign w8279 = ~w8218 & w8245;
assign w8280 = w8248 & ~w8279;
assign w8281 = ~w8224 & w8280;
assign w8282 = w8218 & w8224;
assign w8283 = ~w8279 & ~w8282;
assign w8284 = w8246 & ~w8283;
assign w8285 = ~w8253 & w8284;
assign w8286 = ~w8245 & ~w8271;
assign w8287 = w8254 & w8263;
assign w8288 = ~w8281 & ~w8287;
assign w8289 = ~w8285 & w8288;
assign w8290 = ~w8286 & w8289;
assign w8291 = w8212 & ~w8290;
assign w8292 = ~w8274 & ~w8278;
assign w8293 = ~w8262 & w8292;
assign w8294 = ~w8291 & w8293;
assign w8295 = pi0485 & ~w8294;
assign w8296 = ~pi0485 & w8294;
assign w8297 = ~w8295 & ~w8296;
assign w8298 = w7978 & ~w7983;
assign w8299 = (w7918 & ~w7954) | (w7918 & w63597) | (~w7954 & w63597);
assign w8300 = ~w7973 & w8299;
assign w8301 = ~w8298 & ~w8300;
assign w8302 = w7967 & w7971;
assign w8303 = ~w7924 & w8302;
assign w8304 = ~w7931 & ~w7958;
assign w8305 = ~w7967 & ~w7977;
assign w8306 = ~w8304 & w8305;
assign w8307 = (~w7918 & ~w8302) | (~w7918 & w63598) | (~w8302 & w63598);
assign w8308 = ~w8306 & w8307;
assign w8309 = (w7918 & ~w7958) | (w7918 & w64804) | (~w7958 & w64804);
assign w8310 = ~w7977 & ~w7987;
assign w8311 = w8309 & w8310;
assign w8312 = w7924 & w7931;
assign w8313 = ~w7938 & w7951;
assign w8314 = ~w8312 & w8313;
assign w8315 = (w8314 & w8308) | (w8314 & w63599) | (w8308 & w63599);
assign w8316 = (~w7945 & w8315) | (~w7945 & w64805) | (w8315 & w64805);
assign w8317 = w7952 & w7962;
assign w8318 = ~w7968 & ~w8317;
assign w8319 = w7918 & ~w8318;
assign w8320 = ~w8308 & w64806;
assign w8321 = w7952 & w7971;
assign w8322 = ~w7924 & w8321;
assign w8323 = w7975 & ~w8298;
assign w8324 = ~w8319 & ~w8322;
assign w8325 = ~w8323 & w8324;
assign w8326 = ~w8320 & w8325;
assign w8327 = ~w8316 & w8326;
assign w8328 = pi0496 & ~w8327;
assign w8329 = ~pi0496 & w8327;
assign w8330 = ~w8328 & ~w8329;
assign w8331 = ~pi3384 & pi9040;
assign w8332 = ~pi3394 & ~pi9040;
assign w8333 = ~w8331 & ~w8332;
assign w8334 = pi0478 & ~w8333;
assign w8335 = ~pi0478 & w8333;
assign w8336 = ~w8334 & ~w8335;
assign w8337 = ~pi3416 & pi9040;
assign w8338 = ~pi3389 & ~pi9040;
assign w8339 = ~w8337 & ~w8338;
assign w8340 = pi0448 & ~w8339;
assign w8341 = ~pi0448 & w8339;
assign w8342 = ~w8340 & ~w8341;
assign w8343 = ~pi3365 & pi9040;
assign w8344 = ~pi3452 & ~pi9040;
assign w8345 = ~w8343 & ~w8344;
assign w8346 = pi0474 & ~w8345;
assign w8347 = ~pi0474 & w8345;
assign w8348 = ~w8346 & ~w8347;
assign w8349 = ~w8342 & w8348;
assign w8350 = ~pi3456 & pi9040;
assign w8351 = ~pi3365 & ~pi9040;
assign w8352 = ~w8350 & ~w8351;
assign w8353 = pi0455 & ~w8352;
assign w8354 = ~pi0455 & w8352;
assign w8355 = ~w8353 & ~w8354;
assign w8356 = w8349 & ~w8355;
assign w8357 = ~w8342 & w8355;
assign w8358 = ~pi3369 & pi9040;
assign w8359 = ~pi3408 & ~pi9040;
assign w8360 = ~w8358 & ~w8359;
assign w8361 = pi0466 & ~w8360;
assign w8362 = ~pi0466 & w8360;
assign w8363 = ~w8361 & ~w8362;
assign w8364 = ~w8357 & ~w8363;
assign w8365 = w8357 & w8363;
assign w8366 = ~w8364 & ~w8365;
assign w8367 = ~pi3388 & pi9040;
assign w8368 = ~pi3390 & ~pi9040;
assign w8369 = ~w8367 & ~w8368;
assign w8370 = pi0460 & ~w8369;
assign w8371 = ~pi0460 & w8369;
assign w8372 = ~w8370 & ~w8371;
assign w8373 = ~w8356 & ~w8372;
assign w8374 = w8366 & w8373;
assign w8375 = w8348 & w8363;
assign w8376 = w8342 & ~w8355;
assign w8377 = w8375 & w8376;
assign w8378 = w8349 & ~w8363;
assign w8379 = ~w8377 & ~w8378;
assign w8380 = ~w8374 & w8379;
assign w8381 = ~w8336 & ~w8380;
assign w8382 = w8355 & w8378;
assign w8383 = (~w8336 & ~w8357) | (~w8336 & w64807) | (~w8357 & w64807);
assign w8384 = ~w8348 & w8363;
assign w8385 = ~w8383 & w8384;
assign w8386 = w8355 & w8363;
assign w8387 = w8336 & w8342;
assign w8388 = w8386 & w8387;
assign w8389 = w8348 & ~w8363;
assign w8390 = w8387 & ~w8389;
assign w8391 = w8348 & ~w8355;
assign w8392 = w8364 & ~w8391;
assign w8393 = ~w8336 & ~w8392;
assign w8394 = ~w8355 & w8363;
assign w8395 = w8336 & ~w8394;
assign w8396 = ~w8376 & w8395;
assign w8397 = ~w8390 & ~w8396;
assign w8398 = ~w8393 & w8397;
assign w8399 = w8372 & ~w8388;
assign w8400 = ~w8382 & w8399;
assign w8401 = ~w8385 & w8400;
assign w8402 = ~w8398 & w8401;
assign w8403 = ~w8355 & w8378;
assign w8404 = ~w8357 & ~w8376;
assign w8405 = w8375 & ~w8404;
assign w8406 = w8336 & w8392;
assign w8407 = ~w8372 & ~w8403;
assign w8408 = ~w8405 & w8407;
assign w8409 = ~w8406 & w8408;
assign w8410 = ~w8402 & ~w8409;
assign w8411 = ~w8381 & ~w8410;
assign w8412 = pi0482 & w8411;
assign w8413 = ~pi0482 & ~w8411;
assign w8414 = ~w8412 & ~w8413;
assign w8415 = ~w8143 & w64808;
assign w8416 = w8097 & w8415;
assign w8417 = w8117 & ~w8144;
assign w8418 = w8096 & ~w8110;
assign w8419 = ~w8417 & w8418;
assign w8420 = ~w8097 & w8117;
assign w8421 = w8124 & ~w8142;
assign w8422 = w8420 & w8421;
assign w8423 = w8103 & w8117;
assign w8424 = w8142 & w8423;
assign w8425 = ~w8096 & w8103;
assign w8426 = ~w8117 & w8425;
assign w8427 = w8425 & w64809;
assign w8428 = ~w8111 & ~w8131;
assign w8429 = (~w8140 & ~w8428) | (~w8140 & w64810) | (~w8428 & w64810);
assign w8430 = ~w8424 & ~w8427;
assign w8431 = ~w8422 & w64811;
assign w8432 = ~w8419 & w8431;
assign w8433 = w8110 & w8163;
assign w8434 = ~w8110 & w8117;
assign w8435 = ~w8141 & w8434;
assign w8436 = ~w8426 & ~w8435;
assign w8437 = w8421 & ~w8436;
assign w8438 = w8140 & ~w8149;
assign w8439 = ~w8415 & w8438;
assign w8440 = ~w8433 & ~w8437;
assign w8441 = w8439 & w8440;
assign w8442 = ~w8432 & ~w8441;
assign w8443 = ~w8103 & w8141;
assign w8444 = w8119 & w8131;
assign w8445 = ~w8443 & ~w8444;
assign w8446 = w8154 & ~w8445;
assign w8447 = ~w8103 & w8149;
assign w8448 = ~w8446 & ~w8447;
assign w8449 = ~w8416 & w8448;
assign w8450 = ~w8442 & w8449;
assign w8451 = pi0487 & ~w8450;
assign w8452 = ~pi0487 & w8450;
assign w8453 = ~w8451 & ~w8452;
assign w8454 = w8342 & ~w8348;
assign w8455 = w8363 & w8454;
assign w8456 = ~w8403 & ~w8455;
assign w8457 = w8336 & ~w8456;
assign w8458 = ~w8386 & ~w8404;
assign w8459 = ~w8404 & w64812;
assign w8460 = ~w8336 & w8357;
assign w8461 = w8355 & ~w8363;
assign w8462 = w8342 & w8461;
assign w8463 = ~w8460 & ~w8462;
assign w8464 = ~w8349 & ~w8454;
assign w8465 = ~w8463 & w8464;
assign w8466 = ~w8336 & ~w8384;
assign w8467 = w8366 & w8466;
assign w8468 = ~w8372 & ~w8467;
assign w8469 = w8396 & w8405;
assign w8470 = ~w8459 & ~w8465;
assign w8471 = ~w8469 & w8470;
assign w8472 = w8468 & w8471;
assign w8473 = w8454 & w8386;
assign w8474 = ~w8366 & ~w8384;
assign w8475 = w8393 & w8474;
assign w8476 = ~w8342 & ~w8355;
assign w8477 = ~w8375 & w8476;
assign w8478 = ~w8395 & w8477;
assign w8479 = ~w8363 & ~w8387;
assign w8480 = w8464 & w8479;
assign w8481 = ~w8463 & w8480;
assign w8482 = w8372 & ~w8390;
assign w8483 = ~w8473 & w8482;
assign w8484 = ~w8478 & w8483;
assign w8485 = ~w8481 & w8484;
assign w8486 = ~w8475 & w8485;
assign w8487 = ~w8472 & ~w8486;
assign w8488 = ~w8487 & w64813;
assign w8489 = (pi0492 & w8487) | (pi0492 & w64814) | (w8487 & w64814);
assign w8490 = ~w8488 & ~w8489;
assign w8491 = w8133 & ~w8143;
assign w8492 = w8420 & w8491;
assign w8493 = w8096 & w8103;
assign w8494 = w8143 & w8493;
assign w8495 = ~w8120 & ~w8494;
assign w8496 = ~w8492 & w8495;
assign w8497 = w8496 & w64815;
assign w8498 = (~w8103 & w8121) | (~w8103 & w64816) | (w8121 & w64816);
assign w8499 = ~w8420 & w8498;
assign w8500 = w8090 & ~w8155;
assign w8501 = w8429 & ~w8499;
assign w8502 = ~w8156 & w8501;
assign w8503 = ~w8500 & w8502;
assign w8504 = ~w8497 & ~w8503;
assign w8505 = ~w8443 & ~w8494;
assign w8506 = w8118 & ~w8505;
assign w8507 = ~w8424 & ~w8447;
assign w8508 = ~w8506 & w8507;
assign w8509 = ~w8504 & w8508;
assign w8510 = ~pi0504 & w8509;
assign w8511 = pi0504 & ~w8509;
assign w8512 = ~w8510 & ~w8511;
assign w8513 = ~w8176 & w8184;
assign w8514 = w8012 & ~w8027;
assign w8515 = (~w8012 & w8194) | (~w8012 & w64817) | (w8194 & w64817);
assign w8516 = ~w7999 & ~w8515;
assign w8517 = w8176 & w8516;
assign w8518 = w8030 & w8058;
assign w8519 = ~w8514 & ~w8518;
assign w8520 = ~w8513 & w8519;
assign w8521 = (w8055 & ~w8520) | (w8055 & w64818) | (~w8520 & w64818);
assign w8522 = ~w7999 & ~w8035;
assign w8523 = w8012 & w8026;
assign w8524 = w8190 & ~w8523;
assign w8525 = ~w8522 & ~w8524;
assign w8526 = ~w8028 & ~w8035;
assign w8527 = w8516 & w8526;
assign w8528 = (~w8055 & w8176) | (~w8055 & w64819) | (w8176 & w64819);
assign w8529 = ~w8527 & w8528;
assign w8530 = ~w8525 & ~w8529;
assign w8531 = ~w8521 & w8530;
assign w8532 = pi0511 & ~w8531;
assign w8533 = ~pi0511 & w8531;
assign w8534 = ~w8532 & ~w8533;
assign w8535 = ~w8265 & ~w8280;
assign w8536 = w8253 & ~w8535;
assign w8537 = ~w8224 & ~w8250;
assign w8538 = w8239 & w8245;
assign w8539 = ~w8231 & w8269;
assign w8540 = ~w8252 & ~w8539;
assign w8541 = w8218 & ~w8540;
assign w8542 = ~w8212 & ~w8538;
assign w8543 = ~w8536 & w8542;
assign w8544 = ~w8537 & ~w8541;
assign w8545 = w8543 & w8544;
assign w8546 = ~w8255 & ~w8263;
assign w8547 = ~w8266 & w8546;
assign w8548 = ~w8245 & ~w8547;
assign w8549 = w8246 & w8253;
assign w8550 = w8248 & ~w8283;
assign w8551 = ~w8225 & w8238;
assign w8552 = ~w8282 & w8551;
assign w8553 = w8212 & ~w8287;
assign w8554 = ~w8549 & w8553;
assign w8555 = ~w8550 & ~w8552;
assign w8556 = w8554 & w8555;
assign w8557 = ~w8548 & w8556;
assign w8558 = ~w8545 & ~w8557;
assign w8559 = ~pi0481 & w8558;
assign w8560 = pi0481 & ~w8558;
assign w8561 = ~w8559 & ~w8560;
assign w8562 = w7924 & w7952;
assign w8563 = ~w7954 & ~w8562;
assign w8564 = w7937 & w8312;
assign w8565 = (~w8309 & w8563) | (~w8309 & w64820) | (w8563 & w64820);
assign w8566 = ~w7983 & w8299;
assign w8567 = ~w8563 & w8566;
assign w8568 = (~w7945 & w8567) | (~w7945 & w64821) | (w8567 & w64821);
assign w8569 = w7931 & w8563;
assign w8570 = ~w7918 & ~w7956;
assign w8571 = ~w8566 & ~w8570;
assign w8572 = w7937 & w7973;
assign w8573 = ~w7962 & ~w8572;
assign w8574 = ~w7958 & ~w8573;
assign w8575 = ~w8569 & ~w8574;
assign w8576 = ~w8571 & w8575;
assign w8577 = w7945 & ~w8576;
assign w8578 = ~w8303 & ~w8323;
assign w8579 = ~w8568 & w8578;
assign w8580 = ~w8577 & w8579;
assign w8581 = pi0503 & ~w8580;
assign w8582 = ~pi0503 & w8580;
assign w8583 = ~w8581 & ~w8582;
assign w8584 = ~w7844 & w7878;
assign w8585 = w7836 & w7844;
assign w8586 = w7850 & w8585;
assign w8587 = ~w8584 & ~w8586;
assign w8588 = ~w7885 & ~w8587;
assign w8589 = ~w7835 & w7870;
assign w8590 = w7862 & ~w8589;
assign w8591 = ~w7854 & ~w8590;
assign w8592 = w7861 & w8591;
assign w8593 = w7853 & ~w7888;
assign w8594 = w7878 & ~w8593;
assign w8595 = w8587 & w8594;
assign w8596 = (w7870 & ~w7860) | (w7870 & w64822) | (~w7860 & w64822);
assign w8597 = ~w7906 & w8596;
assign w8598 = ~w8592 & w8597;
assign w8599 = ~w8595 & w8598;
assign w8600 = w7850 & ~w8584;
assign w8601 = ~w7838 & w8600;
assign w8602 = ~w7844 & w7888;
assign w8603 = ~w7882 & ~w8602;
assign w8604 = w7878 & ~w8603;
assign w8605 = w7853 & w7880;
assign w8606 = ~w7870 & ~w8605;
assign w8607 = w7858 & ~w7863;
assign w8608 = ~w8601 & w8606;
assign w8609 = w8607 & w8608;
assign w8610 = ~w8604 & w8609;
assign w8611 = ~w8599 & ~w8610;
assign w8612 = ~w8588 & ~w8611;
assign w8613 = ~pi0493 & w8612;
assign w8614 = pi0493 & ~w8612;
assign w8615 = ~w8613 & ~w8614;
assign w8616 = ~pi3397 & pi9040;
assign w8617 = ~pi3366 & ~pi9040;
assign w8618 = ~w8616 & ~w8617;
assign w8619 = pi0446 & ~w8618;
assign w8620 = ~pi0446 & w8618;
assign w8621 = ~w8619 & ~w8620;
assign w8622 = ~pi3362 & pi9040;
assign w8623 = ~pi3416 & ~pi9040;
assign w8624 = ~w8622 & ~w8623;
assign w8625 = pi0460 & ~w8624;
assign w8626 = ~pi0460 & w8624;
assign w8627 = ~w8625 & ~w8626;
assign w8628 = w8621 & ~w8627;
assign w8629 = ~pi3382 & pi9040;
assign w8630 = ~pi3457 & ~pi9040;
assign w8631 = ~w8629 & ~w8630;
assign w8632 = pi0455 & ~w8631;
assign w8633 = ~pi0455 & w8631;
assign w8634 = ~w8632 & ~w8633;
assign w8635 = ~pi3455 & pi9040;
assign w8636 = ~pi3391 & ~pi9040;
assign w8637 = ~w8635 & ~w8636;
assign w8638 = pi0464 & ~w8637;
assign w8639 = ~pi0464 & w8637;
assign w8640 = ~w8638 & ~w8639;
assign w8641 = ~w8627 & ~w8640;
assign w8642 = ~pi3408 & pi9040;
assign w8643 = ~pi3367 & ~pi9040;
assign w8644 = ~w8642 & ~w8643;
assign w8645 = pi0467 & ~w8644;
assign w8646 = ~pi0467 & w8644;
assign w8647 = ~w8645 & ~w8646;
assign w8648 = w8641 & w8647;
assign w8649 = w8627 & w8640;
assign w8650 = ~w8634 & w8649;
assign w8651 = ~w8648 & ~w8650;
assign w8652 = ~w8641 & ~w8647;
assign w8653 = (~w8634 & w8641) | (~w8634 & w8675) | (w8641 & w8675);
assign w8654 = w8651 & w8653;
assign w8655 = w8651 & w63365;
assign w8656 = ~pi3390 & pi9040;
assign w8657 = ~pi3369 & ~pi9040;
assign w8658 = ~w8656 & ~w8657;
assign w8659 = pi0472 & ~w8658;
assign w8660 = ~pi0472 & w8658;
assign w8661 = ~w8659 & ~w8660;
assign w8662 = w8634 & w8640;
assign w8663 = ~w8634 & ~w8640;
assign w8664 = ~w8662 & ~w8663;
assign w8665 = w8627 & w8647;
assign w8666 = ~w8627 & ~w8647;
assign w8667 = ~w8665 & ~w8666;
assign w8668 = ~w8628 & w8667;
assign w8669 = ~w8634 & w8667;
assign w8670 = ~w8668 & ~w8669;
assign w8671 = w8664 & ~w8670;
assign w8672 = ~w8664 & ~w8668;
assign w8673 = ~w8661 & ~w8672;
assign w8674 = ~w8671 & w8673;
assign w8675 = ~w8634 & w8647;
assign w8676 = w8634 & ~w8647;
assign w8677 = ~w8649 & ~w8676;
assign w8678 = w8662 & ~w8665;
assign w8679 = w8621 & ~w8678;
assign w8680 = ~w8677 & w8679;
assign w8681 = w8679 & w64823;
assign w8682 = ~w8627 & ~w8634;
assign w8683 = ~w8676 & ~w8682;
assign w8684 = ~w8675 & w8683;
assign w8685 = w8621 & ~w8666;
assign w8686 = (w8685 & ~w8684) | (w8685 & w64824) | (~w8684 & w64824);
assign w8687 = w8684 & w64825;
assign w8688 = w8640 & w8666;
assign w8689 = w8634 & w8688;
assign w8690 = ~w8686 & ~w8689;
assign w8691 = ~w8687 & w8690;
assign w8692 = w8661 & ~w8691;
assign w8693 = ~w8655 & ~w8681;
assign w8694 = ~w8674 & w8693;
assign w8695 = ~w8692 & w8694;
assign w8696 = ~pi0500 & w8695;
assign w8697 = pi0500 & ~w8695;
assign w8698 = ~w8696 & ~w8697;
assign w8699 = (w8651 & w8655) | (w8651 & w63600) | (w8655 & w63600);
assign w8700 = w8634 & ~w8640;
assign w8701 = w8667 & w63601;
assign w8702 = ~w8621 & ~w8663;
assign w8703 = ~w8667 & w8702;
assign w8704 = ~w8701 & ~w8703;
assign w8705 = (w8704 & ~w8699) | (w8704 & w64826) | (~w8699 & w64826);
assign w8706 = w8661 & ~w8705;
assign w8707 = w8662 & w8687;
assign w8708 = ~w8666 & ~w8682;
assign w8709 = ~w8648 & ~w8688;
assign w8710 = ~w8701 & w8709;
assign w8711 = w8621 & w8708;
assign w8712 = ~w8710 & w8711;
assign w8713 = ~w8621 & ~w8650;
assign w8714 = ~w8710 & w8713;
assign w8715 = ~w8661 & ~w8703;
assign w8716 = ~w8714 & w8715;
assign w8717 = ~w8699 & w8716;
assign w8718 = ~w8707 & ~w8712;
assign w8719 = ~w8717 & w8718;
assign w8720 = (pi0501 & ~w8719) | (pi0501 & w64827) | (~w8719 & w64827);
assign w8721 = w8719 & w64828;
assign w8722 = ~w8720 & ~w8721;
assign w8723 = w8661 & ~w8681;
assign w8724 = ~w8621 & ~w8649;
assign w8725 = w8683 & w8724;
assign w8726 = ~w8654 & ~w8725;
assign w8727 = ~w8680 & w8726;
assign w8728 = w8634 & w8666;
assign w8729 = ~w8678 & w8724;
assign w8730 = ~w8728 & w8729;
assign w8731 = w8679 & w8710;
assign w8732 = w8661 & ~w8730;
assign w8733 = ~w8731 & w8732;
assign w8734 = ~w8621 & ~w8647;
assign w8735 = w8662 & w8734;
assign w8736 = (~w8735 & w8727) | (~w8735 & w64829) | (w8727 & w64829);
assign w8737 = ~w8733 & w8736;
assign w8738 = pi0508 & w8737;
assign w8739 = ~pi0508 & ~w8737;
assign w8740 = ~w8738 & ~w8739;
assign w8741 = ~pi3389 & pi9040;
assign w8742 = ~pi3456 & ~pi9040;
assign w8743 = ~w8741 & ~w8742;
assign w8744 = pi0448 & ~w8743;
assign w8745 = ~pi0448 & w8743;
assign w8746 = ~w8744 & ~w8745;
assign w8747 = ~pi3391 & pi9040;
assign w8748 = ~pi3378 & ~pi9040;
assign w8749 = ~w8747 & ~w8748;
assign w8750 = pi0473 & ~w8749;
assign w8751 = ~pi0473 & w8749;
assign w8752 = ~w8750 & ~w8751;
assign w8753 = ~w8746 & w8752;
assign w8754 = ~pi3394 & pi9040;
assign w8755 = ~pi3410 & ~pi9040;
assign w8756 = ~w8754 & ~w8755;
assign w8757 = pi0451 & ~w8756;
assign w8758 = ~pi0451 & w8756;
assign w8759 = ~w8757 & ~w8758;
assign w8760 = ~pi3457 & pi9040;
assign w8761 = ~pi3374 & ~pi9040;
assign w8762 = ~w8760 & ~w8761;
assign w8763 = pi0470 & ~w8762;
assign w8764 = ~pi0470 & w8762;
assign w8765 = ~w8763 & ~w8764;
assign w8766 = ~w8759 & ~w8765;
assign w8767 = w8753 & w8766;
assign w8768 = ~pi3420 & pi9040;
assign w8769 = ~pi3382 & ~pi9040;
assign w8770 = ~w8768 & ~w8769;
assign w8771 = pi0479 & ~w8770;
assign w8772 = ~pi0479 & w8770;
assign w8773 = ~w8771 & ~w8772;
assign w8774 = ~w8765 & w8773;
assign w8775 = w8746 & ~w8752;
assign w8776 = ~w8774 & w8775;
assign w8777 = w8752 & w8774;
assign w8778 = ~w8746 & ~w8773;
assign w8779 = w8746 & w8773;
assign w8780 = ~w8778 & ~w8779;
assign w8781 = ~w8765 & ~w8773;
assign w8782 = ~w8753 & ~w8781;
assign w8783 = w8780 & w8782;
assign w8784 = ~w8759 & w8783;
assign w8785 = w8759 & w8765;
assign w8786 = w8778 & w8785;
assign w8787 = ~w8776 & ~w8777;
assign w8788 = ~w8786 & w8787;
assign w8789 = ~w8784 & w8788;
assign w8790 = ~pi3374 & pi9040;
assign w8791 = ~pi3384 & ~pi9040;
assign w8792 = ~w8790 & ~w8791;
assign w8793 = pi0466 & ~w8792;
assign w8794 = ~pi0466 & w8792;
assign w8795 = ~w8793 & ~w8794;
assign w8796 = ~w8789 & w8795;
assign w8797 = ~w8752 & ~w8759;
assign w8798 = w8752 & w8759;
assign w8799 = ~w8797 & ~w8798;
assign w8800 = ~w8780 & w8799;
assign w8801 = ~w8765 & ~w8775;
assign w8802 = ~w8779 & w8801;
assign w8803 = ~w8800 & ~w8802;
assign w8804 = w8773 & w8803;
assign w8805 = ~w8789 & w8804;
assign w8806 = ~w8746 & w8797;
assign w8807 = ~w8777 & ~w8780;
assign w8808 = ~w8775 & w8781;
assign w8809 = (~w8808 & ~w8807) | (~w8808 & w64830) | (~w8807 & w64830);
assign w8810 = ~w8759 & ~w8809;
assign w8811 = ~w8773 & ~w8797;
assign w8812 = ~w8759 & w8773;
assign w8813 = ~w8765 & ~w8812;
assign w8814 = ~w8811 & w8813;
assign w8815 = w8746 & w8798;
assign w8816 = w8753 & w8812;
assign w8817 = ~w8815 & ~w8816;
assign w8818 = ~w8814 & w8817;
assign w8819 = w8783 & ~w8818;
assign w8820 = w8765 & w8773;
assign w8821 = ~w8753 & ~w8775;
assign w8822 = w8780 & ~w8821;
assign w8823 = w8759 & w8822;
assign w8824 = w8822 & w64831;
assign w8825 = ~w8819 & ~w8824;
assign w8826 = (~w8795 & ~w8825) | (~w8795 & w64832) | (~w8825 & w64832);
assign w8827 = w8781 & ~w8821;
assign w8828 = ~w8753 & w8786;
assign w8829 = ~w8827 & ~w8828;
assign w8830 = ~w8773 & w8795;
assign w8831 = ~w8752 & w8759;
assign w8832 = (w8831 & ~w8829) | (w8831 & w64833) | (~w8829 & w64833);
assign w8833 = ~w8767 & ~w8796;
assign w8834 = ~w8805 & ~w8832;
assign w8835 = w8833 & w8834;
assign w8836 = (pi0484 & ~w8835) | (pi0484 & w64834) | (~w8835 & w64834);
assign w8837 = w8835 & w64835;
assign w8838 = ~w8836 & ~w8837;
assign w8839 = w8752 & ~w8773;
assign w8840 = ~w8789 & w8839;
assign w8841 = w8820 & w8821;
assign w8842 = ~w8765 & ~w8798;
assign w8843 = w8807 & w8842;
assign w8844 = ~w8795 & ~w8841;
assign w8845 = ~w8823 & w8844;
assign w8846 = ~w8843 & w8845;
assign w8847 = w8779 & w8797;
assign w8848 = ~w8811 & ~w8847;
assign w8849 = w8765 & ~w8848;
assign w8850 = w8795 & w8818;
assign w8851 = ~w8849 & w8850;
assign w8852 = ~w8846 & ~w8851;
assign w8853 = ~w8840 & ~w8852;
assign w8854 = ~pi0486 & w8853;
assign w8855 = pi0486 & ~w8853;
assign w8856 = ~w8854 & ~w8855;
assign w8857 = (~w8572 & ~w7960) | (~w8572 & w64836) | (~w7960 & w64836);
assign w8858 = ~w7945 & ~w8857;
assign w8859 = ~w7956 & ~w7973;
assign w8860 = (w8859 & ~w7976) | (w8859 & w63602) | (~w7976 & w63602);
assign w8861 = (w7918 & w8860) | (w7918 & w64837) | (w8860 & w64837);
assign w8862 = w7931 & ~w7960;
assign w8863 = (~w7945 & w7955) | (~w7945 & w64838) | (w7955 & w64838);
assign w8864 = ~w8862 & ~w8863;
assign w8865 = ~w7918 & ~w8864;
assign w8866 = ~w7987 & ~w8302;
assign w8867 = ~w7945 & ~w8866;
assign w8868 = w7966 & w7967;
assign w8869 = ~w7956 & w7972;
assign w8870 = ~w8317 & ~w8564;
assign w8871 = ~w8868 & w8870;
assign w8872 = (w7945 & ~w8871) | (w7945 & w64839) | (~w8871 & w64839);
assign w8873 = ~w8321 & ~w8867;
assign w8874 = ~w8872 & w8873;
assign w8875 = ~w8865 & w8874;
assign w8876 = ~w8861 & w8875;
assign w8877 = pi0502 & ~w8876;
assign w8878 = ~pi0502 & w8876;
assign w8879 = ~w8877 & ~w8878;
assign w8880 = (w8423 & ~w8496) | (w8423 & w64840) | (~w8496 & w64840);
assign w8881 = w8122 & w8140;
assign w8882 = ~w8426 & ~w8881;
assign w8883 = w8143 & ~w8882;
assign w8884 = ~w8425 & w8435;
assign w8885 = w8127 & ~w8147;
assign w8886 = w8140 & ~w8884;
assign w8887 = ~w8885 & w8886;
assign w8888 = w8111 & w8119;
assign w8889 = w8117 & w8445;
assign w8890 = ~w8126 & ~w8889;
assign w8891 = ~w8140 & ~w8888;
assign w8892 = ~w8433 & w8891;
assign w8893 = ~w8890 & w8892;
assign w8894 = ~w8887 & ~w8893;
assign w8895 = ~w8880 & ~w8883;
assign w8896 = ~w8894 & w8895;
assign w8897 = pi0505 & ~w8896;
assign w8898 = ~pi0505 & w8896;
assign w8899 = ~w8897 & ~w8898;
assign w8900 = ~w7859 & ~w7892;
assign w8901 = w7861 & w8584;
assign w8902 = w7835 & w7850;
assign w8903 = ~w7855 & ~w7904;
assign w8904 = w8902 & ~w8903;
assign w8905 = ~w7851 & w7878;
assign w8906 = ~w8902 & w8905;
assign w8907 = ~w8593 & w8906;
assign w8908 = w8606 & ~w8904;
assign w8909 = ~w8907 & w8908;
assign w8910 = ~w7829 & w7887;
assign w8911 = w7884 & ~w8910;
assign w8912 = (~w7878 & ~w7884) | (~w7878 & w64841) | (~w7884 & w64841);
assign w8913 = (w7844 & w7856) | (w7844 & w64842) | (w7856 & w64842);
assign w8914 = w7885 & w8913;
assign w8915 = w7864 & w7900;
assign w8916 = ~w8912 & w8915;
assign w8917 = ~w8914 & w8916;
assign w8918 = ~w8909 & ~w8917;
assign w8919 = ~w7907 & ~w8901;
assign w8920 = ~w8900 & w8919;
assign w8921 = ~w8918 & w8920;
assign w8922 = pi0499 & ~w8921;
assign w8923 = ~pi0499 & w8921;
assign w8924 = ~w8922 & ~w8923;
assign w8925 = w8191 & w64843;
assign w8926 = ~w8040 & w8174;
assign w8927 = (~w8523 & w8926) | (~w8523 & w64844) | (w8926 & w64844);
assign w8928 = ~w8177 & w8927;
assign w8929 = ~w7999 & ~w8928;
assign w8930 = w8011 & ~w8066;
assign w8931 = (~w8055 & w8186) | (~w8055 & w64845) | (w8186 & w64845);
assign w8932 = ~w8024 & w8193;
assign w8933 = ~w8012 & ~w8026;
assign w8934 = w8172 & ~w8933;
assign w8935 = ~w8064 & ~w8197;
assign w8936 = ~w8518 & w8935;
assign w8937 = ~w8934 & w8936;
assign w8938 = w8055 & ~w8937;
assign w8939 = ~w8931 & ~w8932;
assign w8940 = ~w8938 & w8939;
assign w8941 = ~w8925 & ~w8929;
assign w8942 = w8940 & w8941;
assign w8943 = pi0522 & ~w8942;
assign w8944 = ~pi0522 & w8942;
assign w8945 = ~w8943 & ~w8944;
assign w8946 = w8683 & w63603;
assign w8947 = w8708 & ~w8946;
assign w8948 = ~w8946 & w8711;
assign w8949 = w8663 & w8666;
assign w8950 = w8652 & w8724;
assign w8951 = w8713 & ~w8950;
assign w8952 = ~w8947 & w8951;
assign w8953 = ~w8948 & ~w8949;
assign w8954 = ~w8952 & w8953;
assign w8955 = ~w8661 & ~w8954;
assign w8956 = ~w8634 & w8688;
assign w8957 = ~w8628 & ~w8679;
assign w8958 = ~w8956 & ~w8957;
assign w8959 = ~w8713 & ~w8958;
assign w8960 = w8628 & w8676;
assign w8961 = ~w8669 & ~w8960;
assign w8962 = (~w8640 & ~w8961) | (~w8640 & w63604) | (~w8961 & w63604);
assign w8963 = w8678 & w8683;
assign w8964 = ~w8950 & ~w8963;
assign w8965 = (w8661 & w8962) | (w8661 & w64846) | (w8962 & w64846);
assign w8966 = ~w8959 & ~w8965;
assign w8967 = ~w8955 & w8966;
assign w8968 = ~pi0495 & w8967;
assign w8969 = pi0495 & ~w8967;
assign w8970 = ~w8968 & ~w8969;
assign w8971 = w8336 & ~w8461;
assign w8972 = ~w8377 & ~w8473;
assign w8973 = ~w8389 & ~w8476;
assign w8974 = ~w8391 & ~w8973;
assign w8975 = ~w8364 & w8974;
assign w8976 = ~w8363 & w8376;
assign w8977 = w8972 & ~w8976;
assign w8978 = ~w8975 & w8977;
assign w8979 = w8336 & ~w8978;
assign w8980 = (~w8372 & ~w8978) | (~w8372 & w64847) | (~w8978 & w64847);
assign w8981 = ~w8979 & w8980;
assign w8982 = ~w8356 & w8383;
assign w8983 = (w8336 & w8973) | (w8336 & w64848) | (w8973 & w64848);
assign w8984 = ~w8982 & ~w8983;
assign w8985 = w8376 & w64849;
assign w8986 = ~w8465 & w63605;
assign w8987 = (w8372 & ~w8986) | (w8372 & w64850) | (~w8986 & w64850);
assign w8988 = ~w8348 & w8461;
assign w8989 = w8468 & w8988;
assign w8990 = ~w8987 & ~w8989;
assign w8991 = ~w8981 & w8990;
assign w8992 = pi0506 & ~w8991;
assign w8993 = ~pi0506 & w8991;
assign w8994 = ~w8992 & ~w8993;
assign w8995 = w7878 & ~w8911;
assign w8996 = w7850 & w7855;
assign w8997 = ~w8913 & ~w8996;
assign w8998 = ~w7838 & w8591;
assign w8999 = ~w7878 & w8997;
assign w9000 = ~w8998 & w8999;
assign w9001 = ~w8995 & ~w9000;
assign w9002 = ~w8906 & ~w9001;
assign w9003 = w7894 & w8902;
assign w9004 = w7855 & w8905;
assign w9005 = ~w7854 & w7870;
assign w9006 = ~w7905 & ~w8585;
assign w9007 = ~w9003 & w9006;
assign w9008 = ~w9004 & w9005;
assign w9009 = w9007 & w9008;
assign w9010 = w7878 & ~w8997;
assign w9011 = w7856 & w7862;
assign w9012 = ~w7870 & ~w9011;
assign w9013 = ~w9010 & w9012;
assign w9014 = ~w9009 & ~w9013;
assign w9015 = ~w9002 & ~w9014;
assign w9016 = pi0497 & w9015;
assign w9017 = ~pi0497 & ~w9015;
assign w9018 = ~w9016 & ~w9017;
assign w9019 = w8782 & w8839;
assign w9020 = ~w8847 & ~w9019;
assign w9021 = w8829 & w9020;
assign w9022 = (w8795 & ~w8825) | (w8795 & w64851) | (~w8825 & w64851);
assign w9023 = w8759 & w8780;
assign w9024 = ~w8753 & ~w9023;
assign w9025 = w8759 & w8795;
assign w9026 = ~w8848 & w64852;
assign w9027 = ~w9024 & w9026;
assign w9028 = w8766 & w8822;
assign w9029 = w8779 & w8813;
assign w9030 = ~w8777 & ~w8815;
assign w9031 = ~w8806 & ~w9029;
assign w9032 = (~w8795 & ~w9031) | (~w8795 & w64853) | (~w9031 & w64853);
assign w9033 = ~w8805 & ~w9028;
assign w9034 = ~w9027 & ~w9032;
assign w9035 = w9033 & w9034;
assign w9036 = w9035 & w64854;
assign w9037 = (pi0488 & ~w9035) | (pi0488 & w64855) | (~w9035 & w64855);
assign w9038 = ~w9036 & ~w9037;
assign w9039 = ~w8248 & ~w8265;
assign w9040 = w8282 & ~w9039;
assign w9041 = w9039 & w63366;
assign w9042 = ~w9040 & ~w9041;
assign w9043 = w8245 & w9042;
assign w9044 = ~w8245 & w8264;
assign w9045 = w9039 & w9044;
assign w9046 = ~w8270 & ~w9045;
assign w9047 = ~w9043 & w9046;
assign w9048 = w8212 & ~w9047;
assign w9049 = ~w8212 & ~w8263;
assign w9050 = ~w9042 & w9049;
assign w9051 = w8245 & ~w8270;
assign w9052 = ~w9050 & w9051;
assign w9053 = (w8218 & ~w9039) | (w8218 & w8275) | (~w9039 & w8275);
assign w9054 = ~w8225 & ~w8265;
assign w9055 = ~w8254 & ~w9054;
assign w9056 = ~w9053 & ~w9055;
assign w9057 = ~w8212 & ~w9056;
assign w9058 = ~w8245 & ~w8549;
assign w9059 = ~w9040 & w9058;
assign w9060 = ~w9057 & w9059;
assign w9061 = ~w9052 & ~w9060;
assign w9062 = ~w9048 & ~w9061;
assign w9063 = ~pi0507 & w9062;
assign w9064 = pi0507 & ~w9062;
assign w9065 = ~w9063 & ~w9064;
assign w9066 = w8765 & w8806;
assign w9067 = ~w9019 & ~w9023;
assign w9068 = w8799 & ~w9067;
assign w9069 = ~w8780 & w8798;
assign w9070 = ~w8816 & ~w9066;
assign w9071 = ~w9069 & w9070;
assign w9072 = ~w9068 & w9071;
assign w9073 = w8795 & ~w9072;
assign w9074 = w8795 & w9030;
assign w9075 = ~w8753 & ~w8803;
assign w9076 = w8765 & ~w8795;
assign w9077 = ~w8821 & w9076;
assign w9078 = w8817 & w9077;
assign w9079 = ~w9075 & ~w9078;
assign w9080 = ~w9074 & ~w9079;
assign w9081 = ~w9073 & ~w9080;
assign w9082 = pi0483 & ~w9081;
assign w9083 = ~pi0483 & w9081;
assign w9084 = ~w9082 & ~w9083;
assign w9085 = w8336 & w8458;
assign w9086 = ~w8403 & ~w9085;
assign w9087 = w8372 & ~w9086;
assign w9088 = w8348 & w8355;
assign w9089 = ~w8985 & ~w9088;
assign w9090 = w8983 & ~w9089;
assign w9091 = w8363 & w8372;
assign w9092 = ~w8376 & w9091;
assign w9093 = ~w9088 & w9092;
assign w9094 = ~w8462 & ~w9093;
assign w9095 = ~w8336 & ~w9094;
assign w9096 = ~w8348 & w8476;
assign w9097 = ~w8388 & ~w9096;
assign w9098 = ~w8405 & w9097;
assign w9099 = ~w8480 & w9098;
assign w9100 = ~w8372 & ~w9099;
assign w9101 = ~w9090 & ~w9095;
assign w9102 = ~w9087 & w9101;
assign w9103 = ~w9100 & w9102;
assign w9104 = pi0523 & ~w9103;
assign w9105 = ~pi0523 & w9103;
assign w9106 = ~w9104 & ~w9105;
assign w9107 = ~w8287 & ~w8546;
assign w9108 = ~w8245 & w9107;
assign w9109 = w8245 & w8254;
assign w9110 = (w9042 & w64856) | (w9042 & w64857) | (w64856 & w64857);
assign w9111 = ~w8259 & ~w8284;
assign w9112 = ~w9108 & w9111;
assign w9113 = ~w9110 & w9112;
assign w9114 = w8212 & ~w9113;
assign w9115 = w8265 & w8282;
assign w9116 = ~w8248 & w8546;
assign w9117 = w9054 & w9116;
assign w9118 = (~w8245 & w9117) | (~w8245 & w63607) | (w9117 & w63607);
assign w9119 = w8245 & ~w8282;
assign w9120 = (~w9115 & ~w9107) | (~w9115 & w64858) | (~w9107 & w64858);
assign w9121 = (~w8212 & w9118) | (~w8212 & w64859) | (w9118 & w64859);
assign w9122 = w8245 & ~w8259;
assign w9123 = ~w8256 & w8276;
assign w9124 = ~w9122 & ~w9123;
assign w9125 = ~w9121 & ~w9124;
assign w9126 = ~w9114 & w9125;
assign w9127 = ~pi0516 & w9126;
assign w9128 = pi0516 & ~w9126;
assign w9129 = ~w9127 & ~w9128;
assign w9130 = ~pi3473 & pi9040;
assign w9131 = ~pi3453 & ~pi9040;
assign w9132 = ~w9130 & ~w9131;
assign w9133 = pi0542 & ~w9132;
assign w9134 = ~pi0542 & w9132;
assign w9135 = ~w9133 & ~w9134;
assign w9136 = ~pi3440 & pi9040;
assign w9137 = ~pi3508 & ~pi9040;
assign w9138 = ~w9136 & ~w9137;
assign w9139 = pi0535 & ~w9138;
assign w9140 = ~pi0535 & w9138;
assign w9141 = ~w9139 & ~w9140;
assign w9142 = w9135 & w9141;
assign w9143 = ~pi3461 & pi9040;
assign w9144 = ~pi3449 & ~pi9040;
assign w9145 = ~w9143 & ~w9144;
assign w9146 = pi0543 & ~w9145;
assign w9147 = ~pi0543 & w9145;
assign w9148 = ~w9146 & ~w9147;
assign w9149 = w9142 & ~w9148;
assign w9150 = ~pi3459 & pi9040;
assign w9151 = ~pi3476 & ~pi9040;
assign w9152 = ~w9150 & ~w9151;
assign w9153 = pi0519 & ~w9152;
assign w9154 = ~pi0519 & w9152;
assign w9155 = ~w9153 & ~w9154;
assign w9156 = ~pi3445 & pi9040;
assign w9157 = ~pi3474 & ~pi9040;
assign w9158 = ~w9156 & ~w9157;
assign w9159 = pi0494 & ~w9158;
assign w9160 = ~pi0494 & w9158;
assign w9161 = ~w9159 & ~w9160;
assign w9162 = ~w9155 & ~w9161;
assign w9163 = ~w9135 & ~w9141;
assign w9164 = w9135 & ~w9161;
assign w9165 = ~w9135 & w9161;
assign w9166 = ~w9164 & ~w9165;
assign w9167 = ~w9142 & w9148;
assign w9168 = w9166 & w9167;
assign w9169 = (~w9162 & w9168) | (~w9162 & w63608) | (w9168 & w63608);
assign w9170 = ~w9135 & ~w9148;
assign w9171 = ~w9142 & ~w9170;
assign w9172 = ~w9166 & w9171;
assign w9173 = ~w9155 & w9172;
assign w9174 = ~w9169 & ~w9173;
assign w9175 = ~pi3460 & pi9040;
assign w9176 = ~pi3428 & ~pi9040;
assign w9177 = ~w9175 & ~w9176;
assign w9178 = pi0540 & ~w9177;
assign w9179 = ~pi0540 & w9177;
assign w9180 = ~w9178 & ~w9179;
assign w9181 = (w9180 & ~w9174) | (w9180 & w64860) | (~w9174 & w64860);
assign w9182 = ~w9141 & w9166;
assign w9183 = w9141 & ~w9166;
assign w9184 = ~w9182 & ~w9183;
assign w9185 = w9155 & w9184;
assign w9186 = w9141 & w9162;
assign w9187 = (~w9186 & ~w9184) | (~w9186 & w64861) | (~w9184 & w64861);
assign w9188 = ~w9148 & ~w9187;
assign w9189 = ~w9141 & ~w9155;
assign w9190 = w9135 & w9148;
assign w9191 = w9189 & w9190;
assign w9192 = ~w9135 & w9148;
assign w9193 = w9166 & w64862;
assign w9194 = w9192 & w9193;
assign w9195 = ~w9141 & w9161;
assign w9196 = w9135 & ~w9155;
assign w9197 = w9195 & w9196;
assign w9198 = w9141 & ~w9161;
assign w9199 = ~w9195 & ~w9198;
assign w9200 = w9142 & w9162;
assign w9201 = ~w9199 & ~w9200;
assign w9202 = w9148 & w9201;
assign w9203 = w9201 & w63609;
assign w9204 = ~w9197 & ~w9203;
assign w9205 = ~w9135 & ~w9189;
assign w9206 = ~w9148 & ~w9196;
assign w9207 = ~w9205 & w9206;
assign w9208 = w9141 & w9161;
assign w9209 = w9155 & w9208;
assign w9210 = ~w9207 & ~w9209;
assign w9211 = w9172 & ~w9210;
assign w9212 = ~w9170 & ~w9190;
assign w9213 = ~w9198 & w9212;
assign w9214 = ~w9155 & ~w9164;
assign w9215 = ~w9195 & w9214;
assign w9216 = ~w9213 & w9215;
assign w9217 = ~w9211 & ~w9216;
assign w9218 = (~w9180 & ~w9217) | (~w9180 & w63610) | (~w9217 & w63610);
assign w9219 = ~w9191 & ~w9194;
assign w9220 = ~w9181 & w9219;
assign w9221 = ~w9188 & ~w9218;
assign w9222 = (pi0553 & ~w9221) | (pi0553 & w64863) | (~w9221 & w64863);
assign w9223 = w9221 & w64864;
assign w9224 = ~w9222 & ~w9223;
assign w9225 = w9141 & ~w9174;
assign w9226 = w9141 & ~w9162;
assign w9227 = ~w9148 & w9166;
assign w9228 = ~w9226 & w9227;
assign w9229 = ~w9166 & ~w9199;
assign w9230 = w9155 & w9229;
assign w9231 = w9190 & w9199;
assign w9232 = ~w9180 & ~w9231;
assign w9233 = ~w9228 & w9232;
assign w9234 = ~w9230 & w9233;
assign w9235 = ~w9197 & ~w9205;
assign w9236 = w9148 & ~w9235;
assign w9237 = w9180 & ~w9200;
assign w9238 = w9210 & w9237;
assign w9239 = ~w9236 & w9238;
assign w9240 = ~w9234 & ~w9239;
assign w9241 = ~w9225 & ~w9240;
assign w9242 = ~pi0555 & w9241;
assign w9243 = pi0555 & ~w9241;
assign w9244 = ~w9242 & ~w9243;
assign w9245 = ~pi3474 & pi9040;
assign w9246 = ~pi3438 & ~pi9040;
assign w9247 = ~w9245 & ~w9246;
assign w9248 = pi0536 & ~w9247;
assign w9249 = ~pi0536 & w9247;
assign w9250 = ~w9248 & ~w9249;
assign w9251 = ~pi3434 & pi9040;
assign w9252 = ~pi3462 & ~pi9040;
assign w9253 = ~w9251 & ~w9252;
assign w9254 = pi0540 & ~w9253;
assign w9255 = ~pi0540 & w9253;
assign w9256 = ~w9254 & ~w9255;
assign w9257 = ~pi3453 & pi9040;
assign w9258 = ~pi3512 & ~pi9040;
assign w9259 = ~w9257 & ~w9258;
assign w9260 = pi0530 & ~w9259;
assign w9261 = ~pi0530 & w9259;
assign w9262 = ~w9260 & ~w9261;
assign w9263 = ~w9256 & w9262;
assign w9264 = ~pi3443 & pi9040;
assign w9265 = ~pi3460 & ~pi9040;
assign w9266 = ~w9264 & ~w9265;
assign w9267 = pi0494 & ~w9266;
assign w9268 = ~pi0494 & w9266;
assign w9269 = ~w9267 & ~w9268;
assign w9270 = w9263 & ~w9269;
assign w9271 = ~pi3511 & pi9040;
assign w9272 = ~pi3459 & ~pi9040;
assign w9273 = ~w9271 & ~w9272;
assign w9274 = pi0524 & ~w9273;
assign w9275 = ~pi0524 & w9273;
assign w9276 = ~w9274 & ~w9275;
assign w9277 = w9269 & ~w9276;
assign w9278 = w9256 & w9277;
assign w9279 = w9277 & w64865;
assign w9280 = w9269 & w9276;
assign w9281 = ~w9256 & w9280;
assign w9282 = ~w9256 & ~w9276;
assign w9283 = w9256 & w9276;
assign w9284 = ~w9269 & w9283;
assign w9285 = ~w9282 & ~w9284;
assign w9286 = ~w9281 & w9285;
assign w9287 = ~pi3430 & pi9040;
assign w9288 = ~pi3469 & ~pi9040;
assign w9289 = ~w9287 & ~w9288;
assign w9290 = pi0528 & ~w9289;
assign w9291 = ~pi0528 & w9289;
assign w9292 = ~w9290 & ~w9291;
assign w9293 = w9262 & ~w9269;
assign w9294 = ~w9276 & w9293;
assign w9295 = ~w9292 & ~w9294;
assign w9296 = w9286 & w9295;
assign w9297 = ~w9270 & ~w9279;
assign w9298 = ~w9296 & w9297;
assign w9299 = ~w9250 & ~w9298;
assign w9300 = w9263 & w64866;
assign w9301 = (~w9250 & ~w9283) | (~w9250 & w64867) | (~w9283 & w64867);
assign w9302 = w9256 & ~w9262;
assign w9303 = ~w9301 & w9302;
assign w9304 = w9250 & w9269;
assign w9305 = ~w9256 & ~w9304;
assign w9306 = ~w9278 & ~w9305;
assign w9307 = ~w9262 & w9269;
assign w9308 = w9282 & w9307;
assign w9309 = w9250 & ~w9308;
assign w9310 = ~w9276 & w9309;
assign w9311 = w9306 & w9310;
assign w9312 = ~w9262 & w9282;
assign w9313 = ~w9281 & ~w9312;
assign w9314 = ~w9250 & ~w9313;
assign w9315 = w9283 & w9304;
assign w9316 = w9292 & ~w9315;
assign w9317 = ~w9300 & w9316;
assign w9318 = ~w9303 & w9317;
assign w9319 = ~w9314 & w9318;
assign w9320 = ~w9311 & w9319;
assign w9321 = ~w9285 & w9293;
assign w9322 = w9250 & ~w9313;
assign w9323 = ~w9279 & ~w9292;
assign w9324 = ~w9321 & w9323;
assign w9325 = ~w9322 & w9324;
assign w9326 = ~w9320 & ~w9325;
assign w9327 = ~w9326 & w64868;
assign w9328 = (pi0551 & w9326) | (pi0551 & w64869) | (w9326 & w64869);
assign w9329 = ~w9327 & ~w9328;
assign w9330 = ~pi3448 & pi9040;
assign w9331 = ~pi3431 & ~pi9040;
assign w9332 = ~w9330 & ~w9331;
assign w9333 = pi0513 & ~w9332;
assign w9334 = ~pi0513 & w9332;
assign w9335 = ~w9333 & ~w9334;
assign w9336 = ~pi3479 & pi9040;
assign w9337 = ~pi3439 & ~pi9040;
assign w9338 = ~w9336 & ~w9337;
assign w9339 = pi0510 & ~w9338;
assign w9340 = ~pi0510 & w9338;
assign w9341 = ~w9339 & ~w9340;
assign w9342 = ~w9335 & ~w9341;
assign w9343 = ~pi3467 & pi9040;
assign w9344 = ~pi3470 & ~pi9040;
assign w9345 = ~w9343 & ~w9344;
assign w9346 = pi0527 & ~w9345;
assign w9347 = ~pi0527 & w9345;
assign w9348 = ~w9346 & ~w9347;
assign w9349 = w9342 & ~w9348;
assign w9350 = ~pi3463 & pi9040;
assign w9351 = ~pi3468 & ~pi9040;
assign w9352 = ~w9350 & ~w9351;
assign w9353 = pi0517 & ~w9352;
assign w9354 = ~pi0517 & w9352;
assign w9355 = ~w9353 & ~w9354;
assign w9356 = ~w9341 & w9355;
assign w9357 = ~pi3442 & pi9040;
assign w9358 = ~pi3481 & ~pi9040;
assign w9359 = ~w9357 & ~w9358;
assign w9360 = pi0521 & ~w9359;
assign w9361 = ~pi0521 & w9359;
assign w9362 = ~w9360 & ~w9361;
assign w9363 = ~w9348 & ~w9362;
assign w9364 = w9356 & w9363;
assign w9365 = w9348 & ~w9362;
assign w9366 = ~w9348 & w9362;
assign w9367 = ~w9365 & ~w9366;
assign w9368 = ~w9355 & w9367;
assign w9369 = (~w9335 & ~w9367) | (~w9335 & w63611) | (~w9367 & w63611);
assign w9370 = ~w9341 & w9348;
assign w9371 = ~w9355 & ~w9370;
assign w9372 = w9348 & w9356;
assign w9373 = ~w9371 & ~w9372;
assign w9374 = w9369 & ~w9373;
assign w9375 = ~w9364 & ~w9374;
assign w9376 = w9349 & w9375;
assign w9377 = ~pi3447 & pi9040;
assign w9378 = ~pi3510 & ~pi9040;
assign w9379 = ~w9377 & ~w9378;
assign w9380 = pi0531 & ~w9379;
assign w9381 = ~pi0531 & w9379;
assign w9382 = ~w9380 & ~w9381;
assign w9383 = w9342 & w64870;
assign w9384 = ~w9335 & ~w9362;
assign w9385 = ~w9355 & w9365;
assign w9386 = ~w9341 & ~w9355;
assign w9387 = w9335 & ~w9386;
assign w9388 = ~w9385 & w9387;
assign w9389 = w9341 & w9355;
assign w9390 = ~w9386 & ~w9389;
assign w9391 = ~w9335 & ~w9390;
assign w9392 = ~w9388 & ~w9391;
assign w9393 = ~w9362 & w9389;
assign w9394 = w9366 & w9389;
assign w9395 = ~w9341 & w9366;
assign w9396 = (~w9348 & ~w9366) | (~w9348 & w63367) | (~w9366 & w63367);
assign w9397 = ~w9355 & w9362;
assign w9398 = ~w9396 & w9397;
assign w9399 = ~w9394 & ~w9398;
assign w9400 = ~w9367 & ~w9371;
assign w9401 = ~w9370 & w9400;
assign w9402 = w9399 & w9401;
assign w9403 = (~w9392 & w64871) | (~w9392 & w64872) | (w64871 & w64872);
assign w9404 = ~w9402 & w9403;
assign w9405 = ~w9382 & ~w9404;
assign w9406 = w9341 & ~w9362;
assign w9407 = ~w9386 & ~w9406;
assign w9408 = ~w9400 & w9407;
assign w9409 = w9348 & w9389;
assign w9410 = w9365 & w9386;
assign w9411 = ~w9409 & ~w9410;
assign w9412 = (~w9335 & w9408) | (~w9335 & w63613) | (w9408 & w63613);
assign w9413 = (~w9400 & w64873) | (~w9400 & w64874) | (w64873 & w64874);
assign w9414 = ~w9355 & w9395;
assign w9415 = w9411 & ~w9414;
assign w9416 = ~w9413 & w9415;
assign w9417 = ~w9349 & ~w9412;
assign w9418 = ~w9416 & w9417;
assign w9419 = ~w9376 & ~w9418;
assign w9420 = (pi0549 & ~w9419) | (pi0549 & w64875) | (~w9419 & w64875);
assign w9421 = w9419 & w64876;
assign w9422 = ~w9420 & ~w9421;
assign w9423 = ~pi3433 & pi9040;
assign w9424 = ~pi3463 & ~pi9040;
assign w9425 = ~w9423 & ~w9424;
assign w9426 = pi0542 & ~w9425;
assign w9427 = ~pi0542 & w9425;
assign w9428 = ~w9426 & ~w9427;
assign w9429 = ~pi3431 & pi9040;
assign w9430 = ~pi3450 & ~pi9040;
assign w9431 = ~w9429 & ~w9430;
assign w9432 = pi0515 & ~w9431;
assign w9433 = ~pi0515 & w9431;
assign w9434 = ~w9432 & ~w9433;
assign w9435 = ~pi3477 & pi9040;
assign w9436 = ~pi3478 & ~pi9040;
assign w9437 = ~w9435 & ~w9436;
assign w9438 = pi0518 & ~w9437;
assign w9439 = ~pi0518 & w9437;
assign w9440 = ~w9438 & ~w9439;
assign w9441 = w9434 & ~w9440;
assign w9442 = ~pi3432 & pi9040;
assign w9443 = ~pi3479 & ~pi9040;
assign w9444 = ~w9442 & ~w9443;
assign w9445 = pi0539 & ~w9444;
assign w9446 = ~pi0539 & w9444;
assign w9447 = ~w9445 & ~w9446;
assign w9448 = w9441 & w9447;
assign w9449 = ~w9434 & ~w9440;
assign w9450 = ~w9447 & w9449;
assign w9451 = ~w9448 & ~w9450;
assign w9452 = ~pi3471 & pi9040;
assign w9453 = ~pi3466 & ~pi9040;
assign w9454 = ~w9452 & ~w9453;
assign w9455 = pi0509 & ~w9454;
assign w9456 = ~pi0509 & w9454;
assign w9457 = ~w9455 & ~w9456;
assign w9458 = w9434 & ~w9447;
assign w9459 = ~pi3425 & pi9040;
assign w9460 = ~pi3447 & ~pi9040;
assign w9461 = ~w9459 & ~w9460;
assign w9462 = pi0535 & ~w9461;
assign w9463 = ~pi0535 & w9461;
assign w9464 = ~w9462 & ~w9463;
assign w9465 = w9440 & ~w9464;
assign w9466 = ~w9458 & ~w9465;
assign w9467 = ~w9447 & w9465;
assign w9468 = (w9457 & ~w9465) | (w9457 & w64877) | (~w9465 & w64877);
assign w9469 = w9434 & ~w9464;
assign w9470 = w9457 & ~w9469;
assign w9471 = ~w9468 & ~w9470;
assign w9472 = ~w9466 & ~w9471;
assign w9473 = ~w9434 & w9440;
assign w9474 = w9447 & w9473;
assign w9475 = w9473 & w9491;
assign w9476 = (~w9475 & w9451) | (~w9475 & w64878) | (w9451 & w64878);
assign w9477 = ~w9472 & w9476;
assign w9478 = w9428 & ~w9477;
assign w9479 = ~w9447 & w9464;
assign w9480 = ~w9440 & w9479;
assign w9481 = w9473 & w9484;
assign w9482 = ~w9480 & ~w9481;
assign w9483 = ~w9449 & w9482;
assign w9484 = w9447 & ~w9464;
assign w9485 = ~w9479 & ~w9484;
assign w9486 = w9434 & w9440;
assign w9487 = ~w9464 & w9486;
assign w9488 = ~w9449 & ~w9487;
assign w9489 = (w9457 & w9488) | (w9457 & w64879) | (w9488 & w64879);
assign w9490 = ~w9483 & w9489;
assign w9491 = w9447 & w9464;
assign w9492 = w9486 & w9491;
assign w9493 = w9458 & ~w9468;
assign w9494 = w9449 & w9464;
assign w9495 = (w9457 & ~w9449) | (w9457 & w64880) | (~w9449 & w64880);
assign w9496 = w9441 & w9484;
assign w9497 = w9495 & ~w9496;
assign w9498 = w9440 & w9464;
assign w9499 = ~w9434 & w9484;
assign w9500 = ~w9457 & ~w9498;
assign w9501 = ~w9499 & w9500;
assign w9502 = ~w9497 & ~w9501;
assign w9503 = ~w9492 & ~w9493;
assign w9504 = ~w9502 & w9503;
assign w9505 = ~w9428 & ~w9504;
assign w9506 = w9434 & ~w9457;
assign w9507 = w9467 & w9506;
assign w9508 = ~w9490 & ~w9507;
assign w9509 = ~w9478 & w9508;
assign w9510 = ~w9505 & w9509;
assign w9511 = pi0544 & ~w9510;
assign w9512 = ~pi0544 & w9510;
assign w9513 = ~w9511 & ~w9512;
assign w9514 = (~w9363 & w9400) | (~w9363 & w63368) | (w9400 & w63368);
assign w9515 = w9367 & w63614;
assign w9516 = (w9335 & w9514) | (w9335 & w63615) | (w9514 & w63615);
assign w9517 = (~w9335 & ~w9356) | (~w9335 & w64881) | (~w9356 & w64881);
assign w9518 = (w9517 & w9399) | (w9517 & w63616) | (w9399 & w63616);
assign w9519 = ~w9516 & ~w9518;
assign w9520 = ~w9370 & w9385;
assign w9521 = (~w9382 & w9519) | (~w9382 & w64882) | (w9519 & w64882);
assign w9522 = w9335 & w9362;
assign w9523 = w9370 & w9522;
assign w9524 = ~w9355 & w9396;
assign w9525 = ~w9409 & ~w9524;
assign w9526 = (w9406 & w9524) | (w9406 & w63617) | (w9524 & w63617);
assign w9527 = (w9335 & w9398) | (w9335 & w64883) | (w9398 & w64883);
assign w9528 = ~w9383 & ~w9410;
assign w9529 = ~w9526 & w9528;
assign w9530 = (w9382 & ~w9529) | (w9382 & w64884) | (~w9529 & w64884);
assign w9531 = ~w9335 & w9382;
assign w9532 = ~w9525 & w9531;
assign w9533 = ~w9364 & ~w9523;
assign w9534 = ~w9532 & w9533;
assign w9535 = ~w9530 & w9534;
assign w9536 = ~w9521 & w9535;
assign w9537 = pi0547 & w9536;
assign w9538 = ~pi0547 & ~w9536;
assign w9539 = ~w9537 & ~w9538;
assign w9540 = ~w9270 & ~w9307;
assign w9541 = w9250 & w9256;
assign w9542 = ~w9310 & ~w9541;
assign w9543 = ~w9540 & ~w9542;
assign w9544 = ~w9263 & w9304;
assign w9545 = ~w9250 & ~w9269;
assign w9546 = w9282 & w9545;
assign w9547 = ~w9250 & w9262;
assign w9548 = ~w9285 & w9547;
assign w9549 = ~w9262 & w9276;
assign w9550 = w9545 & w9549;
assign w9551 = w9263 & w9280;
assign w9552 = ~w9550 & ~w9551;
assign w9553 = w9305 & ~w9552;
assign w9554 = ~w9269 & ~w9276;
assign w9555 = ~w9280 & ~w9554;
assign w9556 = w9302 & ~w9555;
assign w9557 = w9292 & ~w9544;
assign w9558 = ~w9546 & w9557;
assign w9559 = ~w9556 & w9558;
assign w9560 = ~w9548 & ~w9553;
assign w9561 = w9559 & w9560;
assign w9562 = ~w9292 & w9552;
assign w9563 = ~w9283 & w9555;
assign w9564 = w9555 & w64885;
assign w9565 = w9286 & w9547;
assign w9566 = w9262 & w9284;
assign w9567 = w9250 & w9566;
assign w9568 = w9562 & ~w9564;
assign w9569 = ~w9567 & w9568;
assign w9570 = ~w9565 & w9569;
assign w9571 = (~w9543 & w9570) | (~w9543 & w64886) | (w9570 & w64886);
assign w9572 = pi0563 & w9571;
assign w9573 = ~pi0563 & ~w9571;
assign w9574 = ~w9572 & ~w9573;
assign w9575 = w9192 & w9198;
assign w9576 = ~w9148 & w9229;
assign w9577 = ~w9575 & ~w9576;
assign w9578 = ~w9155 & ~w9577;
assign w9579 = ~w9149 & ~w9209;
assign w9580 = ~w9161 & w9189;
assign w9581 = ~w9575 & ~w9580;
assign w9582 = w9579 & w9581;
assign w9583 = ~w9180 & ~w9582;
assign w9584 = ~w9142 & w9180;
assign w9585 = w9155 & w9161;
assign w9586 = w9212 & w9585;
assign w9587 = ~w9584 & w9586;
assign w9588 = ~w9201 & w9236;
assign w9589 = w9206 & ~w9208;
assign w9590 = w9184 & w9589;
assign w9591 = ~w9588 & ~w9590;
assign w9592 = (w9180 & ~w9591) | (w9180 & w64887) | (~w9591 & w64887);
assign w9593 = ~w9191 & ~w9587;
assign w9594 = ~w9583 & w9593;
assign w9595 = ~w9578 & w9594;
assign w9596 = ~w9592 & w9595;
assign w9597 = pi0565 & w9596;
assign w9598 = ~pi0565 & ~w9596;
assign w9599 = ~w9597 & ~w9598;
assign w9600 = ~w9167 & w9199;
assign w9601 = (w9600 & ~w9184) | (w9600 & w64888) | (~w9184 & w64888);
assign w9602 = ~w9579 & w9601;
assign w9603 = ~w9155 & w9167;
assign w9604 = w9199 & w9603;
assign w9605 = w9237 & ~w9604;
assign w9606 = ~w9185 & w9605;
assign w9607 = ~w9180 & ~w9193;
assign w9608 = ~w9202 & w9607;
assign w9609 = ~w9601 & w9608;
assign w9610 = ~w9606 & ~w9609;
assign w9611 = ~w9602 & ~w9610;
assign w9612 = pi0561 & w9611;
assign w9613 = ~pi0561 & ~w9611;
assign w9614 = ~w9612 & ~w9613;
assign w9615 = ~pi3428 & pi9040;
assign w9616 = ~pi3434 & ~pi9040;
assign w9617 = ~w9615 & ~w9616;
assign w9618 = pi0512 & ~w9617;
assign w9619 = ~pi0512 & w9617;
assign w9620 = ~w9618 & ~w9619;
assign w9621 = ~pi3512 & pi9040;
assign w9622 = ~pi3440 & ~pi9040;
assign w9623 = ~w9621 & ~w9622;
assign w9624 = pi0520 & ~w9623;
assign w9625 = ~pi0520 & w9623;
assign w9626 = ~w9624 & ~w9625;
assign w9627 = w9620 & ~w9626;
assign w9628 = ~pi3437 & pi9040;
assign w9629 = ~pi3443 & ~pi9040;
assign w9630 = ~w9628 & ~w9629;
assign w9631 = pi0541 & ~w9630;
assign w9632 = ~pi0541 & w9630;
assign w9633 = ~w9631 & ~w9632;
assign w9634 = ~pi3438 & pi9040;
assign w9635 = ~pi3509 & ~pi9040;
assign w9636 = ~w9634 & ~w9635;
assign w9637 = pi0532 & ~w9636;
assign w9638 = ~pi0532 & w9636;
assign w9639 = ~w9637 & ~w9638;
assign w9640 = ~w9633 & w9639;
assign w9641 = w9627 & w9640;
assign w9642 = ~pi3444 & pi9040;
assign w9643 = ~pi3430 & ~pi9040;
assign w9644 = ~w9642 & ~w9643;
assign w9645 = pi0526 & ~w9644;
assign w9646 = ~pi0526 & w9644;
assign w9647 = ~w9645 & ~w9646;
assign w9648 = w9620 & ~w9639;
assign w9649 = w9626 & ~w9633;
assign w9650 = w9648 & w9649;
assign w9651 = w9647 & ~w9650;
assign w9652 = ~w9641 & w9651;
assign w9653 = ~w9620 & w9639;
assign w9654 = ~w9626 & ~w9653;
assign w9655 = w9649 & w9653;
assign w9656 = ~w9633 & ~w9648;
assign w9657 = ~w9654 & w9656;
assign w9658 = (~w9647 & ~w9657) | (~w9647 & w64889) | (~w9657 & w64889);
assign w9659 = ~w9652 & ~w9658;
assign w9660 = ~pi3436 & pi9040;
assign w9661 = ~pi3473 & ~pi9040;
assign w9662 = ~w9660 & ~w9661;
assign w9663 = pi0537 & ~w9662;
assign w9664 = ~pi0537 & w9662;
assign w9665 = ~w9663 & ~w9664;
assign w9666 = w9620 & ~w9647;
assign w9667 = ~w9639 & ~w9666;
assign w9668 = w9633 & ~w9647;
assign w9669 = w9620 & w9639;
assign w9670 = ~w9668 & w9669;
assign w9671 = ~w9626 & w9633;
assign w9672 = ~w9649 & ~w9671;
assign w9673 = ~w9667 & ~w9670;
assign w9674 = w9672 & w9673;
assign w9675 = w9620 & ~w9671;
assign w9676 = ~w9639 & ~w9647;
assign w9677 = w9654 & ~w9676;
assign w9678 = ~w9675 & w9677;
assign w9679 = w9665 & ~w9674;
assign w9680 = ~w9678 & w9679;
assign w9681 = ~w9675 & w9676;
assign w9682 = ~w9639 & w9649;
assign w9683 = ~w9620 & w9626;
assign w9684 = ~w9633 & ~w9683;
assign w9685 = w9639 & w9647;
assign w9686 = ~w9684 & w9685;
assign w9687 = ~w9627 & w9686;
assign w9688 = ~w9641 & ~w9665;
assign w9689 = ~w9682 & w9688;
assign w9690 = ~w9681 & w9689;
assign w9691 = ~w9687 & w9690;
assign w9692 = ~w9680 & ~w9691;
assign w9693 = ~w9659 & ~w9692;
assign w9694 = pi0557 & w9693;
assign w9695 = ~pi0557 & ~w9693;
assign w9696 = ~w9694 & ~w9695;
assign w9697 = ~pi3450 & pi9040;
assign w9698 = ~pi3467 & ~pi9040;
assign w9699 = ~w9697 & ~w9698;
assign w9700 = pi0517 & ~w9699;
assign w9701 = ~pi0517 & w9699;
assign w9702 = ~w9700 & ~w9701;
assign w9703 = ~pi3468 & pi9040;
assign w9704 = ~pi3425 & ~pi9040;
assign w9705 = ~w9703 & ~w9704;
assign w9706 = pi0538 & ~w9705;
assign w9707 = ~pi0538 & w9705;
assign w9708 = ~w9706 & ~w9707;
assign w9709 = ~pi3481 & pi9040;
assign w9710 = ~pi3477 & ~pi9040;
assign w9711 = ~w9709 & ~w9710;
assign w9712 = pi0537 & ~w9711;
assign w9713 = ~pi0537 & w9711;
assign w9714 = ~w9712 & ~w9713;
assign w9715 = ~pi3429 & pi9040;
assign w9716 = ~pi3426 & ~pi9040;
assign w9717 = ~w9715 & ~w9716;
assign w9718 = pi0521 & ~w9717;
assign w9719 = ~pi0521 & w9717;
assign w9720 = ~w9718 & ~w9719;
assign w9721 = w9714 & ~w9720;
assign w9722 = ~pi3439 & pi9040;
assign w9723 = ~pi3427 & ~pi9040;
assign w9724 = ~w9722 & ~w9723;
assign w9725 = pi0512 & ~w9724;
assign w9726 = ~pi0512 & w9724;
assign w9727 = ~w9725 & ~w9726;
assign w9728 = w9721 & w63618;
assign w9729 = ~pi3466 & pi9040;
assign w9730 = ~pi3435 & ~pi9040;
assign w9731 = ~w9729 & ~w9730;
assign w9732 = pi0534 & ~w9731;
assign w9733 = ~pi0534 & w9731;
assign w9734 = ~w9732 & ~w9733;
assign w9735 = w9714 & w9720;
assign w9736 = ~w9727 & w9735;
assign w9737 = (~w9734 & ~w9735) | (~w9734 & w64890) | (~w9735 & w64890);
assign w9738 = ~w9708 & ~w9714;
assign w9739 = w9727 & w9738;
assign w9740 = w9737 & ~w9739;
assign w9741 = ~w9720 & ~w9727;
assign w9742 = ~w9708 & w9714;
assign w9743 = w9741 & w9742;
assign w9744 = w9734 & ~w9743;
assign w9745 = w9720 & w9727;
assign w9746 = w9714 & w9745;
assign w9747 = w9744 & ~w9746;
assign w9748 = ~w9714 & ~w9727;
assign w9749 = w9708 & ~w9714;
assign w9750 = ~w9741 & ~w9745;
assign w9751 = w9749 & w9750;
assign w9752 = (~w9748 & ~w9750) | (~w9748 & w64891) | (~w9750 & w64891);
assign w9753 = (~w9740 & ~w9747) | (~w9740 & w64892) | (~w9747 & w64892);
assign w9754 = ~w9708 & w9745;
assign w9755 = ~w9728 & ~w9754;
assign w9756 = ~w9753 & w9755;
assign w9757 = w9702 & ~w9756;
assign w9758 = ~w9714 & ~w9720;
assign w9759 = w9708 & ~w9727;
assign w9760 = w9758 & w9759;
assign w9761 = ~w9728 & ~w9760;
assign w9762 = w9708 & w9720;
assign w9763 = ~w9758 & ~w9762;
assign w9764 = w9748 & w9763;
assign w9765 = w9761 & ~w9764;
assign w9766 = w9734 & ~w9765;
assign w9767 = ~w9734 & w9759;
assign w9768 = ~w9754 & ~w9767;
assign w9769 = w9714 & ~w9768;
assign w9770 = ~w9720 & w9734;
assign w9771 = w9749 & ~w9770;
assign w9772 = (w9727 & ~w9770) | (w9727 & w63618) | (~w9770 & w63618);
assign w9773 = ~w9771 & w9772;
assign w9774 = ~w9714 & ~w9734;
assign w9775 = ~w9708 & w9774;
assign w9776 = w9737 & w9763;
assign w9777 = ~w9727 & ~w9775;
assign w9778 = ~w9776 & w9777;
assign w9779 = ~w9702 & ~w9773;
assign w9780 = ~w9778 & w9779;
assign w9781 = ~w9766 & ~w9769;
assign w9782 = ~w9780 & w9781;
assign w9783 = ~w9757 & w9782;
assign w9784 = pi0556 & ~w9783;
assign w9785 = ~pi0556 & w9783;
assign w9786 = ~w9784 & ~w9785;
assign w9787 = w9392 & w9400;
assign w9788 = w9362 & w9409;
assign w9789 = w9356 & w9362;
assign w9790 = ~w9385 & ~w9789;
assign w9791 = w9335 & ~w9790;
assign w9792 = w9335 & w9368;
assign w9793 = ~w9369 & ~w9791;
assign w9794 = (~w9788 & ~w9793) | (~w9788 & w64893) | (~w9793 & w64893);
assign w9795 = ~w9382 & ~w9794;
assign w9796 = w9355 & w9384;
assign w9797 = ~w9395 & ~w9410;
assign w9798 = ~w9796 & w9797;
assign w9799 = ~w9515 & w9798;
assign w9800 = (w9382 & ~w9799) | (w9382 & w64894) | (~w9799 & w64894);
assign w9801 = ~w9787 & ~w9800;
assign w9802 = ~w9795 & w9801;
assign w9803 = ~pi0559 & w9802;
assign w9804 = pi0559 & ~w9802;
assign w9805 = ~w9803 & ~w9804;
assign w9806 = w9721 & w9759;
assign w9807 = ~w9734 & w9806;
assign w9808 = ~w9714 & w9763;
assign w9809 = w9737 & ~w9808;
assign w9810 = ~w9747 & ~w9809;
assign w9811 = w9745 & w9774;
assign w9812 = ~w9739 & ~w9811;
assign w9813 = w9761 & w9812;
assign w9814 = (~w9702 & w9810) | (~w9702 & w64895) | (w9810 & w64895);
assign w9815 = ~w9720 & w9748;
assign w9816 = w9748 & w64896;
assign w9817 = ~w9736 & ~w9816;
assign w9818 = w9734 & ~w9817;
assign w9819 = ~w9734 & w9742;
assign w9820 = ~w9751 & ~w9819;
assign w9821 = ~w9818 & w9820;
assign w9822 = w9702 & ~w9821;
assign w9823 = w9708 & w9735;
assign w9824 = ~w9739 & ~w9823;
assign w9825 = w9734 & ~w9741;
assign w9826 = ~w9758 & w9825;
assign w9827 = w9824 & w9826;
assign w9828 = w9759 & w9827;
assign w9829 = (~w9807 & ~w9747) | (~w9807 & w64897) | (~w9747 & w64897);
assign w9830 = ~w9828 & w9829;
assign w9831 = ~w9814 & w9830;
assign w9832 = ~w9822 & w9831;
assign w9833 = pi0545 & w9832;
assign w9834 = ~pi0545 & ~w9832;
assign w9835 = ~w9833 & ~w9834;
assign w9836 = ~pi3424 & pi9040;
assign w9837 = ~pi3444 & ~pi9040;
assign w9838 = ~w9836 & ~w9837;
assign w9839 = pi0524 & ~w9838;
assign w9840 = ~pi0524 & w9838;
assign w9841 = ~w9839 & ~w9840;
assign w9842 = ~pi3509 & pi9040;
assign w9843 = ~pi3441 & ~pi9040;
assign w9844 = ~w9842 & ~w9843;
assign w9845 = pi0532 & ~w9844;
assign w9846 = ~pi0532 & w9844;
assign w9847 = ~w9845 & ~w9846;
assign w9848 = w9841 & ~w9847;
assign w9849 = ~w9841 & w9847;
assign w9850 = ~w9848 & ~w9849;
assign w9851 = ~pi3446 & pi9040;
assign w9852 = ~pi3461 & ~pi9040;
assign w9853 = ~w9851 & ~w9852;
assign w9854 = pi0528 & ~w9853;
assign w9855 = ~pi0528 & w9853;
assign w9856 = ~w9854 & ~w9855;
assign w9857 = w9850 & w9856;
assign w9858 = ~pi3462 & pi9040;
assign w9859 = ~pi3445 & ~pi9040;
assign w9860 = ~w9858 & ~w9859;
assign w9861 = pi0525 & ~w9860;
assign w9862 = ~pi0525 & w9860;
assign w9863 = ~w9861 & ~w9862;
assign w9864 = (~w9863 & ~w9850) | (~w9863 & w64898) | (~w9850 & w64898);
assign w9865 = ~pi3472 & pi9040;
assign w9866 = ~pi3437 & ~pi9040;
assign w9867 = ~w9865 & ~w9866;
assign w9868 = pi0520 & ~w9867;
assign w9869 = ~pi0520 & w9867;
assign w9870 = ~w9868 & ~w9869;
assign w9871 = ~w9864 & ~w9870;
assign w9872 = w9848 & ~w9856;
assign w9873 = ~pi3476 & pi9040;
assign w9874 = ~pi3436 & ~pi9040;
assign w9875 = ~w9873 & ~w9874;
assign w9876 = pi0533 & ~w9875;
assign w9877 = ~pi0533 & w9875;
assign w9878 = ~w9876 & ~w9877;
assign w9879 = w9856 & w9878;
assign w9880 = ~w9841 & w9879;
assign w9881 = ~w9847 & ~w9878;
assign w9882 = w9847 & w9878;
assign w9883 = ~w9856 & ~w9881;
assign w9884 = ~w9882 & w9883;
assign w9885 = ~w9872 & ~w9880;
assign w9886 = ~w9884 & w9885;
assign w9887 = w9871 & ~w9886;
assign w9888 = w9856 & w9881;
assign w9889 = ~w9841 & w9888;
assign w9890 = w9863 & w9889;
assign w9891 = ~w9841 & ~w9878;
assign w9892 = ~w9847 & ~w9856;
assign w9893 = w9847 & w9856;
assign w9894 = ~w9892 & ~w9893;
assign w9895 = ~w9856 & w9863;
assign w9896 = w9894 & ~w9895;
assign w9897 = w9891 & w9896;
assign w9898 = ~w9863 & ~w9891;
assign w9899 = ~w9894 & w9898;
assign w9900 = ~w9897 & ~w9899;
assign w9901 = w9870 & ~w9900;
assign w9902 = ~w9863 & w9870;
assign w9903 = w9841 & ~w9878;
assign w9904 = ~w9864 & w9903;
assign w9905 = w9886 & ~w9902;
assign w9906 = w9905 & w64899;
assign w9907 = ~w9863 & ~w9879;
assign w9908 = ~w9872 & w9907;
assign w9909 = (w9863 & ~w9883) | (w9863 & w64900) | (~w9883 & w64900);
assign w9910 = ~w9889 & w9909;
assign w9911 = ~w9908 & ~w9910;
assign w9912 = w9841 & w9847;
assign w9913 = w9911 & w9912;
assign w9914 = ~w9887 & ~w9890;
assign w9915 = ~w9901 & w9914;
assign w9916 = ~w9906 & ~w9913;
assign w9917 = w9915 & w9916;
assign w9918 = pi0574 & ~w9917;
assign w9919 = ~pi0574 & w9917;
assign w9920 = ~w9918 & ~w9919;
assign w9921 = ~pi3475 & pi9040;
assign w9922 = ~pi3442 & ~pi9040;
assign w9923 = ~w9921 & ~w9922;
assign w9924 = pi0514 & ~w9923;
assign w9925 = ~pi0514 & w9923;
assign w9926 = ~w9924 & ~w9925;
assign w9927 = ~pi3465 & pi9040;
assign w9928 = ~pi3448 & ~pi9040;
assign w9929 = ~w9927 & ~w9928;
assign w9930 = pi0531 & ~w9929;
assign w9931 = ~pi0531 & w9929;
assign w9932 = ~w9930 & ~w9931;
assign w9933 = w9926 & ~w9932;
assign w9934 = ~pi3470 & pi9040;
assign w9935 = ~pi3432 & ~pi9040;
assign w9936 = ~w9934 & ~w9935;
assign w9937 = pi0527 & ~w9936;
assign w9938 = ~pi0527 & w9936;
assign w9939 = ~w9937 & ~w9938;
assign w9940 = ~pi3427 & pi9040;
assign w9941 = ~pi3451 & ~pi9040;
assign w9942 = ~w9940 & ~w9941;
assign w9943 = pi0518 & ~w9942;
assign w9944 = ~pi0518 & w9942;
assign w9945 = ~w9943 & ~w9944;
assign w9946 = ~w9939 & ~w9945;
assign w9947 = ~w9933 & w9946;
assign w9948 = w9939 & w9945;
assign w9949 = ~w9946 & ~w9948;
assign w9950 = w9933 & w9949;
assign w9951 = ~w9947 & ~w9950;
assign w9952 = ~pi3426 & pi9040;
assign w9953 = ~pi3433 & ~pi9040;
assign w9954 = ~w9952 & ~w9953;
assign w9955 = pi0529 & ~w9954;
assign w9956 = ~pi0529 & w9954;
assign w9957 = ~w9955 & ~w9956;
assign w9958 = ~w9951 & w9957;
assign w9959 = ~pi3510 & pi9040;
assign w9960 = ~pi3482 & ~pi9040;
assign w9961 = ~w9959 & ~w9960;
assign w9962 = pi0515 & ~w9961;
assign w9963 = ~pi0515 & w9961;
assign w9964 = ~w9962 & ~w9963;
assign w9965 = ~w9932 & w9947;
assign w9966 = ~w9926 & w9932;
assign w9967 = ~w9933 & ~w9966;
assign w9968 = ~w9939 & w9967;
assign w9969 = w9967 & w64901;
assign w9970 = w9948 & w9966;
assign w9971 = ~w9969 & ~w9970;
assign w9972 = w9957 & ~w9971;
assign w9973 = ~w9939 & w9945;
assign w9974 = w9933 & w9973;
assign w9975 = ~w9965 & ~w9974;
assign w9976 = ~w9972 & w9975;
assign w9977 = w9964 & ~w9976;
assign w9978 = ~w9939 & w9957;
assign w9979 = ~w9946 & ~w9978;
assign w9980 = w9966 & ~w9979;
assign w9981 = w9945 & ~w9978;
assign w9982 = w9967 & w9981;
assign w9983 = w9932 & ~w9945;
assign w9984 = ~w9946 & ~w9983;
assign w9985 = ~w9957 & ~w9984;
assign w9986 = w9951 & w9985;
assign w9987 = ~w9980 & ~w9982;
assign w9988 = (~w9964 & w9986) | (~w9964 & w63619) | (w9986 & w63619);
assign w9989 = w9939 & w9967;
assign w9990 = ~w9932 & w9945;
assign w9991 = ~w9983 & ~w9990;
assign w9992 = w9939 & ~w9991;
assign w9993 = w9932 & w9973;
assign w9994 = ~w9992 & ~w9993;
assign w9995 = ~w9926 & w9945;
assign w9996 = w9949 & ~w9995;
assign w9997 = (w9964 & ~w9949) | (w9964 & w64902) | (~w9949 & w64902);
assign w9998 = (~w9989 & w9994) | (~w9989 & w64903) | (w9994 & w64903);
assign w9999 = ~w9957 & ~w9998;
assign w10000 = ~w9958 & ~w9988;
assign w10001 = ~w9999 & w10000;
assign w10002 = w10001 & w64904;
assign w10003 = (pi0548 & ~w10001) | (pi0548 & w64905) | (~w10001 & w64905);
assign w10004 = ~w10002 & ~w10003;
assign w10005 = w9683 & w9685;
assign w10006 = ~w9626 & ~w9639;
assign w10007 = w9626 & w9639;
assign w10008 = ~w10006 & ~w10007;
assign w10009 = ~w9633 & ~w9647;
assign w10010 = w10008 & w10009;
assign w10011 = ~w9648 & ~w9668;
assign w10012 = w9654 & ~w9666;
assign w10013 = ~w10011 & w10012;
assign w10014 = w9669 & w9672;
assign w10015 = w9665 & ~w10005;
assign w10016 = ~w10010 & w10015;
assign w10017 = ~w10014 & w10016;
assign w10018 = ~w10013 & w10017;
assign w10019 = w9672 & ~w10007;
assign w10020 = w9647 & ~w9683;
assign w10021 = ~w10019 & w10020;
assign w10022 = ~w10019 & w64906;
assign w10023 = w9653 & w9671;
assign w10024 = ~w9665 & ~w10023;
assign w10025 = w10006 & w10011;
assign w10026 = ~w9640 & w9683;
assign w10027 = ~w9648 & ~w10026;
assign w10028 = w9658 & ~w10027;
assign w10029 = ~w9650 & w10024;
assign w10030 = ~w10025 & w10029;
assign w10031 = ~w10022 & w10030;
assign w10032 = ~w10028 & w10031;
assign w10033 = ~w10018 & ~w10032;
assign w10034 = ~w9633 & w10005;
assign w10035 = ~w9620 & w9647;
assign w10036 = w10019 & w10035;
assign w10037 = ~w9641 & ~w10036;
assign w10038 = ~w9685 & ~w10037;
assign w10039 = ~w10034 & ~w10038;
assign w10040 = (pi0554 & w10033) | (pi0554 & w64907) | (w10033 & w64907);
assign w10041 = ~w10033 & w64908;
assign w10042 = ~w10040 & ~w10041;
assign w10043 = ~w9672 & w9686;
assign w10044 = w9633 & ~w10008;
assign w10045 = w9620 & w10044;
assign w10046 = ~w9653 & ~w9682;
assign w10047 = w10020 & ~w10046;
assign w10048 = ~w9641 & ~w10026;
assign w10049 = ~w9647 & ~w10048;
assign w10050 = w9665 & ~w10045;
assign w10051 = ~w10047 & ~w10049;
assign w10052 = w10050 & w10051;
assign w10053 = w9649 & ~w9667;
assign w10054 = w9626 & ~w9639;
assign w10055 = w9651 & w10054;
assign w10056 = w10012 & ~w10021;
assign w10057 = w10024 & ~w10053;
assign w10058 = ~w10055 & w10057;
assign w10059 = ~w10056 & w10058;
assign w10060 = ~w10052 & ~w10059;
assign w10061 = ~w10025 & ~w10045;
assign w10062 = ~w9647 & ~w10061;
assign w10063 = ~w10043 & ~w10062;
assign w10064 = ~w10060 & w10063;
assign w10065 = pi0570 & ~w10064;
assign w10066 = ~pi0570 & w10064;
assign w10067 = ~w10065 & ~w10066;
assign w10068 = ~w9742 & ~w9750;
assign w10069 = w9742 & w9750;
assign w10070 = w9702 & ~w9749;
assign w10071 = ~w10068 & ~w10070;
assign w10072 = ~w10069 & w10071;
assign w10073 = ~w9734 & ~w10072;
assign w10074 = w9721 & w63620;
assign w10075 = w9734 & ~w10074;
assign w10076 = ~w9815 & w9824;
assign w10077 = ~w9702 & ~w10076;
assign w10078 = ~w9760 & w10075;
assign w10079 = ~w10077 & w10078;
assign w10080 = ~w10073 & ~w10079;
assign w10081 = ~w9750 & w9775;
assign w10082 = w9737 & w9823;
assign w10083 = ~w9806 & ~w10069;
assign w10084 = ~w10081 & w10083;
assign w10085 = ~w9827 & ~w10082;
assign w10086 = w10084 & w10085;
assign w10087 = w9702 & ~w10086;
assign w10088 = ~w10080 & ~w10087;
assign w10089 = ~pi0550 & w10088;
assign w10090 = pi0550 & ~w10088;
assign w10091 = ~w10089 & ~w10090;
assign w10092 = ~w9365 & w9387;
assign w10093 = (w10092 & ~w9529) | (w10092 & w64909) | (~w9529 & w64909);
assign w10094 = w9373 & w9514;
assign w10095 = w9391 & ~w10094;
assign w10096 = ~w9342 & w9348;
assign w10097 = w9407 & w10096;
assign w10098 = ~w9374 & w64910;
assign w10099 = w9382 & ~w9414;
assign w10100 = ~w10097 & w10099;
assign w10101 = ~w10098 & w10100;
assign w10102 = w9514 & w64911;
assign w10103 = ~w9374 & w64912;
assign w10104 = ~w10102 & w10103;
assign w10105 = ~w10101 & ~w10104;
assign w10106 = ~w10093 & ~w10095;
assign w10107 = ~w10105 & w10106;
assign w10108 = pi0552 & w10107;
assign w10109 = ~pi0552 & ~w10107;
assign w10110 = ~w10108 & ~w10109;
assign w10111 = w9280 & w9302;
assign w10112 = ~w9279 & ~w10111;
assign w10113 = ~w9256 & ~w9549;
assign w10114 = w9555 & w10113;
assign w10115 = ~w9556 & ~w10114;
assign w10116 = (w10112 & w10115) | (w10112 & w64913) | (w10115 & w64913);
assign w10117 = ~w9250 & ~w10116;
assign w10118 = ~w9294 & w9301;
assign w10119 = ~w9262 & w9554;
assign w10120 = (w9250 & ~w9263) | (w9250 & w64914) | (~w9263 & w64914);
assign w10121 = ~w10119 & w10120;
assign w10122 = ~w10118 & ~w10121;
assign w10123 = ~w9308 & w9552;
assign w10124 = w10112 & w10123;
assign w10125 = (w9292 & ~w10124) | (w9292 & w64915) | (~w10124 & w64915);
assign w10126 = ~w9250 & ~w9281;
assign w10127 = w9562 & ~w10126;
assign w10128 = w10116 & w10127;
assign w10129 = ~w10117 & ~w10125;
assign w10130 = ~w10128 & w10129;
assign w10131 = pi0564 & ~w10130;
assign w10132 = ~pi0564 & w10130;
assign w10133 = ~w10131 & ~w10132;
assign w10134 = ~w9863 & ~w9880;
assign w10135 = w9848 & w9879;
assign w10136 = w9863 & ~w10135;
assign w10137 = w9878 & w9892;
assign w10138 = ~w9841 & w10137;
assign w10139 = w10136 & ~w10138;
assign w10140 = ~w10134 & ~w10139;
assign w10141 = w9891 & w9892;
assign w10142 = ~w9841 & ~w9856;
assign w10143 = (~w10142 & w9894) | (~w10142 & w63621) | (w9894 & w63621);
assign w10144 = ~w9857 & w10143;
assign w10145 = w9863 & w10144;
assign w10146 = (~w9863 & ~w9892) | (~w9863 & w64916) | (~w9892 & w64916);
assign w10147 = (~w10141 & w10143) | (~w10141 & w64917) | (w10143 & w64917);
assign w10148 = (~w9870 & w10145) | (~w9870 & w64918) | (w10145 & w64918);
assign w10149 = ~w9888 & ~w10137;
assign w10150 = ~w9863 & ~w10149;
assign w10151 = w9841 & w9878;
assign w10152 = ~w9893 & w10151;
assign w10153 = w9847 & w10152;
assign w10154 = w9841 & w9895;
assign w10155 = w9892 & ~w10154;
assign w10156 = ~w9878 & ~w10155;
assign w10157 = ~w10144 & w10156;
assign w10158 = ~w10150 & ~w10153;
assign w10159 = ~w10157 & w10158;
assign w10160 = w9870 & ~w10159;
assign w10161 = ~w10140 & ~w10148;
assign w10162 = ~w10160 & w10161;
assign w10163 = pi0568 & w10162;
assign w10164 = ~pi0568 & ~w10162;
assign w10165 = ~w10163 & ~w10164;
assign w10166 = w9848 & ~w9878;
assign w10167 = ~w9879 & ~w10166;
assign w10168 = w10136 & ~w10167;
assign w10169 = w9849 & w10168;
assign w10170 = ~w9911 & ~w10152;
assign w10171 = ~w9847 & ~w9863;
assign w10172 = w10151 & w10171;
assign w10173 = ~w9870 & ~w10172;
assign w10174 = ~w10170 & ~w10173;
assign w10175 = ~w9849 & ~w9892;
assign w10176 = w9886 & ~w10175;
assign w10177 = ~w9848 & ~w10142;
assign w10178 = w9907 & w10177;
assign w10179 = ~w10168 & ~w10178;
assign w10180 = ~w10176 & w10179;
assign w10181 = (~w10169 & w10180) | (~w10169 & w64919) | (w10180 & w64919);
assign w10182 = ~w10174 & w10181;
assign w10183 = pi0580 & ~w10182;
assign w10184 = ~pi0580 & w10182;
assign w10185 = ~w10183 & ~w10184;
assign w10186 = w9714 & w9754;
assign w10187 = ~w9728 & ~w9808;
assign w10188 = ~w9741 & ~w9762;
assign w10189 = w10187 & w63622;
assign w10190 = ~w9806 & ~w9811;
assign w10191 = ~w10186 & w10190;
assign w10192 = (w9702 & w10189) | (w9702 & w64920) | (w10189 & w64920);
assign w10193 = ~w9737 & ~w9819;
assign w10194 = ~w9816 & ~w10074;
assign w10195 = ~w10193 & w10194;
assign w10196 = ~w9744 & ~w10195;
assign w10197 = (~w9776 & ~w10187) | (~w9776 & w64921) | (~w10187 & w64921);
assign w10198 = ~w9721 & w9759;
assign w10199 = ~w10197 & ~w10198;
assign w10200 = ~w9702 & ~w10199;
assign w10201 = ~w9828 & ~w10196;
assign w10202 = ~w10192 & w10201;
assign w10203 = ~w10200 & w10202;
assign w10204 = pi0569 & w10203;
assign w10205 = ~pi0569 & ~w10203;
assign w10206 = ~w10204 & ~w10205;
assign w10207 = w9262 & w9283;
assign w10208 = w9309 & ~w10207;
assign w10209 = ~w10126 & ~w10208;
assign w10210 = w9250 & w9563;
assign w10211 = ~w9277 & w9302;
assign w10212 = ~w9294 & ~w10211;
assign w10213 = ~w9541 & ~w10212;
assign w10214 = w9292 & ~w10210;
assign w10215 = ~w10213 & w10214;
assign w10216 = ~w9306 & w9540;
assign w10217 = ~w9292 & ~w9315;
assign w10218 = ~w10119 & w10217;
assign w10219 = ~w9566 & w10218;
assign w10220 = ~w10216 & w10219;
assign w10221 = ~w10215 & ~w10220;
assign w10222 = ~w10209 & ~w10221;
assign w10223 = ~pi0589 & w10222;
assign w10224 = pi0589 & ~w10222;
assign w10225 = ~w10223 & ~w10224;
assign w10226 = (~w9957 & ~w9933) | (~w9957 & w64922) | (~w9933 & w64922);
assign w10227 = (w9995 & w9992) | (w9995 & w63623) | (w9992 & w63623);
assign w10228 = w9990 & ~w10226;
assign w10229 = ~w10227 & w10228;
assign w10230 = w9973 & w64923;
assign w10231 = ~w9926 & ~w9990;
assign w10232 = w9991 & ~w9996;
assign w10233 = ~w9992 & ~w10232;
assign w10234 = ~w10232 & w64924;
assign w10235 = ~w9949 & ~w9957;
assign w10236 = (w9926 & w10227) | (w9926 & w64925) | (w10227 & w64925);
assign w10237 = w9933 & w9946;
assign w10238 = w9957 & ~w10237;
assign w10239 = ~w9950 & ~w10238;
assign w10240 = w10236 & w10239;
assign w10241 = ~w9964 & ~w10230;
assign w10242 = ~w10235 & w10241;
assign w10243 = ~w10229 & w10242;
assign w10244 = ~w10234 & w10243;
assign w10245 = ~w10240 & w10244;
assign w10246 = w9932 & w9939;
assign w10247 = ~w9965 & ~w10246;
assign w10248 = w9957 & ~w10247;
assign w10249 = ~w9951 & w10236;
assign w10250 = w9964 & ~w10227;
assign w10251 = ~w10248 & w10250;
assign w10252 = ~w10249 & w10251;
assign w10253 = ~w10245 & w64926;
assign w10254 = (~pi0546 & w10245) | (~pi0546 & w64927) | (w10245 & w64927);
assign w10255 = ~w10253 & ~w10254;
assign w10256 = ~w10023 & ~w10045;
assign w10257 = w9647 & ~w10256;
assign w10258 = ~w9627 & ~w9647;
assign w10259 = ~w9684 & w10258;
assign w10260 = ~w9648 & ~w9682;
assign w10261 = w9647 & w10260;
assign w10262 = w9665 & ~w9676;
assign w10263 = ~w10259 & w10262;
assign w10264 = ~w10261 & w10263;
assign w10265 = ~w9665 & ~w10258;
assign w10266 = ~w9669 & w10044;
assign w10267 = ~w10265 & w10266;
assign w10268 = w10258 & ~w10260;
assign w10269 = ~w9655 & ~w10014;
assign w10270 = ~w10036 & w10269;
assign w10271 = ~w10268 & w10270;
assign w10272 = ~w9665 & ~w10271;
assign w10273 = ~w10264 & ~w10267;
assign w10274 = ~w10257 & w10273;
assign w10275 = ~w10272 & w10274;
assign w10276 = pi0578 & ~w10275;
assign w10277 = ~pi0578 & w10275;
assign w10278 = ~w10276 & ~w10277;
assign w10279 = w9850 & ~w10153;
assign w10280 = (w9870 & w10153) | (w9870 & w64928) | (w10153 & w64928);
assign w10281 = w10137 & w10280;
assign w10282 = ~w9892 & w10280;
assign w10283 = w9849 & w9878;
assign w10284 = ~w10141 & ~w10283;
assign w10285 = ~w10282 & w10284;
assign w10286 = w9863 & ~w10285;
assign w10287 = ~w9891 & ~w10151;
assign w10288 = w9894 & ~w10154;
assign w10289 = w10287 & w10288;
assign w10290 = ~w9896 & ~w10287;
assign w10291 = ~w9870 & ~w10289;
assign w10292 = ~w10290 & w10291;
assign w10293 = w9902 & w10175;
assign w10294 = w10279 & w10293;
assign w10295 = ~w10281 & ~w10294;
assign w10296 = ~w10292 & w10295;
assign w10297 = ~w10286 & w10296;
assign w10298 = pi0573 & ~w10297;
assign w10299 = ~pi0573 & w10297;
assign w10300 = ~w10298 & ~w10299;
assign w10301 = ~w9467 & ~w9486;
assign w10302 = ~w9494 & w10301;
assign w10303 = w9457 & ~w10302;
assign w10304 = ~w9440 & ~w9464;
assign w10305 = w9458 & w10304;
assign w10306 = ~w10303 & ~w10305;
assign w10307 = ~w9428 & ~w10306;
assign w10308 = ~w9434 & w9457;
assign w10309 = ~w9475 & ~w9480;
assign w10310 = w9428 & w10304;
assign w10311 = w10309 & ~w10310;
assign w10312 = w10308 & ~w10311;
assign w10313 = ~w9440 & ~w10308;
assign w10314 = w9491 & w10313;
assign w10315 = (w9440 & w9499) | (w9440 & w64929) | (w9499 & w64929);
assign w10316 = ~w10314 & ~w10315;
assign w10317 = w9428 & ~w10316;
assign w10318 = w9473 & ~w9485;
assign w10319 = w9450 & ~w9464;
assign w10320 = w9428 & ~w9447;
assign w10321 = w9441 & ~w10320;
assign w10322 = ~w10318 & ~w10321;
assign w10323 = ~w10319 & w10322;
assign w10324 = ~w9457 & ~w10323;
assign w10325 = ~w10312 & ~w10317;
assign w10326 = ~w10324 & w10325;
assign w10327 = ~w10307 & w10326;
assign w10328 = ~pi0571 & ~w10327;
assign w10329 = pi0571 & w10327;
assign w10330 = ~w10328 & ~w10329;
assign w10331 = w9479 & w9506;
assign w10332 = ~w9450 & ~w10331;
assign w10333 = ~w10313 & ~w10332;
assign w10334 = ~w9448 & ~w9487;
assign w10335 = w9457 & ~w10334;
assign w10336 = ~w9486 & ~w9506;
assign w10337 = w9479 & ~w10336;
assign w10338 = ~w9465 & ~w9491;
assign w10339 = ~w9434 & ~w9457;
assign w10340 = ~w10338 & w10339;
assign w10341 = ~w10337 & ~w10340;
assign w10342 = ~w9428 & ~w9474;
assign w10343 = ~w9496 & w10342;
assign w10344 = ~w10319 & w10343;
assign w10345 = ~w10335 & w10341;
assign w10346 = w10344 & w10345;
assign w10347 = w9485 & ~w9498;
assign w10348 = (w9457 & ~w9485) | (w9457 & w64930) | (~w9485 & w64930);
assign w10349 = ~w10304 & ~w10315;
assign w10350 = w10348 & w10349;
assign w10351 = w9506 & w10347;
assign w10352 = (w9428 & w9488) | (w9428 & w64931) | (w9488 & w64931);
assign w10353 = ~w10351 & w10352;
assign w10354 = ~w10350 & w10353;
assign w10355 = ~w10346 & ~w10354;
assign w10356 = ~w10333 & ~w10355;
assign w10357 = ~pi0562 & w10356;
assign w10358 = pi0562 & ~w10356;
assign w10359 = ~w10357 & ~w10358;
assign w10360 = w10304 & w10348;
assign w10361 = ~w9434 & w9498;
assign w10362 = ~w9450 & ~w9487;
assign w10363 = ~w10361 & w10362;
assign w10364 = ~w9457 & ~w10363;
assign w10365 = w9470 & ~w10301;
assign w10366 = ~w9496 & w10309;
assign w10367 = ~w10365 & w10366;
assign w10368 = ~w10364 & w10367;
assign w10369 = w9428 & ~w10368;
assign w10370 = w9468 & ~w9491;
assign w10371 = w9482 & w10370;
assign w10372 = ~w9495 & ~w10338;
assign w10373 = w10363 & w10372;
assign w10374 = (~w9428 & w10373) | (~w9428 & w64932) | (w10373 & w64932);
assign w10375 = ~w9482 & ~w10341;
assign w10376 = ~w9507 & ~w10360;
assign w10377 = ~w10375 & w10376;
assign w10378 = ~w10374 & w10377;
assign w10379 = ~w10369 & w10378;
assign w10380 = pi0566 & w10379;
assign w10381 = ~pi0566 & ~w10379;
assign w10382 = ~w10380 & ~w10381;
assign w10383 = (w9926 & w9992) | (w9926 & w10230) | (w9992 & w10230);
assign w10384 = w9984 & w10231;
assign w10385 = w9957 & ~w10384;
assign w10386 = ~w10383 & w10385;
assign w10387 = ~w9965 & w10386;
assign w10388 = ~w9957 & w10384;
assign w10389 = ~w10237 & ~w10388;
assign w10390 = (~w9964 & w10387) | (~w9964 & w64933) | (w10387 & w64933);
assign w10391 = ~w9957 & ~w10383;
assign w10392 = ~w10238 & ~w10391;
assign w10393 = ~w9968 & ~w9992;
assign w10394 = (w9964 & ~w10393) | (w9964 & w64934) | (~w10393 & w64934);
assign w10395 = ~w10386 & w10394;
assign w10396 = ~w10392 & ~w10395;
assign w10397 = ~w10390 & w10396;
assign w10398 = pi0560 & w10397;
assign w10399 = ~pi0560 & ~w10397;
assign w10400 = ~w10398 & ~w10399;
assign w10401 = ~w9966 & ~w9984;
assign w10402 = ~w9926 & w9948;
assign w10403 = ~w10401 & ~w10402;
assign w10404 = ~w10235 & ~w10403;
assign w10405 = w9926 & ~w9991;
assign w10406 = ~w9957 & ~w10405;
assign w10407 = w10233 & w10406;
assign w10408 = w9957 & ~w9974;
assign w10409 = ~w9970 & w10226;
assign w10410 = ~w10408 & ~w10409;
assign w10411 = ~w10235 & ~w10246;
assign w10412 = ~w10407 & w63369;
assign w10413 = ~w9926 & w9983;
assign w10414 = ~w9993 & ~w10413;
assign w10415 = w9957 & ~w10414;
assign w10416 = ~w9950 & ~w10415;
assign w10417 = (~w9964 & w10412) | (~w9964 & w63625) | (w10412 & w63625);
assign w10418 = (~w10407 & w64935) | (~w10407 & w64936) | (w64935 & w64936);
assign w10419 = ~w10417 & w64937;
assign w10420 = (pi0567 & w10417) | (pi0567 & w64938) | (w10417 & w64938);
assign w10421 = ~w10419 & ~w10420;
assign w10422 = ~pi3526 & pi9040;
assign w10423 = ~pi3532 & ~pi9040;
assign w10424 = ~w10422 & ~w10423;
assign w10425 = pi0581 & ~w10424;
assign w10426 = ~pi0581 & w10424;
assign w10427 = ~w10425 & ~w10426;
assign w10428 = ~pi3501 & pi9040;
assign w10429 = ~pi3519 & ~pi9040;
assign w10430 = ~w10428 & ~w10429;
assign w10431 = pi0604 & ~w10430;
assign w10432 = ~pi0604 & w10430;
assign w10433 = ~w10431 & ~w10432;
assign w10434 = ~pi3536 & pi9040;
assign w10435 = ~pi3531 & ~pi9040;
assign w10436 = ~w10434 & ~w10435;
assign w10437 = pi0572 & ~w10436;
assign w10438 = ~pi0572 & w10436;
assign w10439 = ~w10437 & ~w10438;
assign w10440 = w10433 & ~w10439;
assign w10441 = ~pi3521 & pi9040;
assign w10442 = ~pi3523 & ~pi9040;
assign w10443 = ~w10441 & ~w10442;
assign w10444 = pi0584 & ~w10443;
assign w10445 = ~pi0584 & w10443;
assign w10446 = ~w10444 & ~w10445;
assign w10447 = w10440 & ~w10446;
assign w10448 = ~pi3529 & pi9040;
assign w10449 = ~pi3488 & ~pi9040;
assign w10450 = ~w10448 & ~w10449;
assign w10451 = pi0607 & ~w10450;
assign w10452 = ~pi0607 & w10450;
assign w10453 = ~w10451 & ~w10452;
assign w10454 = w10440 & w63626;
assign w10455 = ~w10433 & w10439;
assign w10456 = w10446 & ~w10453;
assign w10457 = ~w10455 & ~w10456;
assign w10458 = w10439 & w10453;
assign w10459 = ~w10433 & w10446;
assign w10460 = w10458 & ~w10459;
assign w10461 = ~w10440 & ~w10460;
assign w10462 = ~w10457 & ~w10461;
assign w10463 = ~w10439 & ~w10453;
assign w10464 = ~w10433 & ~w10446;
assign w10465 = w10463 & w10464;
assign w10466 = ~w10454 & ~w10465;
assign w10467 = ~w10462 & w10466;
assign w10468 = w10427 & ~w10467;
assign w10469 = w10446 & ~w10455;
assign w10470 = ~w10427 & ~w10469;
assign w10471 = ~w10458 & ~w10463;
assign w10472 = ~w10433 & w10453;
assign w10473 = w10446 & ~w10472;
assign w10474 = w10471 & w10473;
assign w10475 = w10470 & w10474;
assign w10476 = w10446 & w10453;
assign w10477 = ~w10446 & ~w10453;
assign w10478 = ~w10476 & ~w10477;
assign w10479 = ~w10439 & ~w10478;
assign w10480 = ~w10427 & w10479;
assign w10481 = ~w10453 & w10455;
assign w10482 = (w10427 & ~w10455) | (w10427 & w64939) | (~w10455 & w64939);
assign w10483 = w10427 & ~w10459;
assign w10484 = ~w10482 & ~w10483;
assign w10485 = ~w10457 & ~w10484;
assign w10486 = ~w10446 & w10458;
assign w10487 = w10433 & w10486;
assign w10488 = ~pi3499 & pi9040;
assign w10489 = ~pi3515 & ~pi9040;
assign w10490 = ~w10488 & ~w10489;
assign w10491 = pi0599 & ~w10490;
assign w10492 = ~pi0599 & w10490;
assign w10493 = ~w10491 & ~w10492;
assign w10494 = ~w10487 & w10493;
assign w10495 = ~w10480 & w10494;
assign w10496 = ~w10485 & w10495;
assign w10497 = w10456 & ~w10482;
assign w10498 = w10433 & w10439;
assign w10499 = ~w10427 & ~w10498;
assign w10500 = w10453 & w10464;
assign w10501 = w10499 & ~w10500;
assign w10502 = ~w10439 & w10446;
assign w10503 = w10472 & w10502;
assign w10504 = (w10427 & ~w10440) | (w10427 & w11131) | (~w10440 & w11131);
assign w10505 = ~w10503 & w10504;
assign w10506 = ~w10501 & ~w10505;
assign w10507 = w10476 & w10498;
assign w10508 = ~w10493 & ~w10507;
assign w10509 = ~w10497 & w10508;
assign w10510 = ~w10506 & w10509;
assign w10511 = ~w10496 & ~w10510;
assign w10512 = ~w10468 & ~w10475;
assign w10513 = ~w10511 & w10512;
assign w10514 = pi0608 & w10513;
assign w10515 = ~pi0608 & ~w10513;
assign w10516 = ~w10514 & ~w10515;
assign w10517 = ~pi3498 & pi9040;
assign w10518 = ~pi3514 & ~pi9040;
assign w10519 = ~w10517 & ~w10518;
assign w10520 = pi0592 & ~w10519;
assign w10521 = ~pi0592 & w10519;
assign w10522 = ~w10520 & ~w10521;
assign w10523 = ~pi3527 & pi9040;
assign w10524 = ~pi3491 & ~pi9040;
assign w10525 = ~w10523 & ~w10524;
assign w10526 = pi0591 & ~w10525;
assign w10527 = ~pi0591 & w10525;
assign w10528 = ~w10526 & ~w10527;
assign w10529 = ~pi3528 & pi9040;
assign w10530 = ~pi3492 & ~pi9040;
assign w10531 = ~w10529 & ~w10530;
assign w10532 = pi0558 & ~w10531;
assign w10533 = ~pi0558 & w10531;
assign w10534 = ~w10532 & ~w10533;
assign w10535 = ~w10528 & ~w10534;
assign w10536 = ~pi3494 & pi9040;
assign w10537 = ~pi3525 & ~pi9040;
assign w10538 = ~w10536 & ~w10537;
assign w10539 = pi0599 & ~w10538;
assign w10540 = ~pi0599 & w10538;
assign w10541 = ~w10539 & ~w10540;
assign w10542 = ~pi3495 & pi9040;
assign w10543 = ~pi3507 & ~pi9040;
assign w10544 = ~w10542 & ~w10543;
assign w10545 = pi0595 & ~w10544;
assign w10546 = ~pi0595 & w10544;
assign w10547 = ~w10545 & ~w10546;
assign w10548 = w10541 & ~w10547;
assign w10549 = ~w10535 & ~w10548;
assign w10550 = w10534 & w10541;
assign w10551 = ~w10534 & ~w10541;
assign w10552 = ~w10550 & ~w10551;
assign w10553 = ~pi3562 & pi9040;
assign w10554 = ~pi3504 & ~pi9040;
assign w10555 = ~w10553 & ~w10554;
assign w10556 = pi0604 & ~w10555;
assign w10557 = ~pi0604 & w10555;
assign w10558 = ~w10556 & ~w10557;
assign w10559 = w10552 & w10558;
assign w10560 = ~w10552 & ~w10558;
assign w10561 = ~w10559 & ~w10560;
assign w10562 = w10528 & w10552;
assign w10563 = (w10541 & ~w10552) | (w10541 & w63627) | (~w10552 & w63627);
assign w10564 = w10561 & w63628;
assign w10565 = ~w10528 & ~w10547;
assign w10566 = w10534 & ~w10558;
assign w10567 = ~w10541 & w10565;
assign w10568 = ~w10566 & w10567;
assign w10569 = ~w10541 & ~w10558;
assign w10570 = ~w10535 & w10569;
assign w10571 = w10548 & w10558;
assign w10572 = ~w10570 & ~w10571;
assign w10573 = ~w10528 & w10550;
assign w10574 = ~w10534 & w10558;
assign w10575 = ~w10566 & ~w10574;
assign w10576 = w10562 & ~w10575;
assign w10577 = (~w10573 & ~w10562) | (~w10573 & w63370) | (~w10562 & w63370);
assign w10578 = w10572 & ~w10577;
assign w10579 = ~w10528 & ~w10558;
assign w10580 = ~w10541 & w10547;
assign w10581 = ~w10579 & w10580;
assign w10582 = w10575 & w10581;
assign w10583 = w10562 & w10582;
assign w10584 = ~w10568 & ~w10583;
assign w10585 = ~w10564 & w10584;
assign w10586 = (~w10522 & ~w10585) | (~w10522 & w64940) | (~w10585 & w64940);
assign w10587 = w10541 & w10558;
assign w10588 = ~w10547 & ~w10587;
assign w10589 = ~w10573 & ~w10588;
assign w10590 = w10575 & ~w10589;
assign w10591 = ~w10552 & w63629;
assign w10592 = ~w10590 & ~w10591;
assign w10593 = ~w10547 & ~w10579;
assign w10594 = w10528 & w10574;
assign w10595 = w10593 & ~w10594;
assign w10596 = ~w10590 & w64941;
assign w10597 = ~w10551 & ~w10566;
assign w10598 = ~w10535 & w10547;
assign w10599 = ~w10597 & w10598;
assign w10600 = w10535 & w10587;
assign w10601 = w10565 & w10569;
assign w10602 = ~w10600 & ~w10601;
assign w10603 = ~w10528 & w10552;
assign w10604 = ~w10593 & w10603;
assign w10605 = w10602 & w10604;
assign w10606 = w10572 & ~w10599;
assign w10607 = (w10522 & w10605) | (w10522 & w64942) | (w10605 & w64942);
assign w10608 = ~w10534 & w10582;
assign w10609 = w10541 & w10547;
assign w10610 = w10579 & w10609;
assign w10611 = ~w10608 & ~w10610;
assign w10612 = ~w10596 & w10611;
assign w10613 = ~w10607 & w10612;
assign w10614 = ~w10586 & w10613;
assign w10615 = ~pi0616 & w10614;
assign w10616 = pi0616 & ~w10614;
assign w10617 = ~w10615 & ~w10616;
assign w10618 = ~pi3500 & pi9040;
assign w10619 = ~pi3537 & ~pi9040;
assign w10620 = ~w10618 & ~w10619;
assign w10621 = pi0601 & ~w10620;
assign w10622 = ~pi0601 & w10620;
assign w10623 = ~w10621 & ~w10622;
assign w10624 = ~pi3518 & pi9040;
assign w10625 = ~pi3534 & ~pi9040;
assign w10626 = ~w10624 & ~w10625;
assign w10627 = pi0586 & ~w10626;
assign w10628 = ~pi0586 & w10626;
assign w10629 = ~w10627 & ~w10628;
assign w10630 = ~w10623 & w10629;
assign w10631 = w10623 & ~w10629;
assign w10632 = ~w10630 & ~w10631;
assign w10633 = ~pi3515 & pi9040;
assign w10634 = ~pi3520 & ~pi9040;
assign w10635 = ~w10633 & ~w10634;
assign w10636 = pi0594 & ~w10635;
assign w10637 = ~pi0594 & w10635;
assign w10638 = ~w10636 & ~w10637;
assign w10639 = ~pi3488 & pi9040;
assign w10640 = ~pi3538 & ~pi9040;
assign w10641 = ~w10639 & ~w10640;
assign w10642 = pi0585 & ~w10641;
assign w10643 = ~pi0585 & w10641;
assign w10644 = ~w10642 & ~w10643;
assign w10645 = ~w10638 & w10644;
assign w10646 = w10632 & w10645;
assign w10647 = w10623 & w10644;
assign w10648 = w10638 & ~w10647;
assign w10649 = ~pi3497 & pi9040;
assign w10650 = ~pi3517 & ~pi9040;
assign w10651 = ~w10649 & ~w10650;
assign w10652 = pi0572 & ~w10651;
assign w10653 = ~pi0572 & w10651;
assign w10654 = ~w10652 & ~w10653;
assign w10655 = w10644 & w10654;
assign w10656 = ~w10644 & ~w10654;
assign w10657 = ~w10655 & ~w10656;
assign w10658 = w10630 & w10657;
assign w10659 = ~w10630 & w10656;
assign w10660 = ~w10658 & ~w10659;
assign w10661 = w10648 & ~w10660;
assign w10662 = ~w10629 & w10654;
assign w10663 = ~w10638 & w10662;
assign w10664 = ~w10655 & ~w10663;
assign w10665 = ~pi3524 & pi9040;
assign w10666 = pi3535 & ~pi9040;
assign w10667 = ~w10665 & ~w10666;
assign w10668 = pi0584 & ~w10667;
assign w10669 = ~pi0584 & w10667;
assign w10670 = ~w10668 & ~w10669;
assign w10671 = ~w10648 & ~w10656;
assign w10672 = w10631 & ~w10671;
assign w10673 = ~w10623 & ~w10654;
assign w10674 = w10623 & w10654;
assign w10675 = ~w10673 & ~w10674;
assign w10676 = ~w10629 & ~w10675;
assign w10677 = (~w10638 & ~w10630) | (~w10638 & w64943) | (~w10630 & w64943);
assign w10678 = ~w10676 & w64944;
assign w10679 = w10660 & w10678;
assign w10680 = (w10670 & w10664) | (w10670 & w64945) | (w10664 & w64945);
assign w10681 = ~w10672 & w10680;
assign w10682 = ~w10679 & w10681;
assign w10683 = ~w10623 & ~w10644;
assign w10684 = ~w10647 & ~w10683;
assign w10685 = ~w10638 & w10684;
assign w10686 = ~w10664 & w10685;
assign w10687 = w10623 & ~w10644;
assign w10688 = w10629 & w10687;
assign w10689 = w10647 & w10662;
assign w10690 = ~w10688 & ~w10689;
assign w10691 = w10638 & ~w10690;
assign w10692 = w10629 & ~w10654;
assign w10693 = ~w10662 & ~w10692;
assign w10694 = w10683 & w10693;
assign w10695 = ~w10670 & ~w10694;
assign w10696 = ~w10686 & w10695;
assign w10697 = ~w10691 & w10696;
assign w10698 = ~w10682 & ~w10697;
assign w10699 = ~w10646 & ~w10661;
assign w10700 = ~w10698 & w10699;
assign w10701 = pi0624 & ~w10700;
assign w10702 = ~pi0624 & w10700;
assign w10703 = ~w10701 & ~w10702;
assign w10704 = ~w10541 & w10558;
assign w10705 = (w10704 & w10605) | (w10704 & w64946) | (w10605 & w64946);
assign w10706 = w10575 & w10609;
assign w10707 = ~w10552 & w10588;
assign w10708 = ~w10594 & w10707;
assign w10709 = ~w10576 & ~w10706;
assign w10710 = ~w10708 & w10709;
assign w10711 = ~w10522 & ~w10710;
assign w10712 = w10534 & w10610;
assign w10713 = w10528 & w10548;
assign w10714 = w10528 & w10534;
assign w10715 = w10558 & w10714;
assign w10716 = ~w10581 & ~w10715;
assign w10717 = w10602 & ~w10713;
assign w10718 = ~w10712 & w10716;
assign w10719 = w10717 & w10718;
assign w10720 = w10522 & ~w10719;
assign w10721 = ~w10705 & ~w10720;
assign w10722 = ~w10711 & w10721;
assign w10723 = pi0617 & w10722;
assign w10724 = ~pi0617 & ~w10722;
assign w10725 = ~w10723 & ~w10724;
assign w10726 = (~w10719 & w63371) | (~w10719 & w63372) | (w63371 & w63372);
assign w10727 = (~w10571 & w10719) | (~w10571 & w63373) | (w10719 & w63373);
assign w10728 = ~w10726 & w10727;
assign w10729 = w10561 & w64947;
assign w10730 = (~w10581 & w10577) | (~w10581 & w63630) | (w10577 & w63630);
assign w10731 = ~w10561 & ~w10730;
assign w10732 = (w10522 & w10731) | (w10522 & w64948) | (w10731 & w64948);
assign w10733 = ~w10572 & ~w10602;
assign w10734 = ~w10549 & ~w10716;
assign w10735 = ~w10610 & ~w10733;
assign w10736 = ~w10734 & w10735;
assign w10737 = (w10736 & w10728) | (w10736 & w63631) | (w10728 & w63631);
assign w10738 = w10737 & w64949;
assign w10739 = (pi0629 & ~w10737) | (pi0629 & w64950) | (~w10737 & w64950);
assign w10740 = ~w10738 & ~w10739;
assign w10741 = ~pi3504 & pi9040;
assign w10742 = ~pi3567 & ~pi9040;
assign w10743 = ~w10741 & ~w10742;
assign w10744 = pi0582 & ~w10743;
assign w10745 = ~pi0582 & w10743;
assign w10746 = ~w10744 & ~w10745;
assign w10747 = ~pi3559 & pi9040;
assign w10748 = ~pi3487 & ~pi9040;
assign w10749 = ~w10747 & ~w10748;
assign w10750 = pi0605 & ~w10749;
assign w10751 = ~pi0605 & w10749;
assign w10752 = ~w10750 & ~w10751;
assign w10753 = ~w10746 & w10752;
assign w10754 = ~pi3489 & pi9040;
assign w10755 = ~pi3498 & ~pi9040;
assign w10756 = ~w10754 & ~w10755;
assign w10757 = pi0583 & ~w10756;
assign w10758 = ~pi0583 & w10756;
assign w10759 = ~w10757 & ~w10758;
assign w10760 = w10752 & w10759;
assign w10761 = ~w10746 & ~w10759;
assign w10762 = ~w10760 & ~w10761;
assign w10763 = ~pi3485 & pi9040;
assign w10764 = ~pi3493 & ~pi9040;
assign w10765 = ~w10763 & ~w10764;
assign w10766 = pi0598 & ~w10765;
assign w10767 = ~pi0598 & w10765;
assign w10768 = ~w10766 & ~w10767;
assign w10769 = (w10768 & w10762) | (w10768 & w64951) | (w10762 & w64951);
assign w10770 = ~w10752 & w10759;
assign w10771 = ~pi3483 & pi9040;
assign w10772 = ~pi3503 & ~pi9040;
assign w10773 = ~w10771 & ~w10772;
assign w10774 = pi0579 & ~w10773;
assign w10775 = ~pi0579 & w10773;
assign w10776 = ~w10774 & ~w10775;
assign w10777 = w10746 & ~w10776;
assign w10778 = w10770 & w10777;
assign w10779 = w10753 & w10759;
assign w10780 = w10753 & w64952;
assign w10781 = ~w10778 & ~w10780;
assign w10782 = w10769 & ~w10781;
assign w10783 = ~pi3525 & pi9040;
assign w10784 = ~pi3513 & ~pi9040;
assign w10785 = ~w10783 & ~w10784;
assign w10786 = pi0606 & ~w10785;
assign w10787 = ~pi0606 & w10785;
assign w10788 = ~w10786 & ~w10787;
assign w10789 = ~w10782 & w10788;
assign w10790 = w10746 & ~w10752;
assign w10791 = ~w10753 & ~w10790;
assign w10792 = ~w10761 & ~w10776;
assign w10793 = ~w10791 & w10792;
assign w10794 = w10752 & w10768;
assign w10795 = w10752 & ~w10776;
assign w10796 = ~w10779 & ~w10795;
assign w10797 = w10794 & w10796;
assign w10798 = ~w10752 & ~w10768;
assign w10799 = ~w10746 & w10776;
assign w10800 = w10759 & ~w10799;
assign w10801 = w10798 & ~w10800;
assign w10802 = w10746 & ~w10759;
assign w10803 = w10794 & w10802;
assign w10804 = ~w10793 & ~w10803;
assign w10805 = ~w10801 & w10804;
assign w10806 = ~w10797 & w10805;
assign w10807 = ~w10789 & ~w10806;
assign w10808 = ~w10746 & ~w10768;
assign w10809 = ~w10790 & ~w10808;
assign w10810 = w10762 & w10809;
assign w10811 = (w10776 & w10810) | (w10776 & w64953) | (w10810 & w64953);
assign w10812 = ~w10777 & ~w10799;
assign w10813 = w10759 & ~w10768;
assign w10814 = ~w10795 & w10813;
assign w10815 = w10812 & w10814;
assign w10816 = ~w10811 & ~w10815;
assign w10817 = w10788 & ~w10816;
assign w10818 = w10752 & w10776;
assign w10819 = w10776 & w10802;
assign w10820 = ~w10768 & ~w10770;
assign w10821 = ~w10819 & w10820;
assign w10822 = w10760 & w10812;
assign w10823 = w10795 & w10802;
assign w10824 = ~w10822 & ~w10823;
assign w10825 = w10821 & w10824;
assign w10826 = w10761 & w10788;
assign w10827 = ~w10825 & ~w10826;
assign w10828 = w10761 & w10798;
assign w10829 = ~w10818 & ~w10828;
assign w10830 = ~w10827 & w10829;
assign w10831 = ~w10807 & ~w10817;
assign w10832 = (pi0621 & ~w10831) | (pi0621 & w64954) | (~w10831 & w64954);
assign w10833 = w10831 & w64955;
assign w10834 = ~w10832 & ~w10833;
assign w10835 = ~pi3567 & pi9040;
assign w10836 = ~pi3494 & ~pi9040;
assign w10837 = ~w10835 & ~w10836;
assign w10838 = pi0600 & ~w10837;
assign w10839 = ~pi0600 & w10837;
assign w10840 = ~w10838 & ~w10839;
assign w10841 = ~pi3514 & pi9040;
assign w10842 = ~pi3483 & ~pi9040;
assign w10843 = ~w10841 & ~w10842;
assign w10844 = pi0558 & ~w10843;
assign w10845 = ~pi0558 & w10843;
assign w10846 = ~w10844 & ~w10845;
assign w10847 = w10840 & ~w10846;
assign w10848 = ~pi3506 & pi9040;
assign w10849 = ~pi3489 & ~pi9040;
assign w10850 = ~w10848 & ~w10849;
assign w10851 = pi0592 & ~w10850;
assign w10852 = ~pi0592 & w10850;
assign w10853 = ~w10851 & ~w10852;
assign w10854 = ~pi3491 & pi9040;
assign w10855 = ~pi3580 & ~pi9040;
assign w10856 = ~w10854 & ~w10855;
assign w10857 = pi0602 & ~w10856;
assign w10858 = ~pi0602 & w10856;
assign w10859 = ~w10857 & ~w10858;
assign w10860 = ~w10853 & w10859;
assign w10861 = w10847 & w10860;
assign w10862 = ~pi3486 & pi9040;
assign w10863 = ~pi3485 & ~pi9040;
assign w10864 = ~w10862 & ~w10863;
assign w10865 = pi0575 & ~w10864;
assign w10866 = ~pi0575 & w10864;
assign w10867 = ~w10865 & ~w10866;
assign w10868 = ~w10846 & ~w10859;
assign w10869 = w10840 & ~w10868;
assign w10870 = w10853 & ~w10869;
assign w10871 = ~w10853 & ~w10859;
assign w10872 = w10846 & w10871;
assign w10873 = ~w10870 & ~w10872;
assign w10874 = w10853 & w10859;
assign w10875 = w10871 & w64956;
assign w10876 = ~pi3487 & pi9040;
assign w10877 = ~pi3528 & ~pi9040;
assign w10878 = ~w10876 & ~w10877;
assign w10879 = pi0588 & ~w10878;
assign w10880 = ~pi0588 & w10878;
assign w10881 = ~w10879 & ~w10880;
assign w10882 = (w10881 & ~w10874) | (w10881 & w64957) | (~w10874 & w64957);
assign w10883 = ~w10875 & w10882;
assign w10884 = ~w10873 & w10883;
assign w10885 = w10840 & ~w10859;
assign w10886 = ~w10846 & w10859;
assign w10887 = ~w10853 & ~w10885;
assign w10888 = ~w10886 & w10887;
assign w10889 = ~w10881 & w10888;
assign w10890 = ~w10840 & ~w10846;
assign w10891 = w10846 & w10881;
assign w10892 = ~w10890 & ~w10891;
assign w10893 = w10874 & ~w10892;
assign w10894 = ~w10861 & w10867;
assign w10895 = ~w10893 & w10894;
assign w10896 = ~w10889 & w10895;
assign w10897 = ~w10884 & w10896;
assign w10898 = w10846 & w10853;
assign w10899 = w10885 & w10898;
assign w10900 = ~w10867 & ~w10899;
assign w10901 = w10881 & w10888;
assign w10902 = ~w10871 & ~w10874;
assign w10903 = w10847 & ~w10902;
assign w10904 = w10900 & ~w10903;
assign w10905 = ~w10901 & w10904;
assign w10906 = ~w10897 & ~w10905;
assign w10907 = w10890 & w10902;
assign w10908 = ~w10898 & ~w10907;
assign w10909 = ~w10867 & ~w10908;
assign w10910 = ~w10846 & ~w10853;
assign w10911 = w10840 & w10910;
assign w10912 = ~w10899 & ~w10911;
assign w10913 = ~w10909 & w10912;
assign w10914 = ~w10881 & ~w10913;
assign w10915 = ~w10906 & ~w10914;
assign w10916 = ~pi0610 & w10915;
assign w10917 = pi0610 & ~w10915;
assign w10918 = ~w10916 & ~w10917;
assign w10919 = ~w10759 & ~w10776;
assign w10920 = w10791 & w10919;
assign w10921 = w10802 & w63632;
assign w10922 = w10768 & ~w10921;
assign w10923 = ~w10920 & w10922;
assign w10924 = ~w10768 & ~w10780;
assign w10925 = ~w10923 & ~w10924;
assign w10926 = ~w10768 & ~w10776;
assign w10927 = ~w10791 & w10926;
assign w10928 = w10791 & w63633;
assign w10929 = w10820 & w10928;
assign w10930 = (~w10752 & w10929) | (~w10752 & w64958) | (w10929 & w64958);
assign w10931 = w10788 & ~w10803;
assign w10932 = ~w10822 & w10931;
assign w10933 = ~w10927 & w10932;
assign w10934 = ~w10930 & w10933;
assign w10935 = ~w10769 & ~w10821;
assign w10936 = w10794 & w10799;
assign w10937 = ~w10746 & w10919;
assign w10938 = w10919 & w64959;
assign w10939 = w10761 & w10818;
assign w10940 = ~w10938 & ~w10939;
assign w10941 = ~w10778 & ~w10788;
assign w10942 = ~w10936 & w10941;
assign w10943 = w10940 & w10942;
assign w10944 = ~w10935 & w10943;
assign w10945 = ~w10934 & ~w10944;
assign w10946 = ~w10925 & ~w10945;
assign w10947 = ~pi0618 & w10946;
assign w10948 = pi0618 & ~w10946;
assign w10949 = ~w10947 & ~w10948;
assign w10950 = ~pi3484 & pi9040;
assign w10951 = ~pi3529 & ~pi9040;
assign w10952 = ~w10950 & ~w10951;
assign w10953 = pi0576 & ~w10952;
assign w10954 = ~pi0576 & w10952;
assign w10955 = ~w10953 & ~w10954;
assign w10956 = ~pi3539 & pi9040;
assign w10957 = ~pi3518 & ~pi9040;
assign w10958 = ~w10956 & ~w10957;
assign w10959 = pi0590 & ~w10958;
assign w10960 = ~pi0590 & w10958;
assign w10961 = ~w10959 & ~w10960;
assign w10962 = ~w10955 & w10961;
assign w10963 = ~pi3523 & pi9040;
assign w10964 = ~pi3500 & ~pi9040;
assign w10965 = ~w10963 & ~w10964;
assign w10966 = pi0593 & ~w10965;
assign w10967 = ~pi0593 & w10965;
assign w10968 = ~w10966 & ~w10967;
assign w10969 = ~pi3538 & pi9040;
assign w10970 = ~pi3530 & ~pi9040;
assign w10971 = ~w10969 & ~w10970;
assign w10972 = pi0585 & ~w10971;
assign w10973 = ~pi0585 & w10971;
assign w10974 = ~w10972 & ~w10973;
assign w10975 = w10968 & w10974;
assign w10976 = w10962 & w10975;
assign w10977 = ~pi3533 & pi9040;
assign w10978 = ~pi3499 & ~pi9040;
assign w10979 = ~w10977 & ~w10978;
assign w10980 = pi0596 & ~w10979;
assign w10981 = ~pi0596 & w10979;
assign w10982 = ~w10980 & ~w10981;
assign w10983 = ~w10974 & w10982;
assign w10984 = ~w10961 & w10983;
assign w10985 = ~w10955 & w10984;
assign w10986 = ~w10974 & ~w10982;
assign w10987 = ~w10962 & w10986;
assign w10988 = w10955 & ~w10961;
assign w10989 = w10987 & ~w10988;
assign w10990 = w10961 & w10982;
assign w10991 = w10974 & w10990;
assign w10992 = ~w10984 & ~w10991;
assign w10993 = ~w10989 & w10992;
assign w10994 = w10968 & ~w10993;
assign w10995 = ~w10961 & ~w10982;
assign w10996 = w10955 & w10974;
assign w10997 = w10995 & w10996;
assign w10998 = w10961 & w10983;
assign w10999 = w10983 & w64960;
assign w11000 = ~w10983 & ~w10995;
assign w11001 = ~w10955 & w11000;
assign w11002 = ~w10999 & ~w11001;
assign w11003 = ~w10968 & ~w11002;
assign w11004 = ~pi3535 & pi9040;
assign w11005 = ~pi3501 & ~pi9040;
assign w11006 = ~w11004 & ~w11005;
assign w11007 = pi0601 & ~w11006;
assign w11008 = ~pi0601 & w11006;
assign w11009 = ~w11007 & ~w11008;
assign w11010 = ~w10997 & ~w11009;
assign w11011 = (w11010 & w10993) | (w11010 & w64961) | (w10993 & w64961);
assign w11012 = ~w11003 & w11011;
assign w11013 = ~w10955 & ~w10974;
assign w11014 = ~w10968 & w10982;
assign w11015 = w11013 & w11014;
assign w11016 = w10982 & w10996;
assign w11017 = w10996 & w63634;
assign w11018 = ~w11015 & ~w11017;
assign w11019 = w10995 & ~w10996;
assign w11020 = ~w11013 & w11019;
assign w11021 = w11018 & ~w11020;
assign w11022 = w10961 & ~w10982;
assign w11023 = ~w10987 & w11022;
assign w11024 = w10968 & ~w10999;
assign w11025 = ~w11023 & w11024;
assign w11026 = ~w10968 & ~w10987;
assign w11027 = ~w11016 & w11026;
assign w11028 = ~w11025 & ~w11027;
assign w11029 = w11009 & w11021;
assign w11030 = ~w11028 & w11029;
assign w11031 = ~w11012 & ~w11030;
assign w11032 = ~w10976 & ~w10985;
assign w11033 = ~w11031 & w11032;
assign w11034 = pi0613 & w11033;
assign w11035 = ~pi0613 & ~w11033;
assign w11036 = ~w11034 & ~w11035;
assign w11037 = ~w10860 & ~w10881;
assign w11038 = ~w10846 & ~w10881;
assign w11039 = ~w11037 & ~w11038;
assign w11040 = ~w10883 & w11039;
assign w11041 = ~w10846 & w11040;
assign w11042 = w10859 & ~w10910;
assign w11043 = ~w10868 & ~w11042;
assign w11044 = ~w10840 & w11043;
assign w11045 = w10840 & w10860;
assign w11046 = w10860 & w64962;
assign w11047 = w10860 & w11038;
assign w11048 = ~w10867 & ~w11047;
assign w11049 = ~w10840 & w10859;
assign w11050 = w11038 & w11049;
assign w11051 = w10840 & w10853;
assign w11052 = ~w10881 & w11051;
assign w11053 = ~w10886 & w11052;
assign w11054 = ~w11046 & ~w11050;
assign w11055 = w11048 & ~w11053;
assign w11056 = w11054 & w11055;
assign w11057 = ~w11044 & w11056;
assign w11058 = ~w11041 & w11057;
assign w11059 = w10898 & w11049;
assign w11060 = w10867 & ~w11059;
assign w11061 = w10840 & ~w10853;
assign w11062 = w10891 & ~w11061;
assign w11063 = ~w10859 & w10890;
assign w11064 = w10890 & w64963;
assign w11065 = ~w10847 & ~w10891;
assign w11066 = ~w10910 & ~w11061;
assign w11067 = w11065 & ~w11066;
assign w11068 = ~w10903 & ~w11067;
assign w11069 = ~w10881 & ~w11068;
assign w11070 = w11060 & ~w11062;
assign w11071 = ~w11064 & w11070;
assign w11072 = ~w11069 & w11071;
assign w11073 = ~w10898 & ~w11061;
assign w11074 = ~w10869 & w10881;
assign w11075 = ~w11073 & w11074;
assign w11076 = (~w11075 & w11058) | (~w11075 & w64964) | (w11058 & w64964);
assign w11077 = ~pi0619 & w11076;
assign w11078 = pi0619 & ~w11076;
assign w11079 = ~w11077 & ~w11078;
assign w11080 = w10629 & w10654;
assign w11081 = w10684 & w11080;
assign w11082 = w10647 & w10692;
assign w11083 = ~w11081 & ~w11082;
assign w11084 = ~w10638 & ~w11083;
assign w11085 = w10684 & ~w10693;
assign w11086 = ~w10629 & ~w10644;
assign w11087 = w10673 & w11086;
assign w11088 = w10648 & ~w11087;
assign w11089 = ~w10684 & ~w11088;
assign w11090 = ~w11085 & ~w11089;
assign w11091 = ~w10638 & ~w10657;
assign w11092 = w10670 & ~w11091;
assign w11093 = ~w11084 & w11092;
assign w11094 = ~w11090 & w11093;
assign w11095 = w10683 & w11080;
assign w11096 = ~w10638 & ~w11095;
assign w11097 = ~w11088 & ~w11096;
assign w11098 = ~w10670 & ~w11085;
assign w11099 = ~w11097 & w11098;
assign w11100 = ~w11094 & ~w11099;
assign w11101 = pi0626 & w11100;
assign w11102 = ~pi0626 & ~w11100;
assign w11103 = ~w11101 & ~w11102;
assign w11104 = w10456 & w10506;
assign w11105 = ~w10478 & w64965;
assign w11106 = ~w10486 & ~w11105;
assign w11107 = w10472 & w11106;
assign w11108 = w10459 & w10463;
assign w11109 = (w10499 & w10474) | (w10499 & w63635) | (w10474 & w63635);
assign w11110 = w10427 & ~w10439;
assign w11111 = w10456 & ~w11110;
assign w11112 = w10433 & w10463;
assign w11113 = ~w11111 & w11112;
assign w11114 = ~w10458 & ~w11110;
assign w11115 = w10464 & ~w11114;
assign w11116 = ~w10474 & ~w11115;
assign w11117 = w10439 & w10482;
assign w11118 = w11116 & w11117;
assign w11119 = ~w11109 & ~w11113;
assign w11120 = ~w11118 & w11119;
assign w11121 = (w10493 & ~w11120) | (w10493 & w64966) | (~w11120 & w64966);
assign w11122 = w10477 & w11110;
assign w11123 = ~w10427 & w10454;
assign w11124 = w10433 & w11111;
assign w11125 = w10427 & ~w10433;
assign w11126 = ~w10427 & w10433;
assign w11127 = ~w10446 & ~w11125;
assign w11128 = ~w11126 & w11127;
assign w11129 = w10455 & w11128;
assign w11130 = ~w10463 & ~w10498;
assign w11131 = w10427 & w10446;
assign w11132 = w11130 & w11131;
assign w11133 = ~w11124 & ~w11132;
assign w11134 = ~w11123 & w11133;
assign w11135 = (~w11134 & w64967) | (~w11134 & w64968) | (w64967 & w64968);
assign w11136 = ~w11104 & ~w11122;
assign w11137 = ~w11135 & w11136;
assign w11138 = ~w11121 & w11137;
assign w11139 = ~pi0628 & w11138;
assign w11140 = pi0628 & ~w11138;
assign w11141 = ~w11139 & ~w11140;
assign w11142 = w10547 & ~w10575;
assign w11143 = ~w10600 & w11142;
assign w11144 = (~w10522 & ~w10592) | (~w10522 & w64969) | (~w10592 & w64969);
assign w11145 = w10528 & w10561;
assign w11146 = ~w10528 & ~w10588;
assign w11147 = w10592 & w63637;
assign w11148 = (w10522 & w11147) | (w10522 & w64970) | (w11147 & w64970);
assign w11149 = w10590 & ~w10727;
assign w11150 = ~w11144 & ~w11149;
assign w11151 = w11150 & w64971;
assign w11152 = (pi0623 & ~w11150) | (pi0623 & w64972) | (~w11150 & w64972);
assign w11153 = ~w11151 & ~w11152;
assign w11154 = ~w10968 & w10986;
assign w11155 = w10986 & w64973;
assign w11156 = ~w10961 & w11155;
assign w11157 = w10955 & ~w11000;
assign w11158 = ~w10955 & w10974;
assign w11159 = ~w10990 & ~w10995;
assign w11160 = w11158 & w11159;
assign w11161 = ~w11157 & ~w11160;
assign w11162 = ~w10968 & w11161;
assign w11163 = w10975 & w10995;
assign w11164 = w10968 & w10982;
assign w11165 = w10988 & w11164;
assign w11166 = ~w11163 & ~w11165;
assign w11167 = ~w10955 & ~w10982;
assign w11168 = ~w10968 & w11167;
assign w11169 = w10961 & w11013;
assign w11170 = ~w11167 & ~w11169;
assign w11171 = ~w11168 & ~w11170;
assign w11172 = w11018 & w11166;
assign w11173 = ~w11171 & w11172;
assign w11174 = (w10968 & ~w11173) | (w10968 & w64974) | (~w11173 & w64974);
assign w11175 = w11009 & ~w11162;
assign w11176 = ~w11174 & w11175;
assign w11177 = ~w11009 & ~w11173;
assign w11178 = ~w11163 & ~w11169;
assign w11179 = ~w11021 & ~w11178;
assign w11180 = w11013 & w11022;
assign w11181 = ~w11016 & ~w11180;
assign w11182 = w10968 & ~w11181;
assign w11183 = ~w10968 & ~w11009;
assign w11184 = ~w10962 & ~w11022;
assign w11185 = ~w11167 & w11183;
assign w11186 = ~w11184 & w11185;
assign w11187 = ~w11156 & ~w11186;
assign w11188 = ~w11182 & w11187;
assign w11189 = ~w11179 & w11188;
assign w11190 = ~w11177 & w11189;
assign w11191 = ~w11176 & w11190;
assign w11192 = ~pi0612 & w11191;
assign w11193 = pi0612 & ~w11191;
assign w11194 = ~w11192 & ~w11193;
assign w11195 = w10439 & w10446;
assign w11196 = ~w10481 & ~w11195;
assign w11197 = ~w10447 & w11196;
assign w11198 = w10427 & ~w11197;
assign w11199 = ~w11108 & ~w11198;
assign w11200 = ~w10493 & ~w11199;
assign w11201 = ~w10453 & w10493;
assign w11202 = w10502 & ~w11201;
assign w11203 = w10477 & w10498;
assign w11204 = ~w11202 & ~w11203;
assign w11205 = ~w10427 & ~w11204;
assign w11206 = ~w10471 & w11128;
assign w11207 = w11116 & ~w11123;
assign w11208 = w10493 & ~w11207;
assign w11209 = ~w11205 & ~w11206;
assign w11210 = ~w11208 & w11209;
assign w11211 = ~w11200 & w11210;
assign w11212 = pi0637 & ~w11211;
assign w11213 = ~pi0637 & w11211;
assign w11214 = ~w11212 & ~w11213;
assign w11215 = ~pi3517 & pi9040;
assign w11216 = ~pi3484 & ~pi9040;
assign w11217 = ~w11215 & ~w11216;
assign w11218 = pi0583 & ~w11217;
assign w11219 = ~pi0583 & w11217;
assign w11220 = ~w11218 & ~w11219;
assign w11221 = ~pi3531 & pi9040;
assign w11222 = ~pi3539 & ~pi9040;
assign w11223 = ~w11221 & ~w11222;
assign w11224 = pi0606 & ~w11223;
assign w11225 = ~pi0606 & w11223;
assign w11226 = ~w11224 & ~w11225;
assign w11227 = ~w11220 & w11226;
assign w11228 = ~pi3520 & pi9040;
assign w11229 = ~pi3522 & ~pi9040;
assign w11230 = ~w11228 & ~w11229;
assign w11231 = pi0590 & ~w11230;
assign w11232 = ~pi0590 & w11230;
assign w11233 = ~w11231 & ~w11232;
assign w11234 = ~pi3516 & pi9040;
assign w11235 = ~pi3526 & ~pi9040;
assign w11236 = ~w11234 & ~w11235;
assign w11237 = pi0587 & ~w11236;
assign w11238 = ~pi0587 & w11236;
assign w11239 = ~w11237 & ~w11238;
assign w11240 = (~w11239 & ~w11227) | (~w11239 & w64975) | (~w11227 & w64975);
assign w11241 = ~pi3519 & pi9040;
assign w11242 = ~pi3533 & ~pi9040;
assign w11243 = ~w11241 & ~w11242;
assign w11244 = pi0603 & ~w11243;
assign w11245 = ~pi0603 & w11243;
assign w11246 = ~w11244 & ~w11245;
assign w11247 = w11220 & ~w11246;
assign w11248 = ~w11226 & w11247;
assign w11249 = w11240 & ~w11248;
assign w11250 = w11220 & w11233;
assign w11251 = w11226 & w11250;
assign w11252 = w11226 & ~w11246;
assign w11253 = ~w11220 & ~w11233;
assign w11254 = w11252 & w11253;
assign w11255 = w11239 & ~w11254;
assign w11256 = ~w11251 & w11255;
assign w11257 = ~w11233 & w11239;
assign w11258 = (w11220 & ~w11257) | (w11220 & w11247) | (~w11257 & w11247);
assign w11259 = ~w11226 & ~w11258;
assign w11260 = (~w11249 & ~w11256) | (~w11249 & w64976) | (~w11256 & w64976);
assign w11261 = w11233 & w11246;
assign w11262 = w11226 & w11246;
assign w11263 = ~w11233 & ~w11262;
assign w11264 = w11220 & ~w11263;
assign w11265 = ~w11261 & w11264;
assign w11266 = ~w11260 & ~w11265;
assign w11267 = ~pi3530 & pi9040;
assign w11268 = ~pi3521 & ~pi9040;
assign w11269 = ~w11267 & ~w11268;
assign w11270 = pi0596 & ~w11269;
assign w11271 = ~pi0596 & w11269;
assign w11272 = ~w11270 & ~w11271;
assign w11273 = ~w11266 & w11272;
assign w11274 = ~w11226 & w11246;
assign w11275 = ~w11220 & ~w11274;
assign w11276 = w11240 & w11275;
assign w11277 = ~w11257 & ~w11274;
assign w11278 = w11258 & ~w11277;
assign w11279 = ~w11276 & ~w11278;
assign w11280 = ~w11272 & ~w11279;
assign w11281 = ~w11239 & w11246;
assign w11282 = w11227 & w11281;
assign w11283 = w11250 & w11252;
assign w11284 = w11226 & ~w11233;
assign w11285 = ~w11220 & w11246;
assign w11286 = ~w11284 & w11285;
assign w11287 = ~w11226 & w11233;
assign w11288 = ~w11284 & ~w11287;
assign w11289 = ~w11261 & ~w11288;
assign w11290 = w11239 & ~w11253;
assign w11291 = (~w11286 & ~w11289) | (~w11286 & w64977) | (~w11289 & w64977);
assign w11292 = ~w11281 & ~w11291;
assign w11293 = ~w11258 & ~w11261;
assign w11294 = w11292 & w11293;
assign w11295 = ~w11282 & ~w11283;
assign w11296 = ~w11280 & w11295;
assign w11297 = ~w11294 & w11296;
assign w11298 = ~w11273 & w11297;
assign w11299 = pi0609 & ~w11298;
assign w11300 = ~pi0609 & w11298;
assign w11301 = ~w11299 & ~w11300;
assign w11302 = w11256 & w11265;
assign w11303 = ~w11250 & ~w11253;
assign w11304 = w11220 & ~w11233;
assign w11305 = ~w11252 & ~w11304;
assign w11306 = w11288 & w11305;
assign w11307 = (w11239 & ~w11247) | (w11239 & w64978) | (~w11247 & w64978);
assign w11308 = ~w11306 & w11307;
assign w11309 = (~w11272 & w11306) | (~w11272 & w64979) | (w11306 & w64979);
assign w11310 = w11274 & w11303;
assign w11311 = ~w11309 & w11310;
assign w11312 = ~w11239 & ~w11252;
assign w11313 = w11272 & ~w11312;
assign w11314 = w11253 & w11262;
assign w11315 = ~w11313 & ~w11314;
assign w11316 = w11272 & w11275;
assign w11317 = w11288 & w11316;
assign w11318 = w11239 & ~w11317;
assign w11319 = ~w11315 & ~w11318;
assign w11320 = ~w11285 & w11287;
assign w11321 = w11240 & ~w11320;
assign w11322 = ~w11264 & ~w11286;
assign w11323 = ~w11233 & ~w11322;
assign w11324 = (~w11248 & w11256) | (~w11248 & w64980) | (w11256 & w64980);
assign w11325 = ~w11323 & w11324;
assign w11326 = ~w11272 & ~w11325;
assign w11327 = ~w11302 & ~w11311;
assign w11328 = ~w11319 & w11327;
assign w11329 = ~w11326 & w11328;
assign w11330 = pi0615 & ~w11329;
assign w11331 = ~pi0615 & w11329;
assign w11332 = ~w11330 & ~w11331;
assign w11333 = ~w10427 & w10462;
assign w11334 = w10472 & w11110;
assign w11335 = ~w10446 & w11130;
assign w11336 = w10470 & ~w11335;
assign w11337 = w10483 & ~w11196;
assign w11338 = ~w10503 & ~w11112;
assign w11339 = w10494 & w11338;
assign w11340 = ~w11336 & ~w11337;
assign w11341 = w11339 & w11340;
assign w11342 = w10476 & w11126;
assign w11343 = w10461 & w10482;
assign w11344 = ~w10493 & ~w11342;
assign w11345 = ~w10454 & w11344;
assign w11346 = ~w11129 & w11345;
assign w11347 = ~w11343 & w11346;
assign w11348 = ~w11341 & ~w11347;
assign w11349 = ~w10475 & ~w11334;
assign w11350 = ~w11333 & w11349;
assign w11351 = ~w11348 & w11350;
assign w11352 = pi0635 & ~w11351;
assign w11353 = ~pi0635 & w11351;
assign w11354 = ~w11352 & ~w11353;
assign w11355 = ~pi3492 & pi9040;
assign w11356 = ~pi3506 & ~pi9040;
assign w11357 = ~w11355 & ~w11356;
assign w11358 = pi0577 & ~w11357;
assign w11359 = ~pi0577 & w11357;
assign w11360 = ~w11358 & ~w11359;
assign w11361 = ~pi3493 & pi9040;
assign w11362 = ~pi3502 & ~pi9040;
assign w11363 = ~w11361 & ~w11362;
assign w11364 = pi0602 & ~w11363;
assign w11365 = ~pi0602 & w11363;
assign w11366 = ~w11364 & ~w11365;
assign w11367 = ~pi3496 & pi9040;
assign w11368 = ~pi3559 & ~pi9040;
assign w11369 = ~w11367 & ~w11368;
assign w11370 = pi0605 & ~w11369;
assign w11371 = ~pi0605 & w11369;
assign w11372 = ~w11370 & ~w11371;
assign w11373 = ~w11366 & w11372;
assign w11374 = ~pi3513 & pi9040;
assign w11375 = ~pi3527 & ~pi9040;
assign w11376 = ~w11374 & ~w11375;
assign w11377 = pi0597 & ~w11376;
assign w11378 = ~pi0597 & w11376;
assign w11379 = ~w11377 & ~w11378;
assign w11380 = w11373 & w11379;
assign w11381 = w11366 & ~w11372;
assign w11382 = ~pi3507 & pi9040;
assign w11383 = ~pi3505 & ~pi9040;
assign w11384 = ~w11382 & ~w11383;
assign w11385 = pi0575 & ~w11384;
assign w11386 = ~pi0575 & w11384;
assign w11387 = ~w11385 & ~w11386;
assign w11388 = w11381 & w11387;
assign w11389 = w11372 & ~w11387;
assign w11390 = w11379 & w11389;
assign w11391 = ~w11388 & ~w11390;
assign w11392 = ~pi3503 & pi9040;
assign w11393 = ~pi3490 & ~pi9040;
assign w11394 = ~w11392 & ~w11393;
assign w11395 = pi0582 & ~w11394;
assign w11396 = ~pi0582 & w11394;
assign w11397 = ~w11395 & ~w11396;
assign w11398 = (w11397 & ~w11391) | (w11397 & w64981) | (~w11391 & w64981);
assign w11399 = ~w11372 & ~w11387;
assign w11400 = ~w11366 & ~w11379;
assign w11401 = w11399 & w11400;
assign w11402 = ~w11380 & ~w11401;
assign w11403 = ~w11398 & w11402;
assign w11404 = w11360 & ~w11403;
assign w11405 = w11372 & w11387;
assign w11406 = ~w11399 & ~w11405;
assign w11407 = ~w11366 & ~w11406;
assign w11408 = ~w11388 & ~w11407;
assign w11409 = w11379 & ~w11408;
assign w11410 = w11360 & ~w11387;
assign w11411 = w11406 & ~w11410;
assign w11412 = w11389 & w11618;
assign w11413 = ~w11400 & ~w11412;
assign w11414 = w11411 & ~w11413;
assign w11415 = w11366 & ~w11379;
assign w11416 = (w11415 & ~w11406) | (w11415 & w64982) | (~w11406 & w64982);
assign w11417 = ~w11414 & ~w11416;
assign w11418 = ~w11409 & w11417;
assign w11419 = ~w11397 & ~w11418;
assign w11420 = ~w11379 & w11399;
assign w11421 = w11397 & ~w11412;
assign w11422 = w11360 & ~w11399;
assign w11423 = ~w11373 & ~w11420;
assign w11424 = ~w11422 & w11423;
assign w11425 = w11408 & w11424;
assign w11426 = w11421 & w11425;
assign w11427 = ~w11404 & ~w11426;
assign w11428 = ~w11419 & w11427;
assign w11429 = ~pi0622 & w11428;
assign w11430 = pi0622 & ~w11428;
assign w11431 = ~w11429 & ~w11430;
assign w11432 = w11360 & ~w11405;
assign w11433 = w11379 & w11387;
assign w11434 = ~w11420 & ~w11433;
assign w11435 = w11391 & w11432;
assign w11436 = w11434 & w11435;
assign w11437 = ~w11417 & w11436;
assign w11438 = w11400 & ~w11406;
assign w11439 = w11391 & ~w11438;
assign w11440 = ~w11360 & ~w11439;
assign w11441 = w11360 & ~w11389;
assign w11442 = (w11400 & w11411) | (w11400 & w63638) | (w11411 & w63638);
assign w11443 = ~w11366 & w11433;
assign w11444 = ~w11399 & w63639;
assign w11445 = ~w11443 & w11444;
assign w11446 = ~w11360 & ~w11400;
assign w11447 = ~w11406 & w11446;
assign w11448 = ~w11445 & ~w11447;
assign w11449 = ~w11442 & w11448;
assign w11450 = ~w11410 & ~w11443;
assign w11451 = w11449 & ~w11450;
assign w11452 = (~w11397 & w11451) | (~w11397 & w64983) | (w11451 & w64983);
assign w11453 = w11397 & ~w11449;
assign w11454 = ~w11366 & ~w11387;
assign w11455 = ~w11360 & ~w11454;
assign w11456 = ~w11399 & ~w11433;
assign w11457 = w11455 & ~w11456;
assign w11458 = w11366 & ~w11405;
assign w11459 = ~w11366 & w11405;
assign w11460 = ~w11458 & ~w11459;
assign w11461 = w11372 & w11460;
assign w11462 = w11457 & w11461;
assign w11463 = ~w11437 & ~w11462;
assign w11464 = ~w11453 & w11463;
assign w11465 = (pi0630 & ~w11464) | (pi0630 & w64984) | (~w11464 & w64984);
assign w11466 = w11464 & w64985;
assign w11467 = ~w11465 & ~w11466;
assign w11468 = ~w10872 & ~w11059;
assign w11469 = ~w11064 & w11468;
assign w11470 = w11468 & w64986;
assign w11471 = ~w11060 & ~w11470;
assign w11472 = ~w10899 & ~w11471;
assign w11473 = ~w10881 & ~w11472;
assign w11474 = ~w11045 & ~w11063;
assign w11475 = w11038 & w11474;
assign w11476 = w10881 & ~w11474;
assign w11477 = ~w10899 & ~w11059;
assign w11478 = w11477 & w64987;
assign w11479 = ~w11475 & ~w11476;
assign w11480 = (w10867 & ~w11479) | (w10867 & w64988) | (~w11479 & w64988);
assign w11481 = ~w10860 & w10881;
assign w11482 = w10900 & w11481;
assign w11483 = w11469 & w11482;
assign w11484 = ~w10840 & w10860;
assign w11485 = w11048 & w11484;
assign w11486 = ~w11483 & ~w11485;
assign w11487 = ~w11480 & w11486;
assign w11488 = ~w11473 & w11487;
assign w11489 = ~pi0627 & w11488;
assign w11490 = pi0627 & ~w11488;
assign w11491 = ~w11489 & ~w11490;
assign w11492 = w10768 & w10823;
assign w11493 = w10791 & w64989;
assign w11494 = ~w10795 & w10802;
assign w11495 = w10924 & ~w11494;
assign w11496 = w10768 & ~w10778;
assign w11497 = w10752 & w10761;
assign w11498 = w11496 & ~w11497;
assign w11499 = ~w11495 & ~w11498;
assign w11500 = ~w11493 & ~w11499;
assign w11501 = w10788 & ~w11500;
assign w11502 = w10777 & w10813;
assign w11503 = w10790 & w11496;
assign w11504 = w10792 & w10809;
assign w11505 = ~w10828 & ~w11502;
assign w11506 = ~w11504 & w11505;
assign w11507 = w10940 & w11506;
assign w11508 = (~w10788 & ~w11507) | (~w10788 & w64990) | (~w11507 & w64990);
assign w11509 = ~w10938 & ~w11493;
assign w11510 = ~w10768 & ~w11509;
assign w11511 = ~w10936 & ~w11492;
assign w11512 = ~w11510 & w11511;
assign w11513 = ~w11508 & w11512;
assign w11514 = ~w11501 & w11513;
assign w11515 = pi0625 & ~w11514;
assign w11516 = ~pi0625 & w11514;
assign w11517 = ~w11515 & ~w11516;
assign w11518 = w11014 & w11158;
assign w11519 = ~w10961 & w11518;
assign w11520 = w10962 & w11164;
assign w11521 = w10961 & w10996;
assign w11522 = ~w11014 & ~w11521;
assign w11523 = ~w10990 & ~w11522;
assign w11524 = w11009 & ~w11520;
assign w11525 = ~w11020 & w11524;
assign w11526 = w11178 & w11525;
assign w11527 = ~w11523 & w11526;
assign w11528 = ~w10975 & w11022;
assign w11529 = ~w11154 & w11528;
assign w11530 = ~w10991 & ~w11164;
assign w11531 = ~w10962 & ~w11530;
assign w11532 = ~w10961 & w11154;
assign w11533 = ~w11009 & ~w11529;
assign w11534 = ~w11532 & w11533;
assign w11535 = ~w11531 & w11534;
assign w11536 = ~w11179 & w11535;
assign w11537 = (~w11519 & w11536) | (~w11519 & w64991) | (w11536 & w64991);
assign w11538 = ~pi0620 & w11537;
assign w11539 = pi0620 & ~w11537;
assign w11540 = ~w11538 & ~w11539;
assign w11541 = w10922 & ~w10937;
assign w11542 = w10922 & w64992;
assign w11543 = (~w10808 & ~w10820) | (~w10808 & w63640) | (~w10820 & w63640);
assign w11544 = ~w10796 & ~w11543;
assign w11545 = ~w10928 & ~w11544;
assign w11546 = (w10788 & ~w11545) | (w10788 & w64993) | (~w11545 & w64993);
assign w11547 = ~w10939 & ~w11493;
assign w11548 = w10768 & ~w11547;
assign w11549 = ~w11541 & w11543;
assign w11550 = w10824 & ~w11549;
assign w11551 = ~w10788 & ~w11550;
assign w11552 = ~w10929 & ~w11548;
assign w11553 = ~w11546 & w11552;
assign w11554 = ~w11551 & w11553;
assign w11555 = pi0633 & ~w11554;
assign w11556 = ~pi0633 & w11554;
assign w11557 = ~w11555 & ~w11556;
assign w11558 = ~w10675 & w64994;
assign w11559 = w10638 & ~w11558;
assign w11560 = w10644 & w10675;
assign w11561 = ~w10683 & ~w10692;
assign w11562 = w10632 & ~w11561;
assign w11563 = w10677 & ~w11560;
assign w11564 = ~w11562 & w11563;
assign w11565 = (w11083 & w11564) | (w11083 & w64995) | (w11564 & w64995);
assign w11566 = ~w10670 & ~w11565;
assign w11567 = w10683 & w10692;
assign w11568 = ~w11558 & ~w11567;
assign w11569 = w10670 & ~w11568;
assign w11570 = ~w10638 & w11083;
assign w11571 = ~w11569 & w11570;
assign w11572 = w10670 & ~w10676;
assign w11573 = w11083 & w11572;
assign w11574 = w10638 & ~w11567;
assign w11575 = ~w11573 & w11574;
assign w11576 = ~w11571 & ~w11575;
assign w11577 = ~w11566 & ~w11576;
assign w11578 = ~pi0641 & w11577;
assign w11579 = pi0641 & ~w11577;
assign w11580 = ~w11578 & ~w11579;
assign w11581 = w11409 & w11432;
assign w11582 = ~w11360 & ~w11372;
assign w11583 = w11434 & w11582;
assign w11584 = ~w11441 & w11458;
assign w11585 = ~w11379 & ~w11584;
assign w11586 = w11408 & w11585;
assign w11587 = w11421 & ~w11583;
assign w11588 = ~w11586 & w11587;
assign w11589 = w11422 & ~w11460;
assign w11590 = (~w11420 & ~w11460) | (~w11420 & w64996) | (~w11460 & w64996);
assign w11591 = ~w11360 & ~w11590;
assign w11592 = ~w11397 & ~w11401;
assign w11593 = ~w11589 & w11592;
assign w11594 = ~w11591 & w11593;
assign w11595 = ~w11588 & ~w11594;
assign w11596 = ~w11360 & w11443;
assign w11597 = ~w11581 & ~w11596;
assign w11598 = ~w11595 & w11597;
assign w11599 = pi0611 & w11598;
assign w11600 = ~pi0611 & ~w11598;
assign w11601 = ~w11599 & ~w11600;
assign w11602 = ~w10859 & w10911;
assign w11603 = w10870 & ~w10881;
assign w11604 = ~w11043 & w11603;
assign w11605 = w10881 & w11043;
assign w11606 = w10867 & ~w11602;
assign w11607 = ~w11605 & w11606;
assign w11608 = ~w11604 & w11607;
assign w11609 = w10874 & ~w11065;
assign w11610 = w10900 & ~w11063;
assign w11611 = ~w11067 & ~w11609;
assign w11612 = w11610 & w11611;
assign w11613 = ~w11608 & ~w11612;
assign w11614 = ~w11040 & ~w11613;
assign w11615 = pi0649 & w11614;
assign w11616 = ~pi0649 & ~w11614;
assign w11617 = ~w11615 & ~w11616;
assign w11618 = w11366 & w11379;
assign w11619 = w11582 & w11618;
assign w11620 = ~w11397 & ~w11619;
assign w11621 = w11379 & w11458;
assign w11622 = ~w11457 & ~w11621;
assign w11623 = (~w11620 & w11436) | (~w11620 & w64997) | (w11436 & w64997);
assign w11624 = ~w11366 & ~w11439;
assign w11625 = ~w11381 & ~w11433;
assign w11626 = w11455 & w11625;
assign w11627 = ~w11624 & ~w11626;
assign w11628 = ~w11397 & ~w11627;
assign w11629 = ~w11397 & ~w11621;
assign w11630 = ~w11373 & ~w11629;
assign w11631 = w11360 & ~w11625;
assign w11632 = ~w11630 & w11631;
assign w11633 = ~w11623 & ~w11632;
assign w11634 = ~w11628 & w11633;
assign w11635 = pi0631 & ~w11634;
assign w11636 = ~pi0631 & w11634;
assign w11637 = ~w11635 & ~w11636;
assign w11638 = (~w10968 & w11169) | (~w10968 & w11168) | (w11169 & w11168);
assign w11639 = w11158 & w11164;
assign w11640 = ~w11180 & ~w11521;
assign w11641 = ~w11639 & w11640;
assign w11642 = (w11009 & ~w11641) | (w11009 & w64998) | (~w11641 & w64998);
assign w11643 = w10961 & w10986;
assign w11644 = ~w10997 & ~w11643;
assign w11645 = w11183 & ~w11644;
assign w11646 = ~w10968 & w10992;
assign w11647 = w10955 & w11166;
assign w11648 = ~w11646 & w11647;
assign w11649 = ~w10994 & w11648;
assign w11650 = w10974 & w11167;
assign w11651 = ~w10998 & ~w11650;
assign w11652 = ~w11017 & w11651;
assign w11653 = w10968 & ~w11652;
assign w11654 = ~w10985 & ~w11518;
assign w11655 = ~w11653 & w11654;
assign w11656 = ~w11009 & ~w11655;
assign w11657 = ~w11155 & ~w11645;
assign w11658 = ~w11642 & w11657;
assign w11659 = ~w11649 & w11658;
assign w11660 = ~w11656 & w11659;
assign w11661 = pi0614 & w11660;
assign w11662 = ~pi0614 & ~w11660;
assign w11663 = ~w11661 & ~w11662;
assign w11664 = ~w11239 & w11303;
assign w11665 = w11274 & w11664;
assign w11666 = w11251 & w11281;
assign w11667 = ~w11252 & w11303;
assign w11668 = ~w11252 & w64999;
assign w11669 = ~w11303 & ~w11314;
assign w11670 = ~w11668 & w11669;
assign w11671 = (~w11666 & w11670) | (~w11666 & w65000) | (w11670 & w65000);
assign w11672 = w11272 & ~w11671;
assign w11673 = w11263 & w11292;
assign w11674 = ~w11312 & ~w11664;
assign w11675 = ~w11667 & ~w11674;
assign w11676 = w11309 & ~w11675;
assign w11677 = w11272 & ~w11314;
assign w11678 = ~w11247 & w11263;
assign w11679 = w11677 & ~w11678;
assign w11680 = w11308 & w11679;
assign w11681 = ~w11665 & ~w11680;
assign w11682 = ~w11676 & w11681;
assign w11683 = w11682 & w65001;
assign w11684 = pi0632 & ~w11683;
assign w11685 = ~pi0632 & w11683;
assign w11686 = ~w11684 & ~w11685;
assign w11687 = w10638 & ~w11095;
assign w11688 = w10677 & ~w10689;
assign w11689 = ~w11687 & ~w11688;
assign w11690 = ~w10644 & ~w10675;
assign w11691 = ~w10673 & ~w11086;
assign w11692 = ~w11690 & ~w11691;
assign w11693 = w10623 & ~w10655;
assign w11694 = ~w10692 & w11693;
assign w11695 = w10638 & ~w11080;
assign w11696 = ~w11694 & w11695;
assign w11697 = ~w11692 & w11696;
assign w11698 = w10687 & w10693;
assign w11699 = (~w10638 & w11692) | (~w10638 & w65002) | (w11692 & w65002);
assign w11700 = ~w10670 & ~w11082;
assign w11701 = ~w11697 & w11700;
assign w11702 = ~w11699 & w11701;
assign w11703 = w10638 & w11694;
assign w11704 = w10647 & w10693;
assign w11705 = w11091 & ~w11694;
assign w11706 = ~w10658 & w10670;
assign w11707 = ~w11704 & w11706;
assign w11708 = ~w11703 & ~w11705;
assign w11709 = w11707 & w11708;
assign w11710 = (~w11689 & w11702) | (~w11689 & w65003) | (w11702 & w65003);
assign w11711 = ~pi0659 & w11710;
assign w11712 = pi0659 & ~w11710;
assign w11713 = ~w11711 & ~w11712;
assign w11714 = w11285 & w11287;
assign w11715 = w11255 & ~w11714;
assign w11716 = w11247 & w11284;
assign w11717 = w11275 & w11306;
assign w11718 = ~w11239 & ~w11716;
assign w11719 = ~w11717 & w11718;
assign w11720 = ~w11715 & ~w11719;
assign w11721 = w11239 & ~w11284;
assign w11722 = ~w11305 & w11721;
assign w11723 = w11250 & ~w11262;
assign w11724 = ~w11256 & w11723;
assign w11725 = w11677 & ~w11722;
assign w11726 = ~w11724 & w11725;
assign w11727 = ~w11289 & ~w11674;
assign w11728 = ~w11272 & w11291;
assign w11729 = ~w11727 & w11728;
assign w11730 = ~w11726 & ~w11729;
assign w11731 = ~w11720 & ~w11730;
assign w11732 = ~pi0640 & w11731;
assign w11733 = pi0640 & ~w11731;
assign w11734 = ~w11732 & ~w11733;
assign w11735 = ~pi3546 & pi9040;
assign w11736 = ~pi3572 & ~pi9040;
assign w11737 = ~w11735 & ~w11736;
assign w11738 = pi0638 & ~w11737;
assign w11739 = ~pi0638 & w11737;
assign w11740 = ~w11738 & ~w11739;
assign w11741 = ~pi3596 & pi9040;
assign w11742 = ~pi3592 & ~pi9040;
assign w11743 = ~w11741 & ~w11742;
assign w11744 = pi0639 & ~w11743;
assign w11745 = ~pi0639 & w11743;
assign w11746 = ~w11744 & ~w11745;
assign w11747 = ~pi3563 & pi9040;
assign w11748 = ~pi3584 & ~pi9040;
assign w11749 = ~w11747 & ~w11748;
assign w11750 = pi0661 & ~w11749;
assign w11751 = ~pi0661 & w11749;
assign w11752 = ~w11750 & ~w11751;
assign w11753 = ~pi3595 & pi9040;
assign w11754 = ~pi3566 & ~pi9040;
assign w11755 = ~w11753 & ~w11754;
assign w11756 = pi0668 & ~w11755;
assign w11757 = ~pi0668 & w11755;
assign w11758 = ~w11756 & ~w11757;
assign w11759 = ~w11752 & ~w11758;
assign w11760 = w11752 & w11758;
assign w11761 = ~w11759 & ~w11760;
assign w11762 = w11740 & w11758;
assign w11763 = ~pi3582 & pi9040;
assign w11764 = ~pi3594 & ~pi9040;
assign w11765 = ~w11763 & ~w11764;
assign w11766 = pi0642 & ~w11765;
assign w11767 = ~pi0642 & w11765;
assign w11768 = ~w11766 & ~w11767;
assign w11769 = ~w11762 & ~w11768;
assign w11770 = w11746 & ~w11761;
assign w11771 = w11769 & w11770;
assign w11772 = w11770 & w65004;
assign w11773 = ~w11740 & ~w11746;
assign w11774 = ~w11752 & w11773;
assign w11775 = ~w11740 & w11752;
assign w11776 = w11746 & w11775;
assign w11777 = ~w11774 & ~w11776;
assign w11778 = w11740 & w11752;
assign w11779 = ~w11746 & w11778;
assign w11780 = w11778 & w65005;
assign w11781 = w11777 & ~w11780;
assign w11782 = ~pi3554 & pi9040;
assign w11783 = ~pi3574 & ~pi9040;
assign w11784 = ~w11782 & ~w11783;
assign w11785 = pi0671 & ~w11784;
assign w11786 = ~pi0671 & w11784;
assign w11787 = ~w11785 & ~w11786;
assign w11788 = ~w11781 & w11787;
assign w11789 = ~w11768 & ~w11788;
assign w11790 = w11740 & ~w11758;
assign w11791 = ~w11746 & w11790;
assign w11792 = (w11768 & ~w11790) | (w11768 & w63641) | (~w11790 & w63641);
assign w11793 = w11746 & w11762;
assign w11794 = w11778 & ~w11793;
assign w11795 = w11746 & ~w11752;
assign w11796 = ~w11790 & w11795;
assign w11797 = w11792 & ~w11796;
assign w11798 = ~w11794 & w11797;
assign w11799 = w11787 & ~w11798;
assign w11800 = ~w11740 & w11758;
assign w11801 = ~w11752 & w11800;
assign w11802 = w11740 & ~w11795;
assign w11803 = ~w11801 & ~w11802;
assign w11804 = ~w11746 & ~w11759;
assign w11805 = ~w11759 & w65006;
assign w11806 = ~w11795 & ~w11805;
assign w11807 = ~w11803 & ~w11806;
assign w11808 = ~w11761 & w11773;
assign w11809 = ~w11807 & ~w11808;
assign w11810 = ~w11799 & w11809;
assign w11811 = ~w11789 & ~w11810;
assign w11812 = w11740 & ~w11761;
assign w11813 = w11768 & ~w11800;
assign w11814 = ~w11779 & w11813;
assign w11815 = ~w11812 & w11814;
assign w11816 = ~w11740 & w11768;
assign w11817 = w11795 & ~w11816;
assign w11818 = ~w11793 & ~w11817;
assign w11819 = ~w11815 & ~w11818;
assign w11820 = w11769 & ~w11805;
assign w11821 = w11775 & w65007;
assign w11822 = w11758 & w11773;
assign w11823 = (w11768 & ~w11773) | (w11768 & w65008) | (~w11773 & w65008);
assign w11824 = ~w11821 & w11823;
assign w11825 = ~w11820 & ~w11824;
assign w11826 = (~w11787 & w11819) | (~w11787 & w65009) | (w11819 & w65009);
assign w11827 = ~w11772 & ~w11826;
assign w11828 = ~w11811 & w11827;
assign w11829 = pi0672 & w11828;
assign w11830 = ~pi0672 & ~w11828;
assign w11831 = ~w11829 & ~w11830;
assign w11832 = ~pi3544 & pi9040;
assign w11833 = ~pi3578 & ~pi9040;
assign w11834 = ~w11832 & ~w11833;
assign w11835 = pi0653 & ~w11834;
assign w11836 = ~pi0653 & w11834;
assign w11837 = ~w11835 & ~w11836;
assign w11838 = ~pi3585 & pi9040;
assign w11839 = ~pi3561 & ~pi9040;
assign w11840 = ~w11838 & ~w11839;
assign w11841 = pi0646 & ~w11840;
assign w11842 = ~pi0646 & w11840;
assign w11843 = ~w11841 & ~w11842;
assign w11844 = w11837 & w11843;
assign w11845 = ~pi3589 & pi9040;
assign w11846 = ~pi3573 & ~pi9040;
assign w11847 = ~w11845 & ~w11846;
assign w11848 = pi0657 & ~w11847;
assign w11849 = ~pi0657 & w11847;
assign w11850 = ~w11848 & ~w11849;
assign w11851 = w11844 & w11850;
assign w11852 = ~pi3555 & pi9040;
assign w11853 = ~pi3596 & ~pi9040;
assign w11854 = ~w11852 & ~w11853;
assign w11855 = pi0652 & ~w11854;
assign w11856 = ~pi0652 & w11854;
assign w11857 = ~w11855 & ~w11856;
assign w11858 = w11850 & ~w11857;
assign w11859 = ~w11843 & ~w11858;
assign w11860 = ~w11843 & w11850;
assign w11861 = w11837 & w11860;
assign w11862 = w11860 & w65010;
assign w11863 = w11843 & ~w11850;
assign w11864 = ~w11837 & ~w11860;
assign w11865 = ~w11863 & w11864;
assign w11866 = w11864 & w65011;
assign w11867 = ~w11862 & ~w11866;
assign w11868 = w11859 & w11867;
assign w11869 = ~w11851 & ~w11868;
assign w11870 = ~pi3584 & pi9040;
assign w11871 = ~pi3589 & ~pi9040;
assign w11872 = ~w11870 & ~w11871;
assign w11873 = pi0658 & ~w11872;
assign w11874 = ~pi0658 & w11872;
assign w11875 = ~w11873 & ~w11874;
assign w11876 = ~pi3557 & pi9040;
assign w11877 = ~pi3591 & ~pi9040;
assign w11878 = ~w11876 & ~w11877;
assign w11879 = pi0660 & ~w11878;
assign w11880 = ~pi0660 & w11878;
assign w11881 = ~w11879 & ~w11880;
assign w11882 = w11875 & ~w11881;
assign w11883 = ~w11869 & w11882;
assign w11884 = ~w11843 & ~w11857;
assign w11885 = w11837 & w11884;
assign w11886 = w11884 & w12527;
assign w11887 = ~w11837 & w11850;
assign w11888 = ~w11844 & ~w11887;
assign w11889 = ~w11857 & ~w11888;
assign w11890 = ~w11862 & ~w11889;
assign w11891 = ~w11875 & ~w11881;
assign w11892 = ~w11890 & w11891;
assign w11893 = w11843 & w11875;
assign w11894 = w11858 & w11893;
assign w11895 = ~w11837 & w11863;
assign w11896 = w11857 & ~w11881;
assign w11897 = w11895 & w11896;
assign w11898 = ~w11850 & w11857;
assign w11899 = w11875 & ~w11898;
assign w11900 = w11844 & w11857;
assign w11901 = ~w11837 & ~w11843;
assign w11902 = ~w11858 & w11901;
assign w11903 = ~w11900 & ~w11902;
assign w11904 = ~w11899 & ~w11903;
assign w11905 = ~w11859 & w11887;
assign w11906 = (w11875 & w11905) | (w11875 & w65012) | (w11905 & w65012);
assign w11907 = ~w11875 & w11885;
assign w11908 = ~w11837 & ~w11857;
assign w11909 = w11863 & w11908;
assign w11910 = ~w11907 & ~w11909;
assign w11911 = ~w11904 & w11910;
assign w11912 = (w11881 & ~w11911) | (w11881 & w65013) | (~w11911 & w65013);
assign w11913 = ~w11886 & ~w11894;
assign w11914 = ~w11897 & w11913;
assign w11915 = ~w11892 & w11914;
assign w11916 = ~w11912 & w11915;
assign w11917 = ~w11883 & w11916;
assign w11918 = pi0685 & ~w11917;
assign w11919 = ~pi0685 & w11917;
assign w11920 = ~w11918 & ~w11919;
assign w11921 = ~pi3574 & pi9040;
assign w11922 = ~pi3551 & ~pi9040;
assign w11923 = ~w11921 & ~w11922;
assign w11924 = pi0643 & ~w11923;
assign w11925 = ~pi0643 & w11923;
assign w11926 = ~w11924 & ~w11925;
assign w11927 = ~pi3594 & pi9040;
assign w11928 = ~pi3547 & ~pi9040;
assign w11929 = ~w11927 & ~w11928;
assign w11930 = pi0665 & ~w11929;
assign w11931 = ~pi0665 & w11929;
assign w11932 = ~w11930 & ~w11931;
assign w11933 = w11926 & w11932;
assign w11934 = ~pi3566 & pi9040;
assign w11935 = ~pi3563 & ~pi9040;
assign w11936 = ~w11934 & ~w11935;
assign w11937 = pi0657 & ~w11936;
assign w11938 = ~pi0657 & w11936;
assign w11939 = ~w11937 & ~w11938;
assign w11940 = w11933 & ~w11939;
assign w11941 = ~pi3592 & pi9040;
assign w11942 = ~pi3582 & ~pi9040;
assign w11943 = ~w11941 & ~w11942;
assign w11944 = pi0651 & ~w11943;
assign w11945 = ~pi0651 & w11943;
assign w11946 = ~w11944 & ~w11945;
assign w11947 = ~w11939 & ~w11946;
assign w11948 = w11932 & w11939;
assign w11949 = ~w11947 & ~w11948;
assign w11950 = ~w11926 & ~w11946;
assign w11951 = w11939 & w11950;
assign w11952 = ~w11940 & ~w11951;
assign w11953 = ~w11949 & ~w11952;
assign w11954 = (~w11940 & w11952) | (~w11940 & w65014) | (w11952 & w65014);
assign w11955 = ~w11926 & w11932;
assign w11956 = w11947 & w11955;
assign w11957 = ~pi3572 & pi9040;
assign w11958 = ~pi3595 & ~pi9040;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = pi0645 & ~w11959;
assign w11961 = ~pi0645 & w11959;
assign w11962 = ~w11960 & ~w11961;
assign w11963 = ~w11956 & w11962;
assign w11964 = ~w11954 & w11963;
assign w11965 = ~w11926 & w11946;
assign w11966 = w11939 & w11965;
assign w11967 = ~w11932 & ~w11939;
assign w11968 = w11950 & w11967;
assign w11969 = ~w11966 & ~w11968;
assign w11970 = w11962 & ~w11969;
assign w11971 = ~w11932 & ~w11962;
assign w11972 = w11946 & w11971;
assign w11973 = (~w11972 & w11952) | (~w11972 & w63642) | (w11952 & w63642);
assign w11974 = ~w11970 & w11973;
assign w11975 = ~pi3551 & pi9040;
assign w11976 = ~pi3546 & ~pi9040;
assign w11977 = ~w11975 & ~w11976;
assign w11978 = pi0653 & ~w11977;
assign w11979 = ~pi0653 & w11977;
assign w11980 = ~w11978 & ~w11979;
assign w11981 = ~w11974 & w11980;
assign w11982 = w11926 & ~w11946;
assign w11983 = ~w11932 & w11982;
assign w11984 = (w11962 & ~w11982) | (w11962 & w65015) | (~w11982 & w65015);
assign w11985 = w11939 & ~w11946;
assign w11986 = ~w11932 & w11985;
assign w11987 = ~w11939 & w11946;
assign w11988 = w11926 & w11987;
assign w11989 = ~w11986 & ~w11988;
assign w11990 = w11962 & ~w11989;
assign w11991 = w11955 & w11987;
assign w11992 = (~w11991 & w11989) | (~w11991 & w65016) | (w11989 & w65016);
assign w11993 = ~w11984 & ~w11992;
assign w11994 = ~w11962 & ~w11966;
assign w11995 = ~w11955 & w11985;
assign w11996 = w11994 & ~w11995;
assign w11997 = w11965 & w11967;
assign w11998 = w11962 & ~w11997;
assign w11999 = w11926 & w11946;
assign w12000 = w11939 & w11999;
assign w12001 = w11998 & ~w12000;
assign w12002 = ~w11996 & ~w12001;
assign w12003 = w11933 & w11987;
assign w12004 = ~w11956 & ~w12003;
assign w12005 = ~w11983 & w12004;
assign w12006 = ~w12002 & w12005;
assign w12007 = ~w11980 & ~w12006;
assign w12008 = ~w11964 & ~w11993;
assign w12009 = ~w11981 & w12008;
assign w12010 = ~w12007 & w12009;
assign w12011 = pi0674 & ~w12010;
assign w12012 = ~pi0674 & w12010;
assign w12013 = ~w12011 & ~w12012;
assign w12014 = ~pi3552 & pi9040;
assign w12015 = ~pi3558 & ~pi9040;
assign w12016 = ~w12014 & ~w12015;
assign w12017 = pi0646 & ~w12016;
assign w12018 = ~pi0646 & w12016;
assign w12019 = ~w12017 & ~w12018;
assign w12020 = ~pi3593 & pi9040;
assign w12021 = ~pi3586 & ~pi9040;
assign w12022 = ~w12020 & ~w12021;
assign w12023 = pi0647 & ~w12022;
assign w12024 = ~pi0647 & w12022;
assign w12025 = ~w12023 & ~w12024;
assign w12026 = ~w12019 & w12025;
assign w12027 = ~pi3558 & pi9040;
assign w12028 = ~pi3593 & ~pi9040;
assign w12029 = ~w12027 & ~w12028;
assign w12030 = pi0660 & ~w12029;
assign w12031 = ~pi0660 & w12029;
assign w12032 = ~w12030 & ~w12031;
assign w12033 = ~pi3578 & pi9040;
assign w12034 = ~pi3585 & ~pi9040;
assign w12035 = ~w12033 & ~w12034;
assign w12036 = pi0638 & ~w12035;
assign w12037 = ~pi0638 & w12035;
assign w12038 = ~w12036 & ~w12037;
assign w12039 = ~w12032 & w12038;
assign w12040 = w12026 & w12039;
assign w12041 = ~w12019 & ~w12038;
assign w12042 = ~w12032 & w12041;
assign w12043 = w12041 & w65017;
assign w12044 = ~w12040 & ~w12043;
assign w12045 = ~w12019 & ~w12032;
assign w12046 = w12019 & w12032;
assign w12047 = ~w12045 & ~w12046;
assign w12048 = ~w12038 & w12047;
assign w12049 = w12044 & ~w12048;
assign w12050 = w12032 & ~w12038;
assign w12051 = ~w12039 & ~w12050;
assign w12052 = ~w12025 & ~w12041;
assign w12053 = w12051 & w12052;
assign w12054 = ~pi3591 & pi9040;
assign w12055 = ~pi3555 & ~pi9040;
assign w12056 = ~w12054 & ~w12055;
assign w12057 = pi0663 & ~w12056;
assign w12058 = ~pi0663 & w12056;
assign w12059 = ~w12057 & ~w12058;
assign w12060 = ~w12053 & w12059;
assign w12061 = ~w12049 & w12060;
assign w12062 = w12019 & w12038;
assign w12063 = ~w12041 & ~w12062;
assign w12064 = ~w12059 & ~w12063;
assign w12065 = (w12050 & w12063) | (w12050 & w63643) | (w12063 & w63643);
assign w12066 = w12041 & w12072;
assign w12067 = (~w12059 & w12065) | (~w12059 & w65018) | (w12065 & w65018);
assign w12068 = ~w12025 & w12032;
assign w12069 = ~w12019 & w12059;
assign w12070 = ~w12041 & ~w12069;
assign w12071 = w12068 & ~w12070;
assign w12072 = w12025 & ~w12032;
assign w12073 = ~w12068 & ~w12072;
assign w12074 = w12038 & ~w12069;
assign w12075 = w12073 & w12074;
assign w12076 = ~w12071 & ~w12075;
assign w12077 = ~w12067 & w12076;
assign w12078 = ~pi3586 & pi9040;
assign w12079 = ~pi3554 & ~pi9040;
assign w12080 = ~w12078 & ~w12079;
assign w12081 = pi0639 & ~w12080;
assign w12082 = ~pi0639 & w12080;
assign w12083 = ~w12081 & ~w12082;
assign w12084 = ~w12077 & ~w12083;
assign w12085 = ~w12025 & w12062;
assign w12086 = (w12032 & w12085) | (w12032 & w65019) | (w12085 & w65019);
assign w12087 = w12059 & ~w12086;
assign w12088 = w12019 & w12025;
assign w12089 = ~w12069 & ~w12088;
assign w12090 = w12039 & ~w12089;
assign w12091 = ~w12025 & w12038;
assign w12092 = w12047 & w12091;
assign w12093 = (~w12059 & w12089) | (~w12059 & w65020) | (w12089 & w65020);
assign w12094 = ~w12092 & w12093;
assign w12095 = ~w12087 & ~w12094;
assign w12096 = w12044 & ~w12095;
assign w12097 = w12083 & ~w12096;
assign w12098 = w12019 & ~w12059;
assign w12099 = w12073 & w12098;
assign w12100 = ~w12061 & ~w12099;
assign w12101 = ~w12084 & w12100;
assign w12102 = ~w12097 & w12101;
assign w12103 = pi0681 & ~w12102;
assign w12104 = ~pi0681 & w12102;
assign w12105 = ~w12103 & ~w12104;
assign w12106 = w11837 & w11898;
assign w12107 = ~w11885 & ~w12106;
assign w12108 = w11857 & w11887;
assign w12109 = (~w11875 & ~w11887) | (~w11875 & w12114) | (~w11887 & w12114);
assign w12110 = ~w11850 & ~w11857;
assign w12111 = ~w11844 & ~w11884;
assign w12112 = ~w12110 & w12111;
assign w12113 = w12109 & w12112;
assign w12114 = ~w11857 & ~w11875;
assign w12115 = w11844 & w12114;
assign w12116 = ~w11850 & w12115;
assign w12117 = ~w11851 & ~w12108;
assign w12118 = (w11875 & ~w12117) | (w11875 & w63644) | (~w12117 & w63644);
assign w12119 = ~w12113 & ~w12116;
assign w12120 = w12119 & w63645;
assign w12121 = w11837 & w11858;
assign w12122 = w12109 & ~w12121;
assign w12123 = w11875 & ~w11908;
assign w12124 = ~w11895 & w12123;
assign w12125 = ~w12122 & ~w12124;
assign w12126 = (~w11881 & w12120) | (~w11881 & w65021) | (w12120 & w65021);
assign w12127 = w11904 & w12110;
assign w12128 = (w11881 & ~w12119) | (w11881 & w65022) | (~w12119 & w65022);
assign w12129 = ~w11910 & ~w12122;
assign w12130 = w11860 & w11908;
assign w12131 = ~w11900 & ~w12130;
assign w12132 = w11875 & ~w12131;
assign w12133 = ~w12127 & ~w12132;
assign w12134 = ~w12129 & w12133;
assign w12135 = ~w12128 & w12134;
assign w12136 = (pi0682 & ~w12135) | (pi0682 & w65023) | (~w12135 & w65023);
assign w12137 = w12135 & w65024;
assign w12138 = ~w12136 & ~w12137;
assign w12139 = ~w11966 & ~w11988;
assign w12140 = ~w11933 & ~w11950;
assign w12141 = ~w11949 & w12140;
assign w12142 = w11999 & w63646;
assign w12143 = ~w11962 & ~w11997;
assign w12144 = w11952 & w12143;
assign w12145 = ~w12141 & ~w12142;
assign w12146 = w12144 & w12145;
assign w12147 = (~w11932 & w12146) | (~w11932 & w63647) | (w12146 & w63647);
assign w12148 = ~w11948 & ~w11950;
assign w12149 = ~w11985 & ~w12148;
assign w12150 = w11984 & ~w12149;
assign w12151 = ~w11939 & ~w11999;
assign w12152 = ~w12149 & w65025;
assign w12153 = w11926 & w11962;
assign w12154 = w11932 & w11946;
assign w12155 = ~w12153 & w12154;
assign w12156 = w12139 & w12155;
assign w12157 = ~w12152 & ~w12156;
assign w12158 = (w11980 & w12147) | (w11980 & w65026) | (w12147 & w65026);
assign w12159 = ~w11953 & ~w11962;
assign w12160 = w11967 & w11999;
assign w12161 = w11963 & ~w12160;
assign w12162 = ~w12159 & ~w12161;
assign w12163 = ~w11980 & ~w12150;
assign w12164 = ~w12146 & w12163;
assign w12165 = ~w12162 & ~w12164;
assign w12166 = ~w12158 & w12165;
assign w12167 = pi0689 & ~w12166;
assign w12168 = ~pi0689 & w12166;
assign w12169 = ~w12167 & ~w12168;
assign w12170 = ~pi3570 & pi9040;
assign w12171 = ~pi3571 & ~pi9040;
assign w12172 = ~w12170 & ~w12171;
assign w12173 = pi0654 & ~w12172;
assign w12174 = ~pi0654 & w12172;
assign w12175 = ~w12173 & ~w12174;
assign w12176 = ~pi3541 & pi9040;
assign w12177 = ~pi3587 & ~pi9040;
assign w12178 = ~w12176 & ~w12177;
assign w12179 = pi0671 & ~w12178;
assign w12180 = ~pi0671 & w12178;
assign w12181 = ~w12179 & ~w12180;
assign w12182 = ~pi3613 & pi9040;
assign w12183 = ~pi3579 & ~pi9040;
assign w12184 = ~w12182 & ~w12183;
assign w12185 = pi0634 & ~w12184;
assign w12186 = ~pi0634 & w12184;
assign w12187 = ~w12185 & ~w12186;
assign w12188 = ~pi3576 & pi9040;
assign w12189 = ~pi3540 & ~pi9040;
assign w12190 = ~w12188 & ~w12189;
assign w12191 = pi0668 & ~w12190;
assign w12192 = ~pi0668 & w12190;
assign w12193 = ~w12191 & ~w12192;
assign w12194 = ~w12187 & ~w12193;
assign w12195 = w12187 & w12193;
assign w12196 = ~w12194 & ~w12195;
assign w12197 = ~pi3571 & pi9040;
assign w12198 = ~pi3543 & ~pi9040;
assign w12199 = ~w12197 & ~w12198;
assign w12200 = pi0669 & ~w12199;
assign w12201 = ~pi0669 & w12199;
assign w12202 = ~w12200 & ~w12201;
assign w12203 = ~w12196 & w12202;
assign w12204 = ~pi3590 & pi9040;
assign w12205 = ~pi3556 & ~pi9040;
assign w12206 = ~w12204 & ~w12205;
assign w12207 = pi0644 & ~w12206;
assign w12208 = ~pi0644 & w12206;
assign w12209 = ~w12207 & ~w12208;
assign w12210 = ~w12187 & ~w12209;
assign w12211 = (w12202 & ~w12210) | (w12202 & w12223) | (~w12210 & w12223);
assign w12212 = w12181 & w12187;
assign w12213 = ~w12196 & ~w12212;
assign w12214 = ~w12211 & ~w12213;
assign w12215 = ~w12203 & ~w12214;
assign w12216 = ~w12181 & ~w12193;
assign w12217 = ~w12210 & w12216;
assign w12218 = w12187 & ~w12193;
assign w12219 = ~w12181 & ~w12187;
assign w12220 = w12209 & w12219;
assign w12221 = (w12202 & w12220) | (w12202 & w63648) | (w12220 & w63648);
assign w12222 = ~w12209 & ~w12219;
assign w12223 = ~w12181 & w12202;
assign w12224 = ~w12194 & ~w12223;
assign w12225 = w12222 & ~w12224;
assign w12226 = ~w12221 & ~w12225;
assign w12227 = w12193 & ~w12202;
assign w12228 = w12181 & w12227;
assign w12229 = ~w12217 & ~w12228;
assign w12230 = w12226 & w12229;
assign w12231 = ~w12214 & w63649;
assign w12232 = w12230 & w12231;
assign w12233 = ~w12181 & w12193;
assign w12234 = w12210 & w12233;
assign w12235 = w12212 & ~w12227;
assign w12236 = ~w12181 & ~w12202;
assign w12237 = ~w12218 & w12236;
assign w12238 = ~w12235 & ~w12237;
assign w12239 = ~w12209 & ~w12238;
assign w12240 = w12193 & w12209;
assign w12241 = w12187 & w12240;
assign w12242 = w12223 & w12241;
assign w12243 = ~w12234 & ~w12242;
assign w12244 = ~w12239 & w12243;
assign w12245 = (~w12175 & w12232) | (~w12175 & w65027) | (w12232 & w65027);
assign w12246 = w12175 & ~w12230;
assign w12247 = ~w12193 & ~w12209;
assign w12248 = w12181 & w12247;
assign w12249 = ~w12181 & ~w12247;
assign w12250 = ~w12248 & ~w12249;
assign w12251 = ~w12181 & w12196;
assign w12252 = w12181 & ~w12196;
assign w12253 = ~w12251 & ~w12252;
assign w12254 = ~w12236 & ~w12250;
assign w12255 = w12253 & w12254;
assign w12256 = ~w12187 & w12255;
assign w12257 = w12210 & w12227;
assign w12258 = ~w12202 & w12209;
assign w12259 = w12187 & w12258;
assign w12260 = ~w12253 & w12259;
assign w12261 = w12202 & w12248;
assign w12262 = ~w12257 & ~w12261;
assign w12263 = ~w12260 & w12262;
assign w12264 = ~w12256 & w12263;
assign w12265 = ~w12246 & w12264;
assign w12266 = w12265 & w65028;
assign w12267 = (~pi0675 & ~w12265) | (~pi0675 & w65029) | (~w12265 & w65029);
assign w12268 = ~w12266 & ~w12267;
assign w12269 = w12038 & ~w12089;
assign w12270 = w12025 & ~w12269;
assign w12271 = ~w12049 & w12270;
assign w12272 = ~w12043 & ~w12046;
assign w12273 = w12059 & ~w12272;
assign w12274 = w12083 & ~w12092;
assign w12275 = ~w12273 & w12274;
assign w12276 = ~w12271 & w12275;
assign w12277 = ~w12019 & ~w12025;
assign w12278 = w12051 & ~w12277;
assign w12279 = w12063 & w12278;
assign w12280 = ~w12051 & ~w12088;
assign w12281 = ~w12072 & ~w12088;
assign w12282 = w12051 & ~w12281;
assign w12283 = ~w12280 & ~w12282;
assign w12284 = w12279 & w12283;
assign w12285 = ~w12066 & ~w12083;
assign w12286 = w12025 & w12059;
assign w12287 = w12032 & ~w12286;
assign w12288 = ~w12052 & w12287;
assign w12289 = ~w12064 & ~w12090;
assign w12290 = ~w12288 & w12289;
assign w12291 = w12285 & w12290;
assign w12292 = ~w12284 & w12291;
assign w12293 = ~w12276 & ~w12292;
assign w12294 = ~pi0677 & w12293;
assign w12295 = pi0677 & ~w12293;
assign w12296 = ~w12294 & ~w12295;
assign w12297 = ~w12226 & w12233;
assign w12298 = w12202 & w12252;
assign w12299 = ~w12194 & ~w12212;
assign w12300 = (~w12234 & w12252) | (~w12234 & w65030) | (w12252 & w65030);
assign w12301 = ~w12202 & ~w12300;
assign w12302 = w12209 & ~w12233;
assign w12303 = w12299 & w12302;
assign w12304 = ~w12298 & ~w12303;
assign w12305 = ~w12301 & w12304;
assign w12306 = ~w12175 & ~w12305;
assign w12307 = w12211 & ~w12250;
assign w12308 = w12210 & w65031;
assign w12309 = ~w12236 & ~w12258;
assign w12310 = ~w12249 & ~w12309;
assign w12311 = ~w12241 & ~w12308;
assign w12312 = ~w12310 & w12311;
assign w12313 = ~w12307 & w12312;
assign w12314 = w12175 & ~w12313;
assign w12315 = ~w12297 & ~w12314;
assign w12316 = ~w12306 & w12315;
assign w12317 = ~pi0678 & w12316;
assign w12318 = pi0678 & ~w12316;
assign w12319 = ~w12317 & ~w12318;
assign w12320 = ~pi3556 & pi9040;
assign w12321 = ~pi3570 & ~pi9040;
assign w12322 = ~w12320 & ~w12321;
assign w12323 = pi0670 & ~w12322;
assign w12324 = ~pi0670 & w12322;
assign w12325 = ~w12323 & ~w12324;
assign w12326 = ~pi3579 & pi9040;
assign w12327 = ~pi3568 & ~pi9040;
assign w12328 = ~w12326 & ~w12327;
assign w12329 = pi0634 & ~w12328;
assign w12330 = ~pi0634 & w12328;
assign w12331 = ~w12329 & ~w12330;
assign w12332 = ~pi3542 & pi9040;
assign w12333 = ~pi3613 & ~pi9040;
assign w12334 = ~w12332 & ~w12333;
assign w12335 = pi0664 & ~w12334;
assign w12336 = ~pi0664 & w12334;
assign w12337 = ~w12335 & ~w12336;
assign w12338 = ~w12331 & w12337;
assign w12339 = ~pi3583 & pi9040;
assign w12340 = ~pi3569 & ~pi9040;
assign w12341 = ~w12339 & ~w12340;
assign w12342 = pi0654 & ~w12341;
assign w12343 = ~pi0654 & w12341;
assign w12344 = ~w12342 & ~w12343;
assign w12345 = w12338 & w12344;
assign w12346 = (~w12325 & ~w12338) | (~w12325 & w65032) | (~w12338 & w65032);
assign w12347 = ~pi3616 & pi9040;
assign w12348 = ~pi3542 & ~pi9040;
assign w12349 = ~w12347 & ~w12348;
assign w12350 = pi0650 & ~w12349;
assign w12351 = ~pi0650 & w12349;
assign w12352 = ~w12350 & ~w12351;
assign w12353 = w12344 & w12352;
assign w12354 = ~w12331 & ~w12337;
assign w12355 = w12331 & w12337;
assign w12356 = ~w12354 & ~w12355;
assign w12357 = w12353 & w12356;
assign w12358 = ~w12344 & w12352;
assign w12359 = w12354 & w12358;
assign w12360 = ~w12357 & ~w12359;
assign w12361 = w12337 & w12358;
assign w12362 = w12358 & w12338;
assign w12363 = w12360 & ~w12362;
assign w12364 = w12346 & ~w12363;
assign w12365 = ~pi3550 & pi9040;
assign w12366 = ~pi3548 & ~pi9040;
assign w12367 = ~w12365 & ~w12366;
assign w12368 = pi0648 & ~w12367;
assign w12369 = ~pi0648 & w12367;
assign w12370 = ~w12368 & ~w12369;
assign w12371 = ~w12337 & ~w12344;
assign w12372 = ~w12352 & w12371;
assign w12373 = ~w12344 & w12355;
assign w12374 = ~w12372 & ~w12373;
assign w12375 = w12325 & ~w12374;
assign w12376 = ~w12331 & w12352;
assign w12377 = ~w12337 & w12376;
assign w12378 = w12346 & ~w12377;
assign w12379 = (~w12325 & ~w12355) | (~w12325 & w65033) | (~w12355 & w65033);
assign w12380 = ~w12371 & w12379;
assign w12381 = w12378 & w12380;
assign w12382 = w12360 & ~w12375;
assign w12383 = (~w12370 & ~w12382) | (~w12370 & w65034) | (~w12382 & w65034);
assign w12384 = w12344 & ~w12352;
assign w12385 = ~w12346 & w12384;
assign w12386 = w12344 & w12354;
assign w12387 = w12331 & w12371;
assign w12388 = ~w12386 & ~w12387;
assign w12389 = w12337 & w12344;
assign w12390 = w12352 & w12389;
assign w12391 = w12331 & w12372;
assign w12392 = w12325 & ~w12390;
assign w12393 = ~w12391 & w12392;
assign w12394 = ~w12388 & w12393;
assign w12395 = w12325 & w12331;
assign w12396 = w12389 & w12395;
assign w12397 = ~w12325 & ~w12374;
assign w12398 = ~w12362 & ~w12396;
assign w12399 = ~w12385 & w12398;
assign w12400 = ~w12397 & w12399;
assign w12401 = ~w12394 & w12400;
assign w12402 = w12370 & ~w12401;
assign w12403 = ~w12364 & ~w12383;
assign w12404 = ~w12402 & w12403;
assign w12405 = ~pi0673 & w12404;
assign w12406 = pi0673 & ~w12404;
assign w12407 = ~w12405 & ~w12406;
assign w12408 = ~w11983 & w11994;
assign w12409 = w11998 & w63650;
assign w12410 = w11973 & w12409;
assign w12411 = w11926 & ~w11967;
assign w12412 = w11949 & w12411;
assign w12413 = (~w12412 & w12410) | (~w12412 & w65035) | (w12410 & w65035);
assign w12414 = w11980 & ~w12413;
assign w12415 = ~w11986 & w12004;
assign w12416 = w11984 & ~w12415;
assign w12417 = w11980 & ~w12142;
assign w12418 = ~w11971 & ~w11982;
assign w12419 = ~w12148 & ~w12418;
assign w12420 = w11967 & w12153;
assign w12421 = ~w12142 & ~w12420;
assign w12422 = ~w12419 & w12421;
assign w12423 = ~w12417 & ~w12422;
assign w12424 = ~w11933 & ~w11987;
assign w12425 = ~w11980 & ~w12424;
assign w12426 = ~w12154 & ~w12425;
assign w12427 = ~w11962 & ~w11999;
assign w12428 = ~w12426 & w12427;
assign w12429 = ~w12416 & ~w12428;
assign w12430 = ~w12423 & w12429;
assign w12431 = ~w12414 & w12430;
assign w12432 = pi0684 & ~w12431;
assign w12433 = ~pi0684 & w12431;
assign w12434 = ~w12432 & ~w12433;
assign w12435 = ~pi3615 & pi9040;
assign w12436 = ~pi3560 & ~pi9040;
assign w12437 = ~w12435 & ~w12436;
assign w12438 = pi0655 & ~w12437;
assign w12439 = ~pi0655 & w12437;
assign w12440 = ~w12438 & ~w12439;
assign w12441 = ~pi3548 & pi9040;
assign w12442 = ~pi3590 & ~pi9040;
assign w12443 = ~w12441 & ~w12442;
assign w12444 = pi0666 & ~w12443;
assign w12445 = ~pi0666 & w12443;
assign w12446 = ~w12444 & ~w12445;
assign w12447 = w12440 & ~w12446;
assign w12448 = ~w12440 & w12446;
assign w12449 = ~w12447 & ~w12448;
assign w12450 = ~pi3564 & pi9040;
assign w12451 = ~pi3565 & ~pi9040;
assign w12452 = ~w12450 & ~w12451;
assign w12453 = pi0662 & ~w12452;
assign w12454 = ~pi0662 & w12452;
assign w12455 = ~w12453 & ~w12454;
assign w12456 = ~pi3560 & pi9040;
assign w12457 = ~pi3553 & ~pi9040;
assign w12458 = ~w12456 & ~w12457;
assign w12459 = pi0643 & ~w12458;
assign w12460 = ~pi0643 & w12458;
assign w12461 = ~w12459 & ~w12460;
assign w12462 = ~w12455 & w12461;
assign w12463 = ~pi3577 & pi9040;
assign w12464 = ~pi3616 & ~pi9040;
assign w12465 = ~w12463 & ~w12464;
assign w12466 = pi0667 & ~w12465;
assign w12467 = ~pi0667 & w12465;
assign w12468 = ~w12466 & ~w12467;
assign w12469 = w12462 & w12468;
assign w12470 = ~w12449 & w12469;
assign w12471 = ~w12455 & ~w12468;
assign w12472 = ~w12446 & ~w12461;
assign w12473 = ~w12455 & w12472;
assign w12474 = ~w12440 & w12473;
assign w12475 = ~w12440 & w12468;
assign w12476 = w12440 & ~w12468;
assign w12477 = ~w12475 & ~w12476;
assign w12478 = ~w12446 & w12468;
assign w12479 = w12461 & ~w12478;
assign w12480 = w12477 & w12479;
assign w12481 = ~w12474 & ~w12480;
assign w12482 = w12447 & w12462;
assign w12483 = w12455 & w12461;
assign w12484 = w12449 & w12483;
assign w12485 = w12449 & w63651;
assign w12486 = ~w12482 & ~w12485;
assign w12487 = w12440 & ~w12455;
assign w12488 = w12446 & ~w12461;
assign w12489 = w12487 & w12488;
assign w12490 = ~w12485 & w65036;
assign w12491 = w12481 & w12490;
assign w12492 = ~w12440 & w12461;
assign w12493 = ~pi3588 & pi9040;
assign w12494 = ~pi3545 & ~pi9040;
assign w12495 = ~w12493 & ~w12494;
assign w12496 = pi0651 & ~w12495;
assign w12497 = ~pi0651 & w12495;
assign w12498 = ~w12496 & ~w12497;
assign w12499 = ~w12446 & w12498;
assign w12500 = w12492 & w12499;
assign w12501 = ~w12491 & ~w12500;
assign w12502 = w12471 & ~w12501;
assign w12503 = ~w12475 & ~w12487;
assign w12504 = w12472 & ~w12503;
assign w12505 = w12446 & ~w12468;
assign w12506 = ~w12447 & ~w12505;
assign w12507 = w12483 & ~w12506;
assign w12508 = ~w12504 & ~w12507;
assign w12509 = ~w12448 & ~w12472;
assign w12510 = ~w12479 & w12509;
assign w12511 = w12455 & w12510;
assign w12512 = w12508 & ~w12511;
assign w12513 = w12448 & ~w12455;
assign w12514 = ~w12462 & w12477;
assign w12515 = ~w12482 & ~w12513;
assign w12516 = (w12515 & ~w12508) | (w12515 & w65037) | (~w12508 & w65037);
assign w12517 = ~w12498 & ~w12516;
assign w12518 = (~w12470 & w12512) | (~w12470 & w65038) | (w12512 & w65038);
assign w12519 = ~w12517 & w12518;
assign w12520 = ~w12502 & w12519;
assign w12521 = pi0690 & w12520;
assign w12522 = ~pi0690 & ~w12520;
assign w12523 = ~w12521 & ~w12522;
assign w12524 = ~w11864 & w11882;
assign w12525 = ~w12121 & w12524;
assign w12526 = w11865 & w11891;
assign w12527 = w11837 & ~w11850;
assign w12528 = ~w11875 & w12527;
assign w12529 = ~w11857 & w11860;
assign w12530 = ~w11895 & ~w12121;
assign w12531 = w11875 & ~w12530;
assign w12532 = ~w11909 & ~w12528;
assign w12533 = ~w12529 & w12532;
assign w12534 = ~w11866 & w12533;
assign w12535 = ~w12531 & w12534;
assign w12536 = w11881 & ~w12535;
assign w12537 = w11851 & w11896;
assign w12538 = ~w12116 & ~w12537;
assign w12539 = ~w12525 & w12538;
assign w12540 = ~w12526 & w12539;
assign w12541 = ~w12129 & w12540;
assign w12542 = ~w12536 & w12541;
assign w12543 = pi0692 & w12542;
assign w12544 = ~pi0692 & ~w12542;
assign w12545 = ~w12543 & ~w12544;
assign w12546 = (~w12066 & w12283) | (~w12066 & w65039) | (w12283 & w65039);
assign w12547 = w12059 & ~w12546;
assign w12548 = w12025 & w12283;
assign w12549 = w12083 & ~w12548;
assign w12550 = ~w12041 & ~w12059;
assign w12551 = w12283 & w12550;
assign w12552 = w12285 & ~w12551;
assign w12553 = ~w12549 & ~w12552;
assign w12554 = ~w12019 & ~w12073;
assign w12555 = ~w12278 & ~w12554;
assign w12556 = w12019 & w12072;
assign w12557 = ~w12059 & ~w12556;
assign w12558 = ~w12555 & w12557;
assign w12559 = ~w12060 & w12083;
assign w12560 = ~w12558 & w12559;
assign w12561 = ~w12547 & ~w12560;
assign w12562 = ~w12553 & w12561;
assign w12563 = pi0700 & ~w12562;
assign w12564 = ~pi0700 & w12562;
assign w12565 = ~w12563 & ~w12564;
assign w12566 = w11790 & w65040;
assign w12567 = w11773 & w11760;
assign w12568 = ~w12566 & ~w12567;
assign w12569 = ~w11768 & ~w12568;
assign w12570 = w11746 & w11790;
assign w12571 = ~w11776 & ~w12570;
assign w12572 = w11768 & ~w12571;
assign w12573 = (~w11779 & w11777) | (~w11779 & w63652) | (w11777 & w63652);
assign w12574 = ~w12572 & w12573;
assign w12575 = (~w11787 & ~w12574) | (~w11787 & w65041) | (~w12574 & w65041);
assign w12576 = w11768 & w11774;
assign w12577 = w11792 & ~w11803;
assign w12578 = ~w11773 & ~w12570;
assign w12579 = ~w11771 & ~w12577;
assign w12580 = ~w11780 & ~w11801;
assign w12581 = ~w11821 & w12580;
assign w12582 = ~w11791 & ~w11793;
assign w12583 = w11814 & ~w12582;
assign w12584 = ~w11740 & w11746;
assign w12585 = ~w11768 & ~w11775;
assign w12586 = ~w12584 & w12585;
assign w12587 = w12582 & w12586;
assign w12588 = ~w12583 & ~w12587;
assign w12589 = (w11787 & ~w12588) | (w11787 & w65042) | (~w12588 & w65042);
assign w12590 = w11758 & w11817;
assign w12591 = ~w12589 & w12590;
assign w12592 = (w12579 & w65043) | (w12579 & w65044) | (w65043 & w65044);
assign w12593 = ~w12575 & w12592;
assign w12594 = ~w12591 & w12593;
assign w12595 = pi0697 & ~w12594;
assign w12596 = ~pi0697 & w12594;
assign w12597 = ~w12595 & ~w12596;
assign w12598 = w12325 & w12352;
assign w12599 = w12331 & ~w12352;
assign w12600 = ~w12598 & ~w12599;
assign w12601 = ~w12344 & w12600;
assign w12602 = w12331 & ~w12358;
assign w12603 = (w12325 & ~w12358) | (w12325 & w63654) | (~w12358 & w63654);
assign w12604 = w12337 & ~w12376;
assign w12605 = ~w12602 & w12604;
assign w12606 = ~w12603 & w12605;
assign w12607 = w12601 & w12606;
assign w12608 = w12356 & ~w12389;
assign w12609 = w12356 & w65045;
assign w12610 = ~w12370 & ~w12606;
assign w12611 = ~w12338 & ~w12353;
assign w12612 = w12346 & ~w12611;
assign w12613 = w12345 & w12598;
assign w12614 = ~w12609 & ~w12613;
assign w12615 = ~w12612 & w12614;
assign w12616 = w12610 & w12615;
assign w12617 = ~w12358 & w12395;
assign w12618 = ~w12356 & w12384;
assign w12619 = ~w12371 & ~w12390;
assign w12620 = ~w12325 & ~w12602;
assign w12621 = ~w12619 & w12620;
assign w12622 = w12370 & ~w12617;
assign w12623 = ~w12618 & w12622;
assign w12624 = ~w12621 & w12623;
assign w12625 = ~w12616 & ~w12624;
assign w12626 = ~w12359 & ~w12385;
assign w12627 = ~w12600 & ~w12626;
assign w12628 = ~w12607 & ~w12627;
assign w12629 = ~w12625 & w12628;
assign w12630 = pi0679 & w12629;
assign w12631 = ~pi0679 & ~w12629;
assign w12632 = ~w12630 & ~w12631;
assign w12633 = ~w11867 & w11875;
assign w12634 = w11843 & ~w11898;
assign w12635 = ~w11908 & ~w12114;
assign w12636 = w12634 & w12635;
assign w12637 = ~w11886 & ~w12115;
assign w12638 = w12114 & w12637;
assign w12639 = w11881 & ~w12130;
assign w12640 = ~w12636 & w12639;
assign w12641 = ~w12638 & w12640;
assign w12642 = w11861 & w11875;
assign w12643 = ~w11881 & ~w12642;
assign w12644 = w12637 & w12643;
assign w12645 = ~w12641 & ~w12644;
assign w12646 = ~w11881 & w11901;
assign w12647 = ~w11900 & ~w12646;
assign w12648 = w11850 & ~w12647;
assign w12649 = ~w11897 & ~w12648;
assign w12650 = ~w11875 & ~w12649;
assign w12651 = w11843 & ~w11882;
assign w12652 = ~w11908 & ~w12106;
assign w12653 = ~w11843 & w11875;
assign w12654 = ~w12651 & ~w12653;
assign w12655 = ~w12652 & w12654;
assign w12656 = ~w12633 & ~w12655;
assign w12657 = ~w12650 & w12656;
assign w12658 = ~w12645 & w12657;
assign w12659 = pi0686 & ~w12658;
assign w12660 = ~pi0686 & w12658;
assign w12661 = ~w12659 & ~w12660;
assign w12662 = w12196 & w12236;
assign w12663 = ~w12255 & ~w12662;
assign w12664 = ~w12232 & w12663;
assign w12665 = w12175 & ~w12664;
assign w12666 = w12202 & w12234;
assign w12667 = ~w12240 & ~w12247;
assign w12668 = (~w12667 & w12260) | (~w12667 & w63655) | (w12260 & w63655);
assign w12669 = (w12222 & w12662) | (w12222 & w65046) | (w12662 & w65046);
assign w12670 = ~w12228 & ~w12241;
assign w12671 = ~w12210 & ~w12259;
assign w12672 = ~w12299 & ~w12671;
assign w12673 = ~w12222 & w12223;
assign w12674 = w12299 & w12673;
assign w12675 = w12670 & ~w12672;
assign w12676 = (~w12175 & ~w12675) | (~w12175 & w65047) | (~w12675 & w65047);
assign w12677 = ~w12666 & ~w12669;
assign w12678 = ~w12668 & w12677;
assign w12679 = ~w12676 & w12678;
assign w12680 = ~w12665 & w12679;
assign w12681 = pi0688 & ~w12680;
assign w12682 = ~pi0688 & w12680;
assign w12683 = ~w12681 & ~w12682;
assign w12684 = w11746 & ~w11787;
assign w12685 = w11760 & w12684;
assign w12686 = ~w11807 & ~w12685;
assign w12687 = ~w11768 & ~w12686;
assign w12688 = (~w11787 & w11815) | (~w11787 & w65048) | (w11815 & w65048);
assign w12689 = w11775 & w11813;
assign w12690 = ~w11772 & ~w12689;
assign w12691 = ~w12688 & w12690;
assign w12692 = ~w12589 & w12691;
assign w12693 = ~w12687 & w12692;
assign w12694 = pi0698 & ~w12693;
assign w12695 = ~pi0698 & w12693;
assign w12696 = ~w12694 & ~w12695;
assign w12697 = ~w11926 & w11964;
assign w12698 = ~w11969 & ~w12148;
assign w12699 = ~w11962 & ~w12160;
assign w12700 = ~w12698 & w12699;
assign w12701 = ~w11998 & ~w12700;
assign w12702 = w11982 & w12146;
assign w12703 = w11989 & w12148;
assign w12704 = w11998 & w12703;
assign w12705 = ~w11991 & w12417;
assign w12706 = ~w12704 & w12705;
assign w12707 = ~w12702 & w12706;
assign w12708 = w11949 & ~w11966;
assign w12709 = ~w11962 & ~w12708;
assign w12710 = w11955 & ~w11987;
assign w12711 = ~w11980 & ~w12710;
assign w12712 = ~w11990 & w12711;
assign w12713 = ~w12709 & w12712;
assign w12714 = ~w12707 & ~w12713;
assign w12715 = ~w12697 & ~w12701;
assign w12716 = (pi0693 & w12714) | (pi0693 & w65049) | (w12714 & w65049);
assign w12717 = ~w12714 & w65050;
assign w12718 = ~w12716 & ~w12717;
assign w12719 = w12455 & ~w12461;
assign w12720 = w12448 & w12719;
assign w12721 = ~w12473 & ~w12720;
assign w12722 = w12468 & ~w12721;
assign w12723 = ~w12440 & w12722;
assign w12724 = w12490 & ~w12498;
assign w12725 = w12506 & w12510;
assign w12726 = ~w12449 & w12471;
assign w12727 = ~w12725 & ~w12726;
assign w12728 = ~w12724 & ~w12727;
assign w12729 = w12478 & ~w12487;
assign w12730 = ~w12492 & w12729;
assign w12731 = w12448 & w12469;
assign w12732 = ~w12506 & w12719;
assign w12733 = (~w12498 & ~w12729) | (~w12498 & w65051) | (~w12729 & w65051);
assign w12734 = ~w12731 & ~w12732;
assign w12735 = w12733 & w12734;
assign w12736 = w12481 & w12735;
assign w12737 = w12449 & w12455;
assign w12738 = w12472 & w12503;
assign w12739 = w12737 & w12738;
assign w12740 = w12498 & ~w12739;
assign w12741 = w12486 & w12740;
assign w12742 = ~w12736 & ~w12741;
assign w12743 = ~w12742 & w65052;
assign w12744 = pi0676 & ~w12743;
assign w12745 = ~pi0676 & w12743;
assign w12746 = ~w12744 & ~w12745;
assign w12747 = w12440 & w12468;
assign w12748 = w12472 & w12747;
assign w12749 = ~w12484 & ~w12748;
assign w12750 = (w12498 & ~w12749) | (w12498 & w65053) | (~w12749 & w65053);
assign w12751 = ~w12487 & w12488;
assign w12752 = ~w12482 & ~w12751;
assign w12753 = w12498 & ~w12752;
assign w12754 = ~w12474 & ~w12484;
assign w12755 = ~w12753 & w12754;
assign w12756 = ~w12468 & ~w12755;
assign w12757 = ~w12489 & ~w12730;
assign w12758 = w12747 & ~w12757;
assign w12759 = w12449 & ~w12492;
assign w12760 = ~w12478 & ~w12505;
assign w12761 = w12461 & ~w12760;
assign w12762 = ~w12759 & ~w12761;
assign w12763 = ~w12455 & ~w12762;
assign w12764 = w12446 & ~w12462;
assign w12765 = w12475 & w12764;
assign w12766 = ~w12738 & ~w12765;
assign w12767 = ~w12763 & w12766;
assign w12768 = ~w12498 & ~w12767;
assign w12769 = ~w12750 & ~w12758;
assign w12770 = ~w12756 & w12769;
assign w12771 = ~w12768 & w12770;
assign w12772 = pi0683 & ~w12771;
assign w12773 = ~pi0683 & w12771;
assign w12774 = ~w12772 & ~w12773;
assign w12775 = ~w11746 & w11768;
assign w12776 = ~w12581 & w12775;
assign w12777 = w11740 & ~w11804;
assign w12778 = ~w11822 & ~w12777;
assign w12779 = w11768 & ~w12778;
assign w12780 = w11759 & w12584;
assign w12781 = ~w11787 & ~w12780;
assign w12782 = ~w12779 & w12781;
assign w12783 = ~w11760 & ~w12775;
assign w12784 = w11758 & w12775;
assign w12785 = ~w11740 & ~w12783;
assign w12786 = ~w12784 & w12785;
assign w12787 = w11740 & ~w11806;
assign w12788 = w11787 & ~w12786;
assign w12789 = ~w12787 & w12788;
assign w12790 = ~w12782 & ~w12789;
assign w12791 = w12586 & ~w12777;
assign w12792 = w12581 & w12791;
assign w12793 = ~w11752 & w11787;
assign w12794 = ~w11768 & w12584;
assign w12795 = ~w12793 & w12794;
assign w12796 = ~w12776 & ~w12795;
assign w12797 = ~w12792 & w12796;
assign w12798 = ~w12790 & w12797;
assign w12799 = pi0695 & ~w12798;
assign w12800 = ~pi0695 & w12798;
assign w12801 = ~w12799 & ~w12800;
assign w12802 = ~w12040 & w12059;
assign w12803 = w12032 & w12085;
assign w12804 = w12557 & ~w12803;
assign w12805 = ~w12802 & ~w12804;
assign w12806 = ~w12051 & w12277;
assign w12807 = (~w12059 & w12279) | (~w12059 & w65054) | (w12279 & w65054);
assign w12808 = ~w12042 & ~w12085;
assign w12809 = w12025 & w12065;
assign w12810 = (w12083 & w12808) | (w12083 & w65055) | (w12808 & w65055);
assign w12811 = ~w12809 & w12810;
assign w12812 = ~w12807 & w12811;
assign w12813 = ~w12025 & w12065;
assign w12814 = ~w12089 & w65056;
assign w12815 = w12064 & ~w12806;
assign w12816 = (~w12083 & ~w12063) | (~w12083 & w65057) | (~w12063 & w65057);
assign w12817 = ~w12814 & w12816;
assign w12818 = ~w12815 & w12817;
assign w12819 = ~w12813 & w12818;
assign w12820 = ~w12812 & ~w12819;
assign w12821 = ~w12805 & ~w12820;
assign w12822 = ~pi0699 & w12821;
assign w12823 = pi0699 & ~w12821;
assign w12824 = ~w12822 & ~w12823;
assign w12825 = ~pi3568 & pi9040;
assign w12826 = ~pi3575 & ~pi9040;
assign w12827 = ~w12825 & ~w12826;
assign w12828 = pi0648 & ~w12827;
assign w12829 = ~pi0648 & w12827;
assign w12830 = ~w12828 & ~w12829;
assign w12831 = ~pi3549 & pi9040;
assign w12832 = ~pi3564 & ~pi9040;
assign w12833 = ~w12831 & ~w12832;
assign w12834 = pi0636 & ~w12833;
assign w12835 = ~pi0636 & w12833;
assign w12836 = ~w12834 & ~w12835;
assign w12837 = ~w12830 & w12836;
assign w12838 = ~pi3543 & pi9040;
assign w12839 = ~pi3541 & ~pi9040;
assign w12840 = ~w12838 & ~w12839;
assign w12841 = pi0664 & ~w12840;
assign w12842 = ~pi0664 & w12840;
assign w12843 = ~w12841 & ~w12842;
assign w12844 = ~pi3545 & pi9040;
assign w12845 = ~pi3583 & ~pi9040;
assign w12846 = ~w12844 & ~w12845;
assign w12847 = pi0655 & ~w12846;
assign w12848 = ~pi0655 & w12846;
assign w12849 = ~w12847 & ~w12848;
assign w12850 = ~w12830 & ~w12849;
assign w12851 = w12830 & w12849;
assign w12852 = ~w12850 & ~w12851;
assign w12853 = ~pi3540 & pi9040;
assign w12854 = ~pi3615 & ~pi9040;
assign w12855 = ~w12853 & ~w12854;
assign w12856 = pi0656 & ~w12855;
assign w12857 = ~pi0656 & w12855;
assign w12858 = ~w12856 & ~w12857;
assign w12859 = ~w12843 & ~w12858;
assign w12860 = ~w12852 & w12859;
assign w12861 = w12830 & ~w12843;
assign w12862 = ~w12830 & ~w12858;
assign w12863 = ~w12861 & ~w12862;
assign w12864 = w12852 & w12863;
assign w12865 = ~w12860 & ~w12864;
assign w12866 = ~w12843 & ~w12865;
assign w12867 = w12837 & w12866;
assign w12868 = w12843 & ~w12849;
assign w12869 = ~w12830 & ~w12843;
assign w12870 = ~w12868 & ~w12869;
assign w12871 = ~w12843 & w12849;
assign w12872 = ~w12864 & ~w12871;
assign w12873 = ~pi3569 & pi9040;
assign w12874 = ~pi3550 & ~pi9040;
assign w12875 = ~w12873 & ~w12874;
assign w12876 = pi0666 & ~w12875;
assign w12877 = ~pi0666 & w12875;
assign w12878 = ~w12876 & ~w12877;
assign w12879 = ~w12836 & w12878;
assign w12880 = w12870 & w12879;
assign w12881 = w12872 & w12880;
assign w12882 = ~w12843 & w12858;
assign w12883 = w12836 & ~w12850;
assign w12884 = ~w12843 & w12851;
assign w12885 = w12843 & ~w12851;
assign w12886 = ~w12884 & ~w12885;
assign w12887 = w12883 & ~w12886;
assign w12888 = w12882 & w12887;
assign w12889 = w12843 & w12858;
assign w12890 = w12850 & w12889;
assign w12891 = w12836 & ~w12872;
assign w12892 = w12878 & ~w12890;
assign w12893 = ~w12891 & w12892;
assign w12894 = ~w12852 & w12882;
assign w12895 = w12830 & w12858;
assign w12896 = w12868 & w12895;
assign w12897 = ~w12894 & ~w12896;
assign w12898 = ~w12830 & w12849;
assign w12899 = w12889 & w12898;
assign w12900 = ~w12836 & w12899;
assign w12901 = ~w12837 & w12852;
assign w12902 = w12843 & ~w12858;
assign w12903 = ~w12901 & w12902;
assign w12904 = w12852 & w65058;
assign w12905 = ~w12878 & ~w12900;
assign w12906 = w12897 & w12905;
assign w12907 = ~w12903 & ~w12904;
assign w12908 = w12906 & w12907;
assign w12909 = ~w12893 & ~w12908;
assign w12910 = ~w12881 & ~w12888;
assign w12911 = ~w12867 & w12910;
assign w12912 = ~w12909 & w12911;
assign w12913 = pi0714 & ~w12912;
assign w12914 = ~pi0714 & w12912;
assign w12915 = ~w12913 & ~w12914;
assign w12916 = ~w12850 & w12886;
assign w12917 = (~w12862 & ~w12886) | (~w12862 & w63656) | (~w12886 & w63656);
assign w12918 = ~w12851 & w12870;
assign w12919 = (~w12836 & ~w12870) | (~w12836 & w65059) | (~w12870 & w65059);
assign w12920 = ~w12917 & w12919;
assign w12921 = ~w12917 & w65060;
assign w12922 = ~w12843 & w12895;
assign w12923 = ~w12837 & ~w12922;
assign w12924 = w12858 & ~w12861;
assign w12925 = w12883 & w12924;
assign w12926 = w12836 & w12859;
assign w12927 = ~w12898 & w12926;
assign w12928 = ~w12836 & ~w12859;
assign w12929 = ~w12852 & w12928;
assign w12930 = ~w12925 & ~w12927;
assign w12931 = ~w12929 & w12930;
assign w12932 = w12930 & w65061;
assign w12933 = w12931 & w63657;
assign w12934 = ~w12836 & ~w12865;
assign w12935 = (~w12878 & w12933) | (~w12878 & w65062) | (w12933 & w65062);
assign w12936 = w12878 & ~w12932;
assign w12937 = ~w12868 & w12895;
assign w12938 = w12836 & ~w12937;
assign w12939 = ~w12849 & w12902;
assign w12940 = w12938 & ~w12939;
assign w12941 = w12865 & w12940;
assign w12942 = w12918 & w12941;
assign w12943 = ~w12921 & ~w12942;
assign w12944 = ~w12936 & w12943;
assign w12945 = w12944 & w65063;
assign w12946 = (~pi0702 & ~w12944) | (~pi0702 & w65064) | (~w12944 & w65064);
assign w12947 = ~w12945 & ~w12946;
assign w12948 = ~w12212 & ~w12220;
assign w12949 = w12667 & ~w12948;
assign w12950 = ~w12215 & ~w12949;
assign w12951 = ~w12235 & ~w12670;
assign w12952 = w12175 & ~w12951;
assign w12953 = ~w12950 & ~w12952;
assign w12954 = w12209 & ~w12253;
assign w12955 = ~w12209 & ~w12212;
assign w12956 = w12203 & w12955;
assign w12957 = ~w12308 & ~w12956;
assign w12958 = ~w12954 & w12957;
assign w12959 = w12175 & ~w12958;
assign w12960 = ~w12953 & ~w12959;
assign w12961 = ~pi0680 & w12960;
assign w12962 = pi0680 & ~w12960;
assign w12963 = ~w12961 & ~w12962;
assign w12964 = ~w12378 & w12608;
assign w12965 = ~w12359 & ~w12964;
assign w12966 = w12370 & ~w12965;
assign w12967 = ~w12352 & w12389;
assign w12968 = ~w12386 & ~w12967;
assign w12969 = w12370 & ~w12968;
assign w12970 = w12379 & ~w12969;
assign w12971 = ~w12393 & ~w12970;
assign w12972 = ~w12376 & w12601;
assign w12973 = ~w12352 & w12354;
assign w12974 = ~w12396 & ~w12973;
assign w12975 = ~w12357 & w12974;
assign w12976 = ~w12972 & w12975;
assign w12977 = ~w12370 & ~w12976;
assign w12978 = ~w12971 & ~w12977;
assign w12979 = ~w12966 & w12978;
assign w12980 = ~pi0694 & w12979;
assign w12981 = pi0694 & ~w12979;
assign w12982 = ~w12980 & ~w12981;
assign w12983 = ~w12492 & ~w12513;
assign w12984 = ~w12506 & ~w12983;
assign w12985 = ~w12722 & ~w12984;
assign w12986 = w12490 & w12985;
assign w12987 = (~w12498 & ~w12985) | (~w12498 & w65065) | (~w12985 & w65065);
assign w12988 = w12498 & ~w12719;
assign w12989 = ~w12764 & w12988;
assign w12990 = (w12476 & w12989) | (w12476 & w65066) | (w12989 & w65066);
assign w12991 = w12455 & w12468;
assign w12992 = (w12991 & ~w12749) | (w12991 & w65067) | (~w12749 & w65067);
assign w12993 = ~w12475 & ~w12737;
assign w12994 = w12498 & ~w12993;
assign w12995 = w12986 & w12994;
assign w12996 = ~w12739 & ~w12990;
assign w12997 = ~w12992 & w12996;
assign w12998 = ~w12987 & w12997;
assign w12999 = ~w12995 & w12998;
assign w13000 = pi0696 & ~w12999;
assign w13001 = ~pi0696 & w12999;
assign w13002 = ~w13000 & ~w13001;
assign w13003 = ~w12357 & ~w12618;
assign w13004 = w12331 & ~w13003;
assign w13005 = ~w12376 & ~w12388;
assign w13006 = (~w12370 & w13005) | (~w12370 & w63658) | (w13005 & w63658);
assign w13007 = ~w13004 & ~w13006;
assign w13008 = ~w12325 & ~w13007;
assign w13009 = w12603 & ~w12973;
assign w13010 = ~w12391 & ~w12606;
assign w13011 = ~w13004 & w13010;
assign w13012 = (w12370 & ~w13011) | (w12370 & w63659) | (~w13011 & w63659);
assign w13013 = ~w12379 & w12610;
assign w13014 = w13007 & w13013;
assign w13015 = ~w13008 & ~w13012;
assign w13016 = (pi0687 & ~w13015) | (pi0687 & w65068) | (~w13015 & w65068);
assign w13017 = w13015 & w65069;
assign w13018 = ~w13016 & ~w13017;
assign w13019 = ~w12836 & w12922;
assign w13020 = ~w12897 & w12938;
assign w13021 = ~w12830 & w12868;
assign w13022 = w12836 & w13021;
assign w13023 = (~w12858 & w12916) | (~w12858 & w65070) | (w12916 & w65070);
assign w13024 = ~w12836 & ~w12849;
assign w13025 = ~w12862 & ~w12895;
assign w13026 = w13024 & w13025;
assign w13027 = w12878 & ~w12899;
assign w13028 = ~w13026 & w13027;
assign w13029 = ~w13023 & w13028;
assign w13030 = w12850 & w12859;
assign w13031 = ~w12878 & ~w13030;
assign w13032 = ~w12887 & w13031;
assign w13033 = ~w12920 & w13032;
assign w13034 = ~w13029 & ~w13033;
assign w13035 = ~w13019 & ~w13020;
assign w13036 = ~w13034 & w13035;
assign w13037 = pi0701 & w13036;
assign w13038 = ~pi0701 & ~w13036;
assign w13039 = ~w13037 & ~w13038;
assign w13040 = (~w12836 & ~w12870) | (~w12836 & w65071) | (~w12870 & w65071);
assign w13041 = ~w12940 & ~w13040;
assign w13042 = ~w12866 & ~w13041;
assign w13043 = ~w12878 & ~w13042;
assign w13044 = ~w12895 & ~w13021;
assign w13045 = w12879 & ~w13044;
assign w13046 = w12889 & w13024;
assign w13047 = ~w12889 & ~w12941;
assign w13048 = ~w12851 & w12878;
assign w13049 = ~w13047 & w13048;
assign w13050 = ~w13045 & ~w13046;
assign w13051 = ~w12888 & w13050;
assign w13052 = ~w13043 & w13051;
assign w13053 = (~pi0707 & ~w13052) | (~pi0707 & w65072) | (~w13052 & w65072);
assign w13054 = w13052 & w65073;
assign w13055 = ~w13053 & ~w13054;
assign w13056 = ~pi3605 & pi9040;
assign w13057 = ~pi3624 & ~pi9040;
assign w13058 = ~w13056 & ~w13057;
assign w13059 = pi0732 & ~w13058;
assign w13060 = ~pi0732 & w13058;
assign w13061 = ~w13059 & ~w13060;
assign w13062 = ~pi3648 & pi9040;
assign w13063 = ~pi3652 & ~pi9040;
assign w13064 = ~w13062 & ~w13063;
assign w13065 = pi0703 & ~w13064;
assign w13066 = ~pi0703 & w13064;
assign w13067 = ~w13065 & ~w13066;
assign w13068 = ~w13061 & w13067;
assign w13069 = w13061 & ~w13067;
assign w13070 = ~w13068 & ~w13069;
assign w13071 = ~pi3647 & pi9040;
assign w13072 = ~pi3607 & ~pi9040;
assign w13073 = ~w13071 & ~w13072;
assign w13074 = pi0726 & ~w13073;
assign w13075 = ~pi0726 & w13073;
assign w13076 = ~w13074 & ~w13075;
assign w13077 = w13070 & ~w13076;
assign w13078 = ~pi3614 & pi9040;
assign w13079 = ~pi3603 & ~pi9040;
assign w13080 = ~w13078 & ~w13079;
assign w13081 = pi0713 & ~w13080;
assign w13082 = ~pi0713 & w13080;
assign w13083 = ~w13081 & ~w13082;
assign w13084 = w13076 & ~w13083;
assign w13085 = ~w13068 & w13084;
assign w13086 = ~pi3642 & pi9040;
assign w13087 = ~pi3601 & ~pi9040;
assign w13088 = ~w13086 & ~w13087;
assign w13089 = pi0704 & ~w13088;
assign w13090 = ~pi0704 & w13088;
assign w13091 = ~w13089 & ~w13090;
assign w13092 = (~w13091 & w13077) | (~w13091 & w63660) | (w13077 & w63660);
assign w13093 = w13061 & ~w13083;
assign w13094 = w13067 & w13093;
assign w13095 = w13093 & w65074;
assign w13096 = ~w13067 & ~w13083;
assign w13097 = w13076 & w13096;
assign w13098 = (w13091 & ~w13096) | (w13091 & w65075) | (~w13096 & w65075);
assign w13099 = ~w13095 & w13098;
assign w13100 = w13061 & w13076;
assign w13101 = ~w13061 & ~w13076;
assign w13102 = ~w13100 & ~w13101;
assign w13103 = w13067 & w13083;
assign w13104 = ~w13102 & w13103;
assign w13105 = (~w13104 & w13092) | (~w13104 & w65076) | (w13092 & w65076);
assign w13106 = ~pi3640 & pi9040;
assign w13107 = ~pi3619 & ~pi9040;
assign w13108 = ~w13106 & ~w13107;
assign w13109 = pi0731 & ~w13108;
assign w13110 = ~pi0731 & w13108;
assign w13111 = ~w13109 & ~w13110;
assign w13112 = ~w13105 & ~w13111;
assign w13113 = w13067 & ~w13091;
assign w13114 = w13083 & w13101;
assign w13115 = w13113 & w13114;
assign w13116 = w13096 & ~w13102;
assign w13117 = w13068 & w13084;
assign w13118 = ~w13076 & w13083;
assign w13119 = ~w13067 & w13118;
assign w13120 = w13118 & w13069;
assign w13121 = ~w13117 & ~w13120;
assign w13122 = ~w13116 & w13121;
assign w13123 = w13091 & ~w13122;
assign w13124 = w13069 & w13083;
assign w13125 = (w13091 & ~w13069) | (w13091 & w65077) | (~w13069 & w65077);
assign w13126 = w13061 & w13103;
assign w13127 = w13103 & w65078;
assign w13128 = w13125 & ~w13127;
assign w13129 = w13068 & ~w13118;
assign w13130 = ~w13119 & ~w13129;
assign w13131 = w13128 & w13130;
assign w13132 = w13111 & ~w13131;
assign w13133 = ~w13123 & ~w13132;
assign w13134 = ~w13091 & ~w13094;
assign w13135 = ~w13084 & ~w13100;
assign w13136 = ~w13067 & ~w13093;
assign w13137 = ~w13135 & w13136;
assign w13138 = ~w13061 & w13096;
assign w13139 = w13134 & ~w13138;
assign w13140 = ~w13137 & w13139;
assign w13141 = ~w13133 & ~w13140;
assign w13142 = ~w13112 & ~w13115;
assign w13143 = ~w13141 & w13142;
assign w13144 = ~pi0736 & w13143;
assign w13145 = pi0736 & ~w13143;
assign w13146 = ~w13144 & ~w13145;
assign w13147 = ~pi3617 & pi9040;
assign w13148 = ~pi3642 & ~pi9040;
assign w13149 = ~w13147 & ~w13148;
assign w13150 = pi0716 & ~w13149;
assign w13151 = ~pi0716 & w13149;
assign w13152 = ~w13150 & ~w13151;
assign w13153 = ~pi3607 & pi9040;
assign w13154 = ~pi3614 & ~pi9040;
assign w13155 = ~w13153 & ~w13154;
assign w13156 = pi0708 & ~w13155;
assign w13157 = ~pi0708 & w13155;
assign w13158 = ~w13156 & ~w13157;
assign w13159 = ~w13152 & ~w13158;
assign w13160 = ~pi3643 & pi9040;
assign w13161 = ~pi3599 & ~pi9040;
assign w13162 = ~w13160 & ~w13161;
assign w13163 = pi0710 & ~w13162;
assign w13164 = ~pi0710 & w13162;
assign w13165 = ~w13163 & ~w13164;
assign w13166 = ~pi3619 & pi9040;
assign w13167 = ~pi3646 & ~pi9040;
assign w13168 = ~w13166 & ~w13167;
assign w13169 = pi0712 & ~w13168;
assign w13170 = ~pi0712 & w13168;
assign w13171 = ~w13169 & ~w13170;
assign w13172 = ~w13165 & ~w13171;
assign w13173 = ~pi3631 & pi9040;
assign w13174 = ~pi3608 & ~pi9040;
assign w13175 = ~w13173 & ~w13174;
assign w13176 = pi0727 & ~w13175;
assign w13177 = ~pi0727 & w13175;
assign w13178 = ~w13176 & ~w13177;
assign w13179 = w13172 & ~w13178;
assign w13180 = w13165 & ~w13171;
assign w13181 = w13178 & w13180;
assign w13182 = ~w13179 & ~w13181;
assign w13183 = w13159 & ~w13182;
assign w13184 = ~w13152 & w13158;
assign w13185 = ~w13165 & w13178;
assign w13186 = w13165 & w13171;
assign w13187 = ~w13185 & ~w13186;
assign w13188 = ~pi3603 & pi9040;
assign w13189 = ~pi3600 & ~pi9040;
assign w13190 = ~w13188 & ~w13189;
assign w13191 = pi0735 & ~w13190;
assign w13192 = ~pi0735 & w13190;
assign w13193 = ~w13191 & ~w13192;
assign w13194 = ~w13178 & w13186;
assign w13195 = w13159 & ~w13194;
assign w13196 = w13171 & w13185;
assign w13197 = w13195 & ~w13196;
assign w13198 = ~w13158 & ~w13165;
assign w13199 = w13158 & ~w13178;
assign w13200 = ~w13198 & ~w13199;
assign w13201 = ~w13181 & ~w13194;
assign w13202 = (w13152 & ~w13201) | (w13152 & w65079) | (~w13201 & w65079);
assign w13203 = (w13193 & w13187) | (w13193 & w65080) | (w13187 & w65080);
assign w13204 = ~w13197 & w13203;
assign w13205 = ~w13165 & w13171;
assign w13206 = w13199 & w13205;
assign w13207 = ~w13198 & ~w13206;
assign w13208 = w13152 & ~w13207;
assign w13209 = w13159 & w13180;
assign w13210 = w13158 & w13186;
assign w13211 = w13186 & w13199;
assign w13212 = ~w13209 & ~w13211;
assign w13213 = ~w13158 & w13178;
assign w13214 = ~w13199 & ~w13213;
assign w13215 = w13180 & ~w13184;
assign w13216 = ~w13214 & w13215;
assign w13217 = ~w13185 & ~w13213;
assign w13218 = ~w13152 & ~w13198;
assign w13219 = ~w13217 & w13218;
assign w13220 = ~w13216 & ~w13219;
assign w13221 = ~w13208 & w13220;
assign w13222 = w13212 & w13221;
assign w13223 = ~w13193 & ~w13222;
assign w13224 = ~w13198 & ~w13210;
assign w13225 = ~w13179 & ~w13196;
assign w13226 = w13152 & w13225;
assign w13227 = w13225 & w65081;
assign w13228 = ~w13224 & w13227;
assign w13229 = (~w13183 & ~w13204) | (~w13183 & w65082) | (~w13204 & w65082);
assign w13230 = ~w13228 & w13229;
assign w13231 = ~w13223 & w13230;
assign w13232 = pi0748 & w13231;
assign w13233 = ~pi0748 & ~w13231;
assign w13234 = ~w13232 & ~w13233;
assign w13235 = w13201 & w65083;
assign w13236 = ~w13159 & w13171;
assign w13237 = w13213 & w13236;
assign w13238 = ~w13205 & ~w13213;
assign w13239 = ~w13185 & ~w13238;
assign w13240 = w13226 & ~w13239;
assign w13241 = (w13226 & w65084) | (w13226 & w65085) | (w65084 & w65085);
assign w13242 = w13172 & ~w13213;
assign w13243 = ~w13210 & ~w13242;
assign w13244 = (w13152 & w13243) | (w13152 & w63662) | (w13243 & w63662);
assign w13245 = (w13243 & w65086) | (w13243 & w65087) | (w65086 & w65087);
assign w13246 = ~w13152 & ~w13243;
assign w13247 = ~w13158 & w13205;
assign w13248 = w13205 & w63663;
assign w13249 = w13193 & ~w13248;
assign w13250 = w13212 & w13249;
assign w13251 = ~w13246 & w13250;
assign w13252 = ~w13245 & w13251;
assign w13253 = ~w13241 & w13252;
assign w13254 = ~w13181 & w13184;
assign w13255 = w13159 & w13187;
assign w13256 = w13165 & w13201;
assign w13257 = w13244 & ~w13256;
assign w13258 = ~w13254 & ~w13255;
assign w13259 = ~w13193 & ~w13206;
assign w13260 = (w13259 & w13257) | (w13259 & w65088) | (w13257 & w65088);
assign w13261 = ~w13235 & ~w13237;
assign w13262 = (w13261 & w13253) | (w13261 & w65089) | (w13253 & w65089);
assign w13263 = pi0739 & w13262;
assign w13264 = ~pi0739 & ~w13262;
assign w13265 = ~w13263 & ~w13264;
assign w13266 = ~pi3629 & pi9040;
assign w13267 = ~pi3635 & ~pi9040;
assign w13268 = ~w13266 & ~w13267;
assign w13269 = pi0691 & ~w13268;
assign w13270 = ~pi0691 & w13268;
assign w13271 = ~w13269 & ~w13270;
assign w13272 = ~pi3621 & pi9040;
assign w13273 = ~pi3649 & ~pi9040;
assign w13274 = ~w13272 & ~w13273;
assign w13275 = pi0723 & ~w13274;
assign w13276 = ~pi0723 & w13274;
assign w13277 = ~w13275 & ~w13276;
assign w13278 = ~w13271 & w13277;
assign w13279 = ~pi3626 & pi9040;
assign w13280 = ~pi3622 & ~pi9040;
assign w13281 = ~w13279 & ~w13280;
assign w13282 = pi0733 & ~w13281;
assign w13283 = ~pi0733 & w13281;
assign w13284 = ~w13282 & ~w13283;
assign w13285 = ~w13277 & w13284;
assign w13286 = ~w13278 & ~w13285;
assign w13287 = ~pi3654 & pi9040;
assign w13288 = ~pi3628 & ~pi9040;
assign w13289 = ~w13287 & ~w13288;
assign w13290 = pi0728 & ~w13289;
assign w13291 = ~pi0728 & w13289;
assign w13292 = ~w13290 & ~w13291;
assign w13293 = w13286 & ~w13292;
assign w13294 = ~pi3622 & pi9040;
assign w13295 = ~pi3597 & ~pi9040;
assign w13296 = ~w13294 & ~w13295;
assign w13297 = pi0730 & ~w13296;
assign w13298 = ~pi0730 & w13296;
assign w13299 = ~w13297 & ~w13298;
assign w13300 = w13293 & w13299;
assign w13301 = ~w13271 & w13284;
assign w13302 = ~w13292 & w13301;
assign w13303 = ~w13277 & w13302;
assign w13304 = w13277 & w13292;
assign w13305 = w13284 & w13304;
assign w13306 = w13304 & w13301;
assign w13307 = w13271 & w13292;
assign w13308 = w13285 & w13307;
assign w13309 = ~pi3630 & pi9040;
assign w13310 = ~pi3609 & ~pi9040;
assign w13311 = ~w13309 & ~w13310;
assign w13312 = pi0717 & ~w13311;
assign w13313 = ~pi0717 & w13311;
assign w13314 = ~w13312 & ~w13313;
assign w13315 = ~w13308 & ~w13314;
assign w13316 = ~w13306 & w13315;
assign w13317 = ~w13303 & w13316;
assign w13318 = ~w13300 & w13317;
assign w13319 = ~w13278 & w13292;
assign w13320 = w13271 & ~w13277;
assign w13321 = w13299 & ~w13320;
assign w13322 = w13319 & w13321;
assign w13323 = ~w13284 & w13292;
assign w13324 = ~w13292 & w13320;
assign w13325 = ~w13323 & ~w13324;
assign w13326 = ~w13284 & w13324;
assign w13327 = w13299 & ~w13305;
assign w13328 = ~w13326 & w13327;
assign w13329 = ~w13325 & w13328;
assign w13330 = w13293 & ~w13299;
assign w13331 = w13284 & ~w13292;
assign w13332 = ~w13323 & ~w13331;
assign w13333 = w13278 & ~w13332;
assign w13334 = w13314 & ~w13322;
assign w13335 = ~w13333 & w13334;
assign w13336 = ~w13330 & w13335;
assign w13337 = ~w13329 & w13336;
assign w13338 = ~w13318 & ~w13337;
assign w13339 = w13277 & ~w13292;
assign w13340 = ~w13271 & w13339;
assign w13341 = ~w13271 & ~w13277;
assign w13342 = w13292 & w13341;
assign w13343 = w13341 & w13323;
assign w13344 = ~w13307 & ~w13340;
assign w13345 = ~w13343 & w13344;
assign w13346 = ~w13314 & ~w13345;
assign w13347 = ~w13302 & ~w13308;
assign w13348 = ~w13346 & w13347;
assign w13349 = ~w13299 & ~w13348;
assign w13350 = ~w13338 & w65090;
assign w13351 = (pi0740 & w13338) | (pi0740 & w65091) | (w13338 & w65091);
assign w13352 = ~w13350 & ~w13351;
assign w13353 = ~pi3698 & pi9040;
assign w13354 = ~pi3612 & ~pi9040;
assign w13355 = ~w13353 & ~w13354;
assign w13356 = pi0691 & ~w13355;
assign w13357 = ~pi0691 & w13355;
assign w13358 = ~w13356 & ~w13357;
assign w13359 = ~pi3612 & pi9040;
assign w13360 = ~pi3626 & ~pi9040;
assign w13361 = ~w13359 & ~w13360;
assign w13362 = pi0722 & ~w13361;
assign w13363 = ~pi0722 & w13361;
assign w13364 = ~w13362 & ~w13363;
assign w13365 = w13358 & ~w13364;
assign w13366 = ~pi3627 & pi9040;
assign w13367 = ~pi3620 & ~pi9040;
assign w13368 = ~w13366 & ~w13367;
assign w13369 = pi0726 & ~w13368;
assign w13370 = ~pi0726 & w13368;
assign w13371 = ~w13369 & ~w13370;
assign w13372 = ~w13358 & w13371;
assign w13373 = w13358 & ~w13371;
assign w13374 = ~w13372 & ~w13373;
assign w13375 = ~pi3625 & pi9040;
assign w13376 = ~pi3698 & ~pi9040;
assign w13377 = ~w13375 & ~w13376;
assign w13378 = pi0731 & ~w13377;
assign w13379 = ~pi0731 & w13377;
assign w13380 = ~w13378 & ~w13379;
assign w13381 = w13374 & w13380;
assign w13382 = ~w13374 & ~w13380;
assign w13383 = ~w13381 & ~w13382;
assign w13384 = ~pi3653 & pi9040;
assign w13385 = ~pi3604 & ~pi9040;
assign w13386 = ~w13384 & ~w13385;
assign w13387 = pi0706 & ~w13386;
assign w13388 = ~pi0706 & w13386;
assign w13389 = ~w13387 & ~w13388;
assign w13390 = ~w13383 & w13389;
assign w13391 = w13365 & w13390;
assign w13392 = w13364 & ~w13380;
assign w13393 = ~w13371 & ~w13392;
assign w13394 = w13364 & ~w13393;
assign w13395 = ~w13364 & ~w13372;
assign w13396 = ~w13389 & ~w13395;
assign w13397 = ~w13394 & w13396;
assign w13398 = ~w13358 & ~w13380;
assign w13399 = w13364 & w13389;
assign w13400 = w13398 & w13399;
assign w13401 = ~w13371 & w13400;
assign w13402 = ~w13371 & ~w13389;
assign w13403 = ~w13380 & ~w13402;
assign w13404 = ~w13364 & w13380;
assign w13405 = w13358 & ~w13404;
assign w13406 = ~w13403 & ~w13405;
assign w13407 = ~w13371 & ~w13406;
assign w13408 = w13371 & w13404;
assign w13409 = ~pi3649 & pi9040;
assign w13410 = ~pi3602 & ~pi9040;
assign w13411 = ~w13409 & ~w13410;
assign w13412 = pi0728 & ~w13411;
assign w13413 = ~pi0728 & w13411;
assign w13414 = ~w13412 & ~w13413;
assign w13415 = ~w13408 & w13414;
assign w13416 = w13358 & w13380;
assign w13417 = ~w13398 & ~w13416;
assign w13418 = ~w13365 & ~w13389;
assign w13419 = ~w13372 & w13418;
assign w13420 = w13417 & w13419;
assign w13421 = ~w13400 & ~w13420;
assign w13422 = ~w13407 & w13415;
assign w13423 = w13421 & w13422;
assign w13424 = w13364 & ~w13389;
assign w13425 = ~w13416 & w13424;
assign w13426 = w13371 & w13392;
assign w13427 = w13392 & w63664;
assign w13428 = w13402 & w13416;
assign w13429 = ~w13427 & ~w13428;
assign w13430 = ~w13424 & w13429;
assign w13431 = ~w13425 & ~w13430;
assign w13432 = ~w13364 & ~w13416;
assign w13433 = w13374 & w13432;
assign w13434 = ~w13372 & ~w13433;
assign w13435 = ~w13380 & ~w13389;
assign w13436 = w13358 & w13389;
assign w13437 = ~w13404 & ~w13436;
assign w13438 = ~w13393 & ~w13437;
assign w13439 = w13389 & ~w13398;
assign w13440 = ~w13438 & w13439;
assign w13441 = ~w13434 & w13440;
assign w13442 = (~w13433 & w65092) | (~w13433 & w65093) | (w65092 & w65093);
assign w13443 = ~w13441 & w13442;
assign w13444 = ~w13431 & w13443;
assign w13445 = ~w13423 & ~w13444;
assign w13446 = ~w13397 & ~w13401;
assign w13447 = ~w13391 & w13446;
assign w13448 = (pi0742 & w13445) | (pi0742 & w65094) | (w13445 & w65094);
assign w13449 = ~w13445 & w65095;
assign w13450 = ~w13448 & ~w13449;
assign w13451 = ~w13421 & w13426;
assign w13452 = w13371 & ~w13435;
assign w13453 = ~w13364 & ~w13417;
assign w13454 = ~w13452 & w13453;
assign w13455 = w13364 & w13381;
assign w13456 = ~w13374 & w13389;
assign w13457 = w13417 & w13456;
assign w13458 = ~w13414 & ~w13454;
assign w13459 = ~w13455 & ~w13457;
assign w13460 = w13458 & w13459;
assign w13461 = w13380 & ~w13389;
assign w13462 = w13372 & w13461;
assign w13463 = w13371 & w13436;
assign w13464 = ~w13403 & ~w13428;
assign w13465 = w13364 & ~w13464;
assign w13466 = ~w13364 & ~w13461;
assign w13467 = ~w13403 & w13466;
assign w13468 = w13414 & ~w13462;
assign w13469 = ~w13463 & w13468;
assign w13470 = ~w13467 & w13469;
assign w13471 = ~w13465 & w13470;
assign w13472 = ~w13460 & ~w13471;
assign w13473 = ~w13451 & ~w13472;
assign w13474 = ~pi0749 & w13473;
assign w13475 = pi0749 & ~w13473;
assign w13476 = ~w13474 & ~w13475;
assign w13477 = ~w13284 & w13307;
assign w13478 = ~w13303 & ~w13477;
assign w13479 = w13299 & ~w13478;
assign w13480 = w13284 & ~w13299;
assign w13481 = ~w13339 & w13480;
assign w13482 = ~w13319 & w13481;
assign w13483 = ~w13306 & ~w13481;
assign w13484 = ~w13482 & ~w13483;
assign w13485 = ~w13320 & ~w13340;
assign w13486 = ~w13284 & ~w13485;
assign w13487 = ~w13286 & ~w13299;
assign w13488 = (~w13284 & w13286) | (~w13284 & w63666) | (w13286 & w63666);
assign w13489 = w13271 & w13339;
assign w13490 = (w13284 & ~w13339) | (w13284 & w13301) | (~w13339 & w13301);
assign w13491 = ~w13488 & ~w13490;
assign w13492 = ~w13299 & w13340;
assign w13493 = ~w13314 & ~w13492;
assign w13494 = ~w13491 & w13493;
assign w13495 = ~w13484 & ~w13486;
assign w13496 = w13494 & w13495;
assign w13497 = ~w13284 & w13304;
assign w13498 = ~w13299 & ~w13497;
assign w13499 = w13271 & ~w13331;
assign w13500 = ~w13498 & w13499;
assign w13501 = w13271 & ~w13480;
assign w13502 = ~w13292 & ~w13301;
assign w13503 = ~w13501 & w13502;
assign w13504 = ~w13299 & w13503;
assign w13505 = w13314 & ~w13343;
assign w13506 = ~w13482 & w13505;
assign w13507 = ~w13500 & ~w13504;
assign w13508 = w13506 & w13507;
assign w13509 = ~w13496 & ~w13508;
assign w13510 = ~w13479 & ~w13509;
assign w13511 = ~pi0750 & w13510;
assign w13512 = pi0750 & ~w13510;
assign w13513 = ~w13511 & ~w13512;
assign w13514 = ~w13152 & w13201;
assign w13515 = ~w13159 & ~w13248;
assign w13516 = ~w13514 & ~w13515;
assign w13517 = ~w13171 & w13213;
assign w13518 = w13158 & ~w13225;
assign w13519 = w13152 & w13239;
assign w13520 = ~w13152 & w13165;
assign w13521 = ~w13178 & w13520;
assign w13522 = ~w13517 & ~w13521;
assign w13523 = ~w13248 & w13522;
assign w13524 = ~w13518 & w13523;
assign w13525 = (w13193 & ~w13524) | (w13193 & w65096) | (~w13524 & w65096);
assign w13526 = ~w13152 & ~w13225;
assign w13527 = w13178 & w13210;
assign w13528 = ~w13526 & ~w13527;
assign w13529 = ~w13240 & w13528;
assign w13530 = ~w13193 & ~w13529;
assign w13531 = ~w13516 & ~w13525;
assign w13532 = ~w13530 & w13531;
assign w13533 = pi0746 & w13532;
assign w13534 = ~pi0746 & ~w13532;
assign w13535 = ~w13533 & ~w13534;
assign w13536 = ~pi3608 & pi9040;
assign w13537 = ~pi3605 & ~pi9040;
assign w13538 = ~w13536 & ~w13537;
assign w13539 = pi0724 & ~w13538;
assign w13540 = ~pi0724 & w13538;
assign w13541 = ~w13539 & ~w13540;
assign w13542 = ~pi3601 & pi9040;
assign w13543 = ~pi3648 & ~pi9040;
assign w13544 = ~w13542 & ~w13543;
assign w13545 = pi0727 & ~w13544;
assign w13546 = ~pi0727 & w13544;
assign w13547 = ~w13545 & ~w13546;
assign w13548 = ~pi3600 & pi9040;
assign w13549 = ~pi3651 & ~pi9040;
assign w13550 = ~w13548 & ~w13549;
assign w13551 = pi0705 & ~w13550;
assign w13552 = ~pi0705 & w13550;
assign w13553 = ~w13551 & ~w13552;
assign w13554 = w13547 & w13553;
assign w13555 = ~pi3624 & pi9040;
assign w13556 = ~pi3647 & ~pi9040;
assign w13557 = ~w13555 & ~w13556;
assign w13558 = pi0734 & ~w13557;
assign w13559 = ~pi0734 & w13557;
assign w13560 = ~w13558 & ~w13559;
assign w13561 = w13554 & w13560;
assign w13562 = ~w13541 & w13561;
assign w13563 = ~w13547 & w13560;
assign w13564 = w13541 & ~w13553;
assign w13565 = ~w13563 & w13564;
assign w13566 = ~pi3652 & pi9040;
assign w13567 = ~pi3610 & ~pi9040;
assign w13568 = ~w13566 & ~w13567;
assign w13569 = pi0721 & ~w13568;
assign w13570 = ~pi0721 & w13568;
assign w13571 = ~w13569 & ~w13570;
assign w13572 = ~w13563 & w13571;
assign w13573 = ~w13541 & w13553;
assign w13574 = w13541 & w13560;
assign w13575 = ~w13547 & ~w13574;
assign w13576 = ~w13573 & w13575;
assign w13577 = w13547 & ~w13560;
assign w13578 = ~w13553 & ~w13560;
assign w13579 = w13541 & w13547;
assign w13580 = ~w13578 & ~w13579;
assign w13581 = ~w13577 & ~w13580;
assign w13582 = ~w13560 & w13573;
assign w13583 = (w13571 & ~w13573) | (w13571 & w63322) | (~w13573 & w63322);
assign w13584 = ~w13581 & w13583;
assign w13585 = ~w13576 & w13584;
assign w13586 = (~w13572 & ~w13584) | (~w13572 & w63323) | (~w13584 & w63323);
assign w13587 = w13553 & w13560;
assign w13588 = ~w13541 & w13577;
assign w13589 = ~w13587 & ~w13588;
assign w13590 = (~w13565 & w13586) | (~w13565 & w63667) | (w13586 & w63667);
assign w13591 = w13541 & ~w13571;
assign w13592 = ~w13573 & ~w13579;
assign w13593 = ~w13591 & w13592;
assign w13594 = ~w13590 & w13593;
assign w13595 = ~pi3636 & pi9040;
assign w13596 = ~pi3606 & ~pi9040;
assign w13597 = ~w13595 & ~w13596;
assign w13598 = pi0710 & ~w13597;
assign w13599 = ~pi0710 & w13597;
assign w13600 = ~w13598 & ~w13599;
assign w13601 = w13541 & ~w13560;
assign w13602 = ~w13563 & ~w13571;
assign w13603 = ~w13601 & w13602;
assign w13604 = ~w13561 & ~w13578;
assign w13605 = ~w13576 & w13604;
assign w13606 = w13571 & ~w13605;
assign w13607 = (w13553 & w13574) | (w13553 & w13554) | (w13574 & w13554);
assign w13608 = ~w13579 & w13607;
assign w13609 = (~w13608 & ~w13605) | (~w13608 & w65097) | (~w13605 & w65097);
assign w13610 = (w13600 & ~w13609) | (w13600 & w63668) | (~w13609 & w63668);
assign w13611 = ~w13553 & w13560;
assign w13612 = (~w13571 & ~w13611) | (~w13571 & w65098) | (~w13611 & w65098);
assign w13613 = ~w13553 & ~w13601;
assign w13614 = w13612 & w13613;
assign w13615 = ~w13547 & w13571;
assign w13616 = ~w13601 & ~w13615;
assign w13617 = w13553 & ~w13616;
assign w13618 = ~w13593 & w13617;
assign w13619 = (~w13600 & w13618) | (~w13600 & w65099) | (w13618 & w65099);
assign w13620 = w13591 & w13611;
assign w13621 = ~w13562 & ~w13620;
assign w13622 = ~w13619 & w13621;
assign w13623 = ~w13610 & w13622;
assign w13624 = w13623 & w65100;
assign w13625 = (pi0756 & ~w13623) | (pi0756 & w65101) | (~w13623 & w65101);
assign w13626 = ~w13624 & ~w13625;
assign w13627 = ~pi3650 & pi9040;
assign w13628 = ~pi3633 & ~pi9040;
assign w13629 = ~w13627 & ~w13628;
assign w13630 = pi0715 & ~w13629;
assign w13631 = ~pi0715 & w13629;
assign w13632 = ~w13630 & ~w13631;
assign w13633 = ~pi3632 & pi9040;
assign w13634 = ~pi3650 & ~pi9040;
assign w13635 = ~w13633 & ~w13634;
assign w13636 = pi0718 & ~w13635;
assign w13637 = ~pi0718 & w13635;
assign w13638 = ~w13636 & ~w13637;
assign w13639 = ~w13632 & w13638;
assign w13640 = ~pi3637 & pi9040;
assign w13641 = ~pi3623 & ~pi9040;
assign w13642 = ~w13640 & ~w13641;
assign w13643 = pi0719 & ~w13642;
assign w13644 = ~pi0719 & w13642;
assign w13645 = ~w13643 & ~w13644;
assign w13646 = w13639 & ~w13645;
assign w13647 = ~w13638 & w13645;
assign w13648 = ~pi3604 & pi9040;
assign w13649 = ~pi3630 & ~pi9040;
assign w13650 = ~w13648 & ~w13649;
assign w13651 = pi0705 & ~w13650;
assign w13652 = ~pi0705 & w13650;
assign w13653 = ~w13651 & ~w13652;
assign w13654 = ~w13647 & w13653;
assign w13655 = w13632 & ~w13638;
assign w13656 = w13654 & w13655;
assign w13657 = ~w13646 & ~w13656;
assign w13658 = ~pi3602 & pi9040;
assign w13659 = ~pi3653 & ~pi9040;
assign w13660 = ~w13658 & ~w13659;
assign w13661 = pi0725 & ~w13660;
assign w13662 = ~pi0725 & w13660;
assign w13663 = ~w13661 & ~w13662;
assign w13664 = w13653 & w13663;
assign w13665 = ~w13657 & w13664;
assign w13666 = ~pi3644 & pi9040;
assign w13667 = ~pi3618 & ~pi9040;
assign w13668 = ~w13666 & ~w13667;
assign w13669 = pi0734 & ~w13668;
assign w13670 = ~pi0734 & w13668;
assign w13671 = ~w13669 & ~w13670;
assign w13672 = w13638 & ~w13653;
assign w13673 = w13632 & w13645;
assign w13674 = w13672 & w13673;
assign w13675 = ~w13645 & ~w13672;
assign w13676 = w13639 & w13663;
assign w13677 = ~w13675 & w13676;
assign w13678 = ~w13638 & ~w13653;
assign w13679 = ~w13632 & ~w13663;
assign w13680 = ~w13673 & ~w13679;
assign w13681 = w13678 & ~w13680;
assign w13682 = ~w13638 & ~w13664;
assign w13683 = ~w13639 & ~w13645;
assign w13684 = ~w13682 & w13683;
assign w13685 = ~w13677 & ~w13681;
assign w13686 = ~w13684 & w13685;
assign w13687 = w13645 & w13672;
assign w13688 = ~w13638 & w13653;
assign w13689 = ~w13675 & ~w13688;
assign w13690 = w13632 & w13663;
assign w13691 = ~w13675 & w65102;
assign w13692 = ~w13654 & w13679;
assign w13693 = w13657 & ~w13692;
assign w13694 = w13657 & w65103;
assign w13695 = w13685 & w63669;
assign w13696 = (~w63670 & w65104) | (~w63670 & w65105) | (w65104 & w65105);
assign w13697 = ~w13671 & ~w13694;
assign w13698 = ~w13639 & ~w13655;
assign w13699 = ~w13653 & ~w13698;
assign w13700 = w13638 & w13653;
assign w13701 = w13632 & w13700;
assign w13702 = ~w13699 & ~w13701;
assign w13703 = ~w13645 & ~w13663;
assign w13704 = ~w13702 & w13703;
assign w13705 = ~w13665 & ~w13704;
assign w13706 = ~w13697 & w13705;
assign w13707 = ~w13696 & w13706;
assign w13708 = pi0757 & ~w13707;
assign w13709 = ~pi0757 & w13707;
assign w13710 = ~w13708 & ~w13709;
assign w13711 = ~w13547 & ~w13553;
assign w13712 = ~w13554 & ~w13711;
assign w13713 = w13601 & w13712;
assign w13714 = ~w13608 & ~w13713;
assign w13715 = ~w13586 & w65106;
assign w13716 = ~w13541 & w13560;
assign w13717 = w13600 & w13716;
assign w13718 = w13563 & w13564;
assign w13719 = ~w13717 & ~w13718;
assign w13720 = ~w13571 & ~w13719;
assign w13721 = w13572 & ~w13577;
assign w13722 = w13613 & w13721;
assign w13723 = (w13600 & w13722) | (w13600 & w65107) | (w13722 & w65107);
assign w13724 = ~w13564 & w13577;
assign w13725 = w13612 & ~w13724;
assign w13726 = (~w13725 & w13586) | (~w13725 & w63671) | (w13586 & w63671);
assign w13727 = ~w13565 & ~w13607;
assign w13728 = ~w13547 & ~w13727;
assign w13729 = ~w13582 & ~w13728;
assign w13730 = (~w13600 & w13726) | (~w13600 & w65108) | (w13726 & w65108);
assign w13731 = ~w13720 & ~w13723;
assign w13732 = ~w13715 & w13731;
assign w13733 = ~w13730 & w13732;
assign w13734 = pi0752 & w13733;
assign w13735 = ~pi0752 & ~w13733;
assign w13736 = ~w13734 & ~w13735;
assign w13737 = ~pi3618 & pi9040;
assign w13738 = ~pi3634 & ~pi9040;
assign w13739 = ~w13737 & ~w13738;
assign w13740 = pi0709 & ~w13739;
assign w13741 = ~pi0709 & w13739;
assign w13742 = ~w13740 & ~w13741;
assign w13743 = ~pi3620 & pi9040;
assign w13744 = ~pi3637 & ~pi9040;
assign w13745 = ~w13743 & ~w13744;
assign w13746 = pi0715 & ~w13745;
assign w13747 = ~pi0715 & w13745;
assign w13748 = ~w13746 & ~w13747;
assign w13749 = ~pi3635 & pi9040;
assign w13750 = ~pi3621 & ~pi9040;
assign w13751 = ~w13749 & ~w13750;
assign w13752 = pi0723 & ~w13751;
assign w13753 = ~pi0723 & w13751;
assign w13754 = ~w13752 & ~w13753;
assign w13755 = w13748 & ~w13754;
assign w13756 = ~pi3609 & pi9040;
assign w13757 = ~pi3654 & ~pi9040;
assign w13758 = ~w13756 & ~w13757;
assign w13759 = pi0711 & ~w13758;
assign w13760 = ~pi0711 & w13758;
assign w13761 = ~w13759 & ~w13760;
assign w13762 = w13755 & w13761;
assign w13763 = ~pi3634 & pi9040;
assign w13764 = ~pi3625 & ~pi9040;
assign w13765 = ~w13763 & ~w13764;
assign w13766 = pi0717 & ~w13765;
assign w13767 = ~pi0717 & w13765;
assign w13768 = ~w13766 & ~w13767;
assign w13769 = ~w13748 & ~w13768;
assign w13770 = ~w13748 & w13754;
assign w13771 = w13761 & ~w13768;
assign w13772 = ~w13770 & ~w13771;
assign w13773 = ~w13769 & ~w13772;
assign w13774 = (~w13755 & w13772) | (~w13755 & w65109) | (w13772 & w65109);
assign w13775 = ~pi3633 & pi9040;
assign w13776 = ~pi3627 & ~pi9040;
assign w13777 = ~w13775 & ~w13776;
assign w13778 = pi0718 & ~w13777;
assign w13779 = ~pi0718 & w13777;
assign w13780 = ~w13778 & ~w13779;
assign w13781 = ~w13774 & w13780;
assign w13782 = ~w13754 & ~w13761;
assign w13783 = w13769 & w13782;
assign w13784 = ~w13762 & ~w13783;
assign w13785 = ~w13781 & w13784;
assign w13786 = w13742 & ~w13785;
assign w13787 = ~w13742 & ~w13769;
assign w13788 = w13774 & w13787;
assign w13789 = w13754 & w13769;
assign w13790 = w13761 & w13789;
assign w13791 = w13780 & ~w13790;
assign w13792 = ~w13788 & w13791;
assign w13793 = w13754 & w13761;
assign w13794 = ~w13782 & ~w13793;
assign w13795 = w13748 & w13768;
assign w13796 = ~w13769 & ~w13795;
assign w13797 = ~w13761 & ~w13768;
assign w13798 = w13742 & w13797;
assign w13799 = w13796 & ~w13798;
assign w13800 = w13794 & ~w13799;
assign w13801 = w13742 & ~w13768;
assign w13802 = ~w13794 & ~w13801;
assign w13803 = w13796 & w13802;
assign w13804 = ~w13780 & ~w13800;
assign w13805 = ~w13803 & w13804;
assign w13806 = ~w13792 & ~w13805;
assign w13807 = ~w13786 & ~w13806;
assign w13808 = ~pi0759 & w13807;
assign w13809 = pi0759 & ~w13807;
assign w13810 = ~w13808 & ~w13809;
assign w13811 = w13761 & w13768;
assign w13812 = ~w13754 & w13811;
assign w13813 = ~w13742 & ~w13812;
assign w13814 = ~w13770 & ~w13811;
assign w13815 = w13742 & ~w13814;
assign w13816 = w13742 & ~w13769;
assign w13817 = ~w13798 & ~w13816;
assign w13818 = ~w13815 & w13817;
assign w13819 = w13761 & w13770;
assign w13820 = w13768 & w13819;
assign w13821 = ~w13818 & ~w13820;
assign w13822 = ~w13813 & ~w13821;
assign w13823 = w13754 & ~w13795;
assign w13824 = ~w13754 & w13795;
assign w13825 = ~w13823 & ~w13824;
assign w13826 = ~w13761 & ~w13769;
assign w13827 = w13825 & w13826;
assign w13828 = ~w13748 & ~w13797;
assign w13829 = ~w13742 & ~w13811;
assign w13830 = w13828 & w13829;
assign w13831 = w13748 & ~w13825;
assign w13832 = (~w13798 & w13825) | (~w13798 & w65110) | (w13825 & w65110);
assign w13833 = ~w13772 & ~w13832;
assign w13834 = w13780 & ~w13830;
assign w13835 = ~w13827 & w13834;
assign w13836 = ~w13833 & w13835;
assign w13837 = ~w13742 & ~w13828;
assign w13838 = ~w13831 & w13837;
assign w13839 = w13816 & ~w13825;
assign w13840 = ~w13780 & ~w13783;
assign w13841 = ~w13839 & w13840;
assign w13842 = ~w13838 & w13841;
assign w13843 = ~w13836 & ~w13842;
assign w13844 = ~w13822 & ~w13843;
assign w13845 = ~pi0753 & w13844;
assign w13846 = pi0753 & ~w13844;
assign w13847 = ~w13845 & ~w13846;
assign w13848 = ~pi3599 & pi9040;
assign w13849 = ~pi3631 & ~pi9040;
assign w13850 = ~w13848 & ~w13849;
assign w13851 = pi0712 & ~w13850;
assign w13852 = ~pi0712 & w13850;
assign w13853 = ~w13851 & ~w13852;
assign w13854 = ~pi3610 & pi9040;
assign w13855 = ~pi3636 & ~pi9040;
assign w13856 = ~w13854 & ~w13855;
assign w13857 = pi0729 & ~w13856;
assign w13858 = ~pi0729 & w13856;
assign w13859 = ~w13857 & ~w13858;
assign w13860 = w13853 & ~w13859;
assign w13861 = ~pi3645 & pi9040;
assign w13862 = ~pi3638 & ~pi9040;
assign w13863 = ~w13861 & ~w13862;
assign w13864 = pi0735 & ~w13863;
assign w13865 = ~pi0735 & w13863;
assign w13866 = ~w13864 & ~w13865;
assign w13867 = ~pi3646 & pi9040;
assign w13868 = ~pi3643 & ~pi9040;
assign w13869 = ~w13867 & ~w13868;
assign w13870 = pi0720 & ~w13869;
assign w13871 = ~pi0720 & w13869;
assign w13872 = ~w13870 & ~w13871;
assign w13873 = ~w13866 & w13872;
assign w13874 = w13866 & ~w13872;
assign w13875 = ~w13873 & ~w13874;
assign w13876 = w13860 & w13875;
assign w13877 = ~pi3598 & pi9040;
assign w13878 = ~pi3645 & ~pi9040;
assign w13879 = ~w13877 & ~w13878;
assign w13880 = pi0713 & ~w13879;
assign w13881 = ~pi0713 & w13879;
assign w13882 = ~w13880 & ~w13881;
assign w13883 = ~w13853 & ~w13882;
assign w13884 = w13859 & ~w13873;
assign w13885 = w13883 & w13884;
assign w13886 = ~w13866 & w13882;
assign w13887 = ~w13853 & w13872;
assign w13888 = ~w13860 & ~w13887;
assign w13889 = w13886 & ~w13888;
assign w13890 = w13866 & ~w13882;
assign w13891 = ~w13886 & ~w13890;
assign w13892 = ~w13853 & ~w13872;
assign w13893 = w13859 & w13866;
assign w13894 = w13892 & ~w13893;
assign w13895 = w13891 & w13894;
assign w13896 = w13853 & ~w13872;
assign w13897 = w13882 & w13896;
assign w13898 = ~w13887 & ~w13897;
assign w13899 = w13893 & ~w13898;
assign w13900 = ~pi3641 & pi9040;
assign w13901 = ~pi3598 & ~pi9040;
assign w13902 = ~w13900 & ~w13901;
assign w13903 = pi0703 & ~w13902;
assign w13904 = ~pi0703 & w13902;
assign w13905 = ~w13903 & ~w13904;
assign w13906 = ~w13889 & w13905;
assign w13907 = ~w13895 & w13906;
assign w13908 = ~w13899 & w13907;
assign w13909 = w13853 & w13882;
assign w13910 = w13875 & w13909;
assign w13911 = ~w13853 & w13893;
assign w13912 = ~w13859 & w13886;
assign w13913 = ~w13911 & ~w13912;
assign w13914 = ~w13872 & ~w13913;
assign w13915 = w13866 & w13882;
assign w13916 = ~w13866 & w13883;
assign w13917 = ~w13915 & ~w13916;
assign w13918 = ~w13859 & w13872;
assign w13919 = ~w13917 & w13918;
assign w13920 = w13874 & w13883;
assign w13921 = ~w13905 & ~w13920;
assign w13922 = w13860 & w13890;
assign w13923 = ~w13910 & ~w13922;
assign w13924 = w13921 & w13923;
assign w13925 = ~w13914 & ~w13919;
assign w13926 = w13924 & w13925;
assign w13927 = ~w13908 & ~w13926;
assign w13928 = ~w13883 & ~w13909;
assign w13929 = w13859 & w13873;
assign w13930 = w13928 & w13929;
assign w13931 = ~w13876 & ~w13885;
assign w13932 = ~w13930 & w13931;
assign w13933 = ~w13927 & w13932;
assign w13934 = ~pi0738 & ~w13933;
assign w13935 = pi0738 & w13933;
assign w13936 = ~w13934 & ~w13935;
assign w13937 = w13647 & w13690;
assign w13938 = ~w13632 & w13653;
assign w13939 = ~w13663 & ~w13938;
assign w13940 = ~w13687 & w13939;
assign w13941 = ~w13632 & w13678;
assign w13942 = (w13663 & ~w13700) | (w13663 & w63672) | (~w13700 & w63672);
assign w13943 = ~w13941 & w13942;
assign w13944 = ~w13940 & ~w13943;
assign w13945 = w13678 & w63673;
assign w13946 = w13639 & w63674;
assign w13947 = ~w13945 & ~w13946;
assign w13948 = w13673 & w13678;
assign w13949 = ~w13937 & ~w13948;
assign w13950 = w13947 & w13949;
assign w13951 = ~w13944 & w13950;
assign w13952 = ~w13653 & w13663;
assign w13953 = ~w13647 & w13952;
assign w13954 = (~w13656 & ~w13693) | (~w13656 & w63675) | (~w13693 & w63675);
assign w13955 = ~w13690 & ~w13954;
assign w13956 = w13698 & w63676;
assign w13957 = w13939 & w13956;
assign w13958 = w13956 & w65111;
assign w13959 = w13680 & w13688;
assign w13960 = ~w13698 & w13703;
assign w13961 = ~w13680 & w13700;
assign w13962 = ~w13691 & ~w13961;
assign w13963 = w13698 & ~w13962;
assign w13964 = ~w13959 & ~w13960;
assign w13965 = ~w13958 & w13964;
assign w13966 = ~w13963 & w13965;
assign w13967 = w13671 & ~w13966;
assign w13968 = ~w13645 & w13672;
assign w13969 = ~w13676 & w13968;
assign w13970 = w13663 & w13969;
assign w13971 = (~w13970 & w13951) | (~w13970 & w65112) | (w13951 & w65112);
assign w13972 = ~w13955 & w13971;
assign w13973 = w13972 & w65113;
assign w13974 = (~pi0743 & ~w13972) | (~pi0743 & w65114) | (~w13972 & w65114);
assign w13975 = ~w13973 & ~w13974;
assign w13976 = ~w13152 & ~w13256;
assign w13977 = w13158 & ~w13227;
assign w13978 = ~w13976 & w13977;
assign w13979 = w13159 & w13172;
assign w13980 = w13159 & w13186;
assign w13981 = ~w13171 & w13178;
assign w13982 = ~w13206 & ~w13981;
assign w13983 = w13514 & ~w13982;
assign w13984 = ~w13181 & ~w13247;
assign w13985 = (w13152 & ~w13984) | (w13152 & w65115) | (~w13984 & w65115);
assign w13986 = ~w13193 & ~w13980;
assign w13987 = ~w13235 & w13986;
assign w13988 = ~w13983 & ~w13985;
assign w13989 = w13987 & w13988;
assign w13990 = ~w13165 & w13517;
assign w13991 = w13200 & w13236;
assign w13992 = w13195 & ~w13256;
assign w13993 = w13193 & ~w13990;
assign w13994 = ~w13991 & w13993;
assign w13995 = ~w13992 & w13994;
assign w13996 = ~w13989 & ~w13995;
assign w13997 = ~w13978 & ~w13979;
assign w13998 = ~w13996 & w65116;
assign w13999 = (pi0741 & w13996) | (pi0741 & w65117) | (w13996 & w65117);
assign w14000 = ~w13998 & ~w13999;
assign w14001 = w13299 & ~w13314;
assign w14002 = w13304 & w65118;
assign w14003 = ~w13308 & ~w14002;
assign w14004 = ~w13324 & ~w13343;
assign w14005 = ~w13302 & w14004;
assign w14006 = ~w13331 & ~w13341;
assign w14007 = ~w13285 & w13299;
assign w14008 = ~w14006 & w14007;
assign w14009 = w14003 & ~w14008;
assign w14010 = (w14009 & ~w13317) | (w14009 & w65119) | (~w13317 & w65119);
assign w14011 = ~w14001 & ~w14010;
assign w14012 = w13485 & w13487;
assign w14013 = ~w13326 & ~w14012;
assign w14014 = (w13314 & ~w14013) | (w13314 & w63677) | (~w14013 & w63677);
assign w14015 = ~w13339 & w14001;
assign w14016 = w14003 & w14015;
assign w14017 = w14004 & w14016;
assign w14018 = ~w13301 & w13339;
assign w14019 = w13494 & w14018;
assign w14020 = ~w14014 & ~w14017;
assign w14021 = ~w14019 & w14020;
assign w14022 = (~pi0765 & ~w14021) | (~pi0765 & w65120) | (~w14021 & w65120);
assign w14023 = w14021 & w65121;
assign w14024 = ~w14022 & ~w14023;
assign w14025 = w13698 & w65122;
assign w14026 = (w13939 & ~w13657) | (w13939 & w65123) | (~w13657 & w65123);
assign w14027 = ~w13678 & ~w13946;
assign w14028 = w13943 & ~w14027;
assign w14029 = ~w14025 & ~w14028;
assign w14030 = ~w14026 & w14029;
assign w14031 = w13671 & ~w14030;
assign w14032 = ~w13945 & ~w14025;
assign w14033 = ~w13663 & ~w14032;
assign w14034 = ~w13676 & ~w13947;
assign w14035 = (~w13671 & ~w13686) | (~w13671 & w65124) | (~w13686 & w65124);
assign w14036 = ~w13937 & ~w13970;
assign w14037 = ~w14033 & w14036;
assign w14038 = ~w14035 & w14037;
assign w14039 = ~w14031 & w14038;
assign w14040 = ~pi0763 & w14039;
assign w14041 = pi0763 & ~w14039;
assign w14042 = ~w14040 & ~w14041;
assign w14043 = w13076 & w13103;
assign w14044 = w13103 & w63678;
assign w14045 = ~w13138 & ~w14044;
assign w14046 = ~w13119 & ~w14043;
assign w14047 = w13128 & ~w14046;
assign w14048 = ~w13118 & ~w13136;
assign w14049 = ~w13091 & ~w13119;
assign w14050 = ~w14048 & w14049;
assign w14051 = ~w14047 & ~w14050;
assign w14052 = ~w14045 & w14051;
assign w14053 = ~w13093 & ~w13103;
assign w14054 = w13076 & w14053;
assign w14055 = (w13091 & w14054) | (w13091 & w65125) | (w14054 & w65125);
assign w14056 = ~w13096 & ~w13126;
assign w14057 = w13076 & w13094;
assign w14058 = w13067 & w13101;
assign w14059 = ~w14057 & ~w14058;
assign w14060 = ~w13091 & ~w14059;
assign w14061 = (w13111 & w14056) | (w13111 & w65126) | (w14056 & w65126);
assign w14062 = ~w14055 & w14061;
assign w14063 = ~w14060 & w14062;
assign w14064 = w13070 & w65127;
assign w14065 = ~w13070 & w13076;
assign w14066 = (~w13091 & w14065) | (~w13091 & w14171) | (w14065 & w14171);
assign w14067 = ~w13124 & ~w14044;
assign w14068 = ~w14066 & w14067;
assign w14069 = ~w13096 & ~w13113;
assign w14070 = ~w14053 & w14069;
assign w14071 = w14046 & w14070;
assign w14072 = ~w13111 & ~w14064;
assign w14073 = ~w14071 & w14072;
assign w14074 = w14068 & w14073;
assign w14075 = ~w14063 & ~w14074;
assign w14076 = ~w14052 & ~w14075;
assign w14077 = ~pi0744 & w14076;
assign w14078 = pi0744 & ~w14076;
assign w14079 = ~w14077 & ~w14078;
assign w14080 = ~w13374 & w65128;
assign w14081 = ~w13397 & ~w14080;
assign w14082 = ~w13403 & ~w14081;
assign w14083 = ~w13401 & w13429;
assign w14084 = ~w14080 & w14083;
assign w14085 = ~w13441 & w14084;
assign w14086 = w13414 & ~w14085;
assign w14087 = w13404 & w13436;
assign w14088 = (~w13358 & w13426) | (~w13358 & w65129) | (w13426 & w65129);
assign w14089 = ~w14087 & ~w14088;
assign w14090 = w13371 & ~w13399;
assign w14091 = ~w14089 & w14090;
assign w14092 = w13414 & ~w14091;
assign w14093 = ~w13438 & w14089;
assign w14094 = ~w14092 & ~w14093;
assign w14095 = ~w14082 & ~w14086;
assign w14096 = (pi0755 & ~w14095) | (pi0755 & w65130) | (~w14095 & w65130);
assign w14097 = w14095 & w65131;
assign w14098 = ~w14096 & ~w14097;
assign w14099 = ~w13761 & ~w13770;
assign w14100 = w13796 & w14099;
assign w14101 = w13802 & w14100;
assign w14102 = w13782 & ~w13796;
assign w14103 = ~w13742 & ~w13796;
assign w14104 = ~w14102 & ~w14103;
assign w14105 = ~w13773 & ~w14102;
assign w14106 = w13742 & ~w14105;
assign w14107 = w13812 & ~w14103;
assign w14108 = ~w13801 & w14105;
assign w14109 = ~w14107 & w14108;
assign w14110 = (~w14104 & w14109) | (~w14104 & w63375) | (w14109 & w63375);
assign w14111 = ~w13771 & ~w13793;
assign w14112 = w13816 & ~w14111;
assign w14113 = ~w14101 & ~w14112;
assign w14114 = (w13780 & w14110) | (w13780 & w63679) | (w14110 & w63679);
assign w14115 = ~w13754 & ~w13768;
assign w14116 = w13742 & w14100;
assign w14117 = ~w14115 & w14116;
assign w14118 = ~w14109 & w63680;
assign w14119 = w13788 & w13793;
assign w14120 = ~w14117 & ~w14119;
assign w14121 = ~w14118 & w14120;
assign w14122 = ~w14114 & w14121;
assign w14123 = pi0761 & w14122;
assign w14124 = ~pi0761 & ~w14122;
assign w14125 = ~w14123 & ~w14124;
assign w14126 = w13795 & w14107;
assign w14127 = ~w13742 & w13819;
assign w14128 = w13815 & ~w13819;
assign w14129 = ~w13754 & ~w14105;
assign w14130 = ~w13742 & ~w14115;
assign w14131 = w13814 & w14130;
assign w14132 = ~w13780 & ~w14131;
assign w14133 = ~w14128 & w14132;
assign w14134 = ~w14129 & w14133;
assign w14135 = w13761 & w13823;
assign w14136 = ~w13789 & w13829;
assign w14137 = w13817 & ~w14136;
assign w14138 = w13780 & ~w14135;
assign w14139 = ~w14116 & w14138;
assign w14140 = ~w14137 & w14139;
assign w14141 = ~w14134 & ~w14140;
assign w14142 = ~w14126 & ~w14127;
assign w14143 = ~w14141 & w14142;
assign w14144 = ~pi0769 & w14143;
assign w14145 = pi0769 & ~w14143;
assign w14146 = ~w14144 & ~w14145;
assign w14147 = ~w13571 & w13713;
assign w14148 = ~w13712 & ~w13716;
assign w14149 = w13603 & w14148;
assign w14150 = w13712 & w13716;
assign w14151 = ~w13718 & ~w14150;
assign w14152 = ~w14149 & w14151;
assign w14153 = ~w13585 & w14152;
assign w14154 = w13600 & ~w14153;
assign w14155 = ~w14148 & ~w14150;
assign w14156 = ~w13571 & ~w14155;
assign w14157 = (~w13600 & w13581) | (~w13600 & w65132) | (w13581 & w65132);
assign w14158 = w13575 & ~w13591;
assign w14159 = ~w13590 & w14158;
assign w14160 = (~w14147 & w14156) | (~w14147 & w65133) | (w14156 & w65133);
assign w14161 = ~w14154 & w14160;
assign w14162 = (pi0754 & ~w14161) | (pi0754 & w65134) | (~w14161 & w65134);
assign w14163 = w14161 & w65135;
assign w14164 = ~w14162 & ~w14163;
assign w14165 = ~w13114 & w13135;
assign w14166 = ~w13093 & w13111;
assign w14167 = w13125 & ~w14166;
assign w14168 = w14165 & w14167;
assign w14169 = ~w13091 & ~w13121;
assign w14170 = w13100 & ~w14069;
assign w14171 = w13118 & w63681;
assign w14172 = ~w13111 & ~w14170;
assign w14173 = ~w14171 & w14172;
assign w14174 = ~w13135 & w14053;
assign w14175 = ~w13095 & w13111;
assign w14176 = ~w14174 & w14175;
assign w14177 = w14051 & w14176;
assign w14178 = ~w14173 & ~w14177;
assign w14179 = ~w13115 & ~w14168;
assign w14180 = ~w14169 & w14179;
assign w14181 = ~w14178 & w14180;
assign w14182 = pi0758 & ~w14181;
assign w14183 = ~pi0758 & w14181;
assign w14184 = ~w14182 & ~w14183;
assign w14185 = w13374 & w13425;
assign w14186 = ~w13462 & ~w14185;
assign w14187 = ~w13390 & w14186;
assign w14188 = w13414 & ~w14187;
assign w14189 = w13415 & ~w13463;
assign w14190 = w13371 & ~w13461;
assign w14191 = ~w13402 & ~w13417;
assign w14192 = ~w14190 & w14191;
assign w14193 = ~w13433 & ~w14192;
assign w14194 = ~w14189 & ~w14193;
assign w14195 = w13364 & ~w13414;
assign w14196 = ~w13374 & w14195;
assign w14197 = ~w13462 & w14196;
assign w14198 = ~w14194 & ~w14197;
assign w14199 = ~w14188 & w14198;
assign w14200 = pi0747 & ~w14199;
assign w14201 = ~pi0747 & w14199;
assign w14202 = ~w14200 & ~w14201;
assign w14203 = ~w13299 & ~w13489;
assign w14204 = ~w13328 & ~w14203;
assign w14205 = w13307 & w13321;
assign w14206 = ~w13343 & ~w13503;
assign w14207 = ~w14205 & w14206;
assign w14208 = w13316 & w14207;
assign w14209 = ~w13342 & w13498;
assign w14210 = w13321 & ~w13340;
assign w14211 = ~w14209 & ~w14210;
assign w14212 = ~w13303 & w13314;
assign w14213 = ~w14211 & w14212;
assign w14214 = ~w14208 & ~w14213;
assign w14215 = ~w14204 & ~w14214;
assign w14216 = ~pi0768 & w14215;
assign w14217 = pi0768 & ~w14215;
assign w14218 = ~w14216 & ~w14217;
assign w14219 = w13873 & w13883;
assign w14220 = w13853 & w13872;
assign w14221 = (~w13859 & ~w14220) | (~w13859 & w65136) | (~w14220 & w65136);
assign w14222 = w13886 & ~w13896;
assign w14223 = ~w14221 & w14222;
assign w14224 = ~w13891 & ~w14220;
assign w14225 = ~w13873 & ~w14220;
assign w14226 = w13891 & ~w14225;
assign w14227 = ~w14224 & ~w14226;
assign w14228 = w13872 & w14227;
assign w14229 = w14227 & w13918;
assign w14230 = ~w13896 & ~w13915;
assign w14231 = ~w13866 & ~w13882;
assign w14232 = ~w13892 & ~w14231;
assign w14233 = w13887 & w13915;
assign w14234 = (~w14233 & ~w13917) | (~w14233 & w65137) | (~w13917 & w65137);
assign w14235 = ~w14230 & ~w14234;
assign w14236 = ~w13859 & ~w13928;
assign w14237 = w13921 & ~w14219;
assign w14238 = w14237 & w65138;
assign w14239 = ~w14229 & w14238;
assign w14240 = ~w14235 & w14239;
assign w14241 = ~w13875 & w13891;
assign w14242 = w13928 & w14241;
assign w14243 = w13872 & w13890;
assign w14244 = ~w13897 & ~w13916;
assign w14245 = ~w14243 & w14244;
assign w14246 = w14224 & ~w14245;
assign w14247 = ~w13885 & ~w13893;
assign w14248 = w13913 & ~w14247;
assign w14249 = w13886 & w13887;
assign w14250 = ~w13859 & w14249;
assign w14251 = w13905 & ~w14250;
assign w14252 = ~w14242 & w14251;
assign w14253 = ~w14246 & w14252;
assign w14254 = ~w14248 & w14253;
assign w14255 = ~w14240 & ~w14254;
assign w14256 = ~pi0737 & w14255;
assign w14257 = pi0737 & ~w14255;
assign w14258 = ~w14256 & ~w14257;
assign w14259 = w13091 & ~w13137;
assign w14260 = w13136 & w14165;
assign w14261 = w13134 & ~w14260;
assign w14262 = ~w14259 & ~w14261;
assign w14263 = ~w13113 & ~w14058;
assign w14264 = ~w13083 & ~w14263;
assign w14265 = ~w13097 & ~w13103;
assign w14266 = ~w13114 & w14265;
assign w14267 = w13091 & ~w14266;
assign w14268 = ~w13111 & ~w14264;
assign w14269 = ~w14267 & w14268;
assign w14270 = w13096 & w13098;
assign w14271 = w13111 & ~w13120;
assign w14272 = ~w14270 & w14271;
assign w14273 = (w14068 & w65139) | (w14068 & w65140) | (w65139 & w65140);
assign w14274 = ~w14269 & ~w14273;
assign w14275 = ~w14262 & ~w14274;
assign w14276 = ~pi0751 & w14275;
assign w14277 = pi0751 & ~w14275;
assign w14278 = ~w14276 & ~w14277;
assign w14279 = ~w13961 & ~w13969;
assign w14280 = (~w13671 & ~w13954) | (~w13671 & w65141) | (~w13954 & w65141);
assign w14281 = w13632 & ~w13663;
assign w14282 = (w14281 & w13675) | (w14281 & w65142) | (w13675 & w65142);
assign w14283 = ~w13956 & ~w14282;
assign w14284 = w13671 & ~w14283;
assign w14285 = ~w13646 & ~w13938;
assign w14286 = w13671 & ~w14285;
assign w14287 = ~w13948 & ~w14025;
assign w14288 = ~w14286 & w14287;
assign w14289 = w13663 & ~w14288;
assign w14290 = ~w13957 & ~w14284;
assign w14291 = ~w14289 & w14290;
assign w14292 = ~w14280 & w14291;
assign w14293 = ~pi0764 & w14292;
assign w14294 = pi0764 & ~w14292;
assign w14295 = ~w14293 & ~w14294;
assign w14296 = w13578 & w13579;
assign w14297 = ~w13586 & ~w14296;
assign w14298 = w13581 & w13613;
assign w14299 = w13563 & w13573;
assign w14300 = ~w13571 & ~w14299;
assign w14301 = ~w14298 & w14300;
assign w14302 = ~w14297 & ~w14301;
assign w14303 = ~w13588 & w13602;
assign w14304 = ~w13562 & w14303;
assign w14305 = ~w13600 & ~w14304;
assign w14306 = w13590 & w14305;
assign w14307 = ~w13572 & ~w13712;
assign w14308 = w13605 & w14307;
assign w14309 = w13580 & w13721;
assign w14310 = ~w13562 & w13600;
assign w14311 = ~w14309 & w14310;
assign w14312 = ~w14308 & w14311;
assign w14313 = ~w14306 & ~w14312;
assign w14314 = ~w14313 & w65143;
assign w14315 = (pi0770 & w14313) | (pi0770 & w65144) | (w14313 & w65144);
assign w14316 = ~w14314 & ~w14315;
assign w14317 = ~w13872 & ~w13883;
assign w14318 = w13891 & w14317;
assign w14319 = w13859 & ~w14318;
assign w14320 = w13853 & ~w13891;
assign w14321 = w13875 & w14230;
assign w14322 = w14221 & ~w14320;
assign w14323 = ~w14321 & w14322;
assign w14324 = ~w14319 & ~w14323;
assign w14325 = (w13905 & w14324) | (w13905 & w65145) | (w14324 & w65145);
assign w14326 = w13859 & ~w14227;
assign w14327 = ~w13859 & w14318;
assign w14328 = (~w13905 & w14326) | (~w13905 & w65146) | (w14326 & w65146);
assign w14329 = ~w13859 & w13905;
assign w14330 = w14219 & ~w14329;
assign w14331 = ~w14229 & ~w14330;
assign w14332 = ~w14328 & w14331;
assign w14333 = ~w14325 & w14332;
assign w14334 = pi0760 & ~w14333;
assign w14335 = ~pi0760 & w14333;
assign w14336 = ~w14334 & ~w14335;
assign w14337 = w13859 & ~w14249;
assign w14338 = w13866 & w13897;
assign w14339 = w14221 & ~w14338;
assign w14340 = ~w14337 & ~w14339;
assign w14341 = w13890 & w14220;
assign w14342 = ~w13859 & ~w14234;
assign w14343 = (w13859 & ~w14244) | (w13859 & w65147) | (~w14244 & w65147);
assign w14344 = w13905 & ~w14341;
assign w14345 = ~w14343 & w14344;
assign w14346 = ~w14342 & w14345;
assign w14347 = ~w13859 & w13920;
assign w14348 = ~w13872 & w13890;
assign w14349 = (~w13883 & w14226) | (~w13883 & w63683) | (w14226 & w63683);
assign w14350 = ~w14236 & ~w14348;
assign w14351 = ~w14349 & w14350;
assign w14352 = ~w13905 & ~w14249;
assign w14353 = (w14352 & w14351) | (w14352 & w65148) | (w14351 & w65148);
assign w14354 = ~w14346 & ~w14353;
assign w14355 = ~w14340 & ~w14354;
assign w14356 = ~pi0767 & w14355;
assign w14357 = pi0767 & ~w14355;
assign w14358 = ~w14356 & ~w14357;
assign w14359 = ~pi3672 & pi9040;
assign w14360 = ~pi3702 & ~pi9040;
assign w14361 = ~w14359 & ~w14360;
assign w14362 = pi0798 & ~w14361;
assign w14363 = ~pi0798 & w14361;
assign w14364 = ~w14362 & ~w14363;
assign w14365 = ~pi3657 & pi9040;
assign w14366 = ~pi3658 & ~pi9040;
assign w14367 = ~w14365 & ~w14366;
assign w14368 = pi0795 & ~w14367;
assign w14369 = ~pi0795 & w14367;
assign w14370 = ~w14368 & ~w14369;
assign w14371 = ~w14364 & ~w14370;
assign w14372 = w14364 & w14370;
assign w14373 = ~w14371 & ~w14372;
assign w14374 = ~pi3690 & pi9040;
assign w14375 = ~pi3684 & ~pi9040;
assign w14376 = ~w14374 & ~w14375;
assign w14377 = pi0774 & ~w14376;
assign w14378 = ~pi0774 & w14376;
assign w14379 = ~w14377 & ~w14378;
assign w14380 = ~pi3701 & pi9040;
assign w14381 = ~pi3668 & ~pi9040;
assign w14382 = ~w14380 & ~w14381;
assign w14383 = pi0766 & ~w14382;
assign w14384 = ~pi0766 & w14382;
assign w14385 = ~w14383 & ~w14384;
assign w14386 = w14379 & w14385;
assign w14387 = ~w14373 & w14386;
assign w14388 = ~w14370 & w14385;
assign w14389 = ~w14364 & w14379;
assign w14390 = ~w14388 & ~w14389;
assign w14391 = ~w14387 & ~w14390;
assign w14392 = w14370 & ~w14385;
assign w14393 = ~w14372 & ~w14392;
assign w14394 = ~w14379 & w14385;
assign w14395 = w14364 & w14394;
assign w14396 = w14393 & ~w14395;
assign w14397 = w14391 & ~w14396;
assign w14398 = ~w14379 & ~w14385;
assign w14399 = ~w14373 & w14398;
assign w14400 = ~w14397 & ~w14399;
assign w14401 = ~pi3677 & pi9040;
assign w14402 = ~pi3682 & ~pi9040;
assign w14403 = ~w14401 & ~w14402;
assign w14404 = pi0771 & ~w14403;
assign w14405 = ~pi0771 & w14403;
assign w14406 = ~w14404 & ~w14405;
assign w14407 = ~w14400 & w14406;
assign w14408 = ~pi3668 & pi9040;
assign w14409 = ~pi3705 & ~pi9040;
assign w14410 = ~w14408 & ~w14409;
assign w14411 = pi0796 & ~w14410;
assign w14412 = ~pi0796 & w14410;
assign w14413 = ~w14411 & ~w14412;
assign w14414 = ~w14370 & w14379;
assign w14415 = ~w14371 & ~w14406;
assign w14416 = ~w14392 & ~w14414;
assign w14417 = w14415 & w14416;
assign w14418 = w14389 & ~w14406;
assign w14419 = ~w14370 & ~w14385;
assign w14420 = w14364 & w14419;
assign w14421 = w14419 & w65149;
assign w14422 = w14370 & w14398;
assign w14423 = ~w14421 & ~w14422;
assign w14424 = w14406 & ~w14423;
assign w14425 = ~w14413 & ~w14418;
assign w14426 = ~w14387 & w14425;
assign w14427 = ~w14417 & w14426;
assign w14428 = ~w14424 & w14427;
assign w14429 = w14379 & ~w14406;
assign w14430 = w14371 & w14385;
assign w14431 = w14429 & w14430;
assign w14432 = w14379 & ~w14385;
assign w14433 = w14364 & w14432;
assign w14434 = ~w14406 & ~w14433;
assign w14435 = ~w14364 & w14398;
assign w14436 = w14434 & ~w14435;
assign w14437 = (w14406 & w14387) | (w14406 & w65150) | (w14387 & w65150);
assign w14438 = ~w14436 & ~w14437;
assign w14439 = w14394 & w14372;
assign w14440 = w14413 & ~w14439;
assign w14441 = ~w14431 & w14440;
assign w14442 = ~w14438 & w14441;
assign w14443 = ~w14428 & ~w14442;
assign w14444 = ~w14407 & ~w14443;
assign w14445 = ~pi0800 & w14444;
assign w14446 = pi0800 & ~w14444;
assign w14447 = ~w14445 & ~w14446;
assign w14448 = ~pi3660 & pi9040;
assign w14449 = ~pi3656 & ~pi9040;
assign w14450 = ~w14448 & ~w14449;
assign w14451 = pi0790 & ~w14450;
assign w14452 = ~pi0790 & w14450;
assign w14453 = ~w14451 & ~w14452;
assign w14454 = ~pi3656 & pi9040;
assign w14455 = ~pi3661 & ~pi9040;
assign w14456 = ~w14454 & ~w14455;
assign w14457 = pi0782 & ~w14456;
assign w14458 = ~pi0782 & w14456;
assign w14459 = ~w14457 & ~w14458;
assign w14460 = ~pi3673 & pi9040;
assign w14461 = ~pi3678 & ~pi9040;
assign w14462 = ~w14460 & ~w14461;
assign w14463 = pi0745 & ~w14462;
assign w14464 = ~pi0745 & w14462;
assign w14465 = ~w14463 & ~w14464;
assign w14466 = ~pi3696 & pi9040;
assign w14467 = ~pi3686 & ~pi9040;
assign w14468 = ~w14466 & ~w14467;
assign w14469 = pi0791 & ~w14468;
assign w14470 = ~pi0791 & w14468;
assign w14471 = ~w14469 & ~w14470;
assign w14472 = ~w14465 & w14471;
assign w14473 = ~pi3678 & pi9040;
assign w14474 = ~pi3669 & ~pi9040;
assign w14475 = ~w14473 & ~w14474;
assign w14476 = pi0789 & ~w14475;
assign w14477 = ~pi0789 & w14475;
assign w14478 = ~w14476 & ~w14477;
assign w14479 = ~w14471 & w14478;
assign w14480 = ~w14472 & ~w14479;
assign w14481 = ~w14465 & ~w14471;
assign w14482 = ~pi3752 & pi9040;
assign w14483 = ~pi3692 & ~pi9040;
assign w14484 = ~w14482 & ~w14483;
assign w14485 = pi0781 & ~w14484;
assign w14486 = ~pi0781 & w14484;
assign w14487 = ~w14485 & ~w14486;
assign w14488 = ~w14465 & ~w14487;
assign w14489 = w14471 & ~w14488;
assign w14490 = ~w14481 & ~w14489;
assign w14491 = ~w14480 & ~w14490;
assign w14492 = ~w14472 & ~w14487;
assign w14493 = ~w14459 & ~w14492;
assign w14494 = ~w14491 & w14493;
assign w14495 = ~w14471 & w14487;
assign w14496 = w14465 & w14478;
assign w14497 = w14495 & w14496;
assign w14498 = w14478 & w14488;
assign w14499 = ~w14497 & ~w14498;
assign w14500 = ~w14494 & w14499;
assign w14501 = ~w14453 & ~w14500;
assign w14502 = w14453 & ~w14479;
assign w14503 = w14492 & w14502;
assign w14504 = ~w14459 & ~w14497;
assign w14505 = w14471 & ~w14487;
assign w14506 = ~w14495 & ~w14505;
assign w14507 = ~w14465 & w14478;
assign w14508 = w14506 & w14507;
assign w14509 = ~w14503 & w14504;
assign w14510 = ~w14508 & w14509;
assign w14511 = ~w14478 & w14487;
assign w14512 = ~w14453 & ~w14472;
assign w14513 = w14511 & ~w14512;
assign w14514 = w14505 & w14507;
assign w14515 = ~w14453 & ~w14487;
assign w14516 = w14480 & w14515;
assign w14517 = w14496 & w14506;
assign w14518 = w14465 & ~w14478;
assign w14519 = w14487 & w14518;
assign w14520 = w14518 & w15330;
assign w14521 = w14481 & w14487;
assign w14522 = ~w14520 & ~w14521;
assign w14523 = ~w14517 & w14522;
assign w14524 = w14453 & ~w14523;
assign w14525 = w14459 & ~w14514;
assign w14526 = ~w14513 & w14525;
assign w14527 = ~w14516 & w14526;
assign w14528 = ~w14524 & w14527;
assign w14529 = ~w14510 & ~w14528;
assign w14530 = ~w14501 & ~w14529;
assign w14531 = ~pi0804 & w14530;
assign w14532 = pi0804 & ~w14530;
assign w14533 = ~w14531 & ~w14532;
assign w14534 = ~pi3699 & pi9040;
assign w14535 = ~pi3708 & ~pi9040;
assign w14536 = ~w14534 & ~w14535;
assign w14537 = pi0799 & ~w14536;
assign w14538 = ~pi0799 & w14536;
assign w14539 = ~w14537 & ~w14538;
assign w14540 = ~pi3680 & pi9040;
assign w14541 = ~pi3665 & ~pi9040;
assign w14542 = ~w14540 & ~w14541;
assign w14543 = pi0795 & ~w14542;
assign w14544 = ~pi0795 & w14542;
assign w14545 = ~w14543 & ~w14544;
assign w14546 = ~w14539 & w14545;
assign w14547 = ~pi3703 & pi9040;
assign w14548 = ~pi3683 & ~pi9040;
assign w14549 = ~w14547 & ~w14548;
assign w14550 = pi0745 & ~w14549;
assign w14551 = ~pi0745 & w14549;
assign w14552 = ~w14550 & ~w14551;
assign w14553 = ~pi3697 & pi9040;
assign w14554 = ~pi3755 & ~pi9040;
assign w14555 = ~w14553 & ~w14554;
assign w14556 = pi0796 & ~w14555;
assign w14557 = ~pi0796 & w14555;
assign w14558 = ~w14556 & ~w14557;
assign w14559 = ~w14552 & w14558;
assign w14560 = w14552 & ~w14558;
assign w14561 = ~w14559 & ~w14560;
assign w14562 = ~pi3708 & pi9040;
assign w14563 = ~pi3679 & ~pi9040;
assign w14564 = ~w14562 & ~w14563;
assign w14565 = pi0779 & ~w14564;
assign w14566 = ~pi0779 & w14564;
assign w14567 = ~w14565 & ~w14566;
assign w14568 = w14545 & ~w14552;
assign w14569 = (~w14567 & ~w14568) | (~w14567 & w63324) | (~w14568 & w63324);
assign w14570 = ~w14561 & w14569;
assign w14571 = ~w14546 & ~w14570;
assign w14572 = ~w14561 & w14567;
assign w14573 = ~w14561 & w63684;
assign w14574 = ~w14539 & w14559;
assign w14575 = ~w14573 & ~w14574;
assign w14576 = w14571 & ~w14575;
assign w14577 = w14558 & ~w14567;
assign w14578 = w14545 & w14577;
assign w14579 = ~w14545 & w14552;
assign w14580 = ~w14568 & ~w14579;
assign w14581 = ~w14539 & ~w14558;
assign w14582 = ~w14574 & ~w14581;
assign w14583 = w14582 & w63685;
assign w14584 = w14569 & ~w14583;
assign w14585 = w14539 & w14558;
assign w14586 = (~w14581 & w14570) | (~w14581 & w63376) | (w14570 & w63376);
assign w14587 = ~w14539 & w14558;
assign w14588 = ~w14552 & w14567;
assign w14589 = ~w14579 & ~w14588;
assign w14590 = ~w14546 & ~w14559;
assign w14591 = ~w14587 & w14590;
assign w14592 = ~w14589 & w14591;
assign w14593 = ~w14586 & ~w14592;
assign w14594 = ~w14585 & ~w14593;
assign w14595 = (~w14576 & w14594) | (~w14576 & w63686) | (w14594 & w63686);
assign w14596 = ~pi3755 & pi9040;
assign w14597 = ~pi3662 & ~pi9040;
assign w14598 = ~w14596 & ~w14597;
assign w14599 = pi0781 & ~w14598;
assign w14600 = ~pi0781 & w14598;
assign w14601 = ~w14599 & ~w14600;
assign w14602 = ~w14595 & ~w14601;
assign w14603 = ~w14539 & w14583;
assign w14604 = ~w14545 & ~w14567;
assign w14605 = w14585 & w14604;
assign w14606 = ~w14552 & ~w14567;
assign w14607 = w14546 & w14606;
assign w14608 = ~w14605 & ~w14607;
assign w14609 = ~w14593 & w14601;
assign w14610 = ~w14545 & w14567;
assign w14611 = ~w14580 & w14581;
assign w14612 = ~w14558 & ~w14604;
assign w14613 = w14582 & w63687;
assign w14614 = ~w14611 & ~w14613;
assign w14615 = (w14610 & w14613) | (w14610 & w65151) | (w14613 & w65151);
assign w14616 = (w14608 & ~w14583) | (w14608 & w65152) | (~w14583 & w65152);
assign w14617 = ~w14615 & w14616;
assign w14618 = ~w14609 & w14617;
assign w14619 = ~w14602 & w65153;
assign w14620 = (pi0811 & w14602) | (pi0811 & w65154) | (w14602 & w65154);
assign w14621 = ~w14619 & ~w14620;
assign w14622 = w14539 & w14545;
assign w14623 = ~w14593 & w14622;
assign w14624 = ~w14539 & ~w14577;
assign w14625 = ~w14612 & w14624;
assign w14626 = w14577 & w14579;
assign w14627 = ~w14612 & ~w14626;
assign w14628 = w14539 & ~w14627;
assign w14629 = ~w14569 & w14589;
assign w14630 = w14601 & ~w14625;
assign w14631 = ~w14628 & w14630;
assign w14632 = ~w14629 & w14631;
assign w14633 = w14545 & ~w14606;
assign w14634 = ~w14539 & w14561;
assign w14635 = ~w14633 & w14634;
assign w14636 = w14580 & ~w14585;
assign w14637 = ~w14572 & ~w14580;
assign w14638 = ~w14636 & ~w14637;
assign w14639 = ~w14601 & ~w14635;
assign w14640 = ~w14638 & w14639;
assign w14641 = ~w14632 & ~w14640;
assign w14642 = ~w14623 & ~w14641;
assign w14643 = pi0818 & w14642;
assign w14644 = ~pi0818 & ~w14642;
assign w14645 = ~w14643 & ~w14644;
assign w14646 = w14478 & ~w14487;
assign w14647 = ~w14453 & ~w14465;
assign w14648 = ~w14646 & ~w14647;
assign w14649 = w14471 & ~w14507;
assign w14650 = ~w14648 & w14649;
assign w14651 = w14515 & w14650;
assign w14652 = w14478 & ~w14647;
assign w14653 = w14490 & ~w14652;
assign w14654 = w14453 & w14465;
assign w14655 = ~w14646 & w14654;
assign w14656 = w14506 & ~w14511;
assign w14657 = ~w14453 & ~w14480;
assign w14658 = w14656 & w14657;
assign w14659 = ~w14655 & ~w14658;
assign w14660 = ~w14511 & ~w14515;
assign w14661 = ~w14481 & ~w14646;
assign w14662 = ~w14488 & w14661;
assign w14663 = w14656 & w14662;
assign w14664 = w14453 & ~w14663;
assign w14665 = ~w14658 & w63688;
assign w14666 = ~w14664 & w14665;
assign w14667 = ~w14650 & ~w14653;
assign w14668 = (~w14459 & w14666) | (~w14459 & w65155) | (w14666 & w65155);
assign w14669 = w14481 & w14646;
assign w14670 = ~w14519 & ~w14669;
assign w14671 = w14453 & ~w14670;
assign w14672 = w14481 & ~w14660;
assign w14673 = ~w14520 & ~w14672;
assign w14674 = (w14459 & ~w14659) | (w14459 & w65156) | (~w14659 & w65156);
assign w14675 = ~w14651 & ~w14671;
assign w14676 = ~w14674 & w14675;
assign w14677 = ~w14668 & w14676;
assign w14678 = pi0813 & ~w14677;
assign w14679 = ~pi0813 & w14677;
assign w14680 = ~w14678 & ~w14679;
assign w14681 = ~pi3689 & pi9040;
assign w14682 = pi3675 & ~pi9040;
assign w14683 = ~w14681 & ~w14682;
assign w14684 = pi0774 & ~w14683;
assign w14685 = ~pi0774 & w14683;
assign w14686 = ~w14684 & ~w14685;
assign w14687 = ~pi3705 & pi9040;
assign w14688 = ~pi3664 & ~pi9040;
assign w14689 = ~w14687 & ~w14688;
assign w14690 = pi0792 & ~w14689;
assign w14691 = ~pi0792 & w14689;
assign w14692 = ~w14690 & ~w14691;
assign w14693 = ~pi3695 & pi9040;
assign w14694 = ~pi3671 & ~pi9040;
assign w14695 = ~w14693 & ~w14694;
assign w14696 = pi0787 & ~w14695;
assign w14697 = ~pi0787 & w14695;
assign w14698 = ~w14696 & ~w14697;
assign w14699 = ~w14692 & w14698;
assign w14700 = w14692 & ~w14698;
assign w14701 = ~w14699 & ~w14700;
assign w14702 = ~pi3706 & pi9040;
assign w14703 = ~pi3681 & ~pi9040;
assign w14704 = ~w14702 & ~w14703;
assign w14705 = pi0788 & ~w14704;
assign w14706 = ~pi0788 & w14704;
assign w14707 = ~w14705 & ~w14706;
assign w14708 = ~pi3675 & pi9040;
assign w14709 = ~pi3677 & ~pi9040;
assign w14710 = ~w14708 & ~w14709;
assign w14711 = pi0786 & ~w14710;
assign w14712 = ~pi0786 & w14710;
assign w14713 = ~w14711 & ~w14712;
assign w14714 = w14707 & ~w14713;
assign w14715 = ~pi3670 & pi9040;
assign w14716 = ~pi3663 & ~pi9040;
assign w14717 = ~w14715 & ~w14716;
assign w14718 = pi0766 & ~w14717;
assign w14719 = ~pi0766 & w14717;
assign w14720 = ~w14718 & ~w14719;
assign w14721 = ~w14714 & w14720;
assign w14722 = w14701 & w14721;
assign w14723 = w14713 & ~w14720;
assign w14724 = (~w14707 & ~w14723) | (~w14707 & w63689) | (~w14723 & w63689);
assign w14725 = ~w14713 & ~w14720;
assign w14726 = w14699 & w14725;
assign w14727 = ~w14723 & ~w14726;
assign w14728 = w14724 & ~w14727;
assign w14729 = ~w14714 & ~w14725;
assign w14730 = w14700 & ~w14729;
assign w14731 = ~w14722 & ~w14730;
assign w14732 = ~w14728 & w14731;
assign w14733 = w14686 & ~w14732;
assign w14734 = w14700 & w14720;
assign w14735 = (~w14713 & ~w14700) | (~w14713 & w14725) | (~w14700 & w14725);
assign w14736 = w14692 & w14713;
assign w14737 = w14724 & ~w14736;
assign w14738 = ~w14735 & w14737;
assign w14739 = ~w14713 & w14720;
assign w14740 = w14699 & w14739;
assign w14741 = ~w14692 & ~w14720;
assign w14742 = ~w14698 & ~w14713;
assign w14743 = w14741 & w14742;
assign w14744 = ~w14698 & w14713;
assign w14745 = w14741 & w14744;
assign w14746 = ~w14734 & ~w14745;
assign w14747 = w14707 & ~w14746;
assign w14748 = (~w14714 & w14746) | (~w14714 & w65157) | (w14746 & w65157);
assign w14749 = w14692 & w14732;
assign w14750 = ~w14740 & ~w14743;
assign w14751 = ~w14738 & w14750;
assign w14752 = (w14751 & ~w14749) | (w14751 & w63690) | (~w14749 & w63690);
assign w14753 = ~w14686 & ~w14752;
assign w14754 = ~w14707 & ~w14713;
assign w14755 = ~w14701 & ~w14707;
assign w14756 = w14707 & ~w14740;
assign w14757 = ~w14699 & w14725;
assign w14758 = w14699 & w14723;
assign w14759 = ~w14757 & ~w14758;
assign w14760 = w14756 & w14759;
assign w14761 = ~w14754 & ~w14755;
assign w14762 = ~w14760 & w14761;
assign w14763 = ~w14733 & ~w14762;
assign w14764 = ~w14753 & w65158;
assign w14765 = (pi0805 & w14753) | (pi0805 & w65159) | (w14753 & w65159);
assign w14766 = ~w14764 & ~w14765;
assign w14767 = ~pi3674 & pi9040;
assign w14768 = ~pi3657 & ~pi9040;
assign w14769 = ~w14767 & ~w14768;
assign w14770 = pi0785 & ~w14769;
assign w14771 = ~pi0785 & w14769;
assign w14772 = ~w14770 & ~w14771;
assign w14773 = ~pi3682 & pi9040;
assign w14774 = ~pi3676 & ~pi9040;
assign w14775 = ~w14773 & ~w14774;
assign w14776 = pi0762 & ~w14775;
assign w14777 = ~pi0762 & w14775;
assign w14778 = ~w14776 & ~w14777;
assign w14779 = ~w14772 & ~w14778;
assign w14780 = ~pi3704 & pi9040;
assign w14781 = ~pi3674 & ~pi9040;
assign w14782 = ~w14780 & ~w14781;
assign w14783 = pi0778 & ~w14782;
assign w14784 = ~pi0778 & w14782;
assign w14785 = ~w14783 & ~w14784;
assign w14786 = ~pi3685 & pi9040;
assign w14787 = ~pi3707 & ~pi9040;
assign w14788 = ~w14786 & ~w14787;
assign w14789 = pi0786 & ~w14788;
assign w14790 = ~pi0786 & w14788;
assign w14791 = ~w14789 & ~w14790;
assign w14792 = w14785 & ~w14791;
assign w14793 = ~pi3663 & pi9040;
assign w14794 = ~pi3655 & ~pi9040;
assign w14795 = ~w14793 & ~w14794;
assign w14796 = pi0773 & ~w14795;
assign w14797 = ~pi0773 & w14795;
assign w14798 = ~w14796 & ~w14797;
assign w14799 = w14792 & w14798;
assign w14800 = ~w14785 & ~w14791;
assign w14801 = ~w14798 & w14800;
assign w14802 = ~w14799 & ~w14801;
assign w14803 = w14779 & ~w14802;
assign w14804 = ~pi3684 & pi9040;
assign w14805 = ~pi3685 & ~pi9040;
assign w14806 = ~w14804 & ~w14805;
assign w14807 = pi0792 & ~w14806;
assign w14808 = ~pi0792 & w14806;
assign w14809 = ~w14807 & ~w14808;
assign w14810 = w14785 & w14791;
assign w14811 = ~w14785 & w14798;
assign w14812 = ~w14810 & ~w14811;
assign w14813 = ~w14772 & w14778;
assign w14814 = ~w14812 & w14813;
assign w14815 = w14791 & w14811;
assign w14816 = w14779 & ~w14815;
assign w14817 = ~w14814 & ~w14816;
assign w14818 = ~w14778 & ~w14812;
assign w14819 = ~w14812 & w65160;
assign w14820 = ~w14817 & ~w14819;
assign w14821 = w14798 & w14810;
assign w14822 = w14792 & ~w14798;
assign w14823 = w14792 & w65160;
assign w14824 = w14778 & w14811;
assign w14825 = (w14772 & ~w14810) | (w14772 & w65161) | (~w14810 & w65161);
assign w14826 = ~w14824 & w14825;
assign w14827 = ~w14823 & w14826;
assign w14828 = (w14809 & w14820) | (w14809 & w65162) | (w14820 & w65162);
assign w14829 = ~w14778 & ~w14785;
assign w14830 = w14772 & ~w14829;
assign w14831 = w14791 & w14812;
assign w14832 = w14830 & ~w14831;
assign w14833 = ~w14778 & w14798;
assign w14834 = w14785 & w14833;
assign w14835 = ~w14772 & ~w14824;
assign w14836 = ~w14834 & w14835;
assign w14837 = ~w14832 & ~w14836;
assign w14838 = w14778 & w14810;
assign w14839 = w14810 & w14843;
assign w14840 = w14779 & w14792;
assign w14841 = ~w14839 & ~w14840;
assign w14842 = ~w14791 & w14833;
assign w14843 = w14778 & ~w14798;
assign w14844 = w14772 & w14843;
assign w14845 = ~w14842 & ~w14844;
assign w14846 = w14785 & ~w14845;
assign w14847 = ~w14809 & w14841;
assign w14848 = ~w14846 & w14847;
assign w14849 = ~w14837 & w14848;
assign w14850 = ~w14828 & ~w14849;
assign w14851 = w14791 & w14829;
assign w14852 = w14829 & w65163;
assign w14853 = w14833 & w14800;
assign w14854 = ~w14838 & ~w14852;
assign w14855 = ~w14853 & w14854;
assign w14856 = w14772 & ~w14855;
assign w14857 = ~w14803 & ~w14856;
assign w14858 = ~w14850 & w14857;
assign w14859 = pi0801 & ~w14858;
assign w14860 = ~pi0801 & w14858;
assign w14861 = ~w14859 & ~w14860;
assign w14862 = ~pi3659 & pi9040;
assign w14863 = ~pi3673 & ~pi9040;
assign w14864 = ~w14862 & ~w14863;
assign w14865 = pi0797 & ~w14864;
assign w14866 = ~pi0797 & w14864;
assign w14867 = ~w14865 & ~w14866;
assign w14868 = ~pi3662 & pi9040;
assign w14869 = ~pi3752 & ~pi9040;
assign w14870 = ~w14868 & ~w14869;
assign w14871 = pi0772 & ~w14870;
assign w14872 = ~pi0772 & w14870;
assign w14873 = ~w14871 & ~w14872;
assign w14874 = ~pi3669 & pi9040;
assign w14875 = ~pi3680 & ~pi9040;
assign w14876 = ~w14874 & ~w14875;
assign w14877 = pi0777 & ~w14876;
assign w14878 = ~pi0777 & w14876;
assign w14879 = ~w14877 & ~w14878;
assign w14880 = w14873 & ~w14879;
assign w14881 = ~pi3683 & pi9040;
assign w14882 = ~pi3687 & ~pi9040;
assign w14883 = ~w14881 & ~w14882;
assign w14884 = pi0780 & ~w14883;
assign w14885 = ~pi0780 & w14883;
assign w14886 = ~w14884 & ~w14885;
assign w14887 = ~pi3700 & pi9040;
assign w14888 = ~pi3697 & ~pi9040;
assign w14889 = ~w14887 & ~w14888;
assign w14890 = pi0784 & ~w14889;
assign w14891 = ~pi0784 & w14889;
assign w14892 = ~w14890 & ~w14891;
assign w14893 = w14873 & ~w14892;
assign w14894 = (~w14886 & ~w14893) | (~w14886 & w65164) | (~w14893 & w65164);
assign w14895 = w14880 & w14894;
assign w14896 = ~w14873 & ~w14879;
assign w14897 = ~pi3687 & pi9040;
assign w14898 = ~pi3694 & ~pi9040;
assign w14899 = ~w14897 & ~w14898;
assign w14900 = pi0793 & ~w14899;
assign w14901 = ~pi0793 & w14899;
assign w14902 = ~w14900 & ~w14901;
assign w14903 = w14886 & ~w14902;
assign w14904 = w14892 & w14902;
assign w14905 = ~w14892 & ~w14902;
assign w14906 = ~w14904 & ~w14905;
assign w14907 = (w14896 & ~w14906) | (w14896 & w63691) | (~w14906 & w63691);
assign w14908 = ~w14886 & ~w14902;
assign w14909 = w14886 & w14902;
assign w14910 = ~w14908 & ~w14909;
assign w14911 = ~w14873 & w14902;
assign w14912 = w14879 & ~w14911;
assign w14913 = ~w14910 & w14912;
assign w14914 = ~w14907 & ~w14913;
assign w14915 = ~w14895 & w14914;
assign w14916 = w14880 & w14909;
assign w14917 = w14892 & w14909;
assign w14918 = ~w14916 & ~w14917;
assign w14919 = w14873 & ~w14902;
assign w14920 = w14892 & ~w14919;
assign w14921 = ~w14911 & w14920;
assign w14922 = ~w14918 & ~w14921;
assign w14923 = w14893 & ~w14902;
assign w14924 = w14893 & w65165;
assign w14925 = ~w14922 & ~w14924;
assign w14926 = w14915 & w14925;
assign w14927 = ~w14867 & ~w14926;
assign w14928 = ~w14873 & w14879;
assign w14929 = ~w14892 & w14902;
assign w14930 = w14928 & w14929;
assign w14931 = ~w14916 & ~w14930;
assign w14932 = w14886 & w14928;
assign w14933 = w14928 & w14903;
assign w14934 = (w14896 & ~w14906) | (w14896 & w63692) | (~w14906 & w63692);
assign w14935 = w14906 & w14934;
assign w14936 = ~w14911 & ~w14919;
assign w14937 = ~w14886 & ~w14892;
assign w14938 = ~w14936 & w14937;
assign w14939 = w14873 & w14879;
assign w14940 = w14904 & w14939;
assign w14941 = w14931 & ~w14940;
assign w14942 = ~w14933 & ~w14938;
assign w14943 = w14941 & w14942;
assign w14944 = (w14867 & ~w14943) | (w14867 & w65166) | (~w14943 & w65166);
assign w14945 = ~w14879 & ~w14893;
assign w14946 = ~w14920 & w14945;
assign w14947 = w14886 & ~w14946;
assign w14948 = ~w14886 & ~w14930;
assign w14949 = ~w14909 & ~w14948;
assign w14950 = ~w14947 & w14949;
assign w14951 = ~w14944 & ~w14950;
assign w14952 = ~w14927 & w14951;
assign w14953 = ~pi0806 & w14952;
assign w14954 = pi0806 & ~w14952;
assign w14955 = ~w14953 & ~w14954;
assign w14956 = w14886 & ~w14924;
assign w14957 = w14919 & w14956;
assign w14958 = w14873 & w14929;
assign w14959 = ~w14886 & w14939;
assign w14960 = ~w14932 & ~w14959;
assign w14961 = ~w14892 & ~w14960;
assign w14962 = ~w14934 & ~w14958;
assign w14963 = ~w14961 & w14962;
assign w14964 = (~w14867 & ~w14963) | (~w14867 & w65167) | (~w14963 & w65167);
assign w14965 = w14896 & w14905;
assign w14966 = w14912 & w14920;
assign w14967 = ~w14965 & ~w14966;
assign w14968 = ~w14886 & ~w14967;
assign w14969 = w14880 & ~w14929;
assign w14970 = w14948 & ~w14969;
assign w14971 = w14896 & w14902;
assign w14972 = w14956 & ~w14971;
assign w14973 = ~w14970 & ~w14972;
assign w14974 = ~w14966 & ~w14973;
assign w14975 = w14867 & ~w14974;
assign w14976 = ~w14922 & ~w14968;
assign w14977 = ~w14964 & w14976;
assign w14978 = ~w14975 & w14977;
assign w14979 = pi0814 & ~w14978;
assign w14980 = ~pi0814 & w14978;
assign w14981 = ~w14979 & ~w14980;
assign w14982 = ~pi3664 & pi9040;
assign w14983 = ~pi3690 & ~pi9040;
assign w14984 = ~w14982 & ~w14983;
assign w14985 = pi0783 & ~w14984;
assign w14986 = ~pi0783 & w14984;
assign w14987 = ~w14985 & ~w14986;
assign w14988 = ~pi3667 & pi9040;
assign w14989 = ~pi3695 & ~pi9040;
assign w14990 = ~w14988 & ~w14989;
assign w14991 = pi0777 & ~w14990;
assign w14992 = ~pi0777 & w14990;
assign w14993 = ~w14991 & ~w14992;
assign w14994 = ~w14987 & w14993;
assign w14995 = ~pi3655 & pi9040;
assign w14996 = ~pi3701 & ~pi9040;
assign w14997 = ~w14995 & ~w14996;
assign w14998 = pi0773 & ~w14997;
assign w14999 = ~pi0773 & w14997;
assign w15000 = ~w14998 & ~w14999;
assign w15001 = ~pi3709 & pi9040;
assign w15002 = ~pi3706 & ~pi9040;
assign w15003 = ~w15001 & ~w15002;
assign w15004 = pi0797 & ~w15003;
assign w15005 = ~pi0797 & w15003;
assign w15006 = ~w15004 & ~w15005;
assign w15007 = w15000 & w15006;
assign w15008 = w14994 & w15007;
assign w15009 = ~w14987 & ~w15000;
assign w15010 = w14987 & w15000;
assign w15011 = ~w15009 & ~w15010;
assign w15012 = w14987 & ~w15006;
assign w15013 = w14993 & ~w15012;
assign w15014 = w15011 & w15013;
assign w15015 = w14994 & ~w15006;
assign w15016 = ~w14993 & w15007;
assign w15017 = ~pi3702 & pi9040;
assign w15018 = ~pi3667 & ~pi9040;
assign w15019 = ~w15017 & ~w15018;
assign w15020 = pi0775 & ~w15019;
assign w15021 = ~pi0775 & w15019;
assign w15022 = ~w15020 & ~w15021;
assign w15023 = (~w15022 & ~w15007) | (~w15022 & w65168) | (~w15007 & w65168);
assign w15024 = ~w15015 & w15023;
assign w15025 = (w15022 & ~w15007) | (w15022 & w65169) | (~w15007 & w65169);
assign w15026 = ~w14993 & ~w15006;
assign w15027 = w14987 & w15006;
assign w15028 = ~w14994 & ~w15000;
assign w15029 = ~w15027 & w15028;
assign w15030 = w15025 & ~w15026;
assign w15031 = ~w15029 & w15030;
assign w15032 = ~w15024 & ~w15031;
assign w15033 = ~w15014 & ~w15032;
assign w15034 = ~pi3658 & pi9040;
assign w15035 = pi3689 & ~pi9040;
assign w15036 = ~w15034 & ~w15035;
assign w15037 = pi0778 & ~w15036;
assign w15038 = ~pi0778 & w15036;
assign w15039 = ~w15037 & ~w15038;
assign w15040 = ~w15033 & w15039;
assign w15041 = ~w14993 & ~w15000;
assign w15042 = w15022 & ~w15041;
assign w15043 = w15009 & w15042;
assign w15044 = w15011 & w15022;
assign w15045 = w14993 & w15012;
assign w15046 = ~w15044 & w15045;
assign w15047 = ~w15043 & ~w15046;
assign w15048 = ~w15039 & ~w15047;
assign w15049 = ~w15022 & w15027;
assign w15050 = ~w15007 & ~w15022;
assign w15051 = ~w15012 & ~w15039;
assign w15052 = w15050 & w15051;
assign w15053 = ~w15049 & ~w15052;
assign w15054 = ~w14993 & ~w15053;
assign w15055 = ~w15000 & w15006;
assign w15056 = w14993 & w15055;
assign w15057 = ~w15026 & ~w15056;
assign w15058 = w15044 & ~w15057;
assign w15059 = ~w15008 & ~w15058;
assign w15060 = ~w15054 & w15059;
assign w15061 = ~w15048 & w15060;
assign w15062 = ~w15040 & w15061;
assign w15063 = ~pi0809 & w15062;
assign w15064 = pi0809 & ~w15062;
assign w15065 = ~w15063 & ~w15064;
assign w15066 = w14778 & w14799;
assign w15067 = ~w14818 & ~w15066;
assign w15068 = ~w14772 & ~w14809;
assign w15069 = ~w15067 & w15068;
assign w15070 = ~w14779 & w14791;
assign w15071 = w14833 & w15070;
assign w15072 = w14778 & ~w14809;
assign w15073 = w14812 & w65170;
assign w15074 = w14772 & ~w14809;
assign w15075 = w14800 & ~w14833;
assign w15076 = ~w14821 & ~w14822;
assign w15077 = ~w15075 & w15076;
assign w15078 = w14800 & w14843;
assign w15079 = w15074 & ~w15078;
assign w15080 = ~w15077 & w15079;
assign w15081 = ~w14815 & ~w14853;
assign w15082 = ~w15066 & w15081;
assign w15083 = w14772 & ~w15082;
assign w15084 = ~w14838 & ~w15075;
assign w15085 = ~w14772 & ~w15084;
assign w15086 = ~w14852 & ~w15078;
assign w15087 = w14841 & w15086;
assign w15088 = ~w15085 & w15087;
assign w15089 = ~w15083 & w15088;
assign w15090 = w14809 & ~w15089;
assign w15091 = ~w14823 & ~w15071;
assign w15092 = ~w15073 & w15091;
assign w15093 = ~w15069 & w15092;
assign w15094 = ~w15080 & w15093;
assign w15095 = ~w15090 & w15094;
assign w15096 = pi0802 & ~w15095;
assign w15097 = ~pi0802 & w15095;
assign w15098 = ~w15096 & ~w15097;
assign w15099 = w14506 & w14518;
assign w15100 = w14502 & ~w14661;
assign w15101 = ~w14497 & ~w14650;
assign w15102 = ~w15099 & ~w15100;
assign w15103 = w15101 & w15102;
assign w15104 = ~w14471 & ~w14488;
assign w15105 = ~w14507 & w15104;
assign w15106 = ~w14519 & w15105;
assign w15107 = ~w14459 & ~w14514;
assign w15108 = ~w14520 & w15107;
assign w15109 = ~w15106 & w15108;
assign w15110 = w14453 & ~w14505;
assign w15111 = w15109 & w15110;
assign w15112 = ~w14459 & w14505;
assign w15113 = w14648 & w15112;
assign w15114 = w14459 & ~w14491;
assign w15115 = ~w14453 & ~w15109;
assign w15116 = ~w15114 & w15115;
assign w15117 = (~w15113 & w15103) | (~w15113 & w65171) | (w15103 & w65171);
assign w15118 = ~w15111 & w15117;
assign w15119 = ~w15116 & w15118;
assign w15120 = pi0807 & ~w15119;
assign w15121 = ~pi0807 & w15119;
assign w15122 = ~w15120 & ~w15121;
assign w15123 = w14608 & ~w14611;
assign w15124 = ~w14612 & ~w15123;
assign w15125 = ~w14558 & w14622;
assign w15126 = w14606 & w15125;
assign w15127 = ~w14604 & ~w15125;
assign w15128 = ~w14552 & ~w15127;
assign w15129 = w14552 & w14567;
assign w15130 = ~w14581 & ~w14585;
assign w15131 = w15129 & w15130;
assign w15132 = ~w14587 & ~w15129;
assign w15133 = w14545 & ~w15132;
assign w15134 = ~w14601 & ~w15131;
assign w15135 = ~w15133 & w15134;
assign w15136 = ~w15128 & w15135;
assign w15137 = w14601 & ~w14626;
assign w15138 = ~w14576 & w15137;
assign w15139 = w14614 & w15138;
assign w15140 = ~w15136 & ~w15139;
assign w15141 = ~w15124 & ~w15126;
assign w15142 = ~w14603 & w15141;
assign w15143 = ~w15140 & w65172;
assign w15144 = (pi0830 & w15140) | (pi0830 & w65173) | (w15140 & w65173);
assign w15145 = ~w15143 & ~w15144;
assign w15146 = w15041 & w15049;
assign w15147 = ~w14987 & w15006;
assign w15148 = ~w15022 & w15147;
assign w15149 = ~w14987 & w15000;
assign w15150 = ~w15055 & ~w15149;
assign w15151 = ~w15012 & w15150;
assign w15152 = w15150 & w65174;
assign w15153 = ~w15016 & ~w15152;
assign w15154 = w15022 & ~w15153;
assign w15155 = w14993 & w15000;
assign w15156 = ~w15041 & ~w15155;
assign w15157 = w15012 & w15156;
assign w15158 = w15039 & ~w15148;
assign w15159 = ~w15157 & w15158;
assign w15160 = ~w15154 & w15159;
assign w15161 = w14987 & w15056;
assign w15162 = w15147 & ~w15156;
assign w15163 = w15025 & ~w15162;
assign w15164 = ~w15006 & w15149;
assign w15165 = w15023 & ~w15164;
assign w15166 = ~w15163 & ~w15165;
assign w15167 = w15012 & w15041;
assign w15168 = ~w15015 & ~w15167;
assign w15169 = w15050 & w15155;
assign w15170 = ~w15039 & ~w15161;
assign w15171 = w15168 & ~w15169;
assign w15172 = w15170 & w15171;
assign w15173 = ~w15166 & w15172;
assign w15174 = ~w15160 & ~w15173;
assign w15175 = ~w15014 & ~w15157;
assign w15176 = w15163 & ~w15175;
assign w15177 = ~w15146 & ~w15176;
assign w15178 = ~w15174 & w15177;
assign w15179 = pi0810 & w15178;
assign w15180 = ~pi0810 & ~w15178;
assign w15181 = ~w15179 & ~w15180;
assign w15182 = w14692 & w14698;
assign w15183 = ~w14720 & ~w15182;
assign w15184 = w14720 & ~w14744;
assign w15185 = ~w15183 & ~w15184;
assign w15186 = ~w14736 & w15185;
assign w15187 = ~w14736 & ~w14743;
assign w15188 = w14707 & ~w15187;
assign w15189 = ~w14701 & ~w14713;
assign w15190 = w14692 & w14720;
assign w15191 = ~w14721 & ~w15190;
assign w15192 = w15189 & ~w15191;
assign w15193 = ~w14686 & ~w14758;
assign w15194 = ~w15186 & w15193;
assign w15195 = ~w15188 & ~w15192;
assign w15196 = w15194 & w15195;
assign w15197 = w14739 & w15182;
assign w15198 = ~w14741 & ~w15190;
assign w15199 = w14698 & w14713;
assign w15200 = w15198 & w15199;
assign w15201 = ~w15197 & ~w15200;
assign w15202 = ~w14707 & ~w15201;
assign w15203 = w14742 & w15198;
assign w15204 = ~w14707 & ~w14723;
assign w15205 = ~w14739 & w15204;
assign w15206 = ~w15203 & w15205;
assign w15207 = ~w14720 & w15189;
assign w15208 = ~w14692 & ~w14754;
assign w15209 = w15184 & w15208;
assign w15210 = w14686 & ~w14745;
assign w15211 = ~w15197 & w15210;
assign w15212 = ~w15209 & w15211;
assign w15213 = ~w15206 & ~w15207;
assign w15214 = w15212 & w15213;
assign w15215 = ~w15202 & w15214;
assign w15216 = ~w15196 & ~w15215;
assign w15217 = ~pi0812 & w15216;
assign w15218 = pi0812 & ~w15216;
assign w15219 = ~w15217 & ~w15218;
assign w15220 = ~w15151 & w15168;
assign w15221 = ~w15029 & w15042;
assign w15222 = w15220 & w15221;
assign w15223 = ~w15147 & w15156;
assign w15224 = ~w15162 & ~w15223;
assign w15225 = w15022 & ~w15220;
assign w15226 = ~w15012 & w15224;
assign w15227 = ~w15225 & w15226;
assign w15228 = w15039 & ~w15222;
assign w15229 = ~w15227 & w15228;
assign w15230 = ~w15022 & ~w15224;
assign w15231 = (~w15039 & w15220) | (~w15039 & w65175) | (w15220 & w65175);
assign w15232 = ~w15230 & w15231;
assign w15233 = w14994 & w15055;
assign w15234 = ~w15167 & ~w15233;
assign w15235 = w15022 & ~w15234;
assign w15236 = ~w15022 & w15157;
assign w15237 = ~w15235 & ~w15236;
assign w15238 = (w15237 & w15229) | (w15237 & w65176) | (w15229 & w65176);
assign w15239 = ~pi0820 & w15238;
assign w15240 = pi0820 & ~w15238;
assign w15241 = ~w15239 & ~w15240;
assign w15242 = w14879 & w14886;
assign w15243 = ~w14923 & w14931;
assign w15244 = w15242 & ~w15243;
assign w15245 = w14880 & w14904;
assign w15246 = ~w14906 & w14928;
assign w15247 = w14960 & ~w15246;
assign w15248 = w14896 & ~w14904;
assign w15249 = ~w14908 & w15248;
assign w15250 = ~w15245 & ~w15249;
assign w15251 = (w15250 & ~w14963) | (w15250 & w65177) | (~w14963 & w65177);
assign w15252 = w14867 & ~w15251;
assign w15253 = ~w14910 & ~w14929;
assign w15254 = w15247 & w15253;
assign w15255 = (~w14867 & w15254) | (~w14867 & w65178) | (w15254 & w65178);
assign w15256 = ~w14896 & w14929;
assign w15257 = ~w14939 & w15256;
assign w15258 = w14937 & ~w15257;
assign w15259 = w14914 & w15258;
assign w15260 = ~w15244 & ~w15259;
assign w15261 = ~w15255 & w15260;
assign w15262 = ~w15252 & w15261;
assign w15263 = ~pi0815 & ~w15262;
assign w15264 = pi0815 & w15262;
assign w15265 = ~w15263 & ~w15264;
assign w15266 = w14821 & w15072;
assign w15267 = ~w14831 & ~w14834;
assign w15268 = w14772 & ~w15267;
assign w15269 = ~w14772 & w14785;
assign w15270 = ~w14798 & w15269;
assign w15271 = ~w14842 & ~w15270;
assign w15272 = ~w15268 & w15271;
assign w15273 = w14809 & ~w15272;
assign w15274 = ~w14801 & ~w14815;
assign w15275 = ~w14778 & w14809;
assign w15276 = ~w15074 & ~w15275;
assign w15277 = ~w15274 & w15276;
assign w15278 = w14779 & w14785;
assign w15279 = w15077 & w15278;
assign w15280 = w14852 & ~w15068;
assign w15281 = w15074 & w15274;
assign w15282 = w15267 & w15281;
assign w15283 = ~w15266 & ~w15277;
assign w15284 = ~w15280 & w15283;
assign w15285 = ~w15279 & ~w15282;
assign w15286 = w15284 & w15285;
assign w15287 = ~w15273 & w15286;
assign w15288 = pi0808 & ~w15287;
assign w15289 = ~pi0808 & w15287;
assign w15290 = ~w15288 & ~w15289;
assign w15291 = w15023 & ~w15150;
assign w15292 = ~w15056 & ~w15164;
assign w15293 = w15022 & w15292;
assign w15294 = w14987 & ~w14993;
assign w15295 = ~w15055 & w15294;
assign w15296 = (~w15295 & w15293) | (~w15295 & w65179) | (w15293 & w65179);
assign w15297 = ~w15039 & ~w15296;
assign w15298 = w15027 & w15041;
assign w15299 = ~w15010 & w15042;
assign w15300 = w15292 & w15299;
assign w15301 = ~w15008 & ~w15298;
assign w15302 = ~w15169 & w15301;
assign w15303 = ~w15300 & w15302;
assign w15304 = w15039 & ~w15303;
assign w15305 = ~w15152 & ~w15233;
assign w15306 = ~w15022 & ~w15305;
assign w15307 = ~w15011 & w15220;
assign w15308 = w15032 & w15307;
assign w15309 = ~w15304 & ~w15306;
assign w15310 = w15309 & w65180;
assign w15311 = pi0833 & ~w15310;
assign w15312 = ~pi0833 & w15310;
assign w15313 = ~w15311 & ~w15312;
assign w15314 = w14601 & ~w15133;
assign w15315 = w14539 & ~w14580;
assign w15316 = ~w14629 & w15315;
assign w15317 = w14580 & ~w14583;
assign w15318 = w14561 & w14610;
assign w15319 = ~w15316 & ~w15318;
assign w15320 = ~w15317 & w15319;
assign w15321 = ~w15314 & ~w15320;
assign w15322 = w14601 & ~w15318;
assign w15323 = ~w14573 & w15322;
assign w15324 = ~w14584 & w15323;
assign w15325 = ~w15321 & ~w15324;
assign w15326 = pi0817 & w15325;
assign w15327 = ~pi0817 & ~w15325;
assign w15328 = ~w15326 & ~w15327;
assign w15329 = ~w14507 & ~w14654;
assign w15330 = w14471 & w14487;
assign w15331 = ~w15329 & w15330;
assign w15332 = ~w14662 & w15329;
assign w15333 = w14504 & ~w15331;
assign w15334 = ~w15332 & w15333;
assign w15335 = ~w14513 & w14522;
assign w15336 = ~w14453 & ~w15335;
assign w15337 = w14453 & w14490;
assign w15338 = w14459 & ~w14669;
assign w15339 = ~w15337 & w15338;
assign w15340 = ~w15336 & w15339;
assign w15341 = ~w15334 & ~w15340;
assign w15342 = ~w14453 & ~w14505;
assign w15343 = ~w14647 & ~w15342;
assign w15344 = ~w14664 & w15343;
assign w15345 = ~w15341 & ~w15344;
assign w15346 = ~pi0846 & w15345;
assign w15347 = pi0846 & ~w15345;
assign w15348 = ~w15346 & ~w15347;
assign w15349 = w14389 & w14419;
assign w15350 = ~w14386 & ~w14430;
assign w15351 = ~w14422 & w15350;
assign w15352 = w14406 & ~w15351;
assign w15353 = ~w14413 & ~w15349;
assign w15354 = ~w15352 & w15353;
assign w15355 = ~w14370 & w14395;
assign w15356 = w14370 & ~w14406;
assign w15357 = ~w14373 & w65181;
assign w15358 = w14385 & w14389;
assign w15359 = w14406 & ~w14414;
assign w15360 = w14419 & w15359;
assign w15361 = w14372 & w14432;
assign w15362 = w14413 & ~w15358;
assign w15363 = ~w15361 & w15362;
assign w15364 = ~w15355 & ~w15360;
assign w15365 = w15363 & w15364;
assign w15366 = ~w15357 & w15365;
assign w15367 = ~w15354 & ~w15366;
assign w15368 = w14370 & w14394;
assign w15369 = ~w14435 & ~w15368;
assign w15370 = w14393 & ~w15369;
assign w15371 = ~w14413 & w14432;
assign w15372 = w14434 & ~w15371;
assign w15373 = ~w15355 & w15372;
assign w15374 = ~w15370 & w15373;
assign w15375 = w14406 & ~w15368;
assign w15376 = w14364 & w14386;
assign w15377 = ~w14398 & ~w15376;
assign w15378 = w14373 & ~w15377;
assign w15379 = w15375 & ~w15378;
assign w15380 = w14406 & ~w14430;
assign w15381 = w14396 & w15380;
assign w15382 = ~w15379 & ~w15381;
assign w15383 = ~w15374 & w15382;
assign w15384 = ~w15367 & ~w15383;
assign w15385 = ~pi0827 & w15384;
assign w15386 = pi0827 & ~w15384;
assign w15387 = ~w15385 & ~w15386;
assign w15388 = w14896 & w14917;
assign w15389 = w14903 & ~w14945;
assign w15390 = w14894 & ~w14921;
assign w15391 = w14867 & ~w15389;
assign w15392 = (w15391 & ~w14915) | (w15391 & w65182) | (~w14915 & w65182);
assign w15393 = w14879 & w14919;
assign w15394 = w14894 & ~w15393;
assign w15395 = ~w14947 & ~w15394;
assign w15396 = ~w14867 & ~w14940;
assign w15397 = ~w15257 & w15396;
assign w15398 = ~w15395 & w15397;
assign w15399 = ~w15392 & ~w15398;
assign w15400 = w14867 & ~w14939;
assign w15401 = ~w14879 & ~w14886;
assign w15402 = ~w15242 & ~w15401;
assign w15403 = ~w15400 & w15402;
assign w15404 = w14921 & ~w15403;
assign w15405 = ~w15388 & ~w15404;
assign w15406 = ~w15399 & w15405;
assign w15407 = pi0821 & w15406;
assign w15408 = ~pi0821 & ~w15406;
assign w15409 = ~w15407 & ~w15408;
assign w15410 = w15356 & w15358;
assign w15411 = w14406 & w14435;
assign w15412 = ~w14370 & w14435;
assign w15413 = ~w14370 & ~w14406;
assign w15414 = w14394 & w15413;
assign w15415 = ~w14413 & ~w15414;
assign w15416 = ~w14370 & w14386;
assign w15417 = ~w14433 & ~w15416;
assign w15418 = w14406 & ~w15417;
assign w15419 = ~w14418 & ~w15358;
assign w15420 = w14370 & ~w15419;
assign w15421 = ~w14395 & ~w14421;
assign w15422 = ~w15412 & w15415;
assign w15423 = w15421 & w15422;
assign w15424 = ~w15357 & ~w15418;
assign w15425 = ~w15420 & w15424;
assign w15426 = w15423 & w15425;
assign w15427 = (~w14406 & ~w14430) | (~w14406 & w65183) | (~w14430 & w65183);
assign w15428 = ~w14373 & w14432;
assign w15429 = w15427 & ~w15428;
assign w15430 = ~w14364 & w14392;
assign w15431 = ~w15376 & ~w15430;
assign w15432 = w15375 & w15431;
assign w15433 = ~w15429 & ~w15432;
assign w15434 = w14413 & ~w15378;
assign w15435 = ~w15433 & w15434;
assign w15436 = ~w15410 & ~w15411;
assign w15437 = (w15436 & w15426) | (w15436 & w65184) | (w15426 & w65184);
assign w15438 = pi0822 & ~w15437;
assign w15439 = ~pi0822 & w15437;
assign w15440 = ~w15438 & ~w15439;
assign w15441 = w14813 & ~w15076;
assign w15442 = ~w14799 & ~w14851;
assign w15443 = (w14772 & ~w15442) | (w14772 & w65185) | (~w15442 & w65185);
assign w15444 = w14779 & w14810;
assign w15445 = ~w14823 & ~w15444;
assign w15446 = ~w14809 & w15445;
assign w15447 = ~w15443 & w15446;
assign w15448 = ~w14829 & ~w14843;
assign w15449 = w15070 & w15448;
assign w15450 = w14809 & ~w14853;
assign w15451 = ~w15449 & w15450;
assign w15452 = ~w15447 & ~w15451;
assign w15453 = w14809 & w15445;
assign w15454 = ~w14800 & ~w15453;
assign w15455 = w14779 & ~w15454;
assign w15456 = ~w14791 & w14811;
assign w15457 = ~w15073 & ~w15456;
assign w15458 = w15068 & ~w15457;
assign w15459 = ~w14801 & w15082;
assign w15460 = w14830 & ~w15459;
assign w15461 = ~w15441 & ~w15458;
assign w15462 = ~w15452 & w15461;
assign w15463 = ~w15455 & ~w15460;
assign w15464 = w15462 & w15463;
assign w15465 = pi0803 & ~w15464;
assign w15466 = ~pi0803 & w15464;
assign w15467 = ~w15465 & ~w15466;
assign w15468 = w14406 & ~w14420;
assign w15469 = ~w14397 & w15427;
assign w15470 = ~w15468 & ~w15469;
assign w15471 = w15369 & ~w15416;
assign w15472 = ~w14406 & ~w15471;
assign w15473 = ~w15350 & w15359;
assign w15474 = ~w14421 & ~w15430;
assign w15475 = w14440 & w15474;
assign w15476 = ~w15473 & w15475;
assign w15477 = ~w15472 & w15476;
assign w15478 = ~w14398 & ~w14429;
assign w15479 = w14372 & ~w15478;
assign w15480 = w15415 & ~w15479;
assign w15481 = ~w15381 & w15480;
assign w15482 = ~w15477 & ~w15481;
assign w15483 = ~w15470 & ~w15482;
assign w15484 = ~pi0823 & w15483;
assign w15485 = pi0823 & ~w15483;
assign w15486 = ~w15484 & ~w15485;
assign w15487 = w14707 & ~w14743;
assign w15488 = (w14746 & ~w15201) | (w14746 & w63693) | (~w15201 & w63693);
assign w15489 = (~w14726 & w15488) | (~w14726 & w65186) | (w15488 & w65186);
assign w15490 = w14686 & ~w15489;
assign w15491 = w14714 & w14741;
assign w15492 = w14698 & w15491;
assign w15493 = ~w14707 & ~w15190;
assign w15494 = ~w14745 & w15493;
assign w15495 = ~w15189 & w15494;
assign w15496 = ~w14747 & w15201;
assign w15497 = (~w14686 & ~w15496) | (~w14686 & w65187) | (~w15496 & w65187);
assign w15498 = ~w15202 & ~w15492;
assign w15499 = ~w15497 & w15498;
assign w15500 = ~w15490 & w15499;
assign w15501 = pi0824 & ~w15500;
assign w15502 = ~pi0824 & w15500;
assign w15503 = ~w15501 & ~w15502;
assign w15504 = w14707 & ~w15185;
assign w15505 = w14724 & ~w15197;
assign w15506 = ~w15203 & w15505;
assign w15507 = ~w15504 & ~w15506;
assign w15508 = w14723 & w15182;
assign w15509 = ~w15491 & ~w15508;
assign w15510 = ~w15507 & w15509;
assign w15511 = ~w14686 & ~w15510;
assign w15512 = w14692 & ~w14754;
assign w15513 = ~w14758 & ~w15512;
assign w15514 = ~w15185 & ~w15513;
assign w15515 = ~w14740 & ~w15206;
assign w15516 = (w14686 & ~w15515) | (w14686 & w65188) | (~w15515 & w65188);
assign w15517 = ~w14699 & ~w14734;
assign w15518 = ~w14754 & ~w14756;
assign w15519 = ~w15517 & w15518;
assign w15520 = ~w15516 & ~w15519;
assign w15521 = ~w15511 & w15520;
assign w15522 = ~pi0829 & w15521;
assign w15523 = pi0829 & ~w15521;
assign w15524 = ~w15522 & ~w15523;
assign w15525 = ~pi3691 & pi9040;
assign w15526 = ~pi3660 & ~pi9040;
assign w15527 = ~w15525 & ~w15526;
assign w15528 = pi0791 & ~w15527;
assign w15529 = ~pi0791 & w15527;
assign w15530 = ~w15528 & ~w15529;
assign w15531 = ~pi3666 & pi9040;
assign w15532 = ~pi3700 & ~pi9040;
assign w15533 = ~w15531 & ~w15532;
assign w15534 = pi0794 & ~w15533;
assign w15535 = ~pi0794 & w15533;
assign w15536 = ~w15534 & ~w15535;
assign w15537 = ~w15530 & w15536;
assign w15538 = ~pi3661 & pi9040;
assign w15539 = ~pi3693 & ~pi9040;
assign w15540 = ~w15538 & ~w15539;
assign w15541 = pi0793 & ~w15540;
assign w15542 = ~pi0793 & w15540;
assign w15543 = ~w15541 & ~w15542;
assign w15544 = ~pi3665 & pi9040;
assign w15545 = ~pi3691 & ~pi9040;
assign w15546 = ~w15544 & ~w15545;
assign w15547 = pi0776 & ~w15546;
assign w15548 = ~pi0776 & w15546;
assign w15549 = ~w15547 & ~w15548;
assign w15550 = w15543 & w15549;
assign w15551 = w15537 & w15550;
assign w15552 = ~pi3693 & pi9040;
assign w15553 = ~pi3696 & ~pi9040;
assign w15554 = ~w15552 & ~w15553;
assign w15555 = pi0782 & ~w15554;
assign w15556 = ~pi0782 & w15554;
assign w15557 = ~w15555 & ~w15556;
assign w15558 = w15551 & w15557;
assign w15559 = w15530 & w15536;
assign w15560 = ~w15530 & ~w15536;
assign w15561 = w15543 & ~w15557;
assign w15562 = ~w15543 & w15557;
assign w15563 = ~w15561 & ~w15562;
assign w15564 = w15560 & w15563;
assign w15565 = w15530 & w15557;
assign w15566 = w15536 & w15561;
assign w15567 = ~w15565 & ~w15566;
assign w15568 = ~w15566 & w63694;
assign w15569 = ~w15564 & w15568;
assign w15570 = ~w15559 & ~w15569;
assign w15571 = w15530 & ~w15543;
assign w15572 = w15536 & w15557;
assign w15573 = ~w15571 & ~w15572;
assign w15574 = ~w15543 & w15559;
assign w15575 = ~w15573 & ~w15574;
assign w15576 = ~pi3679 & pi9040;
assign w15577 = ~pi3659 & ~pi9040;
assign w15578 = ~w15576 & ~w15577;
assign w15579 = pi0772 & ~w15578;
assign w15580 = ~pi0772 & w15578;
assign w15581 = ~w15579 & ~w15580;
assign w15582 = ~w15575 & w15581;
assign w15583 = ~w15570 & w15582;
assign w15584 = ~w15530 & ~w15557;
assign w15585 = ~w15549 & ~w15584;
assign w15586 = ~w15575 & ~w15585;
assign w15587 = ~w15549 & ~w15573;
assign w15588 = ~w15586 & ~w15587;
assign w15589 = ~w15563 & ~w15567;
assign w15590 = (~w15530 & w15589) | (~w15530 & w65189) | (w15589 & w65189);
assign w15591 = ~w15588 & ~w15590;
assign w15592 = ~w15581 & ~w15591;
assign w15593 = ~w15543 & ~w15557;
assign w15594 = w15530 & w15593;
assign w15595 = (w15581 & w15594) | (w15581 & w65190) | (w15594 & w65190);
assign w15596 = ~w15574 & ~w15595;
assign w15597 = ~w15549 & ~w15596;
assign w15598 = ~w15558 & ~w15597;
assign w15599 = ~w15583 & w15598;
assign w15600 = ~w15592 & w15599;
assign w15601 = pi0825 & ~w15600;
assign w15602 = ~pi0825 & w15600;
assign w15603 = ~w15601 & ~w15602;
assign w15604 = w15559 & w15593;
assign w15605 = ~w15530 & w15543;
assign w15606 = (~w15605 & w15567) | (~w15605 & w65191) | (w15567 & w65191);
assign w15607 = ~w15549 & ~w15593;
assign w15608 = w15606 & w15607;
assign w15609 = ~w15604 & ~w15608;
assign w15610 = w15581 & ~w15609;
assign w15611 = ~w15536 & w15593;
assign w15612 = ~w15530 & w15611;
assign w15613 = ~w15581 & ~w15612;
assign w15614 = w15606 & ~w15612;
assign w15615 = w15549 & ~w15613;
assign w15616 = ~w15614 & w15615;
assign w15617 = ~w15550 & ~w15563;
assign w15618 = ~w15559 & ~w15560;
assign w15619 = ~w15566 & w15618;
assign w15620 = ~w15617 & ~w15619;
assign w15621 = w15617 & w15618;
assign w15622 = ~w15581 & ~w15620;
assign w15623 = (~w15551 & ~w15622) | (~w15551 & w65192) | (~w15622 & w65192);
assign w15624 = ~w15616 & w15623;
assign w15625 = ~w15610 & w15624;
assign w15626 = pi0831 & ~w15625;
assign w15627 = ~pi0831 & w15625;
assign w15628 = ~w15626 & ~w15627;
assign w15629 = ~w15565 & ~w15584;
assign w15630 = w15543 & ~w15629;
assign w15631 = ~w15549 & w15562;
assign w15632 = ~w15630 & ~w15631;
assign w15633 = ~w15629 & w15632;
assign w15634 = ~w15570 & w15633;
assign w15635 = ~w15543 & ~w15565;
assign w15636 = (w15549 & w15630) | (w15549 & w65193) | (w15630 & w65193);
assign w15637 = ~w15549 & ~w15611;
assign w15638 = ~w15630 & w15637;
assign w15639 = ~w15636 & ~w15638;
assign w15640 = w15613 & ~w15639;
assign w15641 = w15549 & ~w15561;
assign w15642 = w15536 & ~w15557;
assign w15643 = ~w15605 & w15642;
assign w15644 = ~w15641 & w15643;
assign w15645 = ~w15536 & ~w15632;
assign w15646 = ~w15536 & w15549;
assign w15647 = w15594 & w15646;
assign w15648 = w15560 & w15562;
assign w15649 = w15581 & ~w15648;
assign w15650 = ~w15644 & w15649;
assign w15651 = ~w15647 & w15650;
assign w15652 = ~w15645 & w15651;
assign w15653 = ~w15640 & ~w15652;
assign w15654 = w15537 & w15585;
assign w15655 = ~w15634 & ~w15654;
assign w15656 = ~w15653 & w15655;
assign w15657 = pi0816 & w15656;
assign w15658 = ~pi0816 & ~w15656;
assign w15659 = ~w15657 & ~w15658;
assign w15660 = (~w15549 & w15589) | (~w15549 & w63695) | (w15589 & w63695);
assign w15661 = ~w15568 & ~w15654;
assign w15662 = (~w15560 & ~w15563) | (~w15560 & w63696) | (~w15563 & w63696);
assign w15663 = w15560 & ~w15641;
assign w15664 = ~w15617 & w15663;
assign w15665 = ~w15662 & ~w15664;
assign w15666 = ~w15661 & ~w15665;
assign w15667 = (w15581 & ~w15662) | (w15581 & w65194) | (~w15662 & w65194);
assign w15668 = ~w15666 & w63697;
assign w15669 = (~w15581 & w15666) | (~w15581 & w65195) | (w15666 & w65195);
assign w15670 = w15587 & w15630;
assign w15671 = ~w15563 & w15646;
assign w15672 = w15629 & w15671;
assign w15673 = ~w15670 & ~w15672;
assign w15674 = ~w15668 & w15673;
assign w15675 = (pi0832 & ~w15674) | (pi0832 & w65196) | (~w15674 & w65196);
assign w15676 = w15674 & w65197;
assign w15677 = ~w15675 & ~w15676;
assign w15678 = ~pi3717 & pi9040;
assign w15679 = ~pi3750 & ~pi9040;
assign w15680 = ~w15678 & ~w15679;
assign w15681 = pi0835 & ~w15680;
assign w15682 = ~pi0835 & w15680;
assign w15683 = ~w15681 & ~w15682;
assign w15684 = ~pi3716 & pi9040;
assign w15685 = ~pi3774 & ~pi9040;
assign w15686 = ~w15684 & ~w15685;
assign w15687 = pi0854 & ~w15686;
assign w15688 = ~pi0854 & w15686;
assign w15689 = ~w15687 & ~w15688;
assign w15690 = w15683 & ~w15689;
assign w15691 = ~pi3725 & pi9040;
assign w15692 = ~pi3735 & ~pi9040;
assign w15693 = ~w15691 & ~w15692;
assign w15694 = pi0838 & ~w15693;
assign w15695 = ~pi0838 & w15693;
assign w15696 = ~w15694 & ~w15695;
assign w15697 = ~pi3738 & pi9040;
assign w15698 = ~pi3712 & ~pi9040;
assign w15699 = ~w15697 & ~w15698;
assign w15700 = pi0850 & ~w15699;
assign w15701 = ~pi0850 & w15699;
assign w15702 = ~w15700 & ~w15701;
assign w15703 = ~pi3768 & pi9040;
assign w15704 = ~pi3722 & ~pi9040;
assign w15705 = ~w15703 & ~w15704;
assign w15706 = pi0828 & ~w15705;
assign w15707 = ~pi0828 & w15705;
assign w15708 = ~w15706 & ~w15707;
assign w15709 = ~w15702 & w15708;
assign w15710 = ~w15683 & ~w15696;
assign w15711 = w15709 & w15710;
assign w15712 = w15689 & ~w15708;
assign w15713 = ~w15683 & ~w15712;
assign w15714 = ~w15709 & ~w15713;
assign w15715 = ~w15696 & ~w15711;
assign w15716 = ~w15714 & w15715;
assign w15717 = w15690 & w15716;
assign w15718 = ~w15690 & ~w15709;
assign w15719 = ~w15689 & ~w15702;
assign w15720 = w15683 & ~w15708;
assign w15721 = ~w15683 & w15708;
assign w15722 = ~w15720 & ~w15721;
assign w15723 = ~w15719 & ~w15722;
assign w15724 = ~w15718 & w15723;
assign w15725 = ~w15683 & ~w15708;
assign w15726 = w15689 & w15702;
assign w15727 = w15725 & w15726;
assign w15728 = ~w15711 & ~w15727;
assign w15729 = w15719 & w15725;
assign w15730 = ~w15724 & w65198;
assign w15731 = w15696 & ~w15730;
assign w15732 = ~pi3750 & pi9040;
assign w15733 = ~pi3769 & ~pi9040;
assign w15734 = ~w15732 & ~w15733;
assign w15735 = pi0863 & ~w15734;
assign w15736 = ~pi0863 & w15734;
assign w15737 = ~w15735 & ~w15736;
assign w15738 = w15696 & ~w15709;
assign w15739 = w15690 & ~w15738;
assign w15740 = w15689 & ~w15702;
assign w15741 = w15710 & w15740;
assign w15742 = w15702 & w15725;
assign w15743 = w15683 & w15689;
assign w15744 = ~w15702 & ~w15708;
assign w15745 = w15743 & w15744;
assign w15746 = ~w15742 & ~w15745;
assign w15747 = w15696 & ~w15746;
assign w15748 = w15702 & w15708;
assign w15749 = w15696 & ~w15743;
assign w15750 = w15748 & ~w15749;
assign w15751 = ~w15737 & ~w15741;
assign w15752 = ~w15739 & w15751;
assign w15753 = ~w15750 & w15752;
assign w15754 = ~w15747 & w15753;
assign w15755 = w15721 & w15726;
assign w15756 = ~w15696 & ~w15708;
assign w15757 = ~w15755 & ~w15756;
assign w15758 = ~w15713 & ~w15743;
assign w15759 = ~w15757 & ~w15758;
assign w15760 = w15690 & w15708;
assign w15761 = w15696 & ~w15712;
assign w15762 = ~w15760 & w15761;
assign w15763 = ~w15738 & ~w15762;
assign w15764 = ~w15718 & ~w15763;
assign w15765 = w15737 & ~w15759;
assign w15766 = ~w15764 & w15765;
assign w15767 = ~w15754 & ~w15766;
assign w15768 = ~w15717 & ~w15731;
assign w15769 = ~w15767 & w15768;
assign w15770 = pi0866 & ~w15769;
assign w15771 = ~pi0866 & w15769;
assign w15772 = ~w15770 & ~w15771;
assign w15773 = ~pi3754 & pi9040;
assign w15774 = ~pi3743 & ~pi9040;
assign w15775 = ~w15773 & ~w15774;
assign w15776 = pi0859 & ~w15775;
assign w15777 = ~pi0859 & w15775;
assign w15778 = ~w15776 & ~w15777;
assign w15779 = ~pi3773 & pi9040;
assign w15780 = ~pi3716 & ~pi9040;
assign w15781 = ~w15779 & ~w15780;
assign w15782 = pi0844 & ~w15781;
assign w15783 = ~pi0844 & w15781;
assign w15784 = ~w15782 & ~w15783;
assign w15785 = ~w15778 & w15784;
assign w15786 = w15778 & ~w15784;
assign w15787 = ~w15785 & ~w15786;
assign w15788 = ~pi3749 & pi9040;
assign w15789 = ~pi3738 & ~pi9040;
assign w15790 = ~w15788 & ~w15789;
assign w15791 = pi0837 & ~w15790;
assign w15792 = ~pi0837 & w15790;
assign w15793 = ~w15791 & ~w15792;
assign w15794 = w15787 & w15793;
assign w15795 = ~pi3766 & pi9040;
assign w15796 = ~pi3773 & ~pi9040;
assign w15797 = ~w15795 & ~w15796;
assign w15798 = pi0852 & ~w15797;
assign w15799 = ~pi0852 & w15797;
assign w15800 = ~w15798 & ~w15799;
assign w15801 = w15794 & ~w15800;
assign w15802 = ~pi3726 & pi9040;
assign w15803 = ~pi3758 & ~pi9040;
assign w15804 = ~w15802 & ~w15803;
assign w15805 = pi0835 & ~w15804;
assign w15806 = ~pi0835 & w15804;
assign w15807 = ~w15805 & ~w15806;
assign w15808 = ~pi3722 & pi9040;
assign w15809 = ~pi3725 & ~pi9040;
assign w15810 = ~w15808 & ~w15809;
assign w15811 = pi0828 & ~w15810;
assign w15812 = ~pi0828 & w15810;
assign w15813 = ~w15811 & ~w15812;
assign w15814 = ~w15793 & w15813;
assign w15815 = w15785 & w15814;
assign w15816 = ~w15778 & w15813;
assign w15817 = ~w15793 & w15800;
assign w15818 = w15784 & w15793;
assign w15819 = ~w15817 & ~w15818;
assign w15820 = w15816 & ~w15819;
assign w15821 = ~w15784 & ~w15813;
assign w15822 = ~w15818 & ~w15821;
assign w15823 = ~w15784 & ~w15793;
assign w15824 = w15778 & ~w15813;
assign w15825 = ~w15816 & ~w15824;
assign w15826 = w15823 & w15825;
assign w15827 = ~w15794 & ~w15826;
assign w15828 = w15822 & ~w15827;
assign w15829 = (~w15820 & w15827) | (~w15820 & w63698) | (w15827 & w63698);
assign w15830 = w15778 & w15800;
assign w15831 = ~w15823 & w15830;
assign w15832 = w15822 & w15831;
assign w15833 = ~w15778 & ~w15813;
assign w15834 = w15823 & w15833;
assign w15835 = ~w15815 & ~w15834;
assign w15836 = ~w15832 & w15835;
assign w15837 = (w15836 & w15829) | (w15836 & w65199) | (w15829 & w65199);
assign w15838 = w15807 & ~w15837;
assign w15839 = ~w15793 & ~w15813;
assign w15840 = w15785 & w15839;
assign w15841 = w15787 & w15813;
assign w15842 = (~w15817 & w15841) | (~w15817 & w65200) | (w15841 & w65200);
assign w15843 = ~w15800 & w15822;
assign w15844 = w15778 & ~w15831;
assign w15845 = ~w15843 & w15844;
assign w15846 = ~w15842 & ~w15845;
assign w15847 = ~w15807 & ~w15846;
assign w15848 = w15793 & w15813;
assign w15849 = ~w15839 & ~w15848;
assign w15850 = w15785 & w15849;
assign w15851 = ~w15785 & w15839;
assign w15852 = ~w15850 & ~w15851;
assign w15853 = w15800 & ~w15852;
assign w15854 = ~w15801 & ~w15853;
assign w15855 = ~w15847 & w15854;
assign w15856 = ~w15838 & w15855;
assign w15857 = pi0884 & w15856;
assign w15858 = ~pi0884 & ~w15856;
assign w15859 = ~w15857 & ~w15858;
assign w15860 = ~pi3774 & pi9040;
assign w15861 = ~pi3754 & ~pi9040;
assign w15862 = ~w15860 & ~w15861;
assign w15863 = pi0859 & ~w15862;
assign w15864 = ~pi0859 & w15862;
assign w15865 = ~w15863 & ~w15864;
assign w15866 = ~pi3715 & pi9040;
assign w15867 = ~pi3746 & ~pi9040;
assign w15868 = ~w15866 & ~w15867;
assign w15869 = pi0837 & ~w15868;
assign w15870 = ~pi0837 & w15868;
assign w15871 = ~w15869 & ~w15870;
assign w15872 = ~pi3733 & pi9040;
assign w15873 = ~pi3714 & ~pi9040;
assign w15874 = ~w15872 & ~w15873;
assign w15875 = pi0840 & ~w15874;
assign w15876 = ~pi0840 & w15874;
assign w15877 = ~w15875 & ~w15876;
assign w15878 = ~w15871 & w15877;
assign w15879 = ~pi3769 & pi9040;
assign w15880 = ~pi3747 & ~pi9040;
assign w15881 = ~w15879 & ~w15880;
assign w15882 = pi0851 & ~w15881;
assign w15883 = ~pi0851 & w15881;
assign w15884 = ~w15882 & ~w15883;
assign w15885 = ~pi3747 & pi9040;
assign w15886 = ~pi3726 & ~pi9040;
assign w15887 = ~w15885 & ~w15886;
assign w15888 = pi0834 & ~w15887;
assign w15889 = ~pi0834 & w15887;
assign w15890 = ~w15888 & ~w15889;
assign w15891 = w15884 & ~w15890;
assign w15892 = ~w15871 & ~w15891;
assign w15893 = w15877 & w15890;
assign w15894 = (~w15878 & w15892) | (~w15878 & w63699) | (w15892 & w63699);
assign w15895 = ~w15884 & w15890;
assign w15896 = w15894 & w15895;
assign w15897 = ~pi3758 & pi9040;
assign w15898 = ~pi3766 & ~pi9040;
assign w15899 = ~w15897 & ~w15898;
assign w15900 = pi0856 & ~w15899;
assign w15901 = ~pi0856 & w15899;
assign w15902 = ~w15900 & ~w15901;
assign w15903 = ~w15890 & ~w15902;
assign w15904 = w15878 & w15903;
assign w15905 = ~w15877 & ~w15884;
assign w15906 = w15871 & ~w15890;
assign w15907 = w15905 & w15906;
assign w15908 = ~w15904 & ~w15907;
assign w15909 = ~w15896 & w15908;
assign w15910 = w15871 & w15877;
assign w15911 = w15884 & w15910;
assign w15912 = (w15902 & ~w15910) | (w15902 & w63700) | (~w15910 & w63700);
assign w15913 = w15878 & w15884;
assign w15914 = w15878 & w63701;
assign w15915 = ~w15877 & w15884;
assign w15916 = w15871 & w15915;
assign w15917 = ~w15871 & w15905;
assign w15918 = ~w15916 & ~w15917;
assign w15919 = w15890 & ~w15918;
assign w15920 = (~w15914 & w15918) | (~w15914 & w65201) | (w15918 & w65201);
assign w15921 = (w15912 & w15919) | (w15912 & w63702) | (w15919 & w63702);
assign w15922 = ~w15914 & ~w15915;
assign w15923 = w15921 & ~w15922;
assign w15924 = w15894 & ~w15902;
assign w15925 = w15909 & ~w15924;
assign w15926 = ~w15923 & w15925;
assign w15927 = w15865 & ~w15926;
assign w15928 = w15891 & w15902;
assign w15929 = ~w15865 & w15890;
assign w15930 = w15905 & w15929;
assign w15931 = ~w15928 & ~w15930;
assign w15932 = w15871 & ~w15931;
assign w15933 = w15878 & ~w15884;
assign w15934 = w15878 & w65202;
assign w15935 = ~w15878 & ~w15905;
assign w15936 = ~w15890 & w15935;
assign w15937 = ~w15914 & ~w15936;
assign w15938 = ~w15936 & w65203;
assign w15939 = ~w15865 & ~w15938;
assign w15940 = ~w15921 & w15939;
assign w15941 = ~w15932 & ~w15934;
assign w15942 = ~w15940 & w15941;
assign w15943 = ~w15927 & w65204;
assign w15944 = (~pi0869 & w15927) | (~pi0869 & w65205) | (w15927 & w65205);
assign w15945 = ~w15943 & ~w15944;
assign w15946 = ~pi3728 & pi9040;
assign w15947 = ~pi3729 & ~pi9040;
assign w15948 = ~w15946 & ~w15947;
assign w15949 = pi0819 & ~w15948;
assign w15950 = ~pi0819 & w15948;
assign w15951 = ~w15949 & ~w15950;
assign w15952 = ~pi3721 & pi9040;
assign w15953 = ~pi3772 & ~pi9040;
assign w15954 = ~w15952 & ~w15953;
assign w15955 = pi0863 & ~w15954;
assign w15956 = ~pi0863 & w15954;
assign w15957 = ~w15955 & ~w15956;
assign w15958 = w15951 & w15957;
assign w15959 = ~w15951 & ~w15957;
assign w15960 = ~w15958 & ~w15959;
assign w15961 = ~pi3741 & pi9040;
assign w15962 = ~pi3723 & ~pi9040;
assign w15963 = ~w15961 & ~w15962;
assign w15964 = pi0850 & ~w15963;
assign w15965 = ~pi0850 & w15963;
assign w15966 = ~w15964 & ~w15965;
assign w15967 = ~w15951 & w15966;
assign w15968 = w15951 & ~w15966;
assign w15969 = ~w15967 & ~w15968;
assign w15970 = ~pi3740 & pi9040;
assign w15971 = ~pi3737 & ~pi9040;
assign w15972 = ~w15970 & ~w15971;
assign w15973 = pi0860 & ~w15972;
assign w15974 = ~pi0860 & w15972;
assign w15975 = ~w15973 & ~w15974;
assign w15976 = w15957 & w15975;
assign w15977 = w15969 & ~w15976;
assign w15978 = ~w15960 & ~w15977;
assign w15979 = ~w15957 & ~w15975;
assign w15980 = ~w15968 & w15979;
assign w15981 = ~w15978 & ~w15980;
assign w15982 = ~pi3711 & pi9040;
assign w15983 = ~pi3736 & ~pi9040;
assign w15984 = ~w15982 & ~w15983;
assign w15985 = pi0841 & ~w15984;
assign w15986 = ~pi0841 & w15984;
assign w15987 = ~w15985 & ~w15986;
assign w15988 = w15960 & w15987;
assign w15989 = w15969 & w15975;
assign w15990 = (~w15975 & ~w15969) | (~w15975 & w63378) | (~w15969 & w63378);
assign w15991 = w15966 & w15975;
assign w15992 = ~w15987 & w15991;
assign w15993 = ~w15989 & ~w15992;
assign w15994 = ~w15990 & w15993;
assign w15995 = w15957 & w15988;
assign w15996 = w15994 & w15995;
assign w15997 = ~w15960 & ~w15966;
assign w15998 = w15960 & w15966;
assign w15999 = ~w15997 & ~w15998;
assign w16000 = ~w15966 & ~w15987;
assign w16001 = ~w15957 & ~w16000;
assign w16002 = w15957 & ~w15987;
assign w16003 = w15968 & w16002;
assign w16004 = ~w16001 & ~w16003;
assign w16005 = ~w15979 & ~w16004;
assign w16006 = ~w15999 & w16005;
assign w16007 = (w15988 & w15996) | (w15988 & w63379) | (w15996 & w63379);
assign w16008 = ~pi3775 & pi9040;
assign w16009 = ~pi3718 & ~pi9040;
assign w16010 = ~w16008 & ~w16009;
assign w16011 = pi0842 & ~w16010;
assign w16012 = ~pi0842 & w16010;
assign w16013 = ~w16011 & ~w16012;
assign w16014 = (~w16013 & w16007) | (~w16013 & w63703) | (w16007 & w63703);
assign w16015 = w15966 & ~w15975;
assign w16016 = w15957 & w16015;
assign w16017 = ~w15960 & ~w15975;
assign w16018 = (w15968 & w15960) | (w15968 & w63380) | (w15960 & w63380);
assign w16019 = ~w16016 & ~w16018;
assign w16020 = w15959 & w15991;
assign w16021 = ~w15957 & ~w15966;
assign w16022 = (w15987 & w16020) | (w15987 & w63704) | (w16020 & w63704);
assign w16023 = ~w15967 & ~w15979;
assign w16024 = w15960 & ~w15987;
assign w16025 = w16023 & w16024;
assign w16026 = ~w16022 & ~w16025;
assign w16027 = (w16013 & ~w16026) | (w16013 & w63705) | (~w16026 & w63705);
assign w16028 = w15987 & w15997;
assign w16029 = w15989 & w16028;
assign w16030 = ~w15951 & ~w15987;
assign w16031 = w16015 & w16030;
assign w16032 = w15951 & w15987;
assign w16033 = (~w15975 & w16018) | (~w15975 & w63706) | (w16018 & w63706);
assign w16034 = (w16018 & w65206) | (w16018 & w65207) | (w65206 & w65207);
assign w16035 = w15976 & w16000;
assign w16036 = ~w16031 & ~w16035;
assign w16037 = ~w16034 & w16036;
assign w16038 = ~w16027 & w65208;
assign w16039 = ~w16014 & w65209;
assign w16040 = (~pi0867 & w16014) | (~pi0867 & w65210) | (w16014 & w65210);
assign w16041 = ~w16039 & ~w16040;
assign w16042 = w15833 & w15852;
assign w16043 = w15823 & w15824;
assign w16044 = w15778 & w15784;
assign w16045 = w15849 & ~w16044;
assign w16046 = ~w15800 & ~w16045;
assign w16047 = w15814 & w16044;
assign w16048 = ~w15807 & ~w16043;
assign w16049 = ~w16047 & w16048;
assign w16050 = ~w15820 & w16049;
assign w16051 = ~w16046 & w16050;
assign w16052 = ~w16042 & w16051;
assign w16053 = ~w15814 & ~w15821;
assign w16054 = ~w15852 & w16053;
assign w16055 = ~w15800 & w15807;
assign w16056 = ~w15815 & w16055;
assign w16057 = w15778 & w15793;
assign w16058 = w15800 & w15807;
assign w16059 = ~w16057 & w16058;
assign w16060 = ~w15834 & w16059;
assign w16061 = ~w16056 & ~w16060;
assign w16062 = ~w15828 & ~w16061;
assign w16063 = ~w16054 & w16062;
assign w16064 = ~w16052 & ~w16063;
assign w16065 = pi0879 & w16064;
assign w16066 = ~pi0879 & ~w16064;
assign w16067 = ~w16065 & ~w16066;
assign w16068 = ~w15689 & ~w15708;
assign w16069 = w15696 & ~w16068;
assign w16070 = ~w15683 & w15696;
assign w16071 = w15690 & w15748;
assign w16072 = ~w16070 & ~w16071;
assign w16073 = ~w16069 & ~w16072;
assign w16074 = w15683 & ~w15696;
assign w16075 = ~w15726 & ~w16070;
assign w16076 = ~w15708 & ~w16075;
assign w16077 = ~w15719 & ~w16076;
assign w16078 = w16074 & ~w16077;
assign w16079 = ~w15702 & ~w15743;
assign w16080 = w15702 & w16068;
assign w16081 = ~w15740 & ~w16080;
assign w16082 = w15722 & ~w16081;
assign w16083 = (w15737 & ~w15762) | (w15737 & w65211) | (~w15762 & w65211);
assign w16084 = ~w16082 & w16083;
assign w16085 = ~w16078 & w16084;
assign w16086 = ~w15689 & ~w15744;
assign w16087 = w15713 & ~w16086;
assign w16088 = w15683 & ~w15748;
assign w16089 = w16069 & w16088;
assign w16090 = (~w15696 & w15724) | (~w15696 & w65212) | (w15724 & w65212);
assign w16091 = ~w15737 & ~w15745;
assign w16092 = ~w16071 & w16091;
assign w16093 = ~w16087 & ~w16089;
assign w16094 = w16092 & w16093;
assign w16095 = ~w16090 & w16094;
assign w16096 = ~w16085 & ~w16095;
assign w16097 = ~w16073 & ~w16096;
assign w16098 = ~pi0889 & w16097;
assign w16099 = pi0889 & ~w16097;
assign w16100 = ~w16098 & ~w16099;
assign w16101 = ~pi3732 & pi9040;
assign w16102 = ~pi3741 & ~pi9040;
assign w16103 = ~w16101 & ~w16102;
assign w16104 = pi0853 & ~w16103;
assign w16105 = ~pi0853 & w16103;
assign w16106 = ~w16104 & ~w16105;
assign w16107 = ~pi3723 & pi9040;
assign w16108 = ~pi3711 & ~pi9040;
assign w16109 = ~w16107 & ~w16108;
assign w16110 = pi0819 & ~w16109;
assign w16111 = ~pi0819 & w16109;
assign w16112 = ~w16110 & ~w16111;
assign w16113 = ~pi3756 & pi9040;
assign w16114 = ~pi3713 & ~pi9040;
assign w16115 = ~w16113 & ~w16114;
assign w16116 = pi0861 & ~w16115;
assign w16117 = ~pi0861 & w16115;
assign w16118 = ~w16116 & ~w16117;
assign w16119 = w16112 & ~w16118;
assign w16120 = ~pi3739 & pi9040;
assign w16121 = ~pi3734 & ~pi9040;
assign w16122 = ~w16120 & ~w16121;
assign w16123 = pi0857 & ~w16122;
assign w16124 = ~pi0857 & w16122;
assign w16125 = ~w16123 & ~w16124;
assign w16126 = ~pi3777 & pi9040;
assign w16127 = ~pi3721 & ~pi9040;
assign w16128 = ~w16126 & ~w16127;
assign w16129 = pi0842 & ~w16128;
assign w16130 = ~pi0842 & w16128;
assign w16131 = ~w16129 & ~w16130;
assign w16132 = w16125 & w16131;
assign w16133 = w16119 & w16132;
assign w16134 = ~w16112 & w16125;
assign w16135 = ~w16112 & w16118;
assign w16136 = w16131 & ~w16135;
assign w16137 = ~w16134 & w16136;
assign w16138 = w16118 & ~w16131;
assign w16139 = ~w16112 & w16138;
assign w16140 = ~w16137 & ~w16139;
assign w16141 = ~pi3713 & pi9040;
assign w16142 = ~pi3730 & ~pi9040;
assign w16143 = ~w16141 & ~w16142;
assign w16144 = pi0845 & ~w16143;
assign w16145 = ~pi0845 & w16143;
assign w16146 = ~w16144 & ~w16145;
assign w16147 = ~w16140 & ~w16146;
assign w16148 = w16125 & ~w16131;
assign w16149 = ~w16112 & w16148;
assign w16150 = ~w16133 & ~w16149;
assign w16151 = ~w16147 & w16150;
assign w16152 = ~w16106 & ~w16151;
assign w16153 = ~w16125 & w16131;
assign w16154 = ~w16106 & ~w16135;
assign w16155 = w16153 & ~w16154;
assign w16156 = ~w16112 & ~w16118;
assign w16157 = w16131 & w16156;
assign w16158 = w16119 & ~w16131;
assign w16159 = ~w16157 & ~w16158;
assign w16160 = ~w16125 & w16158;
assign w16161 = w16118 & w16132;
assign w16162 = w16106 & ~w16161;
assign w16163 = ~w16160 & w16162;
assign w16164 = ~w16159 & w16163;
assign w16165 = ~w16106 & ~w16131;
assign w16166 = ~w16118 & ~w16125;
assign w16167 = w16112 & w16138;
assign w16168 = ~w16166 & ~w16167;
assign w16169 = w16165 & ~w16168;
assign w16170 = w16135 & w16148;
assign w16171 = w16112 & w16118;
assign w16172 = w16106 & ~w16138;
assign w16173 = w16171 & w16172;
assign w16174 = w16146 & ~w16170;
assign w16175 = ~w16155 & w16174;
assign w16176 = ~w16173 & w16175;
assign w16177 = ~w16169 & w16176;
assign w16178 = ~w16164 & w16177;
assign w16179 = ~w16112 & w16161;
assign w16180 = ~w16133 & ~w16146;
assign w16181 = ~w16179 & w16180;
assign w16182 = ~w16153 & ~w16165;
assign w16183 = ~w16168 & w16182;
assign w16184 = ~w16118 & w16149;
assign w16185 = w16181 & ~w16184;
assign w16186 = ~w16183 & w16185;
assign w16187 = ~w16178 & ~w16186;
assign w16188 = ~w16187 & w65213;
assign w16189 = (pi0864 & w16187) | (pi0864 & w65214) | (w16187 & w65214);
assign w16190 = ~w16188 & ~w16189;
assign w16191 = w15871 & w15905;
assign w16192 = w15877 & w15891;
assign w16193 = ~w16191 & ~w16192;
assign w16194 = w15902 & ~w16193;
assign w16195 = ~w15871 & w15891;
assign w16196 = ~w15907 & ~w16195;
assign w16197 = ~w15919 & w16196;
assign w16198 = (w15865 & ~w16197) | (w15865 & w65215) | (~w16197 & w65215);
assign w16199 = ~w15877 & ~w15890;
assign w16200 = (w15902 & w16191) | (w15902 & w65216) | (w16191 & w65216);
assign w16201 = ~w15893 & ~w16199;
assign w16202 = w15884 & ~w15902;
assign w16203 = w16201 & w16202;
assign w16204 = ~w16200 & ~w16203;
assign w16205 = ~w15909 & ~w16204;
assign w16206 = ~w15865 & ~w15918;
assign w16207 = ~w15865 & ~w15906;
assign w16208 = w15877 & ~w15884;
assign w16209 = ~w16207 & w16208;
assign w16210 = (~w15902 & w16206) | (~w15902 & w65217) | (w16206 & w65217);
assign w16211 = w15890 & w15911;
assign w16212 = ~w15905 & ~w16192;
assign w16213 = (w15902 & ~w15915) | (w15902 & w65218) | (~w15915 & w65218);
assign w16214 = w16212 & w16213;
assign w16215 = (~w15865 & w16214) | (~w15865 & w65219) | (w16214 & w65219);
assign w16216 = ~w16210 & ~w16215;
assign w16217 = ~w16198 & w16216;
assign w16218 = ~w16205 & w16217;
assign w16219 = pi0870 & ~w16218;
assign w16220 = ~pi0870 & w16218;
assign w16221 = ~w16219 & ~w16220;
assign w16222 = ~w15892 & w15935;
assign w16223 = ~w15906 & w16222;
assign w16224 = w16214 & w16223;
assign w16225 = ~w15890 & w15924;
assign w16226 = w15877 & w15902;
assign w16227 = w15895 & w16226;
assign w16228 = w15895 & w15910;
assign w16229 = ~w15913 & ~w16228;
assign w16230 = w15937 & ~w16229;
assign w16231 = ~w15865 & ~w15904;
assign w16232 = ~w16227 & w16231;
assign w16233 = w16204 & w16232;
assign w16234 = ~w16230 & w16233;
assign w16235 = ~w16192 & w63707;
assign w16236 = (~w15902 & w15935) | (~w15902 & w15903) | (w15935 & w15903);
assign w16237 = ~w16235 & w16236;
assign w16238 = w15890 & w15915;
assign w16239 = w15912 & ~w16238;
assign w16240 = ~w15934 & w16239;
assign w16241 = ~w16237 & ~w16240;
assign w16242 = w15865 & ~w16241;
assign w16243 = ~w16205 & w16242;
assign w16244 = ~w16224 & ~w16225;
assign w16245 = (w16244 & w16243) | (w16244 & w65220) | (w16243 & w65220);
assign w16246 = pi0878 & ~w16245;
assign w16247 = ~pi0878 & w16245;
assign w16248 = ~w16246 & ~w16247;
assign w16249 = w15967 & w16002;
assign w16250 = w16013 & ~w16249;
assign w16251 = ~w15975 & ~w16002;
assign w16252 = ~w16001 & w16251;
assign w16253 = w15975 & ~w16004;
assign w16254 = w15966 & w16032;
assign w16255 = w16250 & ~w16254;
assign w16256 = ~w16252 & w16255;
assign w16257 = ~w16253 & w16256;
assign w16258 = (w15991 & ~w16026) | (w15991 & w65221) | (~w16026 & w65221);
assign w16259 = w15966 & ~w16030;
assign w16260 = w16017 & ~w16259;
assign w16261 = ~w15969 & ~w15988;
assign w16262 = ~w15977 & ~w16261;
assign w16263 = ~w16013 & ~w16260;
assign w16264 = ~w16262 & w16263;
assign w16265 = ~w16258 & w16264;
assign w16266 = ~w16257 & ~w16265;
assign w16267 = ~pi0871 & w16266;
assign w16268 = pi0871 & ~w16266;
assign w16269 = ~w16267 & ~w16268;
assign w16270 = ~pi3745 & pi9040;
assign w16271 = ~pi3751 & ~pi9040;
assign w16272 = ~w16270 & ~w16271;
assign w16273 = pi0847 & ~w16272;
assign w16274 = ~pi0847 & w16272;
assign w16275 = ~w16273 & ~w16274;
assign w16276 = ~pi3729 & pi9040;
assign w16277 = ~pi3816 & ~pi9040;
assign w16278 = ~w16276 & ~w16277;
assign w16279 = pi0839 & ~w16278;
assign w16280 = ~pi0839 & w16278;
assign w16281 = ~w16279 & ~w16280;
assign w16282 = ~w16275 & w16281;
assign w16283 = ~pi3816 & pi9040;
assign w16284 = ~pi3756 & ~pi9040;
assign w16285 = ~w16283 & ~w16284;
assign w16286 = pi0849 & ~w16285;
assign w16287 = ~pi0849 & w16285;
assign w16288 = ~w16286 & ~w16287;
assign w16289 = w16282 & ~w16288;
assign w16290 = ~pi3757 & pi9040;
assign w16291 = ~pi3777 & ~pi9040;
assign w16292 = ~w16290 & ~w16291;
assign w16293 = pi0855 & ~w16292;
assign w16294 = ~pi0855 & w16292;
assign w16295 = ~w16293 & ~w16294;
assign w16296 = w16275 & w16281;
assign w16297 = ~pi3737 & pi9040;
assign w16298 = ~pi3731 & ~pi9040;
assign w16299 = ~w16297 & ~w16298;
assign w16300 = pi0848 & ~w16299;
assign w16301 = ~pi0848 & w16299;
assign w16302 = ~w16300 & ~w16301;
assign w16303 = (~w16295 & ~w16296) | (~w16295 & w65222) | (~w16296 & w65222);
assign w16304 = ~w16289 & w16303;
assign w16305 = ~w16288 & w16302;
assign w16306 = w16275 & ~w16281;
assign w16307 = ~w16295 & ~w16302;
assign w16308 = w16288 & w16306;
assign w16309 = ~w16307 & w16308;
assign w16310 = (~w16305 & ~w16308) | (~w16305 & w65223) | (~w16308 & w65223);
assign w16311 = w16304 & ~w16310;
assign w16312 = w16281 & ~w16302;
assign w16313 = w16275 & ~w16288;
assign w16314 = w16295 & ~w16313;
assign w16315 = w16312 & w16314;
assign w16316 = w16288 & ~w16302;
assign w16317 = ~w16275 & ~w16281;
assign w16318 = ~w16305 & ~w16316;
assign w16319 = w16317 & w16318;
assign w16320 = ~w16315 & ~w16319;
assign w16321 = ~w16311 & w16320;
assign w16322 = ~w16282 & ~w16306;
assign w16323 = w16305 & ~w16322;
assign w16324 = w16295 & ~w16302;
assign w16325 = ~w16288 & w16317;
assign w16326 = w16282 & w16288;
assign w16327 = ~w16325 & ~w16326;
assign w16328 = w16324 & w16327;
assign w16329 = w16295 & w16302;
assign w16330 = ~w16325 & w16329;
assign w16331 = ~w16304 & ~w16330;
assign w16332 = ~w16328 & w16331;
assign w16333 = w16288 & w16296;
assign w16334 = w16302 & w16333;
assign w16335 = ~w16323 & ~w16334;
assign w16336 = ~w16332 & w16335;
assign w16337 = ~w16321 & ~w16336;
assign w16338 = w16307 & w16317;
assign w16339 = w16288 & w16338;
assign w16340 = w16306 & w16324;
assign w16341 = ~pi3751 & pi9040;
assign w16342 = ~pi3740 & ~pi9040;
assign w16343 = ~w16341 & ~w16342;
assign w16344 = pi0858 & ~w16343;
assign w16345 = ~pi0858 & w16343;
assign w16346 = ~w16344 & ~w16345;
assign w16347 = ~w16281 & w16302;
assign w16348 = ~w16312 & ~w16347;
assign w16349 = ~w16288 & ~w16295;
assign w16350 = ~w16348 & w16349;
assign w16351 = w16282 & w16329;
assign w16352 = w16313 & w16347;
assign w16353 = ~w16351 & ~w16352;
assign w16354 = ~w16340 & w16346;
assign w16355 = ~w16334 & w16354;
assign w16356 = ~w16339 & ~w16350;
assign w16357 = w16353 & w16356;
assign w16358 = w16355 & w16357;
assign w16359 = w16281 & w16295;
assign w16360 = ~w16316 & w16359;
assign w16361 = ~w16307 & ~w16360;
assign w16362 = w16275 & ~w16361;
assign w16363 = ~w16295 & w16326;
assign w16364 = w16317 & w16324;
assign w16365 = w16288 & w16348;
assign w16366 = w16314 & ~w16365;
assign w16367 = ~w16331 & w16366;
assign w16368 = ~w16346 & ~w16364;
assign w16369 = ~w16319 & w16368;
assign w16370 = ~w16363 & w16369;
assign w16371 = ~w16362 & w16370;
assign w16372 = ~w16367 & w16371;
assign w16373 = ~w16358 & ~w16372;
assign w16374 = ~w16373 & w65224;
assign w16375 = (pi0868 & w16373) | (pi0868 & w65225) | (w16373 & w65225);
assign w16376 = ~w16374 & ~w16375;
assign w16377 = w16112 & w16153;
assign w16378 = ~w16184 & ~w16377;
assign w16379 = w16106 & ~w16378;
assign w16380 = w16106 & ~w16148;
assign w16381 = w16112 & w16380;
assign w16382 = w16156 & ~w16182;
assign w16383 = w16153 & w16171;
assign w16384 = ~w16106 & w16125;
assign w16385 = ~w16138 & w16384;
assign w16386 = ~w16136 & w16385;
assign w16387 = ~w16106 & ~w16125;
assign w16388 = w16135 & w16387;
assign w16389 = w16148 & w16171;
assign w16390 = ~w16388 & ~w16389;
assign w16391 = w16165 & ~w16390;
assign w16392 = w16146 & ~w16381;
assign w16393 = ~w16382 & ~w16383;
assign w16394 = ~w16386 & w16393;
assign w16395 = ~w16391 & w16392;
assign w16396 = w16394 & w16395;
assign w16397 = ~w16179 & ~w16385;
assign w16398 = ~w16386 & ~w16397;
assign w16399 = ~w16119 & ~w16139;
assign w16400 = ~w16125 & ~w16399;
assign w16401 = w16135 & w16165;
assign w16402 = ~w16146 & ~w16401;
assign w16403 = w16390 & w16402;
assign w16404 = ~w16400 & w16403;
assign w16405 = ~w16398 & w16404;
assign w16406 = ~w16396 & ~w16405;
assign w16407 = ~w16379 & ~w16406;
assign w16408 = ~pi0873 & w16407;
assign w16409 = pi0873 & ~w16407;
assign w16410 = ~w16408 & ~w16409;
assign w16411 = (w15696 & w15722) | (w15696 & w65226) | (w15722 & w65226);
assign w16412 = ~w15744 & w16411;
assign w16413 = w15719 & w15720;
assign w16414 = ~w16412 & ~w16413;
assign w16415 = ~w15737 & ~w16414;
assign w16416 = ~w15748 & w16086;
assign w16417 = w15713 & w16075;
assign w16418 = ~w16416 & w16417;
assign w16419 = ~w15745 & ~w15755;
assign w16420 = ~w16080 & w16419;
assign w16421 = w16070 & ~w16420;
assign w16422 = ~w15689 & w15737;
assign w16423 = ~w15708 & w16074;
assign w16424 = ~w16422 & w16423;
assign w16425 = ~w15747 & w16076;
assign w16426 = w15721 & w15740;
assign w16427 = ~w15760 & ~w16426;
assign w16428 = ~w16425 & w16427;
assign w16429 = w15737 & ~w16428;
assign w16430 = ~w16418 & ~w16424;
assign w16431 = ~w16421 & w16430;
assign w16432 = ~w16415 & w16431;
assign w16433 = ~w16429 & w16432;
assign w16434 = pi0894 & ~w16433;
assign w16435 = ~pi0894 & w16433;
assign w16436 = ~w16434 & ~w16435;
assign w16437 = w15871 & w16199;
assign w16438 = w16229 & ~w16437;
assign w16439 = (~w15865 & ~w16229) | (~w15865 & w65227) | (~w16229 & w65227);
assign w16440 = w15920 & ~w16439;
assign w16441 = w15902 & ~w16440;
assign w16442 = w15903 & w15910;
assign w16443 = ~w15934 & ~w16442;
assign w16444 = ~w15865 & ~w16443;
assign w16445 = w16229 & w65228;
assign w16446 = ~w15877 & w16207;
assign w16447 = w15918 & w16446;
assign w16448 = ~w16445 & ~w16447;
assign w16449 = ~w15902 & ~w16448;
assign w16450 = w15903 & ~w15933;
assign w16451 = (~w16450 & ~w16438) | (~w16450 & w65229) | (~w16438 & w65229);
assign w16452 = w15865 & ~w16442;
assign w16453 = ~w16451 & w16452;
assign w16454 = ~w16441 & ~w16444;
assign w16455 = ~w16449 & ~w16453;
assign w16456 = w16454 & w16455;
assign w16457 = ~pi0865 & ~w16456;
assign w16458 = pi0865 & w16456;
assign w16459 = ~w16457 & ~w16458;
assign w16460 = ~pi3743 & pi9040;
assign w16461 = ~pi3753 & ~pi9040;
assign w16462 = ~w16460 & ~w16461;
assign w16463 = pi0851 & ~w16462;
assign w16464 = ~pi0851 & w16462;
assign w16465 = ~w16463 & ~w16464;
assign w16466 = ~pi3742 & pi9040;
assign w16467 = ~pi3765 & ~pi9040;
assign w16468 = ~w16466 & ~w16467;
assign w16469 = pi0847 & ~w16468;
assign w16470 = ~pi0847 & w16468;
assign w16471 = ~w16469 & ~w16470;
assign w16472 = ~pi3746 & pi9040;
assign w16473 = ~pi3768 & ~pi9040;
assign w16474 = ~w16472 & ~w16473;
assign w16475 = pi0862 & ~w16474;
assign w16476 = ~pi0862 & w16474;
assign w16477 = ~w16475 & ~w16476;
assign w16478 = ~w16471 & w16477;
assign w16479 = w16471 & ~w16477;
assign w16480 = ~w16478 & ~w16479;
assign w16481 = ~pi3714 & pi9040;
assign w16482 = ~pi3742 & ~pi9040;
assign w16483 = ~w16481 & ~w16482;
assign w16484 = pi0858 & ~w16483;
assign w16485 = ~pi0858 & w16483;
assign w16486 = ~w16484 & ~w16485;
assign w16487 = w16465 & w16486;
assign w16488 = ~pi3748 & pi9040;
assign w16489 = ~pi3715 & ~pi9040;
assign w16490 = ~w16488 & ~w16489;
assign w16491 = pi0836 & ~w16490;
assign w16492 = ~pi0836 & w16490;
assign w16493 = ~w16491 & ~w16492;
assign w16494 = w16477 & w16493;
assign w16495 = w16487 & ~w16494;
assign w16496 = ~w16465 & w16486;
assign w16497 = w16471 & w16477;
assign w16498 = ~w16496 & ~w16497;
assign w16499 = w16471 & w16486;
assign w16500 = ~w16493 & ~w16499;
assign w16501 = ~w16498 & w16500;
assign w16502 = (~w16480 & w16501) | (~w16480 & w65230) | (w16501 & w65230);
assign w16503 = ~w16465 & w16502;
assign w16504 = ~pi3735 & pi9040;
assign w16505 = ~pi3733 & ~pi9040;
assign w16506 = ~w16504 & ~w16505;
assign w16507 = pi0840 & ~w16506;
assign w16508 = ~pi0840 & w16506;
assign w16509 = ~w16507 & ~w16508;
assign w16510 = ~w16477 & ~w16486;
assign w16511 = ~w16465 & ~w16510;
assign w16512 = w16480 & w16511;
assign w16513 = ~w16471 & ~w16486;
assign w16514 = w16465 & w16513;
assign w16515 = w16465 & ~w16477;
assign w16516 = ~w16496 & ~w16515;
assign w16517 = (w16516 & w16512) | (w16516 & w63708) | (w16512 & w63708);
assign w16518 = w16465 & ~w16486;
assign w16519 = ~w16511 & ~w16518;
assign w16520 = ~w16511 & w65231;
assign w16521 = w16493 & w16520;
assign w16522 = ~w16477 & ~w16493;
assign w16523 = w16486 & w16522;
assign w16524 = ~w16517 & ~w16523;
assign w16525 = (w16509 & ~w16524) | (w16509 & w65232) | (~w16524 & w65232);
assign w16526 = w16496 & w16497;
assign w16527 = w16465 & w16479;
assign w16528 = ~w16526 & ~w16527;
assign w16529 = ~w16517 & w16528;
assign w16530 = ~w16477 & w16512;
assign w16531 = (w16493 & ~w16512) | (w16493 & w16494) | (~w16512 & w16494);
assign w16532 = w16471 & w16487;
assign w16533 = (~w16512 & w65233) | (~w16512 & w65234) | (w65233 & w65234);
assign w16534 = ~w16529 & w16533;
assign w16535 = ~w16471 & w16487;
assign w16536 = (~w16493 & ~w16487) | (~w16493 & w65235) | (~w16487 & w65235);
assign w16537 = ~w16477 & w16518;
assign w16538 = w16536 & ~w16537;
assign w16539 = ~w16533 & ~w16538;
assign w16540 = w16471 & w16510;
assign w16541 = w16478 & ~w16496;
assign w16542 = ~w16465 & w16541;
assign w16543 = w16471 & w16518;
assign w16544 = ~w16493 & w16543;
assign w16545 = ~w16526 & ~w16540;
assign w16546 = ~w16542 & w16545;
assign w16547 = ~w16544 & w16546;
assign w16548 = ~w16539 & w16547;
assign w16549 = ~w16509 & ~w16548;
assign w16550 = ~w16503 & ~w16534;
assign w16551 = ~w16525 & w16550;
assign w16552 = (~pi0875 & ~w16551) | (~pi0875 & w65236) | (~w16551 & w65236);
assign w16553 = w16551 & w65237;
assign w16554 = ~w16552 & ~w16553;
assign w16555 = ~w16106 & ~w16167;
assign w16556 = ~w16163 & ~w16555;
assign w16557 = w16112 & ~w16384;
assign w16558 = w16131 & ~w16156;
assign w16559 = ~w16134 & ~w16557;
assign w16560 = ~w16558 & w16559;
assign w16561 = ~w16173 & w16181;
assign w16562 = ~w16560 & w16561;
assign w16563 = w16118 & w16153;
assign w16564 = ~w16157 & ~w16563;
assign w16565 = ~w16106 & ~w16564;
assign w16566 = w16106 & ~w16399;
assign w16567 = w16146 & ~w16184;
assign w16568 = ~w16565 & w16567;
assign w16569 = ~w16566 & w16568;
assign w16570 = ~w16562 & ~w16569;
assign w16571 = ~w16556 & ~w16570;
assign w16572 = ~pi0902 & w16571;
assign w16573 = pi0902 & ~w16571;
assign w16574 = ~w16572 & ~w16573;
assign w16575 = w16480 & w16495;
assign w16576 = ~w16480 & w16519;
assign w16577 = ~w16512 & w63709;
assign w16578 = ~w16576 & w16577;
assign w16579 = w16510 & w16578;
assign w16580 = (w16493 & ~w16510) | (w16493 & w65238) | (~w16510 & w65238);
assign w16581 = ~w16465 & w16471;
assign w16582 = ~w16518 & ~w16581;
assign w16583 = w16516 & w16582;
assign w16584 = w16580 & ~w16583;
assign w16585 = ~w16465 & ~w16499;
assign w16586 = ~w16583 & w65239;
assign w16587 = ~w16480 & w16496;
assign w16588 = ~w16575 & ~w16587;
assign w16589 = ~w16586 & w16588;
assign w16590 = (w16509 & w16579) | (w16509 & w65240) | (w16579 & w65240);
assign w16591 = ~w16493 & ~w16517;
assign w16592 = w16479 & w16496;
assign w16593 = w16493 & ~w16592;
assign w16594 = ~w16542 & w16593;
assign w16595 = ~w16591 & ~w16594;
assign w16596 = ~w16509 & ~w16584;
assign w16597 = ~w16578 & w16596;
assign w16598 = ~w16595 & ~w16597;
assign w16599 = ~w16590 & w16598;
assign w16600 = pi0880 & ~w16599;
assign w16601 = ~pi0880 & w16599;
assign w16602 = ~w16600 & ~w16601;
assign w16603 = ~w15958 & ~w15987;
assign w16604 = ~w16020 & ~w16033;
assign w16605 = w16603 & ~w16604;
assign w16606 = w16023 & ~w16037;
assign w16607 = ~w15969 & w15979;
assign w16608 = w16013 & ~w16607;
assign w16609 = ~w15996 & w63710;
assign w16610 = ~w15966 & w16030;
assign w16611 = ~w16013 & ~w16020;
assign w16612 = ~w16016 & ~w16254;
assign w16613 = ~w15976 & ~w15979;
assign w16614 = w16032 & w16613;
assign w16615 = ~w16610 & w16611;
assign w16616 = w16612 & ~w16614;
assign w16617 = w16615 & w16616;
assign w16618 = ~w16609 & ~w16617;
assign w16619 = ~w16605 & ~w16606;
assign w16620 = (pi0882 & w16618) | (pi0882 & w65241) | (w16618 & w65241);
assign w16621 = ~w16618 & w65242;
assign w16622 = ~w16620 & ~w16621;
assign w16623 = ~w16535 & ~w16540;
assign w16624 = ~w16496 & ~w16543;
assign w16625 = w16623 & w16624;
assign w16626 = ~w16530 & ~w16625;
assign w16627 = w16493 & ~w16626;
assign w16628 = ~w16493 & ~w16623;
assign w16629 = w16528 & ~w16628;
assign w16630 = (w16509 & w16627) | (w16509 & w65243) | (w16627 & w65243);
assign w16631 = ~w16522 & ~w16543;
assign w16632 = ~w16497 & ~w16513;
assign w16633 = ~w16631 & ~w16632;
assign w16634 = ~w16477 & w16493;
assign w16635 = w16581 & w16634;
assign w16636 = ~w16501 & ~w16635;
assign w16637 = ~w16633 & w16636;
assign w16638 = w16546 & w65244;
assign w16639 = w16580 & ~w16638;
assign w16640 = (~w16502 & w16637) | (~w16502 & w65245) | (w16637 & w65245);
assign w16641 = ~w16639 & w16640;
assign w16642 = ~w16630 & w16641;
assign w16643 = ~pi0874 & w16642;
assign w16644 = pi0874 & ~w16642;
assign w16645 = ~w16643 & ~w16644;
assign w16646 = w16322 & w16349;
assign w16647 = ~w16327 & w16346;
assign w16648 = w16288 & w16295;
assign w16649 = ~w16306 & ~w16346;
assign w16650 = w16648 & w16649;
assign w16651 = ~w16646 & ~w16650;
assign w16652 = ~w16647 & w16651;
assign w16653 = w16302 & ~w16652;
assign w16654 = ~w16296 & ~w16346;
assign w16655 = ~w16313 & w16654;
assign w16656 = ~w16289 & ~w16655;
assign w16657 = w16307 & ~w16656;
assign w16658 = w16295 & w16313;
assign w16659 = w16346 & ~w16658;
assign w16660 = ~w16288 & w16312;
assign w16661 = w16353 & ~w16660;
assign w16662 = ~w16659 & ~w16661;
assign w16663 = ~w16288 & ~w16302;
assign w16664 = w16306 & w16663;
assign w16665 = ~w16333 & ~w16664;
assign w16666 = ~w16295 & ~w16665;
assign w16667 = ~w16309 & ~w16364;
assign w16668 = ~w16666 & w16667;
assign w16669 = w16346 & ~w16668;
assign w16670 = ~w16657 & ~w16662;
assign w16671 = ~w16653 & w16670;
assign w16672 = ~w16669 & w16671;
assign w16673 = pi0872 & ~w16672;
assign w16674 = ~pi0872 & w16672;
assign w16675 = ~w16673 & ~w16674;
assign w16676 = ~w15696 & w15724;
assign w16677 = ~w15721 & ~w15748;
assign w16678 = w16411 & ~w16677;
assign w16679 = ~w15716 & w16420;
assign w16680 = ~w16678 & w16679;
assign w16681 = w15737 & ~w16680;
assign w16682 = w15726 & w16074;
assign w16683 = w15696 & ~w15726;
assign w16684 = ~w16426 & w16683;
assign w16685 = ~w16416 & w16684;
assign w16686 = w15728 & ~w16682;
assign w16687 = ~w16685 & w16686;
assign w16688 = ~w15737 & ~w16687;
assign w16689 = w15744 & w16069;
assign w16690 = (~w16689 & ~w15716) | (~w16689 & w65246) | (~w15716 & w65246);
assign w16691 = ~w16676 & w16690;
assign w16692 = ~w16688 & w16691;
assign w16693 = ~w16681 & w16692;
assign w16694 = pi0900 & w16693;
assign w16695 = ~pi0900 & ~w16693;
assign w16696 = ~w16694 & ~w16695;
assign w16697 = ~pi3730 & pi9040;
assign w16698 = ~pi3739 & ~pi9040;
assign w16699 = ~w16697 & ~w16698;
assign w16700 = pi0826 & ~w16699;
assign w16701 = ~pi0826 & w16699;
assign w16702 = ~w16700 & ~w16701;
assign w16703 = ~pi3720 & pi9040;
assign w16704 = ~pi3745 & ~pi9040;
assign w16705 = ~w16703 & ~w16704;
assign w16706 = pi0861 & ~w16705;
assign w16707 = ~pi0861 & w16705;
assign w16708 = ~w16706 & ~w16707;
assign w16709 = ~pi3719 & pi9040;
assign w16710 = ~pi3720 & ~pi9040;
assign w16711 = ~w16709 & ~w16710;
assign w16712 = pi0848 & ~w16711;
assign w16713 = ~pi0848 & w16711;
assign w16714 = ~w16712 & ~w16713;
assign w16715 = ~w16708 & w16714;
assign w16716 = ~w16708 & ~w16714;
assign w16717 = ~pi3724 & pi9040;
assign w16718 = ~pi3732 & ~pi9040;
assign w16719 = ~w16717 & ~w16718;
assign w16720 = pi0845 & ~w16719;
assign w16721 = ~pi0845 & w16719;
assign w16722 = ~w16720 & ~w16721;
assign w16723 = ~w16714 & ~w16722;
assign w16724 = w16714 & w16722;
assign w16725 = ~w16723 & ~w16724;
assign w16726 = ~pi3718 & pi9040;
assign w16727 = ~pi3724 & ~pi9040;
assign w16728 = ~w16726 & ~w16727;
assign w16729 = pi0843 & ~w16728;
assign w16730 = ~pi0843 & w16728;
assign w16731 = ~w16729 & ~w16730;
assign w16732 = ~w16722 & ~w16731;
assign w16733 = ~w16716 & ~w16732;
assign w16734 = w16725 & w16733;
assign w16735 = ~w16715 & ~w16734;
assign w16736 = ~pi3734 & pi9040;
assign w16737 = ~pi3744 & ~pi9040;
assign w16738 = ~w16736 & ~w16737;
assign w16739 = pi0839 & ~w16738;
assign w16740 = ~pi0839 & w16738;
assign w16741 = ~w16739 & ~w16740;
assign w16742 = (w16741 & w16734) | (w16741 & w65247) | (w16734 & w65247);
assign w16743 = w16715 & w16731;
assign w16744 = w16716 & w16732;
assign w16745 = ~w16743 & ~w16744;
assign w16746 = ~w16742 & w16745;
assign w16747 = w16702 & ~w16746;
assign w16748 = ~w16708 & ~w16731;
assign w16749 = w16708 & w16731;
assign w16750 = ~w16748 & ~w16749;
assign w16751 = w16702 & ~w16722;
assign w16752 = ~w16743 & w16751;
assign w16753 = ~w16752 & w65248;
assign w16754 = (~w16750 & w16752) | (~w16750 & w65249) | (w16752 & w65249);
assign w16755 = ~w16753 & ~w16754;
assign w16756 = ~w16741 & w16755;
assign w16757 = w16723 & w16741;
assign w16758 = w16749 & w16757;
assign w16759 = ~w16702 & w16741;
assign w16760 = ~w16723 & w16759;
assign w16761 = w16735 & w16760;
assign w16762 = ~w16758 & ~w16761;
assign w16763 = ~w16747 & w16762;
assign w16764 = ~w16756 & w16763;
assign w16765 = pi0886 & ~w16764;
assign w16766 = ~pi0886 & w16764;
assign w16767 = ~w16765 & ~w16766;
assign w16768 = w15817 & w15833;
assign w16769 = w15807 & ~w16768;
assign w16770 = w15840 & ~w16769;
assign w16771 = w15800 & ~w15807;
assign w16772 = (w15793 & ~w15825) | (w15793 & w65250) | (~w15825 & w65250);
assign w16773 = ~w15786 & ~w15793;
assign w16774 = w15784 & ~w15824;
assign w16775 = w16773 & ~w16774;
assign w16776 = ~w16772 & ~w16775;
assign w16777 = w16055 & ~w16776;
assign w16778 = w15818 & ~w15825;
assign w16779 = w15825 & w65251;
assign w16780 = ~w16055 & ~w16773;
assign w16781 = w16779 & w16780;
assign w16782 = ~w16047 & ~w16778;
assign w16783 = ~w16781 & w16782;
assign w16784 = ~w16777 & w16783;
assign w16785 = ~w16771 & ~w16784;
assign w16786 = w16771 & ~w16778;
assign w16787 = ~w16779 & w16786;
assign w16788 = ~w16770 & ~w16787;
assign w16789 = ~w16785 & w16788;
assign w16790 = pi0908 & w16789;
assign w16791 = ~pi0908 & ~w16789;
assign w16792 = ~w16790 & ~w16791;
assign w16793 = w15989 & w16603;
assign w16794 = w15987 & w15999;
assign w16795 = w16250 & ~w16793;
assign w16796 = ~w16794 & w16795;
assign w16797 = w16612 & w16796;
assign w16798 = ~w16611 & ~w16796;
assign w16799 = w16002 & w16259;
assign w16800 = ~w16028 & ~w16799;
assign w16801 = ~w15994 & w16800;
assign w16802 = ~w16798 & w16801;
assign w16803 = ~w16802 & w65252;
assign w16804 = (~pi0877 & w16802) | (~pi0877 & w65253) | (w16802 & w65253);
assign w16805 = ~w16803 & ~w16804;
assign w16806 = w16708 & w16724;
assign w16807 = w16708 & ~w16714;
assign w16808 = w16722 & ~w16731;
assign w16809 = ~w16807 & w16808;
assign w16810 = w16715 & ~w16722;
assign w16811 = ~w16806 & ~w16810;
assign w16812 = ~w16723 & w16811;
assign w16813 = (~w16702 & ~w16811) | (~w16702 & w63711) | (~w16811 & w63711);
assign w16814 = (~w16811 & w65254) | (~w16811 & w65255) | (w65254 & w65255);
assign w16815 = w16806 & w16814;
assign w16816 = ~w16725 & w16748;
assign w16817 = ~w16734 & ~w16816;
assign w16818 = ~w16702 & ~w16817;
assign w16819 = w16722 & w16731;
assign w16820 = ~w16708 & w16819;
assign w16821 = ~w16751 & ~w16820;
assign w16822 = (w16731 & ~w16819) | (w16731 & w16749) | (~w16819 & w16749);
assign w16823 = ~w16723 & w16822;
assign w16824 = ~w16816 & ~w16823;
assign w16825 = w16702 & ~w16824;
assign w16826 = (~w16748 & w16725) | (~w16748 & w63712) | (w16725 & w63712);
assign w16827 = (~w16751 & w16725) | (~w16751 & w65256) | (w16725 & w65256);
assign w16828 = ~w16826 & w16827;
assign w16829 = ~w16825 & ~w16828;
assign w16830 = (w16829 & w65257) | (w16829 & w65258) | (w65257 & w65258);
assign w16831 = w16741 & ~w16829;
assign w16832 = ~w16724 & w16749;
assign w16833 = ~w16807 & ~w16819;
assign w16834 = ~w16832 & ~w16833;
assign w16835 = w16702 & ~w16834;
assign w16836 = ~w16724 & w16817;
assign w16837 = w16836 & w63714;
assign w16838 = ~w16815 & ~w16837;
assign w16839 = ~w16831 & w16838;
assign w16840 = w16839 & w65259;
assign w16841 = (~pi0887 & ~w16839) | (~pi0887 & w65260) | (~w16839 & w65260);
assign w16842 = ~w16840 & ~w16841;
assign w16843 = ~w16133 & ~w16383;
assign w16844 = (~w16170 & w16159) | (~w16170 & w63715) | (w16159 & w63715);
assign w16845 = w16843 & w16844;
assign w16846 = w16390 & ~w16555;
assign w16847 = (~w16146 & ~w16845) | (~w16146 & w65261) | (~w16845 & w65261);
assign w16848 = w16146 & w16843;
assign w16849 = ~w16134 & w16154;
assign w16850 = ~w16172 & ~w16380;
assign w16851 = ~w16125 & w16156;
assign w16852 = ~w16850 & ~w16851;
assign w16853 = ~w16401 & ~w16849;
assign w16854 = ~w16852 & w16853;
assign w16855 = ~w16160 & w16390;
assign w16856 = w16848 & w16855;
assign w16857 = ~w16854 & w16856;
assign w16858 = ~w16847 & ~w16857;
assign w16859 = ~w16106 & ~w16848;
assign w16860 = ~w16845 & w16859;
assign w16861 = ~w16858 & ~w16860;
assign w16862 = pi0885 & w16861;
assign w16863 = ~pi0885 & ~w16861;
assign w16864 = ~w16862 & ~w16863;
assign w16865 = w16353 & w65262;
assign w16866 = w16303 & ~w16865;
assign w16867 = w16317 & w16329;
assign w16868 = w16348 & w65263;
assign w16869 = w16312 & w16658;
assign w16870 = ~w16867 & ~w16869;
assign w16871 = ~w16868 & w16870;
assign w16872 = ~w16866 & w16871;
assign w16873 = w16346 & ~w16872;
assign w16874 = ~w16281 & ~w16658;
assign w16875 = w16313 & ~w16359;
assign w16876 = ~w16305 & ~w16875;
assign w16877 = ~w16874 & ~w16876;
assign w16878 = w16320 & ~w16338;
assign w16879 = (~w16346 & ~w16878) | (~w16346 & w65264) | (~w16878 & w65264);
assign w16880 = ~w16302 & w16325;
assign w16881 = ~w16868 & ~w16880;
assign w16882 = ~w16295 & ~w16881;
assign w16883 = ~w16367 & ~w16882;
assign w16884 = ~w16879 & w16883;
assign w16885 = ~w16873 & w16884;
assign w16886 = pi0881 & w16885;
assign w16887 = ~pi0881 & ~w16885;
assign w16888 = ~w16886 & ~w16887;
assign w16889 = (w16648 & ~w16870) | (w16648 & w65265) | (~w16870 & w65265);
assign w16890 = ~w16311 & ~w16328;
assign w16891 = w16346 & ~w16890;
assign w16892 = ~w16336 & ~w16346;
assign w16893 = ~w16275 & ~w16295;
assign w16894 = ~w16346 & ~w16893;
assign w16895 = ~w16296 & ~w16894;
assign w16896 = w16365 & w16895;
assign w16897 = ~w16889 & ~w16896;
assign w16898 = ~w16891 & w16897;
assign w16899 = ~w16892 & w16898;
assign w16900 = pi0888 & ~w16899;
assign w16901 = ~pi0888 & w16899;
assign w16902 = ~w16900 & ~w16901;
assign w16903 = w15800 & w15815;
assign w16904 = w16053 & ~w16774;
assign w16905 = ~w15843 & w16904;
assign w16906 = w15825 & w15849;
assign w16907 = ~w15823 & ~w16906;
assign w16908 = ~w15800 & ~w15826;
assign w16909 = ~w16907 & w16908;
assign w16910 = w16769 & ~w16905;
assign w16911 = ~w16909 & w16910;
assign w16912 = ~w15830 & ~w16057;
assign w16913 = ~w16904 & ~w16912;
assign w16914 = ~w15800 & ~w15849;
assign w16915 = ~w16043 & w16914;
assign w16916 = ~w15807 & ~w15850;
assign w16917 = ~w16913 & w16916;
assign w16918 = ~w16915 & w16917;
assign w16919 = ~w16911 & ~w16918;
assign w16920 = w15793 & ~w15800;
assign w16921 = ~w15821 & w16920;
assign w16922 = ~w15787 & w16921;
assign w16923 = ~w16903 & ~w16922;
assign w16924 = ~w16919 & w16923;
assign w16925 = pi0913 & ~w16924;
assign w16926 = ~pi0913 & w16924;
assign w16927 = ~w16925 & ~w16926;
assign w16928 = ~w16702 & ~w16714;
assign w16929 = ~w16732 & ~w16819;
assign w16930 = w16928 & w16929;
assign w16931 = (w16731 & ~w16811) | (w16731 & w65266) | (~w16811 & w65266);
assign w16932 = ~w16722 & ~w16807;
assign w16933 = ~w16716 & ~w16751;
assign w16934 = ~w16932 & ~w16933;
assign w16935 = ~w16731 & w16811;
assign w16936 = ~w16934 & w16935;
assign w16937 = w16741 & ~w16930;
assign w16938 = (w16937 & w16936) | (w16937 & w65267) | (w16936 & w65267);
assign w16939 = w16811 & w63716;
assign w16940 = w16811 & w65268;
assign w16941 = ~w16732 & w16811;
assign w16942 = w16813 & ~w16941;
assign w16943 = ~w16741 & ~w16744;
assign w16944 = ~w16940 & w16943;
assign w16945 = ~w16942 & w16944;
assign w16946 = ~w16938 & ~w16945;
assign w16947 = w16702 & w16822;
assign w16948 = w16755 & w16947;
assign w16949 = ~w16702 & w16820;
assign w16950 = ~w16948 & ~w16949;
assign w16951 = ~w16946 & w16950;
assign w16952 = pi0876 & ~w16951;
assign w16953 = ~pi0876 & w16951;
assign w16954 = ~w16952 & ~w16953;
assign w16955 = (w16836 & w65269) | (w16836 & w65270) | (w65269 & w65270);
assign w16956 = ~w16814 & ~w16835;
assign w16957 = ~w16708 & ~w16817;
assign w16958 = ~w16956 & ~w16957;
assign w16959 = ~w16741 & ~w16958;
assign w16960 = w16749 & w16928;
assign w16961 = w16743 & w16939;
assign w16962 = w16759 & ~w16808;
assign w16963 = ~w16932 & w16962;
assign w16964 = ~w16960 & ~w16963;
assign w16965 = ~w16961 & w16964;
assign w16966 = ~w16955 & w16965;
assign w16967 = ~w16959 & w16966;
assign w16968 = pi0883 & w16967;
assign w16969 = ~pi0883 & ~w16967;
assign w16970 = ~w16968 & ~w16969;
assign w16971 = w16494 & w16514;
assign w16972 = w16479 & w16487;
assign w16973 = ~w16486 & w16581;
assign w16974 = ~w16495 & ~w16973;
assign w16975 = w16493 & ~w16974;
assign w16976 = w16478 & w16496;
assign w16977 = w16509 & ~w16972;
assign w16978 = ~w16976 & w16977;
assign w16979 = ~w16544 & w16978;
assign w16980 = ~w16975 & w16979;
assign w16981 = ~w16516 & w16536;
assign w16982 = ~w16516 & ~w16582;
assign w16983 = w16493 & ~w16982;
assign w16984 = ~w16509 & ~w16541;
assign w16985 = (w16984 & w16983) | (w16984 & w65271) | (w16983 & w65271);
assign w16986 = w16520 & w16583;
assign w16987 = ~w16493 & ~w16592;
assign w16988 = ~w16986 & w16987;
assign w16989 = ~w16531 & ~w16988;
assign w16990 = (~w16971 & w16980) | (~w16971 & w65272) | (w16980 & w65272);
assign w16991 = ~w16989 & w16990;
assign w16992 = pi0892 & ~w16991;
assign w16993 = ~pi0892 & w16991;
assign w16994 = ~w16992 & ~w16993;
assign w16995 = ~pi3801 & pi9040;
assign w16996 = ~pi3803 & ~pi9040;
assign w16997 = ~w16995 & ~w16996;
assign w16998 = pi0895 & ~w16997;
assign w16999 = ~pi0895 & w16997;
assign w17000 = ~w16998 & ~w16999;
assign w17001 = ~pi3802 & pi9040;
assign w17002 = ~pi3815 & ~pi9040;
assign w17003 = ~w17001 & ~w17002;
assign w17004 = pi0893 & ~w17003;
assign w17005 = ~pi0893 & w17003;
assign w17006 = ~w17004 & ~w17005;
assign w17007 = ~pi3806 & pi9040;
assign w17008 = ~pi3794 & ~pi9040;
assign w17009 = ~w17007 & ~w17008;
assign w17010 = pi0921 & ~w17009;
assign w17011 = ~pi0921 & w17009;
assign w17012 = ~w17010 & ~w17011;
assign w17013 = ~pi3787 & pi9040;
assign w17014 = ~pi3790 & ~pi9040;
assign w17015 = ~w17013 & ~w17014;
assign w17016 = pi0911 & ~w17015;
assign w17017 = ~pi0911 & w17015;
assign w17018 = ~w17016 & ~w17017;
assign w17019 = ~w17000 & w17018;
assign w17020 = ~pi3830 & pi9040;
assign w17021 = ~pi3835 & ~pi9040;
assign w17022 = ~w17020 & ~w17021;
assign w17023 = pi0891 & ~w17022;
assign w17024 = ~pi0891 & w17022;
assign w17025 = ~w17023 & ~w17024;
assign w17026 = w17019 & w17025;
assign w17027 = w17019 & w65273;
assign w17028 = ~w17018 & w17025;
assign w17029 = ~w17012 & w17028;
assign w17030 = ~w17027 & ~w17029;
assign w17031 = ~w17006 & ~w17030;
assign w17032 = w17000 & w17031;
assign w17033 = (~w17006 & ~w17019) | (~w17006 & w65274) | (~w17019 & w65274);
assign w17034 = ~w17018 & ~w17025;
assign w17035 = ~w17000 & w17034;
assign w17036 = w17018 & ~w17025;
assign w17037 = w17000 & w17012;
assign w17038 = w17036 & w17037;
assign w17039 = ~w17035 & ~w17038;
assign w17040 = w17000 & w17036;
assign w17041 = w17006 & ~w17040;
assign w17042 = w17000 & ~w17012;
assign w17043 = ~w17028 & ~w17042;
assign w17044 = ~w17028 & ~w17036;
assign w17045 = w17042 & ~w17044;
assign w17046 = ~w17043 & ~w17045;
assign w17047 = w17041 & ~w17046;
assign w17048 = ~pi3790 & pi9040;
assign w17049 = ~pi3802 & ~pi9040;
assign w17050 = ~w17048 & ~w17049;
assign w17051 = pi0927 & ~w17050;
assign w17052 = ~pi0927 & w17050;
assign w17053 = ~w17051 & ~w17052;
assign w17054 = (w17053 & ~w17039) | (w17053 & w65275) | (~w17039 & w65275);
assign w17055 = ~w17047 & w17054;
assign w17056 = ~w17012 & ~w17025;
assign w17057 = ~w17006 & w17056;
assign w17058 = w17025 & w17037;
assign w17059 = ~w17057 & ~w17058;
assign w17060 = w17018 & ~w17059;
assign w17061 = w17006 & ~w17042;
assign w17062 = ~w17028 & ~w17037;
assign w17063 = ~w17061 & ~w17062;
assign w17064 = ~w17060 & ~w17063;
assign w17065 = ~w17053 & ~w17064;
assign w17066 = ~w17000 & w17012;
assign w17067 = w17036 & w17066;
assign w17068 = ~w17025 & w17066;
assign w17069 = ~w17012 & w17026;
assign w17070 = ~w17068 & ~w17069;
assign w17071 = ~w17053 & ~w17070;
assign w17072 = ~w17012 & w17035;
assign w17073 = ~w17036 & ~w17066;
assign w17074 = ~w17043 & ~w17073;
assign w17075 = ~w17067 & ~w17072;
assign w17076 = ~w17074 & w17075;
assign w17077 = ~w17071 & w17076;
assign w17078 = w17006 & ~w17077;
assign w17079 = ~w17032 & ~w17055;
assign w17080 = ~w17065 & w17079;
assign w17081 = (pi0928 & ~w17080) | (pi0928 & w65276) | (~w17080 & w65276);
assign w17082 = w17080 & w65277;
assign w17083 = ~w17081 & ~w17082;
assign w17084 = ~pi3797 & pi9040;
assign w17085 = ~pi3859 & ~pi9040;
assign w17086 = ~w17084 & ~w17085;
assign w17087 = pi0917 & ~w17086;
assign w17088 = ~pi0917 & w17086;
assign w17089 = ~w17087 & ~w17088;
assign w17090 = ~pi3805 & pi9040;
assign w17091 = ~pi3854 & ~pi9040;
assign w17092 = ~w17090 & ~w17091;
assign w17093 = pi0904 & ~w17092;
assign w17094 = ~pi0904 & w17092;
assign w17095 = ~w17093 & ~w17094;
assign w17096 = ~pi3859 & pi9040;
assign w17097 = ~pi3832 & ~pi9040;
assign w17098 = ~w17096 & ~w17097;
assign w17099 = pi0922 & ~w17098;
assign w17100 = ~pi0922 & w17098;
assign w17101 = ~w17099 & ~w17100;
assign w17102 = ~w17095 & w17101;
assign w17103 = ~pi3827 & pi9040;
assign w17104 = ~pi3805 & ~pi9040;
assign w17105 = ~w17103 & ~w17104;
assign w17106 = pi0912 & ~w17105;
assign w17107 = ~pi0912 & w17105;
assign w17108 = ~w17106 & ~w17107;
assign w17109 = w17102 & w17108;
assign w17110 = w17095 & ~w17101;
assign w17111 = ~pi3831 & pi9040;
assign w17112 = ~pi3812 & ~pi9040;
assign w17113 = ~w17111 & ~w17112;
assign w17114 = pi0898 & ~w17113;
assign w17115 = ~pi0898 & w17113;
assign w17116 = ~w17114 & ~w17115;
assign w17117 = ~w17108 & ~w17116;
assign w17118 = w17110 & w17117;
assign w17119 = ~w17109 & ~w17118;
assign w17120 = w17095 & w17116;
assign w17121 = w17101 & w17120;
assign w17122 = ~pi3795 & pi9040;
assign w17123 = ~pi3796 & ~pi9040;
assign w17124 = ~w17122 & ~w17123;
assign w17125 = pi0910 & ~w17124;
assign w17126 = ~pi0910 & w17124;
assign w17127 = ~w17125 & ~w17126;
assign w17128 = (w17127 & ~w17120) | (w17127 & w65278) | (~w17120 & w65278);
assign w17129 = w17119 & w17128;
assign w17130 = w17095 & ~w17108;
assign w17131 = ~w17102 & ~w17120;
assign w17132 = w17101 & w17131;
assign w17133 = ~w17095 & ~w17116;
assign w17134 = ~w17102 & ~w17133;
assign w17135 = w17101 & w17133;
assign w17136 = ~w17134 & ~w17135;
assign w17137 = ~w17132 & ~w17136;
assign w17138 = w17108 & ~w17137;
assign w17139 = w17119 & w65279;
assign w17140 = ~w17138 & w17139;
assign w17141 = w17108 & w17131;
assign w17142 = w17108 & w17116;
assign w17143 = w17110 & w17142;
assign w17144 = ~w17132 & ~w17143;
assign w17145 = ~w17141 & ~w17144;
assign w17146 = w17101 & w17130;
assign w17147 = (~w17127 & ~w17119) | (~w17127 & w65280) | (~w17119 & w65280);
assign w17148 = ~w17145 & ~w17147;
assign w17149 = ~w17140 & w17148;
assign w17150 = ~w17089 & ~w17149;
assign w17151 = ~w17108 & ~w17127;
assign w17152 = w17101 & ~w17108;
assign w17153 = w17133 & ~w17152;
assign w17154 = w17151 & w17153;
assign w17155 = ~w17095 & ~w17101;
assign w17156 = w17116 & w17127;
assign w17157 = w17155 & w17156;
assign w17158 = w17101 & w17117;
assign w17159 = ~w17157 & ~w17158;
assign w17160 = ~w17108 & w17116;
assign w17161 = ~w17127 & ~w17160;
assign w17162 = w17130 & w17161;
assign w17163 = ~w17117 & ~w17142;
assign w17164 = w17155 & w17163;
assign w17165 = ~w17143 & ~w17162;
assign w17166 = ~w17164 & w17165;
assign w17167 = (~w17159 & ~w17165) | (~w17159 & w65281) | (~w17165 & w65281);
assign w17168 = w17108 & w17120;
assign w17169 = w17133 & w17152;
assign w17170 = ~w17168 & ~w17169;
assign w17171 = w17127 & ~w17170;
assign w17172 = ~w17102 & ~w17110;
assign w17173 = w17160 & ~w17172;
assign w17174 = ~w17127 & ~w17141;
assign w17175 = ~w17173 & w17174;
assign w17176 = w17089 & ~w17129;
assign w17177 = ~w17175 & w17176;
assign w17178 = ~w17154 & ~w17171;
assign w17179 = ~w17167 & w17178;
assign w17180 = ~w17177 & w17179;
assign w17181 = (pi0947 & w17150) | (pi0947 & w65282) | (w17150 & w65282);
assign w17182 = ~w17150 & w65283;
assign w17183 = ~w17181 & ~w17182;
assign w17184 = w17152 & w17156;
assign w17185 = w17127 & ~w17155;
assign w17186 = ~w17146 & w17185;
assign w17187 = (w17186 & ~w17137) | (w17186 & w65284) | (~w17137 & w65284);
assign w17188 = ~w17153 & ~w17168;
assign w17189 = (w17089 & w17188) | (w17089 & w65285) | (w17188 & w65285);
assign w17190 = w17166 & w17189;
assign w17191 = ~w17187 & w17190;
assign w17192 = w17142 & w17155;
assign w17193 = w17131 & w65286;
assign w17194 = ~w17127 & ~w17193;
assign w17195 = w17110 & ~w17116;
assign w17196 = ~w17141 & w17153;
assign w17197 = w17128 & ~w17195;
assign w17198 = ~w17196 & w17197;
assign w17199 = ~w17131 & w17151;
assign w17200 = ~w17089 & ~w17192;
assign w17201 = ~w17199 & w17200;
assign w17202 = (w17201 & w17198) | (w17201 & w65287) | (w17198 & w65287);
assign w17203 = ~w17118 & ~w17184;
assign w17204 = (w17203 & w17191) | (w17203 & w65288) | (w17191 & w65288);
assign w17205 = pi0943 & ~w17204;
assign w17206 = ~pi0943 & w17204;
assign w17207 = ~w17205 & ~w17206;
assign w17208 = ~pi3794 & pi9040;
assign w17209 = ~pi3830 & ~pi9040;
assign w17210 = ~w17208 & ~w17209;
assign w17211 = pi0899 & ~w17210;
assign w17212 = ~pi0899 & w17210;
assign w17213 = ~w17211 & ~w17212;
assign w17214 = ~pi3799 & pi9040;
assign w17215 = ~pi3827 & ~pi9040;
assign w17216 = ~w17214 & ~w17215;
assign w17217 = pi0917 & ~w17216;
assign w17218 = ~pi0917 & w17216;
assign w17219 = ~w17217 & ~w17218;
assign w17220 = w17213 & ~w17219;
assign w17221 = ~pi3835 & pi9040;
assign w17222 = ~pi3806 & ~pi9040;
assign w17223 = ~w17221 & ~w17222;
assign w17224 = pi0895 & ~w17223;
assign w17225 = ~pi0895 & w17223;
assign w17226 = ~w17224 & ~w17225;
assign w17227 = ~pi3803 & pi9040;
assign w17228 = ~pi3804 & ~pi9040;
assign w17229 = ~w17227 & ~w17228;
assign w17230 = pi0898 & ~w17229;
assign w17231 = ~pi0898 & w17229;
assign w17232 = ~w17230 & ~w17231;
assign w17233 = w17226 & w17232;
assign w17234 = ~w17226 & ~w17232;
assign w17235 = ~w17233 & ~w17234;
assign w17236 = w17220 & w17235;
assign w17237 = ~w17220 & w17234;
assign w17238 = ~w17236 & ~w17237;
assign w17239 = ~pi3804 & pi9040;
assign w17240 = ~pi3817 & ~pi9040;
assign w17241 = ~w17239 & ~w17240;
assign w17242 = pi0925 & ~w17241;
assign w17243 = ~pi0925 & w17241;
assign w17244 = ~w17242 & ~w17243;
assign w17245 = ~w17238 & w17244;
assign w17246 = ~pi3822 & pi9040;
assign w17247 = ~pi3838 & ~pi9040;
assign w17248 = ~w17246 & ~w17247;
assign w17249 = pi0891 & ~w17248;
assign w17250 = ~pi0891 & w17248;
assign w17251 = ~w17249 & ~w17250;
assign w17252 = ~w17219 & ~w17232;
assign w17253 = (w17252 & w17236) | (w17252 & w65289) | (w17236 & w65289);
assign w17254 = w17219 & w17232;
assign w17255 = ~w17252 & ~w17254;
assign w17256 = w17255 & w65290;
assign w17257 = ~w17219 & w17226;
assign w17258 = ~w17232 & w17244;
assign w17259 = w17213 & w17232;
assign w17260 = ~w17258 & ~w17259;
assign w17261 = w17257 & ~w17260;
assign w17262 = ~w17256 & ~w17261;
assign w17263 = ~w17244 & ~w17262;
assign w17264 = w17213 & w17219;
assign w17265 = ~w17232 & w17264;
assign w17266 = ~w17213 & w17219;
assign w17267 = w17233 & w17266;
assign w17268 = ~w17265 & ~w17267;
assign w17269 = w17244 & ~w17268;
assign w17270 = ~w17253 & ~w17269;
assign w17271 = ~w17263 & w17270;
assign w17272 = w17251 & ~w17271;
assign w17273 = ~w17234 & ~w17258;
assign w17274 = w17266 & ~w17273;
assign w17275 = w17219 & ~w17226;
assign w17276 = ~w17234 & ~w17275;
assign w17277 = ~w17244 & ~w17276;
assign w17278 = (~w17274 & ~w17238) | (~w17274 & w65291) | (~w17238 & w65291);
assign w17279 = ~w17251 & ~w17278;
assign w17280 = w17232 & ~w17244;
assign w17281 = w17226 & ~w17251;
assign w17282 = ~w17280 & ~w17281;
assign w17283 = ~w17220 & ~w17258;
assign w17284 = ~w17266 & w17283;
assign w17285 = ~w17282 & w17284;
assign w17286 = ~w17245 & ~w17285;
assign w17287 = ~w17279 & w17286;
assign w17288 = ~w17272 & w17287;
assign w17289 = pi0930 & ~w17288;
assign w17290 = ~pi0930 & w17288;
assign w17291 = ~w17289 & ~w17290;
assign w17292 = ~pi3829 & pi9040;
assign w17293 = ~pi3837 & ~pi9040;
assign w17294 = ~w17292 & ~w17293;
assign w17295 = pi0890 & ~w17294;
assign w17296 = ~pi0890 & w17294;
assign w17297 = ~w17295 & ~w17296;
assign w17298 = ~pi3826 & pi9040;
assign w17299 = ~pi3833 & ~pi9040;
assign w17300 = ~w17298 & ~w17299;
assign w17301 = pi0918 & ~w17300;
assign w17302 = ~pi0918 & w17300;
assign w17303 = ~w17301 & ~w17302;
assign w17304 = ~pi3825 & pi9040;
assign w17305 = ~pi3826 & ~pi9040;
assign w17306 = ~w17304 & ~w17305;
assign w17307 = pi0905 & ~w17306;
assign w17308 = ~pi0905 & w17306;
assign w17309 = ~w17307 & ~w17308;
assign w17310 = ~pi3784 & pi9040;
assign w17311 = ~pi3834 & ~pi9040;
assign w17312 = ~w17310 & ~w17311;
assign w17313 = pi0915 & ~w17312;
assign w17314 = ~pi0915 & w17312;
assign w17315 = ~w17313 & ~w17314;
assign w17316 = w17309 & w17315;
assign w17317 = w17297 & ~w17303;
assign w17318 = w17316 & w17317;
assign w17319 = ~w17297 & w17315;
assign w17320 = ~w17309 & w17319;
assign w17321 = ~w17318 & ~w17320;
assign w17322 = ~pi3792 & pi9040;
assign w17323 = ~pi3836 & ~pi9040;
assign w17324 = ~w17322 & ~w17323;
assign w17325 = pi0926 & ~w17324;
assign w17326 = ~pi0926 & w17324;
assign w17327 = ~w17325 & ~w17326;
assign w17328 = ~w17321 & ~w17327;
assign w17329 = ~w17297 & w17303;
assign w17330 = w17309 & w17329;
assign w17331 = ~w17327 & ~w17330;
assign w17332 = w17309 & ~w17315;
assign w17333 = ~w17331 & w17332;
assign w17334 = w17303 & w17320;
assign w17335 = w17297 & w17303;
assign w17336 = ~w17297 & ~w17303;
assign w17337 = (w17327 & w17336) | (w17327 & w65292) | (w17336 & w65292);
assign w17338 = w17335 & w17337;
assign w17339 = ~pi3818 & pi9040;
assign w17340 = ~pi3829 & ~pi9040;
assign w17341 = ~w17339 & ~w17340;
assign w17342 = pi0909 & ~w17341;
assign w17343 = ~pi0909 & w17341;
assign w17344 = ~w17342 & ~w17343;
assign w17345 = w17309 & w17336;
assign w17346 = ~w17303 & ~w17309;
assign w17347 = w17297 & w17346;
assign w17348 = ~w17345 & ~w17347;
assign w17349 = w17297 & ~w17315;
assign w17350 = w17346 & w17349;
assign w17351 = w17327 & ~w17350;
assign w17352 = ~w17348 & w17351;
assign w17353 = ~w17303 & w17315;
assign w17354 = ~w17309 & ~w17329;
assign w17355 = ~w17353 & w17354;
assign w17356 = ~w17327 & w17355;
assign w17357 = ~w17334 & w17344;
assign w17358 = ~w17333 & w17357;
assign w17359 = ~w17338 & ~w17352;
assign w17360 = ~w17356 & w17359;
assign w17361 = w17358 & w17360;
assign w17362 = ~w17318 & ~w17344;
assign w17363 = w17316 & w17329;
assign w17364 = w17362 & ~w17363;
assign w17365 = w17327 & w17355;
assign w17366 = ~w17303 & w17320;
assign w17367 = w17364 & ~w17366;
assign w17368 = ~w17365 & w17367;
assign w17369 = ~w17303 & w17319;
assign w17370 = ~w17344 & ~w17369;
assign w17371 = w17331 & ~w17354;
assign w17372 = w17370 & w17371;
assign w17373 = ~w17328 & ~w17372;
assign w17374 = (w17373 & w17361) | (w17373 & w65293) | (w17361 & w65293);
assign w17375 = pi0937 & ~w17374;
assign w17376 = ~pi0937 & w17374;
assign w17377 = ~w17375 & ~w17376;
assign w17378 = w17120 & w17151;
assign w17379 = ~w17101 & w17378;
assign w17380 = ~w17136 & w17186;
assign w17381 = w17101 & w17142;
assign w17382 = (~w17128 & w17136) | (~w17128 & w65294) | (w17136 & w65294);
assign w17383 = ~w17089 & ~w17380;
assign w17384 = ~w17382 & w17383;
assign w17385 = ~w17167 & w17384;
assign w17386 = ~w17110 & ~w17185;
assign w17387 = ~w17186 & ~w17386;
assign w17388 = w17102 & w17142;
assign w17389 = w17089 & ~w17388;
assign w17390 = w17159 & w17389;
assign w17391 = ~w17164 & w17390;
assign w17392 = ~w17387 & w17391;
assign w17393 = (~w17379 & w17385) | (~w17379 & w65295) | (w17385 & w65295);
assign w17394 = ~pi0941 & w17393;
assign w17395 = pi0941 & ~w17393;
assign w17396 = ~w17394 & ~w17395;
assign w17397 = ~pi3838 & pi9040;
assign w17398 = ~pi3831 & ~pi9040;
assign w17399 = ~w17397 & ~w17398;
assign w17400 = pi0916 & ~w17399;
assign w17401 = ~pi0916 & w17399;
assign w17402 = ~w17400 & ~w17401;
assign w17403 = ~pi3812 & pi9040;
assign w17404 = ~pi3822 & ~pi9040;
assign w17405 = ~w17403 & ~w17404;
assign w17406 = pi0922 & ~w17405;
assign w17407 = ~pi0922 & w17405;
assign w17408 = ~w17406 & ~w17407;
assign w17409 = ~pi3796 & pi9040;
assign w17410 = ~pi3848 & ~pi9040;
assign w17411 = ~w17409 & ~w17410;
assign w17412 = pi0896 & ~w17411;
assign w17413 = ~pi0896 & w17411;
assign w17414 = ~w17412 & ~w17413;
assign w17415 = w17408 & w17414;
assign w17416 = ~pi3848 & pi9040;
assign w17417 = ~pi3858 & ~pi9040;
assign w17418 = ~w17416 & ~w17417;
assign w17419 = pi0919 & ~w17418;
assign w17420 = ~pi0919 & w17418;
assign w17421 = ~w17419 & ~w17420;
assign w17422 = w17415 & ~w17421;
assign w17423 = w17402 & w17422;
assign w17424 = ~pi3832 & pi9040;
assign w17425 = ~pi3798 & ~pi9040;
assign w17426 = ~w17424 & ~w17425;
assign w17427 = pi0904 & ~w17426;
assign w17428 = ~pi0904 & w17426;
assign w17429 = ~w17427 & ~w17428;
assign w17430 = ~w17402 & w17408;
assign w17431 = ~pi3854 & pi9040;
assign w17432 = ~pi3799 & ~pi9040;
assign w17433 = ~w17431 & ~w17432;
assign w17434 = pi0897 & ~w17433;
assign w17435 = ~pi0897 & w17433;
assign w17436 = ~w17434 & ~w17435;
assign w17437 = ~w17430 & w17436;
assign w17438 = ~w17402 & ~w17414;
assign w17439 = ~w17402 & w17421;
assign w17440 = ~w17408 & ~w17414;
assign w17441 = ~w17439 & ~w17440;
assign w17442 = ~w17438 & ~w17441;
assign w17443 = ~w17437 & w17442;
assign w17444 = w17402 & ~w17421;
assign w17445 = ~w17436 & w17444;
assign w17446 = (~w17421 & ~w17444) | (~w17421 & w65296) | (~w17444 & w65296);
assign w17447 = w17442 & w17446;
assign w17448 = ~w17402 & w17414;
assign w17449 = ~w17421 & w17448;
assign w17450 = (w17436 & ~w17448) | (w17436 & w65297) | (~w17448 & w65297);
assign w17451 = w17415 & w17437;
assign w17452 = (w17402 & ~w17437) | (w17402 & w63718) | (~w17437 & w63718);
assign w17453 = w17450 & ~w17452;
assign w17454 = ~w17447 & ~w17453;
assign w17455 = ~w17443 & ~w17454;
assign w17456 = ~w17436 & ~w17438;
assign w17457 = ~w17414 & ~w17439;
assign w17458 = w17408 & ~w17436;
assign w17459 = w17457 & w17458;
assign w17460 = ~w17449 & ~w17459;
assign w17461 = (w17456 & w17459) | (w17456 & w65298) | (w17459 & w65298);
assign w17462 = ~w17408 & w17414;
assign w17463 = w17402 & w17421;
assign w17464 = w17462 & w17463;
assign w17465 = ~w17422 & ~w17464;
assign w17466 = ~w17461 & w17465;
assign w17467 = (w17429 & w17455) | (w17429 & w65299) | (w17455 & w65299);
assign w17468 = ~w17436 & w17463;
assign w17469 = w17402 & ~w17408;
assign w17470 = ~w17430 & ~w17469;
assign w17471 = w17436 & w17441;
assign w17472 = ~w17470 & w17471;
assign w17473 = (~w17468 & ~w17471) | (~w17468 & w65300) | (~w17471 & w65300);
assign w17474 = ~w17414 & ~w17473;
assign w17475 = w17436 & ~w17462;
assign w17476 = ~w17421 & ~w17456;
assign w17477 = ~w17475 & w17476;
assign w17478 = ~w17443 & ~w17477;
assign w17479 = ~w17429 & ~w17478;
assign w17480 = w17439 & w17440;
assign w17481 = ~w17464 & ~w17480;
assign w17482 = w17436 & ~w17481;
assign w17483 = ~w17423 & ~w17482;
assign w17484 = ~w17474 & w17483;
assign w17485 = ~w17479 & w17484;
assign w17486 = ~w17467 & w17485;
assign w17487 = pi0956 & ~w17486;
assign w17488 = ~pi0956 & w17486;
assign w17489 = ~w17487 & ~w17488;
assign w17490 = ~pi3793 & pi9040;
assign w17491 = ~pi3821 & ~pi9040;
assign w17492 = ~w17490 & ~w17491;
assign w17493 = pi0905 & ~w17492;
assign w17494 = ~pi0905 & w17492;
assign w17495 = ~w17493 & ~w17494;
assign w17496 = ~pi3786 & pi9040;
assign w17497 = ~pi3808 & ~pi9040;
assign w17498 = ~w17496 & ~w17497;
assign w17499 = pi0901 & ~w17498;
assign w17500 = ~pi0901 & w17498;
assign w17501 = ~w17499 & ~w17500;
assign w17502 = ~pi3791 & pi9040;
assign w17503 = ~pi3811 & ~pi9040;
assign w17504 = ~w17502 & ~w17503;
assign w17505 = pi0890 & ~w17504;
assign w17506 = ~pi0890 & w17504;
assign w17507 = ~w17505 & ~w17506;
assign w17508 = ~w17501 & ~w17507;
assign w17509 = ~pi3833 & pi9040;
assign w17510 = ~pi3819 & ~pi9040;
assign w17511 = ~w17509 & ~w17510;
assign w17512 = pi0921 & ~w17511;
assign w17513 = ~pi0921 & w17511;
assign w17514 = ~w17512 & ~w17513;
assign w17515 = ~pi3788 & pi9040;
assign w17516 = ~pi3818 & ~pi9040;
assign w17517 = ~w17515 & ~w17516;
assign w17518 = pi0927 & ~w17517;
assign w17519 = ~pi0927 & w17517;
assign w17520 = ~w17518 & ~w17519;
assign w17521 = w17514 & ~w17520;
assign w17522 = w17508 & w17521;
assign w17523 = w17507 & w17520;
assign w17524 = ~w17507 & ~w17520;
assign w17525 = ~w17523 & ~w17524;
assign w17526 = w17514 & w17525;
assign w17527 = ~w17501 & w17520;
assign w17528 = ~pi3819 & pi9040;
assign w17529 = ~pi3825 & ~pi9040;
assign w17530 = ~w17528 & ~w17529;
assign w17531 = pi0923 & ~w17530;
assign w17532 = ~pi0923 & w17530;
assign w17533 = ~w17531 & ~w17532;
assign w17534 = ~w17527 & w17533;
assign w17535 = w17526 & w17534;
assign w17536 = ~w17520 & ~w17533;
assign w17537 = ~w17507 & w17514;
assign w17538 = ~w17523 & ~w17537;
assign w17539 = ~w17536 & w17538;
assign w17540 = ~w17527 & ~w17533;
assign w17541 = ~w17501 & ~w17514;
assign w17542 = ~w17520 & ~w17541;
assign w17543 = w17540 & ~w17542;
assign w17544 = w17539 & w17543;
assign w17545 = ~w17535 & ~w17544;
assign w17546 = w17501 & ~w17545;
assign w17547 = w17507 & ~w17514;
assign w17548 = ~w17533 & ~w17547;
assign w17549 = ~w17523 & ~w17548;
assign w17550 = ~w17547 & w65301;
assign w17551 = ~w17501 & ~w17550;
assign w17552 = ~w17549 & w17551;
assign w17553 = ~w17522 & ~w17552;
assign w17554 = (~w17495 & w17546) | (~w17495 & w65302) | (w17546 & w65302);
assign w17555 = w17520 & w17533;
assign w17556 = w17541 & w17555;
assign w17557 = w17514 & ~w17533;
assign w17558 = (~w17508 & ~w17540) | (~w17508 & w65303) | (~w17540 & w65303);
assign w17559 = w17557 & ~w17558;
assign w17560 = ~w17556 & ~w17559;
assign w17561 = w17501 & w17525;
assign w17562 = ~w17537 & ~w17547;
assign w17563 = w17536 & ~w17562;
assign w17564 = w17561 & w17563;
assign w17565 = ~w17501 & ~w17524;
assign w17566 = w17539 & w17565;
assign w17567 = ~w17533 & ~w17538;
assign w17568 = w17501 & w17524;
assign w17569 = ~w17547 & ~w17568;
assign w17570 = ~w17567 & ~w17569;
assign w17571 = ~w17566 & ~w17570;
assign w17572 = w17520 & w17557;
assign w17573 = (w17495 & ~w17571) | (w17495 & w65304) | (~w17571 & w65304);
assign w17574 = ~w17520 & w17533;
assign w17575 = ~w17514 & ~w17525;
assign w17576 = ~w17525 & w65305;
assign w17577 = w17574 & w17576;
assign w17578 = ~w17564 & ~w17577;
assign w17579 = w17560 & w17578;
assign w17580 = ~w17573 & w17579;
assign w17581 = ~w17554 & w17580;
assign w17582 = pi0931 & ~w17581;
assign w17583 = ~pi0931 & w17581;
assign w17584 = ~w17582 & ~w17583;
assign w17585 = w17213 & ~w17261;
assign w17586 = ~w17238 & w17585;
assign w17587 = ~w17232 & ~w17237;
assign w17588 = w17244 & ~w17587;
assign w17589 = ~w17255 & w17588;
assign w17590 = w17251 & ~w17256;
assign w17591 = ~w17586 & w17590;
assign w17592 = ~w17589 & w17591;
assign w17593 = w17235 & ~w17264;
assign w17594 = ~w17588 & ~w17593;
assign w17595 = (~w17251 & ~w17255) | (~w17251 & w65306) | (~w17255 & w65306);
assign w17596 = ~w17281 & ~w17595;
assign w17597 = ~w17261 & ~w17594;
assign w17598 = ~w17596 & w17597;
assign w17599 = ~w17592 & ~w17598;
assign w17600 = pi0933 & w17599;
assign w17601 = ~pi0933 & ~w17599;
assign w17602 = ~w17600 & ~w17601;
assign w17603 = ~pi3837 & pi9040;
assign w17604 = ~pi3788 & ~pi9040;
assign w17605 = ~w17603 & ~w17604;
assign w17606 = pi0914 & ~w17605;
assign w17607 = ~pi0914 & w17605;
assign w17608 = ~w17606 & ~w17607;
assign w17609 = ~pi3814 & pi9040;
assign w17610 = ~pi3855 & ~pi9040;
assign w17611 = ~w17609 & ~w17610;
assign w17612 = pi0920 & ~w17611;
assign w17613 = ~pi0920 & w17611;
assign w17614 = ~w17612 & ~w17613;
assign w17615 = w17608 & ~w17614;
assign w17616 = ~pi3850 & pi9040;
assign w17617 = ~pi3792 & ~pi9040;
assign w17618 = ~w17616 & ~w17617;
assign w17619 = pi0906 & ~w17618;
assign w17620 = ~pi0906 & w17618;
assign w17621 = ~w17619 & ~w17620;
assign w17622 = ~pi3813 & pi9040;
assign w17623 = ~pi3785 & ~pi9040;
assign w17624 = ~w17622 & ~w17623;
assign w17625 = pi0896 & ~w17624;
assign w17626 = ~pi0896 & w17624;
assign w17627 = ~w17625 & ~w17626;
assign w17628 = ~w17621 & w17627;
assign w17629 = ~pi3823 & pi9040;
assign w17630 = ~pi3850 & ~pi9040;
assign w17631 = ~w17629 & ~w17630;
assign w17632 = pi0924 & ~w17631;
assign w17633 = ~pi0924 & w17631;
assign w17634 = ~w17632 & ~w17633;
assign w17635 = w17628 & ~w17634;
assign w17636 = w17615 & w17635;
assign w17637 = ~w17614 & ~w17627;
assign w17638 = ~w17608 & ~w17621;
assign w17639 = w17637 & w17638;
assign w17640 = w17621 & ~w17627;
assign w17641 = w17615 & w17640;
assign w17642 = ~w17639 & ~w17641;
assign w17643 = w17608 & w17627;
assign w17644 = ~w17637 & ~w17643;
assign w17645 = ~w17621 & ~w17627;
assign w17646 = ~w17634 & ~w17645;
assign w17647 = w17644 & w17646;
assign w17648 = ~pi3836 & pi9040;
assign w17649 = ~pi3823 & ~pi9040;
assign w17650 = ~w17648 & ~w17649;
assign w17651 = pi0916 & ~w17650;
assign w17652 = ~pi0916 & w17650;
assign w17653 = ~w17651 & ~w17652;
assign w17654 = ~w17608 & w17634;
assign w17655 = w17637 & w17654;
assign w17656 = w17614 & w17627;
assign w17657 = w17608 & w17634;
assign w17658 = ~w17638 & ~w17657;
assign w17659 = w17656 & ~w17658;
assign w17660 = w17621 & w17634;
assign w17661 = w17615 & w17660;
assign w17662 = ~w17653 & ~w17655;
assign w17663 = ~w17661 & w17662;
assign w17664 = w17642 & ~w17647;
assign w17665 = ~w17659 & w17664;
assign w17666 = w17663 & w17665;
assign w17667 = ~w17614 & w17627;
assign w17668 = ~w17621 & ~w17667;
assign w17669 = w17621 & ~w17656;
assign w17670 = ~w17668 & ~w17669;
assign w17671 = w17608 & w17670;
assign w17672 = ~w17608 & ~w17634;
assign w17673 = w17637 & w17672;
assign w17674 = w17621 & w17673;
assign w17675 = ~w17608 & w17614;
assign w17676 = ~w17615 & ~w17675;
assign w17677 = ~w17621 & ~w17676;
assign w17678 = ~w17634 & ~w17677;
assign w17679 = w17644 & ~w17675;
assign w17680 = w17634 & ~w17679;
assign w17681 = ~w17678 & ~w17680;
assign w17682 = w17653 & ~w17674;
assign w17683 = ~w17671 & w17682;
assign w17684 = ~w17681 & w17683;
assign w17685 = ~w17666 & ~w17684;
assign w17686 = ~w17645 & ~w17675;
assign w17687 = w17634 & ~w17686;
assign w17688 = ~w17637 & ~w17640;
assign w17689 = w17687 & ~w17688;
assign w17690 = ~w17608 & w17689;
assign w17691 = w17608 & ~w17621;
assign w17692 = ~w17667 & ~w17691;
assign w17693 = ~w17644 & ~w17692;
assign w17694 = w17657 & ~w17693;
assign w17695 = ~w17693 & w65307;
assign w17696 = ~w17636 & ~w17690;
assign w17697 = ~w17695 & w17696;
assign w17698 = ~w17685 & w17697;
assign w17699 = pi0932 & w17698;
assign w17700 = ~pi0932 & ~w17698;
assign w17701 = ~w17699 & ~w17700;
assign w17702 = ~w17320 & ~w17349;
assign w17703 = w17337 & ~w17702;
assign w17704 = ~w17309 & w17315;
assign w17705 = ~w17297 & ~w17327;
assign w17706 = ~w17704 & ~w17705;
assign w17707 = w17303 & ~w17706;
assign w17708 = ~w17319 & w17707;
assign w17709 = w17297 & w17327;
assign w17710 = ~w17309 & ~w17709;
assign w17711 = w17708 & w17710;
assign w17712 = ~w17316 & ~w17329;
assign w17713 = w17303 & w17332;
assign w17714 = ~w17345 & ~w17713;
assign w17715 = w17712 & ~w17714;
assign w17716 = ~w17704 & w17709;
assign w17717 = ~w17346 & ~w17363;
assign w17718 = ~w17327 & ~w17349;
assign w17719 = ~w17717 & w17718;
assign w17720 = w17344 & ~w17716;
assign w17721 = ~w17715 & w17720;
assign w17722 = ~w17719 & w17721;
assign w17723 = ~w17711 & w17722;
assign w17724 = w17331 & ~w17712;
assign w17725 = w17303 & ~w17309;
assign w17726 = ~w17297 & ~w17725;
assign w17727 = ~w17335 & ~w17726;
assign w17728 = ~w17315 & w17727;
assign w17729 = w17327 & w17363;
assign w17730 = ~w17344 & ~w17729;
assign w17731 = ~w17708 & w17730;
assign w17732 = ~w17724 & ~w17728;
assign w17733 = w17731 & w17732;
assign w17734 = (~w17703 & w17723) | (~w17703 & w65308) | (w17723 & w65308);
assign w17735 = pi0949 & ~w17734;
assign w17736 = ~pi0949 & w17734;
assign w17737 = ~w17735 & ~w17736;
assign w17738 = ~w17095 & w17160;
assign w17739 = ~w17132 & w65309;
assign w17740 = ~w17089 & ~w17739;
assign w17741 = ~w17138 & ~w17740;
assign w17742 = w17127 & ~w17741;
assign w17743 = ~w17118 & ~w17378;
assign w17744 = w17151 & w17743;
assign w17745 = w17130 & w17156;
assign w17746 = ~w17169 & ~w17381;
assign w17747 = ~w17745 & w17746;
assign w17748 = ~w17744 & w17747;
assign w17749 = w17089 & ~w17748;
assign w17750 = ~w17135 & ~w17192;
assign w17751 = ~w17127 & ~w17750;
assign w17752 = w17743 & ~w17751;
assign w17753 = ~w17089 & ~w17752;
assign w17754 = w17108 & ~w17121;
assign w17755 = ~w17195 & w17754;
assign w17756 = ~w17130 & w17161;
assign w17757 = ~w17755 & w17756;
assign w17758 = ~w17749 & ~w17757;
assign w17759 = ~w17753 & w17758;
assign w17760 = (pi0938 & ~w17759) | (pi0938 & w65310) | (~w17759 & w65310);
assign w17761 = w17759 & w65311;
assign w17762 = ~w17760 & ~w17761;
assign w17763 = w17621 & w17676;
assign w17764 = w17676 & w65312;
assign w17765 = ~w17639 & ~w17764;
assign w17766 = ~w17634 & ~w17765;
assign w17767 = ~w17628 & w17654;
assign w17768 = ~w17635 & ~w17691;
assign w17769 = (w17614 & ~w17768) | (w17614 & w65313) | (~w17768 & w65313);
assign w17770 = w17627 & w17634;
assign w17771 = ~w17614 & ~w17621;
assign w17772 = w17770 & w17771;
assign w17773 = ~w17673 & ~w17772;
assign w17774 = w17642 & w17773;
assign w17775 = ~w17769 & w17774;
assign w17776 = ~w17653 & ~w17775;
assign w17777 = ~w17686 & w65314;
assign w17778 = ~w17627 & ~w17634;
assign w17779 = w17614 & ~w17691;
assign w17780 = w17778 & w17779;
assign w17781 = w17637 & w17657;
assign w17782 = ~w17636 & ~w17781;
assign w17783 = ~w17780 & w17782;
assign w17784 = ~w17764 & ~w17777;
assign w17785 = w17783 & w17784;
assign w17786 = w17653 & ~w17785;
assign w17787 = ~w17661 & ~w17695;
assign w17788 = ~w17766 & w17787;
assign w17789 = ~w17776 & w17788;
assign w17790 = ~w17786 & w17789;
assign w17791 = pi0935 & ~w17790;
assign w17792 = ~pi0935 & w17790;
assign w17793 = ~w17791 & ~w17792;
assign w17794 = w17608 & w17614;
assign w17795 = ~w17770 & ~w17794;
assign w17796 = w17669 & ~w17795;
assign w17797 = w17670 & w17678;
assign w17798 = ~w17628 & w17693;
assign w17799 = ~w17655 & ~w17796;
assign w17800 = ~w17798 & w17799;
assign w17801 = ~w17797 & w17800;
assign w17802 = w17653 & ~w17801;
assign w17803 = ~w17634 & w17693;
assign w17804 = (w17668 & w17803) | (w17668 & w65315) | (w17803 & w65315);
assign w17805 = ~w17628 & ~w17656;
assign w17806 = w17672 & w17805;
assign w17807 = (~w17653 & w17694) | (~w17653 & w65316) | (w17694 & w65316);
assign w17808 = ~w17686 & w17688;
assign w17809 = ~w17671 & ~w17808;
assign w17810 = w17653 & ~w17770;
assign w17811 = w17677 & ~w17810;
assign w17812 = ~w17809 & w17811;
assign w17813 = ~w17804 & ~w17807;
assign w17814 = ~w17812 & w17813;
assign w17815 = ~w17802 & w17814;
assign w17816 = pi0934 & ~w17815;
assign w17817 = ~pi0934 & w17815;
assign w17818 = ~w17816 & ~w17817;
assign w17819 = ~w17415 & ~w17440;
assign w17820 = w17439 & w17819;
assign w17821 = ~w17464 & ~w17820;
assign w17822 = w17436 & ~w17821;
assign w17823 = w17457 & w17470;
assign w17824 = w17436 & w17823;
assign w17825 = ~w17445 & ~w17820;
assign w17826 = ~w17824 & w17825;
assign w17827 = w17429 & ~w17826;
assign w17828 = ~w17440 & ~w17448;
assign w17829 = ~w17473 & ~w17828;
assign w17830 = w17448 & w17458;
assign w17831 = ~w17451 & ~w17830;
assign w17832 = w17481 & w17831;
assign w17833 = ~w17447 & w17460;
assign w17834 = w17832 & w17833;
assign w17835 = ~w17429 & ~w17834;
assign w17836 = ~w17827 & w65317;
assign w17837 = ~w17835 & w17836;
assign w17838 = pi0946 & w17837;
assign w17839 = ~pi0946 & ~w17837;
assign w17840 = ~w17838 & ~w17839;
assign w17841 = w17521 & ~w17571;
assign w17842 = w17555 & w17562;
assign w17843 = ~w17522 & ~w17575;
assign w17844 = ~w17533 & ~w17843;
assign w17845 = w17561 & ~w17562;
assign w17846 = ~w17495 & ~w17842;
assign w17847 = ~w17845 & w17846;
assign w17848 = ~w17844 & w17847;
assign w17849 = w17527 & w17537;
assign w17850 = w17495 & ~w17849;
assign w17851 = w17507 & w17514;
assign w17852 = w17501 & w17851;
assign w17853 = w17523 & w17541;
assign w17854 = ~w17542 & ~w17853;
assign w17855 = w17533 & ~w17854;
assign w17856 = ~w17543 & ~w17852;
assign w17857 = w17850 & w17856;
assign w17858 = ~w17855 & w17857;
assign w17859 = ~w17848 & ~w17858;
assign w17860 = ~w17841 & ~w17859;
assign w17861 = ~pi0936 & w17860;
assign w17862 = pi0936 & ~w17860;
assign w17863 = ~w17861 & ~w17862;
assign w17864 = ~w17320 & w17348;
assign w17865 = w17332 & w17335;
assign w17866 = ~w17318 & ~w17865;
assign w17867 = (w17866 & w17864) | (w17866 & w65318) | (w17864 & w65318);
assign w17868 = ~w17327 & ~w17867;
assign w17869 = w17337 & w17362;
assign w17870 = ~w17715 & w17869;
assign w17871 = ~w17344 & w17725;
assign w17872 = w17706 & w17871;
assign w17873 = w17331 & ~w17369;
assign w17874 = ~w17315 & w17336;
assign w17875 = w17327 & ~w17874;
assign w17876 = ~w17707 & w17875;
assign w17877 = ~w17873 & ~w17876;
assign w17878 = ~w17350 & w17866;
assign w17879 = ~w17708 & w17878;
assign w17880 = ~w17877 & w17879;
assign w17881 = w17344 & ~w17880;
assign w17882 = ~w17870 & ~w17872;
assign w17883 = ~w17868 & w17882;
assign w17884 = ~w17881 & w17883;
assign w17885 = pi0957 & ~w17884;
assign w17886 = ~pi0957 & w17884;
assign w17887 = ~w17885 & ~w17886;
assign w17888 = ~w17444 & w17819;
assign w17889 = w17444 & ~w17819;
assign w17890 = ~w17888 & ~w17889;
assign w17891 = w17452 & w17890;
assign w17892 = ~w17436 & w17890;
assign w17893 = w17890 & w65319;
assign w17894 = w17402 & w17414;
assign w17895 = ~w17408 & ~w17894;
assign w17896 = w17408 & ~w17421;
assign w17897 = ~w17448 & ~w17896;
assign w17898 = w17470 & w17897;
assign w17899 = w17450 & ~w17898;
assign w17900 = ~w17898 & w65320;
assign w17901 = ~w17891 & ~w17900;
assign w17902 = (w17429 & ~w17901) | (w17429 & w65321) | (~w17901 & w65321);
assign w17903 = ~w17436 & ~w17820;
assign w17904 = w17444 & w17462;
assign w17905 = w17436 & ~w17480;
assign w17906 = ~w17904 & w17905;
assign w17907 = ~w17903 & ~w17906;
assign w17908 = ~w17429 & ~w17899;
assign w17909 = ~w17892 & w17908;
assign w17910 = ~w17907 & ~w17909;
assign w17911 = ~w17902 & w17910;
assign w17912 = pi0955 & ~w17911;
assign w17913 = ~pi0955 & w17911;
assign w17914 = ~w17912 & ~w17913;
assign w17915 = (w17660 & ~w17783) | (w17660 & w65322) | (~w17783 & w65322);
assign w17916 = w17763 & w17778;
assign w17917 = ~w17653 & ~w17916;
assign w17918 = (~w17654 & w17671) | (~w17654 & w63382) | (w17671 & w63382);
assign w17919 = ~w17689 & ~w17918;
assign w17920 = (~w17654 & ~w17676) | (~w17654 & w65323) | (~w17676 & w65323);
assign w17921 = ~w17918 & w63719;
assign w17922 = (~w17917 & w17921) | (~w17917 & w65324) | (w17921 & w65324);
assign w17923 = ~w17653 & ~w17919;
assign w17924 = ~w17915 & ~w17923;
assign w17925 = (pi0948 & ~w17924) | (pi0948 & w65325) | (~w17924 & w65325);
assign w17926 = w17924 & w65326;
assign w17927 = ~w17925 & ~w17926;
assign w17928 = w17028 & w17037;
assign w17929 = ~w17035 & ~w17928;
assign w17930 = w17006 & ~w17038;
assign w17931 = ~w17018 & w17042;
assign w17932 = w17042 & w17034;
assign w17933 = ~w17058 & ~w17932;
assign w17934 = w17930 & w17933;
assign w17935 = ~w17019 & ~w17025;
assign w17936 = ~w17042 & w17935;
assign w17937 = w17025 & w17042;
assign w17938 = (~w17006 & ~w17042) | (~w17006 & w65274) | (~w17042 & w65274);
assign w17939 = ~w17936 & w17938;
assign w17940 = ~w17934 & ~w17939;
assign w17941 = ~w17929 & ~w17940;
assign w17942 = ~w17026 & ~w17937;
assign w17943 = w17006 & ~w17942;
assign w17944 = ~w17006 & w17012;
assign w17945 = ~w17058 & ~w17944;
assign w17946 = ~w17044 & ~w17945;
assign w17947 = w17000 & w17057;
assign w17948 = ~w17040 & ~w17053;
assign w17949 = ~w17069 & w17948;
assign w17950 = ~w17072 & ~w17947;
assign w17951 = w17949 & w17950;
assign w17952 = ~w17943 & ~w17946;
assign w17953 = w17951 & w17952;
assign w17954 = ~w17068 & ~w17937;
assign w17955 = w17044 & ~w17954;
assign w17956 = w17019 & w17056;
assign w17957 = w17056 & w17061;
assign w17958 = ~w17045 & ~w17928;
assign w17959 = ~w17957 & w17958;
assign w17960 = ~w17012 & ~w17018;
assign w17961 = w17006 & ~w17960;
assign w17962 = ~w17019 & w17961;
assign w17963 = w17958 & w65327;
assign w17964 = w17053 & ~w17956;
assign w17965 = ~w17955 & w17964;
assign w17966 = ~w17031 & w17965;
assign w17967 = ~w17963 & w17966;
assign w17968 = (~w17941 & w17967) | (~w17941 & w65328) | (w17967 & w65328);
assign w17969 = ~pi0942 & w17968;
assign w17970 = pi0942 & ~w17968;
assign w17971 = ~w17969 & ~w17970;
assign w17972 = w17012 & w17018;
assign w17973 = ~w17066 & ~w17972;
assign w17974 = ~w17931 & w17973;
assign w17975 = ~w17019 & w17053;
assign w17976 = w17041 & ~w17975;
assign w17977 = w17974 & w17976;
assign w17978 = ~w17006 & w17074;
assign w17979 = (~w17068 & w17936) | (~w17068 & w65329) | (w17936 & w65329);
assign w17980 = w17972 & ~w17979;
assign w17981 = ~w17053 & ~w17947;
assign w17982 = ~w17980 & w17981;
assign w17983 = ~w17026 & ~w17066;
assign w17984 = ~w17972 & ~w17983;
assign w17985 = w17053 & ~w17984;
assign w17986 = ~w17940 & w17985;
assign w17987 = ~w17982 & ~w17986;
assign w17988 = ~w17977 & ~w17978;
assign w17989 = ~w17032 & w17988;
assign w17990 = ~w17987 & w17989;
assign w17991 = pi0952 & ~w17990;
assign w17992 = ~pi0952 & w17990;
assign w17993 = ~w17991 & ~w17992;
assign w17994 = ~w17257 & ~w17275;
assign w17995 = w17259 & ~w17994;
assign w17996 = ~w17220 & w17994;
assign w17997 = ~w17995 & ~w17996;
assign w17998 = w17244 & ~w17251;
assign w17999 = w17233 & w17264;
assign w18000 = w17998 & ~w17999;
assign w18001 = ~w17997 & w18000;
assign w18002 = w17226 & w17265;
assign w18003 = ~w17244 & w17251;
assign w18004 = w17213 & ~w17226;
assign w18005 = ~w17252 & w17994;
assign w18006 = (~w18004 & ~w17994) | (~w18004 & w65330) | (~w17994 & w65330);
assign w18007 = w17213 & ~w17252;
assign w18008 = ~w18006 & ~w18007;
assign w18009 = ~w18003 & ~w18008;
assign w18010 = ~w17213 & ~w17232;
assign w18011 = ~w17219 & w17259;
assign w18012 = ~w17275 & ~w18011;
assign w18013 = ~w18010 & ~w18012;
assign w18014 = ~w17233 & ~w18010;
assign w18015 = ~w17219 & ~w18014;
assign w18016 = w18003 & ~w18015;
assign w18017 = ~w18013 & w18016;
assign w18018 = ~w18009 & ~w18017;
assign w18019 = ~w17995 & ~w17998;
assign w18020 = ~w18002 & w18019;
assign w18021 = ~w18018 & w18020;
assign w18022 = ~w18001 & ~w18021;
assign w18023 = ~pi0950 & w18022;
assign w18024 = pi0950 & ~w18022;
assign w18025 = ~w18023 & ~w18024;
assign w18026 = ~pi3828 & pi9040;
assign w18027 = ~pi3786 & ~pi9040;
assign w18028 = ~w18026 & ~w18027;
assign w18029 = pi0903 & ~w18028;
assign w18030 = ~pi0903 & w18028;
assign w18031 = ~w18029 & ~w18030;
assign w18032 = ~pi3820 & pi9040;
assign w18033 = ~pi3807 & ~pi9040;
assign w18034 = ~w18032 & ~w18033;
assign w18035 = pi0918 & ~w18034;
assign w18036 = ~pi0918 & w18034;
assign w18037 = ~w18035 & ~w18036;
assign w18038 = ~pi3821 & pi9040;
assign w18039 = ~pi3784 & ~pi9040;
assign w18040 = ~w18038 & ~w18039;
assign w18041 = pi0914 & ~w18040;
assign w18042 = ~pi0914 & w18040;
assign w18043 = ~w18041 & ~w18042;
assign w18044 = w18037 & ~w18043;
assign w18045 = ~pi3811 & pi9040;
assign w18046 = ~pi3820 & ~pi9040;
assign w18047 = ~w18045 & ~w18046;
assign w18048 = pi0907 & ~w18047;
assign w18049 = ~pi0907 & w18047;
assign w18050 = ~w18048 & ~w18049;
assign w18051 = w18044 & w18050;
assign w18052 = ~w18031 & w18051;
assign w18053 = ~pi3807 & pi9040;
assign w18054 = ~pi3791 & ~pi9040;
assign w18055 = ~w18053 & ~w18054;
assign w18056 = pi0920 & ~w18055;
assign w18057 = ~pi0920 & w18055;
assign w18058 = ~w18056 & ~w18057;
assign w18059 = ~w18037 & ~w18050;
assign w18060 = ~pi3855 & pi9040;
assign w18061 = ~pi3813 & ~pi9040;
assign w18062 = ~w18060 & ~w18061;
assign w18063 = pi0909 & ~w18062;
assign w18064 = ~pi0909 & w18062;
assign w18065 = ~w18063 & ~w18064;
assign w18066 = ~w18043 & w18065;
assign w18067 = w18059 & w18066;
assign w18068 = w18037 & w18065;
assign w18069 = w18043 & ~w18065;
assign w18070 = ~w18059 & ~w18069;
assign w18071 = ~w18068 & w18070;
assign w18072 = ~w18050 & ~w18065;
assign w18073 = w18043 & w18072;
assign w18074 = ~w18071 & w63720;
assign w18075 = ~w18037 & w18074;
assign w18076 = ~w18037 & ~w18065;
assign w18077 = w18050 & w18065;
assign w18078 = ~w18044 & ~w18077;
assign w18079 = ~w18051 & ~w18078;
assign w18080 = w18031 & ~w18079;
assign w18081 = ~w18031 & ~w18078;
assign w18082 = (~w18076 & w18078) | (~w18076 & w65331) | (w18078 & w65331);
assign w18083 = ~w18080 & w18082;
assign w18084 = ~w18075 & ~w18083;
assign w18085 = ~w18058 & ~w18084;
assign w18086 = ~w18043 & ~w18065;
assign w18087 = w18031 & w18037;
assign w18088 = w18086 & ~w18087;
assign w18089 = ~w18050 & ~w18088;
assign w18090 = w18081 & ~w18089;
assign w18091 = ~w18074 & w18080;
assign w18092 = w18037 & w18050;
assign w18093 = ~w18079 & w18092;
assign w18094 = ~w18090 & ~w18093;
assign w18095 = ~w18091 & w18094;
assign w18096 = w18058 & ~w18095;
assign w18097 = ~w18068 & ~w18076;
assign w18098 = w18043 & w18097;
assign w18099 = ~w18043 & w18068;
assign w18100 = ~w18098 & ~w18099;
assign w18101 = (w18031 & w18098) | (w18031 & w65332) | (w18098 & w65332);
assign w18102 = w18071 & w18101;
assign w18103 = ~w18052 & ~w18102;
assign w18104 = ~w18085 & w18103;
assign w18105 = (pi0966 & ~w18104) | (pi0966 & w65333) | (~w18104 & w65333);
assign w18106 = w18104 & w65334;
assign w18107 = ~w18105 & ~w18106;
assign w18108 = w17935 & w17974;
assign w18109 = w17033 & ~w18108;
assign w18110 = w17034 & w17066;
assign w18111 = w17930 & ~w18110;
assign w18112 = ~w18109 & ~w18111;
assign w18113 = ~w17000 & w17025;
assign w18114 = ~w17961 & w18113;
assign w18115 = w17933 & w17954;
assign w18116 = w17006 & ~w18115;
assign w18117 = ~w17053 & ~w18114;
assign w18118 = ~w18116 & w18117;
assign w18119 = ~w17006 & w17067;
assign w18120 = ~w17027 & w17053;
assign w18121 = ~w18119 & w18120;
assign w18122 = w17959 & w18121;
assign w18123 = ~w18118 & ~w18122;
assign w18124 = ~w18112 & ~w18123;
assign w18125 = ~pi0940 & w18124;
assign w18126 = pi0940 & ~w18124;
assign w18127 = ~w18125 & ~w18126;
assign w18128 = ~w17495 & ~w17541;
assign w18129 = w17563 & w18128;
assign w18130 = ~w17522 & ~w17563;
assign w18131 = w17560 & w18130;
assign w18132 = ~w18129 & ~w18131;
assign w18133 = ~w17572 & ~w17852;
assign w18134 = ~w17565 & w17574;
assign w18135 = ~w17575 & w18134;
assign w18136 = ~w17514 & ~w17558;
assign w18137 = ~w17495 & w18133;
assign w18138 = ~w18135 & w18137;
assign w18139 = ~w18136 & w18138;
assign w18140 = w17495 & ~w17853;
assign w18141 = w17545 & w65335;
assign w18142 = ~w18139 & ~w18141;
assign w18143 = ~w18132 & ~w18142;
assign w18144 = pi0939 & w18143;
assign w18145 = ~pi0939 & ~w18143;
assign w18146 = ~w18144 & ~w18145;
assign w18147 = (~w18065 & ~w18072) | (~w18065 & w18086) | (~w18072 & w18086);
assign w18148 = ~w18037 & w18043;
assign w18149 = ~w18044 & ~w18148;
assign w18150 = ~w18147 & w18149;
assign w18151 = ~w18031 & w18150;
assign w18152 = w18086 & w18092;
assign w18153 = ~w18151 & ~w18152;
assign w18154 = w18058 & ~w18153;
assign w18155 = w18050 & w18148;
assign w18156 = w18059 & w18086;
assign w18157 = w18058 & ~w18086;
assign w18158 = ~w18150 & w18157;
assign w18159 = ~w18155 & ~w18156;
assign w18160 = ~w18158 & w18159;
assign w18161 = w18031 & ~w18160;
assign w18162 = ~w18031 & ~w18037;
assign w18163 = w18073 & w18162;
assign w18164 = ~w18071 & w63383;
assign w18165 = ~w18150 & w18164;
assign w18166 = (~w18066 & ~w18164) | (~w18066 & w63721) | (~w18164 & w63721);
assign w18167 = w18092 & ~w18166;
assign w18168 = w18072 & w18087;
assign w18169 = ~w18067 & ~w18168;
assign w18170 = ~w18066 & ~w18092;
assign w18171 = w18070 & w18170;
assign w18172 = ~w18163 & w18169;
assign w18173 = ~w18171 & w18172;
assign w18174 = (~w18058 & w18167) | (~w18058 & w65336) | (w18167 & w65336);
assign w18175 = ~w18154 & ~w18161;
assign w18176 = ~w18174 & w18175;
assign w18177 = pi0959 & w18176;
assign w18178 = ~pi0959 & ~w18176;
assign w18179 = ~w18177 & ~w18178;
assign w18180 = w18031 & w18050;
assign w18181 = ~w18043 & w18180;
assign w18182 = ~w18097 & w18181;
assign w18183 = w18077 & w18162;
assign w18184 = w18089 & w18100;
assign w18185 = w18069 & w18092;
assign w18186 = ~w18043 & ~w18072;
assign w18187 = ~w18031 & ~w18077;
assign w18188 = w18186 & w18187;
assign w18189 = w18058 & ~w18185;
assign w18190 = ~w18188 & w18189;
assign w18191 = ~w18184 & w18190;
assign w18192 = ~w18031 & ~w18186;
assign w18193 = ~w18098 & w18192;
assign w18194 = ~w18058 & ~w18156;
assign w18195 = ~w18193 & w18194;
assign w18196 = ~w18101 & w18195;
assign w18197 = ~w18191 & ~w18196;
assign w18198 = ~w18182 & ~w18183;
assign w18199 = ~w18197 & w18198;
assign w18200 = pi0951 & ~w18199;
assign w18201 = ~pi0951 & w18199;
assign w18202 = ~w18200 & ~w18201;
assign w18203 = ~w18071 & w18180;
assign w18204 = ~w18031 & ~w18066;
assign w18205 = (~w18204 & w18071) | (~w18204 & w63722) | (w18071 & w63722);
assign w18206 = ~w18069 & ~w18087;
assign w18207 = ~w18165 & w63723;
assign w18208 = ~w18163 & ~w18203;
assign w18209 = (w18058 & w18207) | (w18058 & w65337) | (w18207 & w65337);
assign w18210 = w18077 & w18193;
assign w18211 = (~w18058 & w18165) | (~w18058 & w65338) | (w18165 & w65338);
assign w18212 = w18080 & ~w18169;
assign w18213 = ~w18210 & ~w18212;
assign w18214 = ~w18211 & w18213;
assign w18215 = ~w18209 & w18214;
assign w18216 = pi0965 & w18215;
assign w18217 = ~pi0965 & ~w18215;
assign w18218 = ~w18216 & ~w18217;
assign w18219 = ~w17414 & w17822;
assign w18220 = ~w17436 & ~w17896;
assign w18221 = ~w17823 & ~w17904;
assign w18222 = w18220 & ~w18221;
assign w18223 = ~w17437 & ~w17894;
assign w18224 = ~w17897 & ~w18223;
assign w18225 = w17440 & w17463;
assign w18226 = w17429 & ~w17830;
assign w18227 = ~w18225 & w18226;
assign w18228 = ~w18224 & w18227;
assign w18229 = ~w17414 & ~w17446;
assign w18230 = ~w18220 & ~w18229;
assign w18231 = ~w17469 & ~w18230;
assign w18232 = ~w17429 & ~w17472;
assign w18233 = ~w18231 & w18232;
assign w18234 = ~w18228 & ~w18233;
assign w18235 = ~w17447 & ~w18222;
assign w18236 = ~w18219 & w18235;
assign w18237 = ~w18234 & w18236;
assign w18238 = ~pi0960 & w18237;
assign w18239 = pi0960 & ~w18237;
assign w18240 = ~w18238 & ~w18239;
assign w18241 = ~w17534 & ~w17556;
assign w18242 = ~w17562 & ~w18241;
assign w18243 = w17539 & w17551;
assign w18244 = ~w18242 & w18243;
assign w18245 = w17538 & w17548;
assign w18246 = w17527 & w17851;
assign w18247 = ~w18245 & ~w18246;
assign w18248 = w17501 & ~w17526;
assign w18249 = ~w17575 & w18248;
assign w18250 = (w17850 & w18247) | (w17850 & w65339) | (w18247 & w65339);
assign w18251 = ~w18249 & w18250;
assign w18252 = ~w18244 & w18251;
assign w18253 = ~w17495 & ~w17576;
assign w18254 = ~w18242 & w18247;
assign w18255 = w18253 & w18254;
assign w18256 = ~w18252 & ~w18255;
assign w18257 = ~pi0929 & w18256;
assign w18258 = pi0929 & ~w18256;
assign w18259 = ~w18257 & ~w18258;
assign w18260 = w17303 & w17316;
assign w18261 = w17351 & ~w18260;
assign w18262 = w17297 & w17725;
assign w18263 = w17344 & ~w17714;
assign w18264 = ~w17327 & ~w18262;
assign w18265 = ~w18263 & w18264;
assign w18266 = ~w18261 & ~w18265;
assign w18267 = w17702 & w17710;
assign w18268 = ~w17338 & ~w17874;
assign w18269 = w17364 & ~w18267;
assign w18270 = w18268 & w18269;
assign w18271 = w17327 & w17727;
assign w18272 = w17344 & ~w17366;
assign w18273 = ~w18271 & w18272;
assign w18274 = ~w18270 & ~w18273;
assign w18275 = ~w18266 & ~w18274;
assign w18276 = ~pi0980 & w18275;
assign w18277 = pi0980 & ~w18275;
assign w18278 = ~w18276 & ~w18277;
assign w18279 = w17261 & w18014;
assign w18280 = ~w17235 & ~w17596;
assign w18281 = ~w17267 & ~w18011;
assign w18282 = ~w18280 & w18281;
assign w18283 = ~w17244 & ~w18282;
assign w18284 = ~w17213 & w17233;
assign w18285 = ~w17232 & ~w17244;
assign w18286 = w17219 & ~w18004;
assign w18287 = ~w18285 & w18286;
assign w18288 = ~w18284 & w18287;
assign w18289 = (~w17251 & w18288) | (~w17251 & w65340) | (w18288 & w65340);
assign w18290 = ~w17266 & ~w17276;
assign w18291 = ~w17244 & ~w17259;
assign w18292 = (~w18291 & w18290) | (~w18291 & w65341) | (w18290 & w65341);
assign w18293 = ~w18005 & ~w18010;
assign w18294 = w17994 & ~w18014;
assign w18295 = ~w17244 & ~w18294;
assign w18296 = ~w18293 & w18295;
assign w18297 = (w17251 & w18296) | (w17251 & w65342) | (w18296 & w65342);
assign w18298 = ~w18279 & ~w18289;
assign w18299 = ~w18297 & w18298;
assign w18300 = ~w18283 & w18299;
assign w18301 = ~pi0944 & ~w18300;
assign w18302 = pi0944 & w18300;
assign w18303 = ~w18301 & ~w18302;
assign w18304 = ~pi3910 & pi9040;
assign w18305 = ~pi3916 & ~pi9040;
assign w18306 = ~w18304 & ~w18305;
assign w18307 = pi0990 & ~w18306;
assign w18308 = ~pi0990 & w18306;
assign w18309 = ~w18307 & ~w18308;
assign w18310 = ~pi3927 & pi9040;
assign w18311 = ~pi3884 & ~pi9040;
assign w18312 = ~w18310 & ~w18311;
assign w18313 = pi0973 & ~w18312;
assign w18314 = ~pi0973 & w18312;
assign w18315 = ~w18313 & ~w18314;
assign w18316 = w18309 & ~w18315;
assign w18317 = ~pi3883 & pi9040;
assign w18318 = ~pi3896 & ~pi9040;
assign w18319 = ~w18317 & ~w18318;
assign w18320 = pi0972 & ~w18319;
assign w18321 = ~pi0972 & w18319;
assign w18322 = ~w18320 & ~w18321;
assign w18323 = w18316 & w18322;
assign w18324 = ~pi3882 & pi9040;
assign w18325 = ~pi3944 & ~pi9040;
assign w18326 = ~w18324 & ~w18325;
assign w18327 = pi0975 & ~w18326;
assign w18328 = ~pi0975 & w18326;
assign w18329 = ~w18327 & ~w18328;
assign w18330 = w18316 & w65343;
assign w18331 = ~w18315 & ~w18322;
assign w18332 = w18329 & w18331;
assign w18333 = ~w18330 & ~w18332;
assign w18334 = ~pi3942 & pi9040;
assign w18335 = ~pi3891 & ~pi9040;
assign w18336 = ~w18334 & ~w18335;
assign w18337 = pi0954 & ~w18336;
assign w18338 = ~pi0954 & w18336;
assign w18339 = ~w18337 & ~w18338;
assign w18340 = ~w18333 & w18339;
assign w18341 = ~pi3885 & pi9040;
assign w18342 = ~pi3882 & ~pi9040;
assign w18343 = ~w18341 & ~w18342;
assign w18344 = pi0985 & ~w18343;
assign w18345 = ~pi0985 & w18343;
assign w18346 = ~w18344 & ~w18345;
assign w18347 = w18329 & ~w18339;
assign w18348 = w18309 & w18329;
assign w18349 = w18322 & w18348;
assign w18350 = ~w18347 & ~w18349;
assign w18351 = ~w18309 & ~w18329;
assign w18352 = w18322 & w18351;
assign w18353 = w18350 & ~w18352;
assign w18354 = w18315 & ~w18353;
assign w18355 = ~w18309 & w18322;
assign w18356 = w18309 & ~w18322;
assign w18357 = ~w18355 & ~w18356;
assign w18358 = w18322 & ~w18339;
assign w18359 = ~w18329 & ~w18339;
assign w18360 = ~w18358 & ~w18359;
assign w18361 = ~w18357 & ~w18360;
assign w18362 = ~w18346 & ~w18361;
assign w18363 = ~w18340 & w18362;
assign w18364 = ~w18354 & w18363;
assign w18365 = ~w18309 & w18331;
assign w18366 = ~w18323 & ~w18339;
assign w18367 = ~w18365 & w18366;
assign w18368 = w18315 & ~w18329;
assign w18369 = ~w18355 & ~w18368;
assign w18370 = w18315 & w18322;
assign w18371 = w18351 & w18370;
assign w18372 = ~w18369 & ~w18371;
assign w18373 = w18339 & ~w18372;
assign w18374 = ~w18367 & ~w18373;
assign w18375 = w18315 & ~w18322;
assign w18376 = w18348 & w18375;
assign w18377 = w18346 & ~w18376;
assign w18378 = ~w18374 & w18377;
assign w18379 = ~w18364 & ~w18378;
assign w18380 = ~w18315 & w18329;
assign w18381 = ~w18357 & w18380;
assign w18382 = w18356 & w18368;
assign w18383 = w18331 & w18351;
assign w18384 = ~w18382 & ~w18383;
assign w18385 = ~w18381 & w18384;
assign w18386 = w18339 & ~w18385;
assign w18387 = ~w18339 & w18371;
assign w18388 = ~w18386 & ~w18387;
assign w18389 = ~w18379 & w18388;
assign w18390 = pi1059 & ~w18389;
assign w18391 = ~pi1059 & w18389;
assign w18392 = ~w18390 & ~w18391;
assign w18393 = ~pi3908 & pi9040;
assign w18394 = ~pi3888 & ~pi9040;
assign w18395 = ~w18393 & ~w18394;
assign w18396 = pi0978 & ~w18395;
assign w18397 = ~pi0978 & w18395;
assign w18398 = ~w18396 & ~w18397;
assign w18399 = ~pi3909 & pi9040;
assign w18400 = ~pi3913 & ~pi9040;
assign w18401 = ~w18399 & ~w18400;
assign w18402 = pi0945 & ~w18401;
assign w18403 = ~pi0945 & w18401;
assign w18404 = ~w18402 & ~w18403;
assign w18405 = ~pi3878 & pi9040;
assign w18406 = ~pi3872 & ~pi9040;
assign w18407 = ~w18405 & ~w18406;
assign w18408 = pi0986 & ~w18407;
assign w18409 = ~pi0986 & w18407;
assign w18410 = ~w18408 & ~w18409;
assign w18411 = ~w18404 & w18410;
assign w18412 = ~pi3913 & pi9040;
assign w18413 = ~pi3908 & ~pi9040;
assign w18414 = ~w18412 & ~w18413;
assign w18415 = pi0977 & ~w18414;
assign w18416 = ~pi0977 & w18414;
assign w18417 = ~w18415 & ~w18416;
assign w18418 = ~pi3877 & pi9040;
assign w18419 = ~pi3906 & ~pi9040;
assign w18420 = ~w18418 & ~w18419;
assign w18421 = pi0967 & ~w18420;
assign w18422 = ~pi0967 & w18420;
assign w18423 = ~w18421 & ~w18422;
assign w18424 = ~w18417 & ~w18423;
assign w18425 = w18411 & w18424;
assign w18426 = ~w18417 & w18423;
assign w18427 = ~w18404 & w18426;
assign w18428 = w18404 & w18417;
assign w18429 = ~w18427 & ~w18428;
assign w18430 = ~w18404 & ~w18423;
assign w18431 = ~w18410 & w18430;
assign w18432 = w18430 & w18457;
assign w18433 = w18429 & ~w18432;
assign w18434 = ~pi3898 & pi9040;
assign w18435 = ~pi3924 & ~pi9040;
assign w18436 = ~w18434 & ~w18435;
assign w18437 = pi0979 & ~w18436;
assign w18438 = ~pi0979 & w18436;
assign w18439 = ~w18437 & ~w18438;
assign w18440 = ~w18433 & ~w18439;
assign w18441 = w18404 & ~w18423;
assign w18442 = w18410 & w18417;
assign w18443 = w18441 & w18442;
assign w18444 = w18426 & w18411;
assign w18445 = ~w18443 & ~w18444;
assign w18446 = ~w18425 & w18445;
assign w18447 = ~w18440 & w18446;
assign w18448 = ~w18398 & ~w18447;
assign w18449 = w18404 & w18426;
assign w18450 = ~w18410 & w18424;
assign w18451 = ~w18449 & ~w18450;
assign w18452 = ~w18398 & ~w18451;
assign w18453 = w18417 & w18423;
assign w18454 = w18398 & w18404;
assign w18455 = w18453 & w18454;
assign w18456 = w18417 & w18430;
assign w18457 = ~w18410 & w18417;
assign w18458 = ~w18456 & ~w18457;
assign w18459 = ~w18417 & w18441;
assign w18460 = w18410 & w18459;
assign w18461 = w18458 & ~w18460;
assign w18462 = w18404 & ~w18410;
assign w18463 = ~w18411 & ~w18462;
assign w18464 = ~w18398 & ~w18404;
assign w18465 = w18410 & w18426;
assign w18466 = ~w18431 & ~w18465;
assign w18467 = ~w18464 & w18466;
assign w18468 = w18423 & w18463;
assign w18469 = (~w18398 & w18467) | (~w18398 & w63724) | (w18467 & w63724);
assign w18470 = ~w18461 & ~w18469;
assign w18471 = w18439 & ~w18455;
assign w18472 = ~w18444 & w18471;
assign w18473 = ~w18452 & w18472;
assign w18474 = ~w18470 & w18473;
assign w18475 = w18411 & w18453;
assign w18476 = ~w18439 & ~w18443;
assign w18477 = ~w18475 & w18476;
assign w18478 = w18398 & ~w18451;
assign w18479 = ~w18425 & w18477;
assign w18480 = ~w18478 & w18479;
assign w18481 = ~w18474 & ~w18480;
assign w18482 = ~w18481 & w65344;
assign w18483 = (pi1061 & w18481) | (pi1061 & w65345) | (w18481 & w65345);
assign w18484 = ~w18482 & ~w18483;
assign w18485 = ~pi3924 & pi9040;
assign w18486 = ~pi3893 & ~pi9040;
assign w18487 = ~w18485 & ~w18486;
assign w18488 = pi0987 & ~w18487;
assign w18489 = ~pi0987 & w18487;
assign w18490 = ~w18488 & ~w18489;
assign w18491 = ~pi3922 & pi9040;
assign w18492 = ~pi3907 & ~pi9040;
assign w18493 = ~w18491 & ~w18492;
assign w18494 = pi0975 & ~w18493;
assign w18495 = ~pi0975 & w18493;
assign w18496 = ~w18494 & ~w18495;
assign w18497 = ~pi3928 & pi9040;
assign w18498 = ~pi3874 & ~pi9040;
assign w18499 = ~w18497 & ~w18498;
assign w18500 = pi0945 & ~w18499;
assign w18501 = ~pi0945 & w18499;
assign w18502 = ~w18500 & ~w18501;
assign w18503 = w18496 & ~w18502;
assign w18504 = ~w18496 & w18502;
assign w18505 = ~w18503 & ~w18504;
assign w18506 = ~pi3900 & pi9040;
assign w18507 = ~pi3922 & ~pi9040;
assign w18508 = ~w18506 & ~w18507;
assign w18509 = pi0985 & ~w18508;
assign w18510 = ~pi0985 & w18508;
assign w18511 = ~w18509 & ~w18510;
assign w18512 = ~pi3899 & pi9040;
assign w18513 = ~pi3900 & ~pi9040;
assign w18514 = ~w18512 & ~w18513;
assign w18515 = pi0976 & ~w18514;
assign w18516 = ~pi0976 & w18514;
assign w18517 = ~w18515 & ~w18516;
assign w18518 = (w18517 & ~w18505) | (w18517 & w65346) | (~w18505 & w65346);
assign w18519 = ~w18505 & ~w18511;
assign w18520 = w18518 & ~w18519;
assign w18521 = ~w18496 & w18520;
assign w18522 = w18496 & w18518;
assign w18523 = w18502 & w18517;
assign w18524 = ~w18503 & ~w18523;
assign w18525 = ~w18490 & ~w18524;
assign w18526 = ~w18522 & w18525;
assign w18527 = ~w18521 & w18526;
assign w18528 = ~w18496 & ~w18517;
assign w18529 = w18490 & w18511;
assign w18530 = w18528 & w18529;
assign w18531 = ~w18511 & ~w18528;
assign w18532 = w18502 & w18511;
assign w18533 = w18528 & w18532;
assign w18534 = ~w18531 & ~w18533;
assign w18535 = w18490 & ~w18534;
assign w18536 = ~w18534 & w65347;
assign w18537 = ~w18502 & w18536;
assign w18538 = w18503 & w18517;
assign w18539 = w18529 & w18538;
assign w18540 = ~w18533 & ~w18539;
assign w18541 = w18496 & w18511;
assign w18542 = ~w18490 & ~w18541;
assign w18543 = w18511 & ~w18517;
assign w18544 = w18496 & w18543;
assign w18545 = ~w18542 & ~w18544;
assign w18546 = w18505 & ~w18545;
assign w18547 = ~pi3920 & pi9040;
assign w18548 = ~pi3894 & ~pi9040;
assign w18549 = ~w18547 & ~w18548;
assign w18550 = pi0977 & ~w18549;
assign w18551 = ~pi0977 & w18549;
assign w18552 = ~w18550 & ~w18551;
assign w18553 = (~w18552 & w18545) | (~w18552 & w63725) | (w18545 & w63725);
assign w18554 = w18505 & w18529;
assign w18555 = ~w18552 & ~w18554;
assign w18556 = ~w18553 & ~w18555;
assign w18557 = ~w18502 & ~w18511;
assign w18558 = ~w18531 & ~w18557;
assign w18559 = (~w18517 & ~w18545) | (~w18517 & w65348) | (~w18545 & w65348);
assign w18560 = ~w18558 & w18559;
assign w18561 = ~w18490 & ~w18543;
assign w18562 = ~w18531 & w18561;
assign w18563 = w18496 & w18523;
assign w18564 = ~w18562 & ~w18563;
assign w18565 = ~w18490 & ~w18511;
assign w18566 = ~w18532 & ~w18557;
assign w18567 = ~w18541 & ~w18565;
assign w18568 = w18566 & w18567;
assign w18569 = ~w18564 & w18568;
assign w18570 = w18540 & ~w18569;
assign w18571 = ~w18556 & w18570;
assign w18572 = w18517 & w18557;
assign w18573 = ~w18504 & ~w18572;
assign w18574 = ~w18503 & ~w18532;
assign w18575 = ~w18490 & ~w18574;
assign w18576 = ~w18573 & ~w18575;
assign w18577 = ~w18517 & w18568;
assign w18578 = ~w18576 & ~w18577;
assign w18579 = ~w18490 & w18541;
assign w18580 = w18552 & ~w18579;
assign w18581 = w18578 & w18580;
assign w18582 = (~w18581 & ~w18571) | (~w18581 & w63726) | (~w18571 & w63726);
assign w18583 = ~w18530 & ~w18537;
assign w18584 = ~w18527 & w18583;
assign w18585 = ~w18582 & w65349;
assign w18586 = (~pi1071 & w18582) | (~pi1071 & w65350) | (w18582 & w65350);
assign w18587 = ~w18585 & ~w18586;
assign w18588 = ~pi3926 & pi9040;
assign w18589 = ~pi3871 & ~pi9040;
assign w18590 = ~w18588 & ~w18589;
assign w18591 = pi0953 & ~w18590;
assign w18592 = ~pi0953 & w18590;
assign w18593 = ~w18591 & ~w18592;
assign w18594 = ~pi3911 & pi9040;
assign w18595 = ~pi3889 & ~pi9040;
assign w18596 = ~w18594 & ~w18595;
assign w18597 = pi0961 & ~w18596;
assign w18598 = ~pi0961 & w18596;
assign w18599 = ~w18597 & ~w18598;
assign w18600 = ~w18593 & w18599;
assign w18601 = ~pi3918 & pi9040;
assign w18602 = ~pi3919 & ~pi9040;
assign w18603 = ~w18601 & ~w18602;
assign w18604 = pi0971 & ~w18603;
assign w18605 = ~pi0971 & w18603;
assign w18606 = ~w18604 & ~w18605;
assign w18607 = ~pi3897 & pi9040;
assign w18608 = ~pi3926 & ~pi9040;
assign w18609 = ~w18607 & ~w18608;
assign w18610 = pi0983 & ~w18609;
assign w18611 = ~pi0983 & w18609;
assign w18612 = ~w18610 & ~w18611;
assign w18613 = ~w18606 & ~w18612;
assign w18614 = w18600 & w18613;
assign w18615 = ~pi3889 & pi9040;
assign w18616 = ~pi3942 & ~pi9040;
assign w18617 = ~w18615 & ~w18616;
assign w18618 = pi0989 & ~w18617;
assign w18619 = ~pi0989 & w18617;
assign w18620 = ~w18618 & ~w18619;
assign w18621 = w18599 & ~w18612;
assign w18622 = ~pi3884 & pi9040;
assign w18623 = ~pi3897 & ~pi9040;
assign w18624 = ~w18622 & ~w18623;
assign w18625 = pi0964 & ~w18624;
assign w18626 = ~pi0964 & w18624;
assign w18627 = ~w18625 & ~w18626;
assign w18628 = ~w18593 & ~w18627;
assign w18629 = w18621 & w18628;
assign w18630 = w18593 & w18612;
assign w18631 = w18599 & w18630;
assign w18632 = w18630 & w65351;
assign w18633 = ~w18629 & ~w18632;
assign w18634 = ~w18600 & w18627;
assign w18635 = ~w18599 & w18606;
assign w18636 = w18630 & w18635;
assign w18637 = ~w18599 & ~w18606;
assign w18638 = ~w18621 & ~w18637;
assign w18639 = ~w18593 & w18638;
assign w18640 = w18593 & w18606;
assign w18641 = w18621 & w18640;
assign w18642 = ~w18639 & ~w18641;
assign w18643 = ~w18639 & w65352;
assign w18644 = w18634 & ~w18643;
assign w18645 = ~w18593 & w18606;
assign w18646 = ~w18599 & ~w18612;
assign w18647 = ~w18645 & w18646;
assign w18648 = ~w18631 & ~w18647;
assign w18649 = ~w18627 & ~w18648;
assign w18650 = w18593 & ~w18599;
assign w18651 = w18613 & w18650;
assign w18652 = ~w18593 & w18612;
assign w18653 = ~w18599 & w18652;
assign w18654 = w18652 & w18637;
assign w18655 = ~w18651 & ~w18654;
assign w18656 = ~w18649 & w65353;
assign w18657 = ~w18644 & w18656;
assign w18658 = w18620 & ~w18657;
assign w18659 = ~w18620 & w18627;
assign w18660 = w18606 & w18612;
assign w18661 = ~w18613 & ~w18660;
assign w18662 = w18599 & ~w18661;
assign w18663 = ~w18647 & ~w18662;
assign w18664 = ~w18651 & w18659;
assign w18665 = ~w18663 & w18664;
assign w18666 = ~w18620 & ~w18627;
assign w18667 = ~w18642 & w18666;
assign w18668 = w18630 & w18637;
assign w18669 = ~w18620 & w18668;
assign w18670 = w18612 & w18627;
assign w18671 = w18645 & w18670;
assign w18672 = ~w18614 & ~w18671;
assign w18673 = ~w18669 & w18672;
assign w18674 = ~w18665 & w18673;
assign w18675 = ~w18667 & w18674;
assign w18676 = ~w18658 & w18675;
assign w18677 = pi1060 & w18676;
assign w18678 = ~pi1060 & ~w18676;
assign w18679 = ~w18677 & ~w18678;
assign w18680 = w18490 & w18496;
assign w18681 = ~w18578 & w18680;
assign w18682 = ~w18538 & w18542;
assign w18683 = ~w18566 & w18682;
assign w18684 = ~w18505 & w18566;
assign w18685 = w18517 & w18684;
assign w18686 = w18555 & ~w18683;
assign w18687 = ~w18685 & w18686;
assign w18688 = ~w18502 & w18544;
assign w18689 = w18552 & ~w18688;
assign w18690 = ~w18535 & w18564;
assign w18691 = w18689 & w18690;
assign w18692 = ~w18687 & ~w18691;
assign w18693 = ~w18681 & ~w18692;
assign w18694 = ~pi1066 & w18693;
assign w18695 = pi1066 & ~w18693;
assign w18696 = ~w18694 & ~w18695;
assign w18697 = ~w18599 & ~w18661;
assign w18698 = w18666 & w18697;
assign w18699 = w18599 & w18627;
assign w18700 = w18612 & ~w18699;
assign w18701 = w18645 & ~w18700;
assign w18702 = w18655 & ~w18701;
assign w18703 = w18599 & ~w18627;
assign w18704 = w18637 & w18670;
assign w18705 = ~w18703 & ~w18704;
assign w18706 = ~w18606 & ~w18705;
assign w18707 = ~w18636 & ~w18706;
assign w18708 = w18702 & w18707;
assign w18709 = w18620 & ~w18708;
assign w18710 = ~w18702 & ~w18705;
assign w18711 = w18606 & w18646;
assign w18712 = w18659 & w18711;
assign w18713 = w18652 & w18703;
assign w18714 = ~w18606 & w18713;
assign w18715 = ~w18627 & ~w18660;
assign w18716 = w18599 & ~w18620;
assign w18717 = ~w18645 & w18716;
assign w18718 = ~w18715 & w18717;
assign w18719 = ~w18712 & ~w18714;
assign w18720 = ~w18718 & w18719;
assign w18721 = ~w18698 & w18720;
assign w18722 = ~w18710 & w18721;
assign w18723 = ~w18709 & w18722;
assign w18724 = ~pi1078 & w18723;
assign w18725 = pi1078 & ~w18723;
assign w18726 = ~w18724 & ~w18725;
assign w18727 = ~pi3868 & pi9040;
assign w18728 = ~pi3880 & ~pi9040;
assign w18729 = ~w18727 & ~w18728;
assign w18730 = pi0988 & ~w18729;
assign w18731 = ~pi0988 & w18729;
assign w18732 = ~w18730 & ~w18731;
assign w18733 = ~pi3905 & pi9040;
assign w18734 = ~pi3879 & ~pi9040;
assign w18735 = ~w18733 & ~w18734;
assign w18736 = pi0963 & ~w18735;
assign w18737 = ~pi0963 & w18735;
assign w18738 = ~w18736 & ~w18737;
assign w18739 = w18732 & w18738;
assign w18740 = ~pi3904 & pi9040;
assign w18741 = ~pi3887 & ~pi9040;
assign w18742 = ~w18740 & ~w18741;
assign w18743 = pi0991 & ~w18742;
assign w18744 = ~pi0991 & w18742;
assign w18745 = ~w18743 & ~w18744;
assign w18746 = ~pi3879 & pi9040;
assign w18747 = ~pi3911 & ~pi9040;
assign w18748 = ~w18746 & ~w18747;
assign w18749 = pi0971 & ~w18748;
assign w18750 = ~pi0971 & w18748;
assign w18751 = ~w18749 & ~w18750;
assign w18752 = ~w18745 & w18751;
assign w18753 = w18739 & w18752;
assign w18754 = ~w18732 & ~w18745;
assign w18755 = w18732 & ~w18751;
assign w18756 = ~w18754 & ~w18755;
assign w18757 = w18745 & ~w18751;
assign w18758 = w18738 & w18757;
assign w18759 = ~w18732 & ~w18738;
assign w18760 = w18751 & w18759;
assign w18761 = ~w18758 & ~w18760;
assign w18762 = w18756 & ~w18761;
assign w18763 = ~pi3890 & pi9040;
assign w18764 = ~pi3918 & ~pi9040;
assign w18765 = ~w18763 & ~w18764;
assign w18766 = pi0970 & ~w18765;
assign w18767 = ~pi0970 & w18765;
assign w18768 = ~w18766 & ~w18767;
assign w18769 = (~w18768 & w18761) | (~w18768 & w63384) | (w18761 & w63384);
assign w18770 = ~w18739 & w18751;
assign w18771 = w18769 & w18770;
assign w18772 = w18738 & w18754;
assign w18773 = w18739 & w18757;
assign w18774 = ~w18772 & ~w18773;
assign w18775 = (w18774 & ~w18769) | (w18774 & w63727) | (~w18769 & w63727);
assign w18776 = ~w18732 & w18738;
assign w18777 = w18751 & w18754;
assign w18778 = (w18768 & ~w18754) | (w18768 & w63728) | (~w18754 & w63728);
assign w18779 = ~w18751 & w18776;
assign w18780 = ~w18752 & ~w18779;
assign w18781 = w18778 & ~w18780;
assign w18782 = w18745 & w18776;
assign w18783 = (w18782 & w18780) | (w18782 & w63729) | (w18780 & w63729);
assign w18784 = ~w18745 & ~w18751;
assign w18785 = (w18768 & ~w18784) | (w18768 & w65354) | (~w18784 & w65354);
assign w18786 = w18738 & ~w18768;
assign w18787 = ~w18756 & ~w18786;
assign w18788 = ~w18785 & w18787;
assign w18789 = ~w18783 & ~w18788;
assign w18790 = ~w18775 & w18789;
assign w18791 = w18732 & ~w18738;
assign w18792 = w18784 & w18791;
assign w18793 = w18739 & w18751;
assign w18794 = ~w18792 & ~w18793;
assign w18795 = ~w18759 & w18794;
assign w18796 = ~w18762 & w18795;
assign w18797 = w18768 & ~w18796;
assign w18798 = ~w18790 & ~w18797;
assign w18799 = ~pi3873 & pi9040;
assign w18800 = ~pi3910 & ~pi9040;
assign w18801 = ~w18799 & ~w18800;
assign w18802 = pi0961 & ~w18801;
assign w18803 = ~pi0961 & w18801;
assign w18804 = ~w18802 & ~w18803;
assign w18805 = ~w18798 & w18804;
assign w18806 = ~w18789 & ~w18804;
assign w18807 = (w18768 & ~w18754) | (w18768 & w65354) | (~w18754 & w65354);
assign w18808 = w18757 & w18759;
assign w18809 = w18774 & w65355;
assign w18810 = w18807 & ~w18809;
assign w18811 = ~w18738 & w18745;
assign w18812 = w18732 & ~w18768;
assign w18813 = w18811 & w18812;
assign w18814 = ~w18753 & ~w18813;
assign w18815 = ~w18810 & w18814;
assign w18816 = ~w18806 & w18815;
assign w18817 = ~w18805 & w65356;
assign w18818 = (~pi1062 & w18805) | (~pi1062 & w65357) | (w18805 & w65357);
assign w18819 = ~w18817 & ~w18818;
assign w18820 = ~pi3907 & pi9040;
assign w18821 = ~pi3941 & ~pi9040;
assign w18822 = ~w18820 & ~w18821;
assign w18823 = pi0969 & ~w18822;
assign w18824 = ~pi0969 & w18822;
assign w18825 = ~w18823 & ~w18824;
assign w18826 = ~pi3869 & pi9040;
assign w18827 = ~pi3928 & ~pi9040;
assign w18828 = ~w18826 & ~w18827;
assign w18829 = pi0963 & ~w18828;
assign w18830 = ~pi0963 & w18828;
assign w18831 = ~w18829 & ~w18830;
assign w18832 = w18825 & w18831;
assign w18833 = ~pi3923 & pi9040;
assign w18834 = ~pi3877 & ~pi9040;
assign w18835 = ~w18833 & ~w18834;
assign w18836 = pi0984 & ~w18835;
assign w18837 = ~pi0984 & w18835;
assign w18838 = ~w18836 & ~w18837;
assign w18839 = ~w18832 & ~w18838;
assign w18840 = ~pi3881 & pi9040;
assign w18841 = ~pi3901 & ~pi9040;
assign w18842 = ~w18840 & ~w18841;
assign w18843 = pi0968 & ~w18842;
assign w18844 = ~pi0968 & w18842;
assign w18845 = ~w18843 & ~w18844;
assign w18846 = ~w18831 & w18845;
assign w18847 = w18831 & ~w18845;
assign w18848 = ~w18846 & ~w18847;
assign w18849 = ~w18839 & ~w18848;
assign w18850 = ~pi3893 & pi9040;
assign w18851 = ~pi3869 & ~pi9040;
assign w18852 = ~w18850 & ~w18851;
assign w18853 = pi0982 & ~w18852;
assign w18854 = ~pi0982 & w18852;
assign w18855 = ~w18853 & ~w18854;
assign w18856 = w18849 & w18855;
assign w18857 = ~w18831 & ~w18845;
assign w18858 = w18838 & ~w18855;
assign w18859 = w18825 & ~w18838;
assign w18860 = ~w18858 & ~w18859;
assign w18861 = w18857 & ~w18860;
assign w18862 = ~pi3906 & pi9040;
assign w18863 = ~pi3881 & ~pi9040;
assign w18864 = ~w18862 & ~w18863;
assign w18865 = pi0988 & ~w18864;
assign w18866 = ~pi0988 & w18864;
assign w18867 = ~w18865 & ~w18866;
assign w18868 = ~w18845 & w18855;
assign w18869 = w18831 & ~w18868;
assign w18870 = ~w18825 & w18838;
assign w18871 = w18831 & w18845;
assign w18872 = ~w18838 & w18855;
assign w18873 = ~w18870 & w18871;
assign w18874 = ~w18872 & w18873;
assign w18875 = w18860 & w18869;
assign w18876 = ~w18874 & w18875;
assign w18877 = ~w18861 & w18867;
assign w18878 = ~w18856 & w18877;
assign w18879 = ~w18876 & w18878;
assign w18880 = w18845 & ~w18855;
assign w18881 = ~w18838 & w18880;
assign w18882 = ~w18845 & w18858;
assign w18883 = w18858 & w18847;
assign w18884 = ~w18881 & ~w18883;
assign w18885 = w18825 & w18838;
assign w18886 = ~w18846 & ~w18855;
assign w18887 = ~w18847 & ~w18886;
assign w18888 = ~w18886 & w65358;
assign w18889 = ~w18867 & w18884;
assign w18890 = ~w18888 & w18889;
assign w18891 = ~w18879 & ~w18890;
assign w18892 = ~w18881 & ~w18882;
assign w18893 = w18832 & ~w18892;
assign w18894 = w18848 & w18858;
assign w18895 = w18867 & ~w18880;
assign w18896 = ~w18838 & ~w18869;
assign w18897 = ~w18895 & w18896;
assign w18898 = ~w18894 & ~w18897;
assign w18899 = ~w18825 & ~w18898;
assign w18900 = ~w18893 & ~w18899;
assign w18901 = ~w18891 & w18900;
assign w18902 = pi1081 & ~w18901;
assign w18903 = ~pi1081 & w18901;
assign w18904 = ~w18902 & ~w18903;
assign w18905 = w18453 & w18462;
assign w18906 = ~w18432 & ~w18905;
assign w18907 = (~w18398 & ~w18426) | (~w18398 & w18464) | (~w18426 & w18464);
assign w18908 = ~w18457 & w18907;
assign w18909 = w18398 & w18475;
assign w18910 = w18429 & ~w18456;
assign w18911 = w18908 & ~w18910;
assign w18912 = ~w18427 & ~w18441;
assign w18913 = (~w18410 & w18427) | (~w18410 & w63730) | (w18427 & w63730);
assign w18914 = ~w18909 & ~w18913;
assign w18915 = ~w18911 & w18914;
assign w18916 = ~w18911 & w63731;
assign w18917 = (w18439 & w18916) | (w18439 & w65359) | (w18916 & w65359);
assign w18918 = ~w18417 & ~w18454;
assign w18919 = w18439 & ~w18918;
assign w18920 = ~w18467 & w65360;
assign w18921 = ~w18439 & ~w18915;
assign w18922 = ~w18428 & ~w18462;
assign w18923 = ~w18439 & ~w18457;
assign w18924 = ~w18922 & ~w18923;
assign w18925 = ~w18425 & ~w18924;
assign w18926 = w18398 & ~w18925;
assign w18927 = ~w18920 & ~w18926;
assign w18928 = ~w18921 & w18927;
assign w18929 = (pi1072 & ~w18928) | (pi1072 & w65361) | (~w18928 & w65361);
assign w18930 = w18928 & w65362;
assign w18931 = ~w18929 & ~w18930;
assign w18932 = w18628 & ~w18648;
assign w18933 = w18634 & ~w18640;
assign w18934 = ~w18651 & w18933;
assign w18935 = ~w18621 & w18627;
assign w18936 = ~w18600 & ~w18650;
assign w18937 = w18606 & ~w18935;
assign w18938 = ~w18936 & w18937;
assign w18939 = w18633 & ~w18934;
assign w18940 = ~w18938 & w18939;
assign w18941 = ~w18620 & ~w18940;
assign w18942 = (w18634 & w18701) | (w18634 & w65363) | (w18701 & w65363);
assign w18943 = w18661 & w18699;
assign w18944 = w18593 & ~w18638;
assign w18945 = w18635 & w18652;
assign w18946 = ~w18627 & ~w18945;
assign w18947 = ~w18714 & w18946;
assign w18948 = ~w18944 & w18947;
assign w18949 = w18620 & ~w18933;
assign w18950 = ~w18943 & w18949;
assign w18951 = ~w18948 & w18950;
assign w18952 = ~w18932 & ~w18942;
assign w18953 = ~w18710 & w18952;
assign w18954 = ~w18951 & w18953;
assign w18955 = ~w18941 & w18954;
assign w18956 = pi1065 & ~w18955;
assign w18957 = ~pi1065 & w18955;
assign w18958 = ~w18956 & ~w18957;
assign w18959 = ~w18859 & ~w18883;
assign w18960 = ~w18855 & w18857;
assign w18961 = w18825 & ~w18960;
assign w18962 = w18846 & w18872;
assign w18963 = w18961 & ~w18962;
assign w18964 = ~w18959 & ~w18963;
assign w18965 = w18857 & w18872;
assign w18966 = (~w18825 & ~w18892) | (~w18825 & w65364) | (~w18892 & w65364);
assign w18967 = w18838 & w18855;
assign w18968 = w18871 & w18967;
assign w18969 = ~w18888 & w18959;
assign w18970 = w18849 & ~w18969;
assign w18971 = w18867 & ~w18968;
assign w18972 = ~w18966 & w18971;
assign w18973 = ~w18970 & w18972;
assign w18974 = ~w18838 & w18960;
assign w18975 = ~w18867 & ~w18974;
assign w18976 = w18846 & ~w18855;
assign w18977 = ~w18868 & ~w18976;
assign w18978 = w18885 & ~w18977;
assign w18979 = ~w18859 & ~w18967;
assign w18980 = w18857 & ~w18979;
assign w18981 = w18831 & ~w18838;
assign w18982 = w18846 & w18855;
assign w18983 = ~w18981 & ~w18982;
assign w18984 = ~w18825 & ~w18983;
assign w18985 = ~w18874 & ~w18980;
assign w18986 = w18975 & w18985;
assign w18987 = ~w18978 & ~w18984;
assign w18988 = w18986 & w18987;
assign w18989 = ~w18973 & ~w18988;
assign w18990 = ~w18964 & ~w18989;
assign w18991 = ~pi1057 & w18990;
assign w18992 = pi1057 & ~w18990;
assign w18993 = ~w18991 & ~w18992;
assign w18994 = ~w18614 & ~w18713;
assign w18995 = w18606 & w18621;
assign w18996 = ~w18697 & ~w18995;
assign w18997 = w18627 & ~w18996;
assign w18998 = w18606 & w18620;
assign w18999 = ~w18703 & ~w18998;
assign w19000 = ~w18661 & ~w18999;
assign w19001 = ~w18997 & ~w19000;
assign w19002 = w18593 & ~w19001;
assign w19003 = w18639 & ~w18700;
assign w19004 = w18628 & w18994;
assign w19005 = ~w19003 & ~w19004;
assign w19006 = w18620 & ~w19005;
assign w19007 = ~w18653 & ~w18995;
assign w19008 = ~w18632 & w19007;
assign w19009 = w18659 & ~w19008;
assign w19010 = ~w18668 & ~w18711;
assign w19011 = w18666 & ~w19010;
assign w19012 = w18628 & w18646;
assign w19013 = (~w19012 & w18994) | (~w19012 & w65365) | (w18994 & w65365);
assign w19014 = ~w19011 & w19013;
assign w19015 = ~w19009 & w19014;
assign w19016 = ~w19006 & w19015;
assign w19017 = ~w19002 & w19016;
assign w19018 = pi1058 & ~w19017;
assign w19019 = ~pi1058 & w19017;
assign w19020 = ~w19018 & ~w19019;
assign w19021 = w18768 & ~w18808;
assign w19022 = w18739 & w18784;
assign w19023 = w19021 & ~w19022;
assign w19024 = ~w18769 & ~w19023;
assign w19025 = (~w18768 & ~w18776) | (~w18768 & w65366) | (~w18776 & w65366);
assign w19026 = ~w18753 & ~w18792;
assign w19027 = w19025 & w19026;
assign w19028 = w18761 & w19027;
assign w19029 = ~w18752 & ~w18755;
assign w19030 = w18732 & w19029;
assign w19031 = ~w18738 & w19030;
assign w19032 = w19028 & ~w19031;
assign w19033 = ~w18751 & w18759;
assign w19034 = ~w19030 & w65367;
assign w19035 = ~w18804 & ~w19034;
assign w19036 = w18752 & w18791;
assign w19037 = ~w18739 & ~w18751;
assign w19038 = ~w19030 & w65368;
assign w19039 = w18754 & w19028;
assign w19040 = w19029 & w65369;
assign w19041 = w18755 & w18811;
assign w19042 = ~w19022 & ~w19036;
assign w19043 = ~w19041 & w19042;
assign w19044 = ~w19040 & w19043;
assign w19045 = ~w19038 & w19044;
assign w19046 = ~w19039 & w19045;
assign w19047 = w18804 & ~w19046;
assign w19048 = (~w19024 & w19032) | (~w19024 & w65370) | (w19032 & w65370);
assign w19049 = (pi1077 & w19047) | (pi1077 & w65371) | (w19047 & w65371);
assign w19050 = ~w19047 & w65372;
assign w19051 = ~w19049 & ~w19050;
assign w19052 = w18847 & w18872;
assign w19053 = ~w18968 & ~w19052;
assign w19054 = ~w18974 & w19053;
assign w19055 = ~w18825 & ~w19054;
assign w19056 = w18825 & ~w18847;
assign w19057 = ~w18825 & ~w18871;
assign w19058 = ~w18855 & ~w19056;
assign w19059 = ~w19057 & w19058;
assign w19060 = w18832 & w18881;
assign w19061 = (~w18857 & w19060) | (~w18857 & w65373) | (w19060 & w65373);
assign w19062 = ~w18845 & ~w18860;
assign w19063 = ~w19061 & ~w19062;
assign w19064 = w18975 & ~w19059;
assign w19065 = ~w19063 & w19064;
assign w19066 = w18857 & w18885;
assign w19067 = w19053 & ~w19066;
assign w19068 = w18884 & ~w18982;
assign w19069 = ~w18870 & ~w19057;
assign w19070 = ~w19068 & ~w19069;
assign w19071 = w18867 & ~w19060;
assign w19072 = w19067 & w19071;
assign w19073 = ~w19070 & w19072;
assign w19074 = ~w19065 & ~w19073;
assign w19075 = ~w18978 & ~w19055;
assign w19076 = ~w19074 & w19075;
assign w19077 = ~pi1086 & w19076;
assign w19078 = pi1086 & ~w19076;
assign w19079 = ~w19077 & ~w19078;
assign w19080 = w18751 & w18791;
assign w19081 = ~w19033 & ~w19080;
assign w19082 = w19021 & ~w19081;
assign w19083 = ~w18745 & w18812;
assign w19084 = w18804 & ~w19083;
assign w19085 = ~w18762 & w19084;
assign w19086 = ~w19082 & w19085;
assign w19087 = w18768 & ~w18794;
assign w19088 = w18774 & w65374;
assign w19089 = ~w19087 & w19088;
assign w19090 = ~w18771 & w19089;
assign w19091 = ~w19086 & ~w19090;
assign w19092 = ~w18762 & w18774;
assign w19093 = w18785 & ~w19092;
assign w19094 = ~w18751 & w18813;
assign w19095 = ~w19093 & ~w19094;
assign w19096 = ~w19091 & w19095;
assign w19097 = pi1063 & ~w19096;
assign w19098 = ~pi1063 & w19096;
assign w19099 = ~w19097 & ~w19098;
assign w19100 = w18523 & w18579;
assign w19101 = w18557 & w18680;
assign w19102 = ~w18490 & w18684;
assign w19103 = ~w19101 & ~w19102;
assign w19104 = ~w18517 & ~w19103;
assign w19105 = ~w18502 & w18528;
assign w19106 = ~w18563 & ~w18579;
assign w19107 = w18523 & ~w18529;
assign w19108 = ~w18565 & w19107;
assign w19109 = ~w18552 & ~w19101;
assign w19110 = ~w19105 & w19109;
assign w19111 = w19106 & ~w19108;
assign w19112 = w19110 & w19111;
assign w19113 = ~w18519 & ~w18568;
assign w19114 = w18561 & ~w19113;
assign w19115 = ~w18539 & w65375;
assign w19116 = ~w18536 & w19115;
assign w19117 = ~w19114 & w19116;
assign w19118 = ~w19112 & ~w19117;
assign w19119 = ~w18530 & ~w19100;
assign w19120 = ~w19104 & w19119;
assign w19121 = ~w19118 & w19120;
assign w19122 = pi1096 & ~w19121;
assign w19123 = ~pi1096 & w19121;
assign w19124 = ~w19122 & ~w19123;
assign w19125 = ~pi3886 & pi9040;
assign w19126 = ~pi3878 & ~pi9040;
assign w19127 = ~w19125 & ~w19126;
assign w19128 = pi0962 & ~w19127;
assign w19129 = ~pi0962 & w19127;
assign w19130 = ~w19128 & ~w19129;
assign w19131 = ~pi3901 & pi9040;
assign w19132 = ~pi3876 & ~pi9040;
assign w19133 = ~w19131 & ~w19132;
assign w19134 = pi0967 & ~w19133;
assign w19135 = ~pi0967 & w19133;
assign w19136 = ~w19134 & ~w19135;
assign w19137 = w19130 & w19136;
assign w19138 = ~pi3894 & pi9040;
assign w19139 = ~pi3923 & ~pi9040;
assign w19140 = ~w19138 & ~w19139;
assign w19141 = pi0974 & ~w19140;
assign w19142 = ~pi0974 & w19140;
assign w19143 = ~w19141 & ~w19142;
assign w19144 = ~pi3874 & pi9040;
assign w19145 = ~pi3899 & ~pi9040;
assign w19146 = ~w19144 & ~w19145;
assign w19147 = pi0984 & ~w19146;
assign w19148 = ~pi0984 & w19146;
assign w19149 = ~w19147 & ~w19148;
assign w19150 = ~w19143 & ~w19149;
assign w19151 = w19137 & w19150;
assign w19152 = w19136 & ~w19149;
assign w19153 = (w19143 & ~w19152) | (w19143 & w65376) | (~w19152 & w65376);
assign w19154 = ~pi3941 & pi9040;
assign w19155 = ~pi3925 & ~pi9040;
assign w19156 = ~w19154 & ~w19155;
assign w19157 = pi0979 & ~w19156;
assign w19158 = ~pi0979 & w19156;
assign w19159 = ~w19157 & ~w19158;
assign w19160 = w19149 & ~w19159;
assign w19161 = ~w19149 & w19159;
assign w19162 = ~w19160 & ~w19161;
assign w19163 = ~w19130 & ~w19162;
assign w19164 = ~w19149 & ~w19159;
assign w19165 = w19130 & w19164;
assign w19166 = (w19153 & w19163) | (w19153 & w65377) | (w19163 & w65377);
assign w19167 = w19130 & w19159;
assign w19168 = ~w19152 & w19167;
assign w19169 = w19137 & ~w19168;
assign w19170 = ~w19166 & ~w19169;
assign w19171 = ~pi3925 & pi9040;
assign w19172 = ~pi3920 & ~pi9040;
assign w19173 = ~w19171 & ~w19172;
assign w19174 = pi0968 & ~w19173;
assign w19175 = ~pi0968 & w19173;
assign w19176 = ~w19174 & ~w19175;
assign w19177 = ~w19170 & w19176;
assign w19178 = ~w19152 & ~w19167;
assign w19179 = ~w19136 & ~w19159;
assign w19180 = w19178 & ~w19179;
assign w19181 = ~w19143 & ~w19180;
assign w19182 = w19153 & ~w19168;
assign w19183 = ~w19181 & ~w19182;
assign w19184 = w19130 & w19160;
assign w19185 = w19152 & w19159;
assign w19186 = ~w19184 & ~w19185;
assign w19187 = ~w19130 & ~w19136;
assign w19188 = w19162 & w19187;
assign w19189 = w19186 & ~w19188;
assign w19190 = ~w19136 & ~w19189;
assign w19191 = ~w19183 & ~w19190;
assign w19192 = ~w19176 & ~w19191;
assign w19193 = ~w19143 & w19176;
assign w19194 = (w19193 & w19162) | (w19193 & w65378) | (w19162 & w65378);
assign w19195 = w19136 & w19159;
assign w19196 = w19143 & w19149;
assign w19197 = ~w19195 & w19196;
assign w19198 = ~w19194 & ~w19197;
assign w19199 = ~w19178 & ~w19198;
assign w19200 = ~w19151 & ~w19199;
assign w19201 = ~w19177 & w19200;
assign w19202 = ~w19192 & w19201;
assign w19203 = pi1093 & ~w19202;
assign w19204 = ~pi1093 & w19202;
assign w19205 = ~w19203 & ~w19204;
assign w19206 = ~pi3880 & pi9040;
assign w19207 = ~pi3873 & ~pi9040;
assign w19208 = ~w19206 & ~w19207;
assign w19209 = pi0989 & ~w19208;
assign w19210 = ~pi0989 & w19208;
assign w19211 = ~w19209 & ~w19210;
assign w19212 = ~pi3891 & pi9040;
assign w19213 = ~pi3927 & ~pi9040;
assign w19214 = ~w19212 & ~w19213;
assign w19215 = pi0958 & ~w19214;
assign w19216 = ~pi0958 & w19214;
assign w19217 = ~w19215 & ~w19216;
assign w19218 = ~w19211 & w19217;
assign w19219 = ~pi3896 & pi9040;
assign w19220 = ~pi3905 & ~pi9040;
assign w19221 = ~w19219 & ~w19220;
assign w19222 = pi0983 & ~w19221;
assign w19223 = ~pi0983 & w19221;
assign w19224 = ~w19222 & ~w19223;
assign w19225 = ~pi3916 & pi9040;
assign w19226 = ~pi3903 & ~pi9040;
assign w19227 = ~w19225 & ~w19226;
assign w19228 = pi0973 & ~w19227;
assign w19229 = ~pi0973 & w19227;
assign w19230 = ~w19228 & ~w19229;
assign w19231 = ~w19224 & ~w19230;
assign w19232 = w19218 & w19231;
assign w19233 = ~pi3903 & pi9040;
assign w19234 = ~pi3904 & ~pi9040;
assign w19235 = ~w19233 & ~w19234;
assign w19236 = pi0981 & ~w19235;
assign w19237 = ~pi0981 & w19235;
assign w19238 = ~w19236 & ~w19237;
assign w19239 = ~w19232 & w19238;
assign w19240 = w19224 & w19230;
assign w19241 = ~w19231 & ~w19240;
assign w19242 = w19218 & w19241;
assign w19243 = ~w19231 & ~w19242;
assign w19244 = w19239 & ~w19243;
assign w19245 = w19211 & ~w19217;
assign w19246 = ~w19224 & w19238;
assign w19247 = ~w19231 & ~w19246;
assign w19248 = w19245 & ~w19247;
assign w19249 = ~w19211 & w19230;
assign w19250 = w19224 & w19249;
assign w19251 = ~w19238 & ~w19250;
assign w19252 = w19211 & ~w19230;
assign w19253 = ~w19249 & ~w19252;
assign w19254 = w19224 & ~w19253;
assign w19255 = ~w19232 & ~w19254;
assign w19256 = w19251 & ~w19255;
assign w19257 = ~pi3887 & pi9040;
assign w19258 = ~pi3890 & ~pi9040;
assign w19259 = ~w19257 & ~w19258;
assign w19260 = pi0972 & ~w19259;
assign w19261 = ~pi0972 & w19259;
assign w19262 = ~w19260 & ~w19261;
assign w19263 = ~w19248 & ~w19262;
assign w19264 = ~w19256 & w19263;
assign w19265 = ~w19217 & ~w19224;
assign w19266 = ~w19252 & ~w19265;
assign w19267 = ~w19245 & w19253;
assign w19268 = ~w19266 & w19267;
assign w19269 = w19230 & w19242;
assign w19270 = w19211 & ~w19224;
assign w19271 = w19230 & w19270;
assign w19272 = ~w19250 & ~w19271;
assign w19273 = ~w19217 & ~w19272;
assign w19274 = w19251 & ~w19273;
assign w19275 = w19240 & w19245;
assign w19276 = w19217 & w19270;
assign w19277 = w19238 & ~w19275;
assign w19278 = ~w19276 & w19277;
assign w19279 = ~w19274 & ~w19278;
assign w19280 = (w19262 & ~w19267) | (w19262 & w65379) | (~w19267 & w65379);
assign w19281 = ~w19269 & w19280;
assign w19282 = ~w19279 & w19281;
assign w19283 = w19224 & ~w19238;
assign w19284 = w19230 & ~w19262;
assign w19285 = ~w19283 & ~w19284;
assign w19286 = ~w19218 & ~w19245;
assign w19287 = ~w19246 & w19286;
assign w19288 = ~w19285 & w19287;
assign w19289 = ~w19244 & ~w19288;
assign w19290 = (w19289 & w19282) | (w19289 & w65380) | (w19282 & w65380);
assign w19291 = pi1076 & ~w19290;
assign w19292 = ~pi1076 & w19290;
assign w19293 = ~w19291 & ~w19292;
assign w19294 = ~w18450 & ~w18465;
assign w19295 = w18404 & ~w19294;
assign w19296 = ~w18398 & ~w18466;
assign w19297 = ~w18467 & ~w19296;
assign w19298 = w18439 & ~w18443;
assign w19299 = ~w18905 & w19298;
assign w19300 = ~w19295 & w19299;
assign w19301 = ~w19297 & w19300;
assign w19302 = w18466 & w65381;
assign w19303 = w18445 & ~w18459;
assign w19304 = w18906 & w19303;
assign w19305 = w18398 & ~w18426;
assign w19306 = w19303 & w65382;
assign w19307 = ~w18439 & ~w19302;
assign w19308 = ~w19306 & w19307;
assign w19309 = ~w19301 & ~w19308;
assign w19310 = ~w18398 & ~w19299;
assign w19311 = ~w19304 & w19310;
assign w19312 = ~w19309 & ~w19311;
assign w19313 = ~pi1087 & w19312;
assign w19314 = pi1087 & ~w19312;
assign w19315 = ~w19313 & ~w19314;
assign w19316 = w19164 & w19187;
assign w19317 = w19176 & ~w19186;
assign w19318 = ~w19130 & ~w19176;
assign w19319 = ~w19136 & w19149;
assign w19320 = ~w19318 & w19319;
assign w19321 = ~w19317 & ~w19320;
assign w19322 = ~w19316 & w19321;
assign w19323 = w19143 & ~w19322;
assign w19324 = w19137 & w19176;
assign w19325 = w19164 & w19324;
assign w19326 = ~w19162 & ~w19196;
assign w19327 = ~w19137 & ~w19187;
assign w19328 = w19326 & ~w19327;
assign w19329 = ~w19184 & w19327;
assign w19330 = ~w19326 & w19329;
assign w19331 = ~w19328 & ~w19330;
assign w19332 = ~w19164 & w19193;
assign w19333 = w19321 & w19332;
assign w19334 = (~w19325 & w19331) | (~w19325 & w65383) | (w19331 & w65383);
assign w19335 = ~w19333 & w19334;
assign w19336 = ~w19323 & w19335;
assign w19337 = pi1084 & ~w19336;
assign w19338 = ~pi1084 & w19336;
assign w19339 = ~w19337 & ~w19338;
assign w19340 = w19136 & w19184;
assign w19341 = (w19150 & w19163) | (w19150 & w65384) | (w19163 & w65384);
assign w19342 = ~w19179 & ~w19195;
assign w19343 = w19143 & w19342;
assign w19344 = (w19164 & ~w19342) | (w19164 & w65385) | (~w19342 & w65385);
assign w19345 = w19149 & w19342;
assign w19346 = ~w19185 & ~w19345;
assign w19347 = ~w19130 & ~w19344;
assign w19348 = w19346 & w19347;
assign w19349 = ~w19340 & ~w19341;
assign w19350 = ~w19348 & w19349;
assign w19351 = w19176 & ~w19350;
assign w19352 = (w19143 & w19345) | (w19143 & w65386) | (w19345 & w65386);
assign w19353 = ~w19143 & ~w19161;
assign w19354 = ~w19165 & w19353;
assign w19355 = ~w19345 & w19354;
assign w19356 = ~w19316 & ~w19355;
assign w19357 = (~w19176 & ~w19356) | (~w19176 & w65387) | (~w19356 & w65387);
assign w19358 = w19130 & w19182;
assign w19359 = ~w19136 & ~w19143;
assign w19360 = w19167 & w19359;
assign w19361 = (~w19360 & w19331) | (~w19360 & w65388) | (w19331 & w65388);
assign w19362 = ~w19357 & w19361;
assign w19363 = ~w19351 & w19362;
assign w19364 = pi1064 & ~w19363;
assign w19365 = ~pi1064 & w19363;
assign w19366 = ~w19364 & ~w19365;
assign w19367 = ~w19143 & ~w19189;
assign w19368 = ~w19160 & w19187;
assign w19369 = ~w19184 & ~w19195;
assign w19370 = ~w19353 & ~w19368;
assign w19371 = w19369 & w19370;
assign w19372 = ~w19367 & ~w19371;
assign w19373 = ~w19143 & ~w19160;
assign w19374 = ~w19130 & w19136;
assign w19375 = ~w19373 & w19374;
assign w19376 = w19176 & ~w19375;
assign w19377 = ~w19367 & w65389;
assign w19378 = ~w19176 & ~w19372;
assign w19379 = w19137 & w19355;
assign w19380 = w19163 & w19343;
assign w19381 = ~w19379 & ~w19380;
assign w19382 = ~w19377 & w19381;
assign w19383 = ~w19378 & w19382;
assign w19384 = ~pi1070 & ~w19383;
assign w19385 = pi1070 & w19383;
assign w19386 = ~w19384 & ~w19385;
assign w19387 = w18546 & ~w19106;
assign w19388 = ~w18520 & ~w18559;
assign w19389 = w18689 & ~w19387;
assign w19390 = ~w19388 & w19389;
assign w19391 = w18490 & ~w18505;
assign w19392 = ~w18544 & w19391;
assign w19393 = w18553 & ~w19392;
assign w19394 = ~w18521 & w19393;
assign w19395 = ~w19390 & ~w19394;
assign w19396 = ~pi1069 & w19395;
assign w19397 = pi1069 & ~w19395;
assign w19398 = ~w19396 & ~w19397;
assign w19399 = ~w18453 & ~w18459;
assign w19400 = w18461 & ~w19399;
assign w19401 = w18398 & ~w19400;
assign w19402 = w18439 & ~w18441;
assign w19403 = ~w18458 & w19402;
assign w19404 = w18907 & ~w19403;
assign w19405 = ~w19401 & ~w19404;
assign w19406 = ~w18430 & ~w18918;
assign w19407 = w18463 & ~w19406;
assign w19408 = ~w18455 & w18477;
assign w19409 = ~w19407 & w19408;
assign w19410 = w18398 & ~w18912;
assign w19411 = ~w18425 & w18439;
assign w19412 = ~w19410 & w19411;
assign w19413 = ~w19409 & ~w19412;
assign w19414 = ~w19405 & ~w19413;
assign w19415 = ~pi1141 & w19414;
assign w19416 = pi1141 & ~w19414;
assign w19417 = ~w19415 & ~w19416;
assign w19418 = w19218 & w19224;
assign w19419 = ~w19276 & ~w19418;
assign w19420 = ~w19230 & ~w19419;
assign w19421 = w19211 & w19224;
assign w19422 = ~w19268 & ~w19421;
assign w19423 = w19238 & ~w19422;
assign w19424 = ~w19238 & w19269;
assign w19425 = (w19262 & w19272) | (w19262 & w65390) | (w19272 & w65390);
assign w19426 = ~w19420 & w19425;
assign w19427 = ~w19424 & w19426;
assign w19428 = ~w19423 & w19427;
assign w19429 = ~w19238 & ~w19241;
assign w19430 = ~w19217 & ~w19231;
assign w19431 = w19217 & w19238;
assign w19432 = w19211 & ~w19431;
assign w19433 = ~w19430 & w19432;
assign w19434 = ~w19429 & ~w19433;
assign w19435 = w19217 & w19224;
assign w19436 = ~w19246 & ~w19435;
assign w19437 = w19249 & ~w19436;
assign w19438 = w19241 & w19267;
assign w19439 = ~w19218 & w19438;
assign w19440 = ~w19232 & ~w19262;
assign w19441 = ~w19437 & w19440;
assign w19442 = w19434 & w19441;
assign w19443 = ~w19439 & w19442;
assign w19444 = ~w19428 & ~w19443;
assign w19445 = pi1056 & w19444;
assign w19446 = ~pi1056 & ~w19444;
assign w19447 = ~w19445 & ~w19446;
assign w19448 = w18961 & ~w19067;
assign w19449 = ~w18976 & ~w19069;
assign w19450 = ~w18963 & ~w19449;
assign w19451 = ~w18848 & w18858;
assign w19452 = ~w18968 & ~w19451;
assign w19453 = ~w19450 & w19452;
assign w19454 = ~w18867 & ~w19453;
assign w19455 = w18825 & ~w18867;
assign w19456 = w18846 & w18967;
assign w19457 = ~w18965 & ~w19456;
assign w19458 = ~w19455 & ~w19457;
assign w19459 = ~w18831 & ~w18880;
assign w19460 = w18859 & ~w19459;
assign w19461 = w18870 & ~w18887;
assign w19462 = ~w19052 & ~w19460;
assign w19463 = ~w19461 & w19462;
assign w19464 = w18867 & ~w19463;
assign w19465 = ~w19448 & ~w19458;
assign w19466 = ~w19464 & w19465;
assign w19467 = ~w19454 & w19466;
assign w19468 = pi1079 & ~w19467;
assign w19469 = ~pi1079 & w19467;
assign w19470 = ~w19468 & ~w19469;
assign w19471 = ~w18309 & w18370;
assign w19472 = w18370 & w65391;
assign w19473 = ~w18339 & w19472;
assign w19474 = (w18316 & w18349) | (w18316 & w65392) | (w18349 & w65392);
assign w19475 = ~w18351 & ~w19474;
assign w19476 = w18358 & ~w19475;
assign w19477 = w18329 & w18375;
assign w19478 = ~w18309 & w18380;
assign w19479 = ~w19477 & ~w19478;
assign w19480 = w18339 & ~w19479;
assign w19481 = w18309 & ~w18347;
assign w19482 = w18370 & w19481;
assign w19483 = w18331 & ~w18348;
assign w19484 = ~w18351 & w19483;
assign w19485 = ~w19482 & ~w19484;
assign w19486 = ~w19480 & w19485;
assign w19487 = ~w19476 & w19486;
assign w19488 = w18346 & ~w19487;
assign w19489 = w18322 & w18368;
assign w19490 = ~w18323 & ~w19489;
assign w19491 = (~w18365 & w19490) | (~w18365 & w65393) | (w19490 & w65393);
assign w19492 = w18339 & ~w19491;
assign w19493 = ~w18330 & ~w18376;
assign w19494 = w18347 & ~w18357;
assign w19495 = w18359 & w18375;
assign w19496 = w18384 & ~w19495;
assign w19497 = ~w19472 & ~w19494;
assign w19498 = w19496 & w19497;
assign w19499 = (~w18346 & ~w19498) | (~w18346 & w65394) | (~w19498 & w65394);
assign w19500 = ~w19473 & ~w19492;
assign w19501 = ~w19499 & w19500;
assign w19502 = ~w19488 & w19501;
assign w19503 = pi1067 & w19502;
assign w19504 = ~pi1067 & ~w19502;
assign w19505 = ~w19503 & ~w19504;
assign w19506 = ~w18760 & ~w18792;
assign w19507 = w18778 & ~w19506;
assign w19508 = ~w18784 & ~w19031;
assign w19509 = w19027 & ~w19508;
assign w19510 = w18768 & ~w18811;
assign w19511 = w19029 & ~w19510;
assign w19512 = ~w18768 & ~w19036;
assign w19513 = w18738 & w18755;
assign w19514 = w18778 & ~w19513;
assign w19515 = ~w19512 & ~w19514;
assign w19516 = ~w18804 & ~w19511;
assign w19517 = ~w19515 & w19516;
assign w19518 = w18776 & w19025;
assign w19519 = ~w18753 & w18804;
assign w19520 = ~w19041 & w19519;
assign w19521 = ~w18781 & w19520;
assign w19522 = ~w19518 & w19521;
assign w19523 = ~w19517 & ~w19522;
assign w19524 = ~w19507 & ~w19509;
assign w19525 = ~w19523 & w19524;
assign w19526 = pi1107 & ~w19525;
assign w19527 = ~pi1107 & w19525;
assign w19528 = ~w19526 & ~w19527;
assign w19529 = ~w19478 & w19493;
assign w19530 = ~w18322 & ~w19529;
assign w19531 = w18339 & ~w19530;
assign w19532 = ~w18309 & w19477;
assign w19533 = w18366 & w18384;
assign w19534 = ~w19532 & w19533;
assign w19535 = ~w19531 & ~w19534;
assign w19536 = w18339 & ~w18380;
assign w19537 = w18331 & w19536;
assign w19538 = w18346 & ~w18382;
assign w19539 = ~w19471 & w19538;
assign w19540 = ~w19537 & w19539;
assign w19541 = ~w19474 & w19540;
assign w19542 = w18315 & w18351;
assign w19543 = ~w18370 & ~w19542;
assign w19544 = ~w18332 & w19543;
assign w19545 = w18339 & ~w19544;
assign w19546 = ~w18352 & ~w18358;
assign w19547 = ~w18315 & ~w19546;
assign w19548 = ~w18346 & ~w19547;
assign w19549 = ~w19545 & w19548;
assign w19550 = ~w19541 & ~w19549;
assign w19551 = ~w19535 & ~w19550;
assign w19552 = ~pi1088 & w19551;
assign w19553 = pi1088 & ~w19551;
assign w19554 = ~w19552 & ~w19553;
assign w19555 = w18361 & ~w18385;
assign w19556 = ~w18346 & ~w18348;
assign w19557 = ~w18356 & w19556;
assign w19558 = ~w18316 & ~w19557;
assign w19559 = w19536 & ~w19542;
assign w19560 = ~w19558 & w19559;
assign w19561 = ~w18331 & w18360;
assign w19562 = ~w18348 & ~w19495;
assign w19563 = ~w18346 & ~w19561;
assign w19564 = ~w19562 & w19563;
assign w19565 = ~w18365 & ~w19477;
assign w19566 = ~w19489 & w19565;
assign w19567 = ~w18339 & ~w19566;
assign w19568 = w18339 & ~w19489;
assign w19569 = ~w19543 & w19568;
assign w19570 = w19529 & ~w19569;
assign w19571 = ~w19567 & w19570;
assign w19572 = w18346 & ~w19571;
assign w19573 = ~w18387 & ~w19555;
assign w19574 = ~w19560 & ~w19564;
assign w19575 = w19573 & w19574;
assign w19576 = ~w19572 & w19575;
assign w19577 = pi1075 & ~w19576;
assign w19578 = ~pi1075 & w19576;
assign w19579 = ~w19577 & ~w19578;
assign w19580 = w19217 & ~w19270;
assign w19581 = w19253 & ~w19580;
assign w19582 = ~w19253 & w19435;
assign w19583 = ~w19581 & ~w19582;
assign w19584 = w19217 & ~w19583;
assign w19585 = w19253 & w19430;
assign w19586 = w19238 & ~w19585;
assign w19587 = (~w19238 & ~w19218) | (~w19238 & w65395) | (~w19218 & w65395);
assign w19588 = ~w19245 & ~w19266;
assign w19589 = ~w19254 & w19587;
assign w19590 = ~w19588 & w19589;
assign w19591 = ~w19586 & ~w19590;
assign w19592 = (w19262 & w19591) | (w19262 & w65396) | (w19591 & w65396);
assign w19593 = (~w19239 & w19584) | (~w19239 & w65397) | (w19584 & w65397);
assign w19594 = w19238 & w19583;
assign w19595 = (~w19232 & ~w19585) | (~w19232 & w19239) | (~w19585 & w19239);
assign w19596 = (~w19262 & w19594) | (~w19262 & w65398) | (w19594 & w65398);
assign w19597 = ~w19593 & ~w19596;
assign w19598 = ~w19592 & w19597;
assign w19599 = ~pi1085 & w19598;
assign w19600 = pi1085 & ~w19598;
assign w19601 = ~w19599 & ~w19600;
assign w19602 = ~w19217 & w19252;
assign w19603 = w19429 & ~w19602;
assign w19604 = ~w19271 & ~w19602;
assign w19605 = w19238 & ~w19604;
assign w19606 = ~w19242 & ~w19603;
assign w19607 = ~w19605 & w19606;
assign w19608 = (~w19262 & ~w19607) | (~w19262 & w63732) | (~w19607 & w63732);
assign w19609 = w19252 & w19435;
assign w19610 = ~w19253 & w19265;
assign w19611 = (~w19238 & w19438) | (~w19238 & w65399) | (w19438 & w65399);
assign w19612 = ~w19241 & ~w19435;
assign w19613 = (~w19609 & ~w19434) | (~w19609 & w65400) | (~w19434 & w65400);
assign w19614 = ~w19611 & w19613;
assign w19615 = w19262 & ~w19614;
assign w19616 = w19238 & ~w19269;
assign w19617 = ~w19275 & w19587;
assign w19618 = ~w19616 & ~w19617;
assign w19619 = ~w19608 & ~w19618;
assign w19620 = w19619 & w65401;
assign w19621 = (~pi1068 & ~w19619) | (~pi1068 & w65402) | (~w19619 & w65402);
assign w19622 = ~w19620 & ~w19621;
assign w19623 = ~pi3974 & pi9040;
assign w19624 = ~pi4005 & ~pi9040;
assign w19625 = ~w19623 & ~w19624;
assign w19626 = pi1104 & ~w19625;
assign w19627 = ~pi1104 & w19625;
assign w19628 = ~w19626 & ~w19627;
assign w19629 = ~pi3996 & pi9040;
assign w19630 = ~pi4012 & ~pi9040;
assign w19631 = ~w19629 & ~w19630;
assign w19632 = pi1133 & ~w19631;
assign w19633 = ~pi1133 & w19631;
assign w19634 = ~w19632 & ~w19633;
assign w19635 = w19628 & w19634;
assign w19636 = ~pi3977 & pi9040;
assign w19637 = ~pi3992 & ~pi9040;
assign w19638 = ~w19636 & ~w19637;
assign w19639 = pi1073 & ~w19638;
assign w19640 = ~pi1073 & w19638;
assign w19641 = ~w19639 & ~w19640;
assign w19642 = ~pi4006 & pi9040;
assign w19643 = ~pi3999 & ~pi9040;
assign w19644 = ~w19642 & ~w19643;
assign w19645 = pi1083 & ~w19644;
assign w19646 = ~pi1083 & w19644;
assign w19647 = ~w19645 & ~w19646;
assign w19648 = ~w19641 & ~w19647;
assign w19649 = ~pi4009 & pi9040;
assign w19650 = ~pi3991 & ~pi9040;
assign w19651 = ~w19649 & ~w19650;
assign w19652 = pi1116 & ~w19651;
assign w19653 = ~pi1116 & w19651;
assign w19654 = ~w19652 & ~w19653;
assign w19655 = w19648 & w19654;
assign w19656 = w19634 & ~w19654;
assign w19657 = ~w19647 & w19656;
assign w19658 = w19641 & w19657;
assign w19659 = ~w19655 & ~w19658;
assign w19660 = w19635 & ~w19659;
assign w19661 = ~w19628 & w19647;
assign w19662 = w19641 & ~w19654;
assign w19663 = ~w19634 & w19662;
assign w19664 = w19661 & w19663;
assign w19665 = w19634 & w19641;
assign w19666 = ~w19647 & w19665;
assign w19667 = w19665 & w65403;
assign w19668 = ~pi3973 & pi9040;
assign w19669 = ~pi3988 & ~pi9040;
assign w19670 = ~w19668 & ~w19669;
assign w19671 = pi1102 & ~w19670;
assign w19672 = ~pi1102 & w19670;
assign w19673 = ~w19671 & ~w19672;
assign w19674 = ~w19667 & w19673;
assign w19675 = w19634 & ~w19641;
assign w19676 = w19647 & w19675;
assign w19677 = ~w19634 & w19648;
assign w19678 = ~w19676 & ~w19677;
assign w19679 = ~w19628 & ~w19678;
assign w19680 = ~w19634 & w19654;
assign w19681 = ~w19656 & ~w19680;
assign w19682 = w19641 & w19647;
assign w19683 = w19681 & w19682;
assign w19684 = ~w19634 & w19647;
assign w19685 = ~w19662 & ~w19684;
assign w19686 = w19628 & ~w19685;
assign w19687 = ~w19683 & w19686;
assign w19688 = w19674 & ~w19679;
assign w19689 = ~w19687 & w19688;
assign w19690 = w19641 & w19654;
assign w19691 = ~w19628 & ~w19690;
assign w19692 = ~w19657 & ~w19684;
assign w19693 = w19691 & w19692;
assign w19694 = w19628 & ~w19655;
assign w19695 = w19675 & w19701;
assign w19696 = w19694 & ~w19695;
assign w19697 = ~w19693 & ~w19696;
assign w19698 = ~w19673 & ~w19683;
assign w19699 = ~w19697 & w19698;
assign w19700 = ~w19689 & ~w19699;
assign w19701 = w19647 & ~w19654;
assign w19702 = w19628 & ~w19701;
assign w19703 = ~w19641 & ~w19654;
assign w19704 = w19628 & ~w19647;
assign w19705 = ~w19641 & ~w19704;
assign w19706 = ~w19703 & ~w19705;
assign w19707 = ~w19634 & w19702;
assign w19708 = ~w19706 & w19707;
assign w19709 = ~w19664 & ~w19708;
assign w19710 = ~w19660 & w19709;
assign w19711 = ~w19700 & w19710;
assign w19712 = pi0994 & ~w19711;
assign w19713 = ~pi0994 & w19711;
assign w19714 = ~w19712 & ~w19713;
assign w19715 = ~pi4033 & pi9040;
assign w19716 = ~pi3984 & ~pi9040;
assign w19717 = ~w19715 & ~w19716;
assign w19718 = pi1117 & ~w19717;
assign w19719 = ~pi1117 & w19717;
assign w19720 = ~w19718 & ~w19719;
assign w19721 = ~pi3994 & pi9040;
assign w19722 = ~pi3993 & ~pi9040;
assign w19723 = ~w19721 & ~w19722;
assign w19724 = pi1103 & ~w19723;
assign w19725 = ~pi1103 & w19723;
assign w19726 = ~w19724 & ~w19725;
assign w19727 = w19720 & w19726;
assign w19728 = ~w19720 & ~w19726;
assign w19729 = ~w19727 & ~w19728;
assign w19730 = ~pi4034 & pi9040;
assign w19731 = ~pi3996 & ~pi9040;
assign w19732 = ~w19730 & ~w19731;
assign w19733 = pi1092 & ~w19732;
assign w19734 = ~pi1092 & w19732;
assign w19735 = ~w19733 & ~w19734;
assign w19736 = ~w19729 & w19735;
assign w19737 = ~pi4019 & pi9040;
assign w19738 = ~pi3973 & ~pi9040;
assign w19739 = ~w19737 & ~w19738;
assign w19740 = pi1109 & ~w19739;
assign w19741 = ~pi1109 & w19739;
assign w19742 = ~w19740 & ~w19741;
assign w19743 = ~w19736 & ~w19742;
assign w19744 = ~pi3982 & pi9040;
assign w19745 = ~pi3981 & ~pi9040;
assign w19746 = ~w19744 & ~w19745;
assign w19747 = pi1073 & ~w19746;
assign w19748 = ~pi1073 & w19746;
assign w19749 = ~w19747 & ~w19748;
assign w19750 = ~w19726 & w19749;
assign w19751 = w19720 & ~w19735;
assign w19752 = w19750 & w19751;
assign w19753 = w19742 & ~w19752;
assign w19754 = ~w19726 & ~w19735;
assign w19755 = w19720 & ~w19749;
assign w19756 = w19754 & w19755;
assign w19757 = ~w19720 & ~w19754;
assign w19758 = w19726 & ~w19749;
assign w19759 = ~w19750 & ~w19758;
assign w19760 = w19757 & w19759;
assign w19761 = ~w19756 & ~w19760;
assign w19762 = w19726 & w19735;
assign w19763 = ~w19749 & ~w19762;
assign w19764 = w19761 & w19763;
assign w19765 = w19753 & ~w19764;
assign w19766 = ~w19743 & ~w19765;
assign w19767 = w19720 & w19735;
assign w19768 = (~w19742 & ~w19767) | (~w19742 & w63325) | (~w19767 & w63325);
assign w19769 = ~w19735 & ~w19749;
assign w19770 = ~w19750 & ~w19769;
assign w19771 = ~w19729 & ~w19770;
assign w19772 = w19768 & ~w19771;
assign w19773 = ~w19735 & w19749;
assign w19774 = w19720 & ~w19773;
assign w19775 = w19759 & ~w19774;
assign w19776 = ~w19759 & w19767;
assign w19777 = ~w19775 & ~w19776;
assign w19778 = w19720 & ~w19777;
assign w19779 = w19742 & ~w19760;
assign w19780 = w19735 & ~w19759;
assign w19781 = w19772 & ~w19780;
assign w19782 = ~w19779 & ~w19781;
assign w19783 = (w19772 & w19782) | (w19772 & w63385) | (w19782 & w63385);
assign w19784 = ~pi4020 & pi9040;
assign w19785 = ~pi3978 & ~pi9040;
assign w19786 = ~w19784 & ~w19785;
assign w19787 = pi1083 & ~w19786;
assign w19788 = ~pi1083 & w19786;
assign w19789 = ~w19787 & ~w19788;
assign w19790 = ~w19742 & w19749;
assign w19791 = ~w19751 & w19790;
assign w19792 = w19735 & w19749;
assign w19793 = ~w19791 & ~w19792;
assign w19794 = ~w19729 & ~w19793;
assign w19795 = ~w19720 & ~w19735;
assign w19796 = w19726 & w19795;
assign w19797 = ~w19790 & w19796;
assign w19798 = ~w19789 & ~w19797;
assign w19799 = ~w19794 & w19798;
assign w19800 = ~w19720 & w19749;
assign w19801 = ~w19755 & ~w19800;
assign w19802 = w19754 & w19801;
assign w19803 = w19726 & w19742;
assign w19804 = w19762 & w19800;
assign w19805 = ~w19751 & ~w19804;
assign w19806 = w19803 & ~w19805;
assign w19807 = ~w19754 & ~w19762;
assign w19808 = w19791 & w19807;
assign w19809 = (w19789 & ~w19801) | (w19789 & w65404) | (~w19801 & w65404);
assign w19810 = ~w19808 & w19809;
assign w19811 = ~w19806 & w19810;
assign w19812 = (~w19811 & w19783) | (~w19811 & w63733) | (w19783 & w63733);
assign w19813 = ~w19812 & w65405;
assign w19814 = (pi0993 & w19812) | (pi0993 & w65406) | (w19812 & w65406);
assign w19815 = ~w19813 & ~w19814;
assign w19816 = ~pi4027 & pi9040;
assign w19817 = ~pi3983 & ~pi9040;
assign w19818 = ~w19816 & ~w19817;
assign w19819 = pi1102 & ~w19818;
assign w19820 = ~pi1102 & w19818;
assign w19821 = ~w19819 & ~w19820;
assign w19822 = ~pi4008 & pi9040;
assign w19823 = ~pi4028 & ~pi9040;
assign w19824 = ~w19822 & ~w19823;
assign w19825 = pi1074 & ~w19824;
assign w19826 = ~pi1074 & w19824;
assign w19827 = ~w19825 & ~w19826;
assign w19828 = w19821 & w19827;
assign w19829 = ~w19821 & ~w19827;
assign w19830 = ~w19828 & ~w19829;
assign w19831 = ~pi4007 & pi9040;
assign w19832 = ~pi4013 & ~pi9040;
assign w19833 = ~w19831 & ~w19832;
assign w19834 = pi1116 & ~w19833;
assign w19835 = ~pi1116 & w19833;
assign w19836 = ~w19834 & ~w19835;
assign w19837 = ~w19830 & ~w19836;
assign w19838 = w19830 & w19836;
assign w19839 = ~w19837 & ~w19838;
assign w19840 = ~pi4017 & pi9040;
assign w19841 = ~pi3985 & ~pi9040;
assign w19842 = ~w19840 & ~w19841;
assign w19843 = pi1105 & ~w19842;
assign w19844 = ~pi1105 & w19842;
assign w19845 = ~w19843 & ~w19844;
assign w19846 = w19839 & w19845;
assign w19847 = w19821 & ~w19845;
assign w19848 = ~pi4014 & pi9040;
assign w19849 = ~pi3995 & ~pi9040;
assign w19850 = ~w19848 & ~w19849;
assign w19851 = pi1150 & ~w19850;
assign w19852 = ~pi1150 & w19850;
assign w19853 = ~w19851 & ~w19852;
assign w19854 = ~w19847 & ~w19853;
assign w19855 = w19827 & w19854;
assign w19856 = w19846 & w19855;
assign w19857 = ~w19836 & ~w19845;
assign w19858 = ~w19821 & ~w19857;
assign w19859 = w19827 & ~w19836;
assign w19860 = w19847 & w19859;
assign w19861 = ~w19858 & ~w19860;
assign w19862 = w19853 & ~w19861;
assign w19863 = w19837 & w19845;
assign w19864 = w19862 & w19863;
assign w19865 = ~w19827 & w19836;
assign w19866 = ~w19845 & ~w19853;
assign w19867 = w19865 & w19866;
assign w19868 = w19821 & w19853;
assign w19869 = w19857 & w19868;
assign w19870 = ~pi3998 & pi9040;
assign w19871 = ~pi4030 & ~pi9040;
assign w19872 = ~w19870 & ~w19871;
assign w19873 = pi1089 & ~w19872;
assign w19874 = ~pi1089 & w19872;
assign w19875 = ~w19873 & ~w19874;
assign w19876 = ~w19827 & w19857;
assign w19877 = w19827 & w19845;
assign w19878 = w19836 & w19877;
assign w19879 = w19821 & w19836;
assign w19880 = ~w19853 & w19879;
assign w19881 = ~w19878 & ~w19880;
assign w19882 = ~w19821 & w19853;
assign w19883 = w19877 & w19882;
assign w19884 = ~w19876 & ~w19883;
assign w19885 = w19881 & w19884;
assign w19886 = ~w19830 & ~w19845;
assign w19887 = w19885 & w19886;
assign w19888 = ~w19821 & ~w19853;
assign w19889 = ~w19845 & ~w19859;
assign w19890 = w19888 & w19889;
assign w19891 = w19836 & w19853;
assign w19892 = ~w19836 & ~w19853;
assign w19893 = ~w19891 & ~w19892;
assign w19894 = w19821 & ~w19827;
assign w19895 = w19845 & w19894;
assign w19896 = ~w19893 & w19895;
assign w19897 = w19878 & w19882;
assign w19898 = ~w19875 & ~w19890;
assign w19899 = ~w19896 & ~w19897;
assign w19900 = w19898 & w19899;
assign w19901 = ~w19887 & w19900;
assign w19902 = ~w19828 & ~w19865;
assign w19903 = ~w19853 & ~w19902;
assign w19904 = w19829 & w19845;
assign w19905 = ~w19859 & ~w19904;
assign w19906 = ~w19903 & ~w19905;
assign w19907 = ~w19845 & ~w19865;
assign w19908 = ~w19888 & w19907;
assign w19909 = w19830 & w19908;
assign w19910 = ~w19906 & ~w19909;
assign w19911 = w19875 & ~w19880;
assign w19912 = w19910 & w19911;
assign w19913 = ~w19901 & ~w19912;
assign w19914 = ~w19867 & ~w19869;
assign w19915 = ~w19864 & w19914;
assign w19916 = ~w19856 & w19915;
assign w19917 = ~w19913 & w19916;
assign w19918 = pi0992 & ~w19917;
assign w19919 = ~pi0992 & w19917;
assign w19920 = ~w19918 & ~w19919;
assign w19921 = ~pi4030 & pi9040;
assign w19922 = ~pi4026 & ~pi9040;
assign w19923 = ~w19921 & ~w19922;
assign w19924 = pi1095 & ~w19923;
assign w19925 = ~pi1095 & w19923;
assign w19926 = ~w19924 & ~w19925;
assign w19927 = ~pi3986 & pi9040;
assign w19928 = ~pi4007 & ~pi9040;
assign w19929 = ~w19927 & ~w19928;
assign w19930 = pi1082 & ~w19929;
assign w19931 = ~pi1082 & w19929;
assign w19932 = ~w19930 & ~w19931;
assign w19933 = ~w19926 & ~w19932;
assign w19934 = ~pi4004 & pi9040;
assign w19935 = ~pi4035 & ~pi9040;
assign w19936 = ~w19934 & ~w19935;
assign w19937 = pi1128 & ~w19936;
assign w19938 = ~pi1128 & w19936;
assign w19939 = ~w19937 & ~w19938;
assign w19940 = ~w19932 & w19939;
assign w19941 = w19932 & ~w19939;
assign w19942 = ~w19940 & ~w19941;
assign w19943 = ~pi4015 & pi9040;
assign w19944 = ~pi3997 & ~pi9040;
assign w19945 = ~w19943 & ~w19944;
assign w19946 = pi1114 & ~w19945;
assign w19947 = ~pi1114 & w19945;
assign w19948 = ~w19946 & ~w19947;
assign w19949 = ~w19942 & w63386;
assign w19950 = ~pi3979 & pi9040;
assign w19951 = ~pi4010 & ~pi9040;
assign w19952 = ~w19950 & ~w19951;
assign w19953 = pi1129 & ~w19952;
assign w19954 = ~pi1129 & w19952;
assign w19955 = ~w19953 & ~w19954;
assign w19956 = w19926 & w19955;
assign w19957 = ~pi3975 & pi9040;
assign w19958 = ~pi4027 & ~pi9040;
assign w19959 = ~w19957 & ~w19958;
assign w19960 = pi1110 & ~w19959;
assign w19961 = ~pi1110 & w19959;
assign w19962 = ~w19960 & ~w19961;
assign w19963 = ~w19956 & w19962;
assign w19964 = w19949 & ~w19963;
assign w19965 = ~w19926 & w19932;
assign w19966 = w19939 & w19965;
assign w19967 = ~w19932 & w19956;
assign w19968 = ~w19966 & ~w19967;
assign w19969 = w19932 & ~w19955;
assign w19970 = ~w19940 & ~w19969;
assign w19971 = w19926 & ~w19970;
assign w19972 = w19968 & ~w19971;
assign w19973 = w19939 & ~w19948;
assign w19974 = w19926 & ~w19948;
assign w19975 = ~w19955 & w19974;
assign w19976 = ~w19939 & w19955;
assign w19977 = ~w19974 & w19976;
assign w19978 = ~w19973 & ~w19975;
assign w19979 = ~w19977 & w19978;
assign w19980 = (~w19932 & ~w19978) | (~w19932 & w63734) | (~w19978 & w63734);
assign w19981 = w19972 & ~w19980;
assign w19982 = (w19962 & w19972) | (w19962 & w63735) | (w19972 & w63735);
assign w19983 = ~w19981 & w19982;
assign w19984 = ~w19926 & w19948;
assign w19985 = ~w19970 & w19984;
assign w19986 = ~w19939 & ~w19955;
assign w19987 = w19926 & w19986;
assign w19988 = w19942 & w19955;
assign w19989 = w19968 & w19988;
assign w19990 = ~w19985 & ~w19987;
assign w19991 = ~w19989 & w19990;
assign w19992 = ~w19941 & w19948;
assign w19993 = ~w19940 & w19992;
assign w19994 = w19992 & w63387;
assign w19995 = ~w19949 & ~w19994;
assign w19996 = w19939 & ~w19995;
assign w19997 = ~w19942 & w65407;
assign w19998 = ~w19975 & ~w19997;
assign w19999 = w19991 & ~w19998;
assign w20000 = ~w19996 & w19999;
assign w20001 = w19932 & ~w19974;
assign w20002 = ~w19984 & ~w20001;
assign w20003 = w19955 & ~w20002;
assign w20004 = (~w20003 & ~w19981) | (~w20003 & w65408) | (~w19981 & w65408);
assign w20005 = ~w19962 & ~w19976;
assign w20006 = ~w20004 & w20005;
assign w20007 = ~w19964 & ~w19983;
assign w20008 = ~w20000 & w20007;
assign w20009 = w20008 & w65409;
assign w20010 = (~pi1027 & ~w20008) | (~pi1027 & w65410) | (~w20008 & w65410);
assign w20011 = ~w20009 & ~w20010;
assign w20012 = ~w19933 & ~w19984;
assign w20013 = ~w19992 & ~w20012;
assign w20014 = w19976 & w20013;
assign w20015 = w19965 & w19973;
assign w20016 = ~w19962 & ~w20015;
assign w20017 = (w20016 & w19995) | (w20016 & w65411) | (w19995 & w65411);
assign w20018 = ~w19939 & w19967;
assign w20019 = (~w19995 & w65412) | (~w19995 & w65413) | (w65412 & w65413);
assign w20020 = ~w19955 & w19984;
assign w20021 = ~w19966 & ~w20020;
assign w20022 = w19970 & ~w20021;
assign w20023 = ~w19997 & ~w20022;
assign w20024 = ~w20019 & w20023;
assign w20025 = ~w20017 & ~w20024;
assign w20026 = w19933 & ~w19939;
assign w20027 = ~w19948 & w20026;
assign w20028 = w19948 & w19955;
assign w20029 = w19940 & w20028;
assign w20030 = w19941 & w19974;
assign w20031 = ~w20029 & ~w20030;
assign w20032 = ~w20027 & w20031;
assign w20033 = (~w19962 & ~w19991) | (~w19962 & w65414) | (~w19991 & w65414);
assign w20034 = ~w20014 & ~w20033;
assign w20035 = ~w20025 & w20034;
assign w20036 = pi1004 & w20035;
assign w20037 = ~pi1004 & ~w20035;
assign w20038 = ~w20036 & ~w20037;
assign w20039 = ~w19967 & ~w20026;
assign w20040 = ~w20028 & ~w20039;
assign w20041 = w19932 & ~w19979;
assign w20042 = w19940 & w19984;
assign w20043 = ~w19962 & ~w20042;
assign w20044 = ~w20040 & w20043;
assign w20045 = ~w20041 & w20044;
assign w20046 = w19932 & w20020;
assign w20047 = ~w19926 & w19940;
assign w20048 = ~w20030 & ~w20047;
assign w20049 = w19955 & ~w20048;
assign w20050 = ~w19994 & ~w20049;
assign w20051 = w19997 & w20048;
assign w20052 = w19962 & ~w20046;
assign w20053 = w20050 & w65415;
assign w20054 = ~w20045 & ~w20053;
assign w20055 = w19973 & w20003;
assign w20056 = ~w19994 & ~w20027;
assign w20057 = ~w19955 & ~w20056;
assign w20058 = ~w20029 & ~w20055;
assign w20059 = ~w20057 & w20058;
assign w20060 = ~w20054 & w20059;
assign w20061 = pi1017 & ~w20060;
assign w20062 = ~pi1017 & w20060;
assign w20063 = ~w20061 & ~w20062;
assign w20064 = w19891 & ~w19910;
assign w20065 = ~w19859 & ~w19865;
assign w20066 = w19853 & w20065;
assign w20067 = w19821 & w20066;
assign w20068 = w19830 & ~w20065;
assign w20069 = w19845 & w20068;
assign w20070 = ~w19867 & ~w19892;
assign w20071 = ~w19830 & ~w20070;
assign w20072 = ~w19875 & ~w20067;
assign w20073 = ~w20069 & ~w20071;
assign w20074 = w20072 & w20073;
assign w20075 = w19854 & ~w19858;
assign w20076 = w19847 & w19865;
assign w20077 = w19875 & ~w20076;
assign w20078 = ~w19878 & ~w20075;
assign w20079 = w20077 & w20078;
assign w20080 = ~w19862 & w20079;
assign w20081 = ~w20074 & ~w20080;
assign w20082 = ~w20064 & ~w20081;
assign w20083 = ~pi0996 & w20082;
assign w20084 = pi0996 & ~w20082;
assign w20085 = ~w20083 & ~w20084;
assign w20086 = w19888 & ~w20065;
assign w20087 = ~w19861 & ~w19888;
assign w20088 = ~w19839 & w20087;
assign w20089 = ~w19896 & ~w20086;
assign w20090 = ~w20088 & w20089;
assign w20091 = w19875 & ~w20090;
assign w20092 = w19866 & w20068;
assign w20093 = ~w19855 & ~w19882;
assign w20094 = w19875 & ~w19905;
assign w20095 = ~w19902 & ~w20093;
assign w20096 = ~w20094 & w20095;
assign w20097 = ~w19875 & ~w19885;
assign w20098 = ~w19869 & ~w20092;
assign w20099 = ~w20097 & w20098;
assign w20100 = ~w20096 & w20099;
assign w20101 = ~w20091 & w20100;
assign w20102 = pi0997 & ~w20101;
assign w20103 = ~pi0997 & w20101;
assign w20104 = ~w20102 & ~w20103;
assign w20105 = w19828 & w19889;
assign w20106 = ~w19888 & ~w20105;
assign w20107 = ~w19881 & ~w20106;
assign w20108 = w19853 & ~w20076;
assign w20109 = ~w19859 & w19902;
assign w20110 = ~w20108 & ~w20109;
assign w20111 = ~w20066 & ~w20110;
assign w20112 = ~w19875 & ~w20105;
assign w20113 = ~w19863 & w20112;
assign w20114 = ~w20111 & w20113;
assign w20115 = w19853 & w19889;
assign w20116 = w19902 & w20115;
assign w20117 = w20077 & ~w20116;
assign w20118 = ~w19846 & w20117;
assign w20119 = ~w20114 & ~w20118;
assign w20120 = ~w20107 & ~w20119;
assign w20121 = ~pi0998 & w20120;
assign w20122 = pi0998 & ~w20120;
assign w20123 = ~w20121 & ~w20122;
assign w20124 = ~w19742 & w19752;
assign w20125 = ~w19801 & w19807;
assign w20126 = ~w19762 & ~w19802;
assign w20127 = w19753 & ~w20126;
assign w20128 = w19789 & ~w20124;
assign w20129 = ~w20125 & w20128;
assign w20130 = ~w20127 & w20129;
assign w20131 = w19742 & ~w19773;
assign w20132 = ~w19769 & ~w19792;
assign w20133 = ~w19727 & w20132;
assign w20134 = ~w20131 & ~w20133;
assign w20135 = w19757 & w19763;
assign w20136 = w19750 & ~w19757;
assign w20137 = ~w19768 & w20136;
assign w20138 = ~w19756 & ~w19789;
assign w20139 = ~w20135 & w20138;
assign w20140 = ~w20134 & w20139;
assign w20141 = ~w20137 & w20140;
assign w20142 = ~w20130 & ~w20141;
assign w20143 = pi1005 & w20142;
assign w20144 = ~pi1005 & ~w20142;
assign w20145 = ~w20143 & ~w20144;
assign w20146 = ~w19663 & ~w19682;
assign w20147 = ~w19655 & w20146;
assign w20148 = w19628 & ~w20147;
assign w20149 = ~w19654 & w19684;
assign w20150 = ~w19661 & ~w20149;
assign w20151 = ~w19641 & ~w20150;
assign w20152 = ~w20148 & ~w20151;
assign w20153 = ~w19673 & ~w20152;
assign w20154 = (w19641 & w19657) | (w19641 & w65416) | (w19657 & w65416);
assign w20155 = ~w19680 & ~w19703;
assign w20156 = ~w19704 & ~w20155;
assign w20157 = ~w19706 & ~w20156;
assign w20158 = (w19673 & w20157) | (w19673 & w65417) | (w20157 & w65417);
assign w20159 = ~w19641 & w19680;
assign w20160 = ~w19667 & ~w20159;
assign w20161 = w19704 & ~w20160;
assign w20162 = ~w19647 & ~w19662;
assign w20163 = ~w19675 & w20162;
assign w20164 = ~w19634 & w19641;
assign w20165 = ~w19701 & ~w19703;
assign w20166 = ~w20164 & w20165;
assign w20167 = w20163 & ~w20166;
assign w20168 = ~w19658 & ~w19676;
assign w20169 = ~w20167 & w20168;
assign w20170 = ~w19628 & ~w20169;
assign w20171 = ~w20158 & ~w20161;
assign w20172 = ~w20170 & w20171;
assign w20173 = ~w20153 & w20172;
assign w20174 = pi1001 & ~w20173;
assign w20175 = ~pi1001 & w20173;
assign w20176 = ~w20174 & ~w20175;
assign w20177 = ~pi3984 & pi9040;
assign w20178 = ~pi4032 & ~pi9040;
assign w20179 = ~w20177 & ~w20178;
assign w20180 = pi1098 & ~w20179;
assign w20181 = ~pi1098 & w20179;
assign w20182 = ~w20180 & ~w20181;
assign w20183 = ~pi3993 & pi9040;
assign w20184 = ~pi4006 & ~pi9040;
assign w20185 = ~w20183 & ~w20184;
assign w20186 = pi1136 & ~w20185;
assign w20187 = ~pi1136 & w20185;
assign w20188 = ~w20186 & ~w20187;
assign w20189 = ~w20182 & ~w20188;
assign w20190 = ~pi3990 & pi9040;
assign w20191 = ~pi4034 & ~pi9040;
assign w20192 = ~w20190 & ~w20191;
assign w20193 = pi1092 & ~w20192;
assign w20194 = ~pi1092 & w20192;
assign w20195 = ~w20193 & ~w20194;
assign w20196 = ~w20182 & w20195;
assign w20197 = ~pi4012 & pi9040;
assign w20198 = ~pi4002 & ~pi9040;
assign w20199 = ~w20197 & ~w20198;
assign w20200 = pi1111 & ~w20199;
assign w20201 = ~pi1111 & w20199;
assign w20202 = ~w20200 & ~w20201;
assign w20203 = ~pi3988 & pi9040;
assign w20204 = ~pi4031 & ~pi9040;
assign w20205 = ~w20203 & ~w20204;
assign w20206 = pi1080 & ~w20205;
assign w20207 = ~pi1080 & w20205;
assign w20208 = ~w20206 & ~w20207;
assign w20209 = ~w20202 & ~w20208;
assign w20210 = w20196 & w20209;
assign w20211 = ~w20188 & ~w20202;
assign w20212 = ~w20195 & w20208;
assign w20213 = w20211 & w20212;
assign w20214 = ~w20210 & ~w20213;
assign w20215 = ~w20189 & ~w20214;
assign w20216 = ~pi3991 & pi9040;
assign w20217 = ~pi4020 & ~pi9040;
assign w20218 = ~w20216 & ~w20217;
assign w20219 = pi1103 & ~w20218;
assign w20220 = ~pi1103 & w20218;
assign w20221 = ~w20219 & ~w20220;
assign w20222 = w20182 & ~w20195;
assign w20223 = ~w20196 & ~w20208;
assign w20224 = ~w20222 & w20223;
assign w20225 = w20223 & w65418;
assign w20226 = ~w20202 & w20222;
assign w20227 = ~w20225 & ~w20226;
assign w20228 = w20189 & w20208;
assign w20229 = w20182 & ~w20202;
assign w20230 = w20208 & ~w20229;
assign w20231 = ~w20223 & ~w20230;
assign w20232 = w20188 & w20231;
assign w20233 = ~w20210 & ~w20228;
assign w20234 = ~w20232 & w20233;
assign w20235 = w20227 & w20234;
assign w20236 = w20221 & ~w20235;
assign w20237 = ~w20188 & w20224;
assign w20238 = w20195 & w20208;
assign w20239 = w20202 & w20238;
assign w20240 = w20182 & w20239;
assign w20241 = ~w20237 & ~w20240;
assign w20242 = ~w20221 & ~w20241;
assign w20243 = w20182 & ~w20208;
assign w20244 = ~w20195 & w20243;
assign w20245 = ~w20230 & ~w20244;
assign w20246 = w20188 & ~w20221;
assign w20247 = w20211 & w20238;
assign w20248 = ~w20246 & ~w20247;
assign w20249 = ~w20245 & ~w20248;
assign w20250 = ~w20215 & ~w20249;
assign w20251 = ~w20242 & w20250;
assign w20252 = ~w20236 & w20251;
assign w20253 = pi1006 & w20252;
assign w20254 = ~pi1006 & ~w20252;
assign w20255 = ~w20253 & ~w20254;
assign w20256 = w19661 & w19680;
assign w20257 = ~w19677 & ~w20256;
assign w20258 = ~w19691 & ~w20257;
assign w20259 = ~w19654 & w19682;
assign w20260 = ~w19648 & ~w20259;
assign w20261 = ~w19665 & ~w19680;
assign w20262 = w19628 & ~w20261;
assign w20263 = ~w20154 & w20262;
assign w20264 = w19647 & w19681;
assign w20265 = w19691 & w20264;
assign w20266 = (w19673 & w20260) | (w19673 & w65419) | (w20260 & w65419);
assign w20267 = ~w20265 & w20266;
assign w20268 = ~w20263 & w20267;
assign w20269 = w19680 & w19682;
assign w20270 = ~w19654 & ~w19678;
assign w20271 = ~w19702 & w20155;
assign w20272 = ~w19676 & ~w20271;
assign w20273 = ~w19661 & ~w20272;
assign w20274 = ~w19666 & ~w20256;
assign w20275 = ~w19673 & ~w20269;
assign w20276 = w20274 & w20275;
assign w20277 = ~w20270 & w20276;
assign w20278 = ~w20273 & w20277;
assign w20279 = ~w20268 & ~w20278;
assign w20280 = ~w20258 & ~w20279;
assign w20281 = ~pi1002 & w20280;
assign w20282 = pi1002 & ~w20280;
assign w20283 = ~w20281 & ~w20282;
assign w20284 = ~pi3976 & pi9040;
assign w20285 = ~pi4017 & ~pi9040;
assign w20286 = ~w20284 & ~w20285;
assign w20287 = pi1122 & ~w20286;
assign w20288 = ~pi1122 & w20286;
assign w20289 = ~w20287 & ~w20288;
assign w20290 = ~pi4026 & pi9040;
assign w20291 = ~pi4000 & ~pi9040;
assign w20292 = ~w20290 & ~w20291;
assign w20293 = pi1089 & ~w20292;
assign w20294 = ~pi1089 & w20292;
assign w20295 = ~w20293 & ~w20294;
assign w20296 = w20289 & w20295;
assign w20297 = ~pi3997 & pi9040;
assign w20298 = ~pi3998 & ~pi9040;
assign w20299 = ~w20297 & ~w20298;
assign w20300 = pi1074 & ~w20299;
assign w20301 = ~pi1074 & w20299;
assign w20302 = ~w20300 & ~w20301;
assign w20303 = ~pi4028 & pi9040;
assign w20304 = ~pi4004 & ~pi9040;
assign w20305 = ~w20303 & ~w20304;
assign w20306 = pi1121 & ~w20305;
assign w20307 = ~pi1121 & w20305;
assign w20308 = ~w20306 & ~w20307;
assign w20309 = (~w20308 & ~w20296) | (~w20308 & w65420) | (~w20296 & w65420);
assign w20310 = ~pi3983 & pi9040;
assign w20311 = ~pi3986 & ~pi9040;
assign w20312 = ~w20310 & ~w20311;
assign w20313 = pi1120 & ~w20312;
assign w20314 = ~pi1120 & w20312;
assign w20315 = ~w20313 & ~w20314;
assign w20316 = w20295 & ~w20315;
assign w20317 = ~w20309 & w20316;
assign w20318 = ~w20289 & w20302;
assign w20319 = ~w20295 & w20315;
assign w20320 = w20318 & w20319;
assign w20321 = ~w20289 & ~w20302;
assign w20322 = w20295 & w20321;
assign w20323 = ~w20320 & ~w20322;
assign w20324 = w20308 & ~w20323;
assign w20325 = w20289 & ~w20295;
assign w20326 = ~w20302 & w20315;
assign w20327 = w20325 & w20326;
assign w20328 = ~pi4010 & pi9040;
assign w20329 = ~pi4011 & ~pi9040;
assign w20330 = ~w20328 & ~w20329;
assign w20331 = pi1099 & ~w20330;
assign w20332 = ~pi1099 & w20330;
assign w20333 = ~w20331 & ~w20332;
assign w20334 = ~w20289 & ~w20295;
assign w20335 = ~w20315 & w20334;
assign w20336 = w20302 & w20325;
assign w20337 = ~w20335 & ~w20336;
assign w20338 = ~w20308 & ~w20337;
assign w20339 = w20302 & w20308;
assign w20340 = w20296 & w20339;
assign w20341 = ~w20327 & w20333;
assign w20342 = ~w20340 & w20341;
assign w20343 = ~w20317 & w20342;
assign w20344 = ~w20324 & ~w20338;
assign w20345 = w20343 & w20344;
assign w20346 = w20295 & w20315;
assign w20347 = w20318 & w20346;
assign w20348 = ~w20333 & ~w20347;
assign w20349 = w20308 & ~w20337;
assign w20350 = w20319 & w20321;
assign w20351 = w20296 & w20315;
assign w20352 = w20296 & w20326;
assign w20353 = ~w20350 & ~w20352;
assign w20354 = w20348 & ~w20349;
assign w20355 = w20353 & w20354;
assign w20356 = ~w20345 & ~w20355;
assign w20357 = w20321 & w20316;
assign w20358 = ~w20302 & w20325;
assign w20359 = w20295 & w20302;
assign w20360 = ~w20358 & ~w20359;
assign w20361 = ~w20357 & w20360;
assign w20362 = ~w20333 & ~w20361;
assign w20363 = ~w20295 & w20326;
assign w20364 = ~w20347 & ~w20363;
assign w20365 = ~w20362 & w20364;
assign w20366 = ~w20308 & ~w20365;
assign w20367 = ~w20356 & ~w20366;
assign w20368 = ~pi1007 & w20367;
assign w20369 = pi1007 & ~w20367;
assign w20370 = ~w20368 & ~w20369;
assign w20371 = w20202 & ~w20238;
assign w20372 = w20196 & w20371;
assign w20373 = w20202 & w20208;
assign w20374 = w20222 & w20373;
assign w20375 = ~w20211 & ~w20374;
assign w20376 = ~w20195 & ~w20208;
assign w20377 = ~w20229 & w20376;
assign w20378 = ~w20239 & ~w20377;
assign w20379 = ~w20182 & w20202;
assign w20380 = w20188 & ~w20379;
assign w20381 = ~w20378 & ~w20380;
assign w20382 = w20243 & ~w20377;
assign w20383 = (w20188 & w20382) | (w20188 & w63737) | (w20382 & w63737);
assign w20384 = w20214 & ~w20381;
assign w20385 = w20384 & w63738;
assign w20386 = (~w20221 & w20385) | (~w20221 & w65421) | (w20385 & w65421);
assign w20387 = ~w20196 & w20246;
assign w20388 = ~w20382 & w65422;
assign w20389 = w20227 & w20388;
assign w20390 = (w20221 & ~w20384) | (w20221 & w65423) | (~w20384 & w65423);
assign w20391 = ~w20196 & ~w20209;
assign w20392 = ~w20379 & w20391;
assign w20393 = w20391 & w65424;
assign w20394 = ~w20182 & w20393;
assign w20395 = w20195 & ~w20211;
assign w20396 = w20229 & w20395;
assign w20397 = ~w20394 & ~w20396;
assign w20398 = ~w20389 & w20397;
assign w20399 = ~w20390 & w20398;
assign w20400 = ~w20386 & w20399;
assign w20401 = pi1008 & ~w20400;
assign w20402 = ~pi1008 & w20400;
assign w20403 = ~w20401 & ~w20402;
assign w20404 = w20211 & w20377;
assign w20405 = ~w20221 & ~w20393;
assign w20406 = ~w20243 & w20371;
assign w20407 = w20195 & ~w20202;
assign w20408 = ~w20231 & w20407;
assign w20409 = w20221 & ~w20406;
assign w20410 = ~w20408 & w20409;
assign w20411 = ~w20188 & ~w20405;
assign w20412 = ~w20410 & w20411;
assign w20413 = w20238 & w20379;
assign w20414 = w20212 & w20229;
assign w20415 = ~w20413 & ~w20414;
assign w20416 = ~w20221 & ~w20415;
assign w20417 = ~w20376 & w20379;
assign w20418 = ~w20209 & ~w20417;
assign w20419 = w20222 & w20209;
assign w20420 = w20221 & ~w20419;
assign w20421 = ~w20418 & ~w20420;
assign w20422 = ~w20209 & ~w20222;
assign w20423 = ~w20376 & ~w20422;
assign w20424 = ~w20413 & ~w20423;
assign w20425 = w20221 & w20392;
assign w20426 = w20424 & w20425;
assign w20427 = ~w20239 & ~w20421;
assign w20428 = ~w20426 & w20427;
assign w20429 = w20188 & ~w20428;
assign w20430 = ~w20215 & ~w20404;
assign w20431 = ~w20416 & w20430;
assign w20432 = ~w20412 & w20431;
assign w20433 = ~w20429 & w20432;
assign w20434 = pi1000 & ~w20433;
assign w20435 = ~pi1000 & w20433;
assign w20436 = ~w20434 & ~w20435;
assign w20437 = w20028 & ~w20050;
assign w20438 = w19942 & w20020;
assign w20439 = w19932 & ~w19984;
assign w20440 = w19986 & w20439;
assign w20441 = w19955 & w20013;
assign w20442 = ~w20440 & ~w20441;
assign w20443 = w20017 & w20442;
assign w20444 = w19939 & ~w19955;
assign w20445 = w20002 & w20444;
assign w20446 = w19993 & ~w20439;
assign w20447 = w19976 & w20012;
assign w20448 = w19962 & ~w20447;
assign w20449 = ~w20445 & w20448;
assign w20450 = ~w20446 & w20449;
assign w20451 = ~w20443 & ~w20450;
assign w20452 = ~w20437 & ~w20438;
assign w20453 = ~w20451 & w20452;
assign w20454 = pi1040 & ~w20453;
assign w20455 = ~pi1040 & w20453;
assign w20456 = ~w20454 & ~w20455;
assign w20457 = ~w20302 & ~w20308;
assign w20458 = ~w20319 & ~w20457;
assign w20459 = w20289 & ~w20458;
assign w20460 = ~w20458 & w65425;
assign w20461 = w20308 & w20352;
assign w20462 = ~w20346 & ~w20358;
assign w20463 = w20309 & ~w20462;
assign w20464 = ~w20318 & ~w20358;
assign w20465 = ~w20315 & ~w20464;
assign w20466 = ~w20333 & ~w20460;
assign w20467 = ~w20461 & ~w20463;
assign w20468 = w20467 & w65426;
assign w20469 = w20334 & w20457;
assign w20470 = w20302 & w20316;
assign w20471 = w20316 & w63739;
assign w20472 = w20333 & ~w20471;
assign w20473 = ~w20320 & w20353;
assign w20474 = ~w20308 & ~w20473;
assign w20475 = ~w20319 & w20339;
assign w20476 = ~w20469 & ~w20475;
assign w20477 = ~w20357 & w20476;
assign w20478 = w20472 & w20477;
assign w20479 = ~w20474 & w20478;
assign w20480 = ~w20468 & ~w20479;
assign w20481 = w20302 & ~w20315;
assign w20482 = ~w20295 & ~w20326;
assign w20483 = ~w20339 & ~w20481;
assign w20484 = w20482 & w20483;
assign w20485 = w20459 & w20484;
assign w20486 = ~w20350 & ~w20470;
assign w20487 = w20308 & ~w20486;
assign w20488 = ~w20485 & ~w20487;
assign w20489 = ~w20480 & w20488;
assign w20490 = ~pi1020 & ~w20489;
assign w20491 = pi1020 & w20489;
assign w20492 = ~w20490 & ~w20491;
assign w20493 = w20211 & ~w20422;
assign w20494 = w20395 & w20418;
assign w20495 = w20420 & ~w20493;
assign w20496 = ~w20494 & w20495;
assign w20497 = (w20188 & w20423) | (w20188 & w65427) | (w20423 & w65427);
assign w20498 = (~w20188 & w20372) | (~w20188 & w65428) | (w20372 & w65428);
assign w20499 = ~w20221 & ~w20247;
assign w20500 = ~w20394 & w20499;
assign w20501 = ~w20497 & ~w20498;
assign w20502 = w20500 & w20501;
assign w20503 = ~w20496 & ~w20502;
assign w20504 = w20188 & ~w20374;
assign w20505 = ~w20225 & w20504;
assign w20506 = ~w20195 & ~w20418;
assign w20507 = ~w20188 & ~w20240;
assign w20508 = ~w20506 & w20507;
assign w20509 = ~w20505 & ~w20508;
assign w20510 = ~w20503 & ~w20509;
assign w20511 = pi1021 & ~w20510;
assign w20512 = ~pi1021 & w20510;
assign w20513 = ~w20511 & ~w20512;
assign w20514 = (w19789 & w19782) | (w19789 & w65429) | (w19782 & w65429);
assign w20515 = ~w19761 & ~w19789;
assign w20516 = (~w19742 & w19777) | (~w19742 & w63740) | (w19777 & w63740);
assign w20517 = ~w20515 & w20516;
assign w20518 = w19777 & ~w19789;
assign w20519 = w19742 & ~w19756;
assign w20520 = ~w20518 & w20519;
assign w20521 = ~w20517 & ~w20520;
assign w20522 = ~w20514 & ~w20521;
assign w20523 = ~pi1012 & w20522;
assign w20524 = pi1012 & ~w20522;
assign w20525 = ~w20523 & ~w20524;
assign w20526 = ~pi4031 & pi9040;
assign w20527 = ~pi4009 & ~pi9040;
assign w20528 = ~w20526 & ~w20527;
assign w20529 = pi1162 & ~w20528;
assign w20530 = ~pi1162 & w20528;
assign w20531 = ~w20529 & ~w20530;
assign w20532 = ~pi4032 & pi9040;
assign w20533 = ~pi3977 & ~pi9040;
assign w20534 = ~w20532 & ~w20533;
assign w20535 = pi1110 & ~w20534;
assign w20536 = ~pi1110 & w20534;
assign w20537 = ~w20535 & ~w20536;
assign w20538 = w20531 & ~w20537;
assign w20539 = ~pi4002 & pi9040;
assign w20540 = ~pi3982 & ~pi9040;
assign w20541 = ~w20539 & ~w20540;
assign w20542 = pi1095 & ~w20541;
assign w20543 = ~pi1095 & w20541;
assign w20544 = ~w20542 & ~w20543;
assign w20545 = ~pi4003 & pi9040;
assign w20546 = ~pi4019 & ~pi9040;
assign w20547 = ~w20545 & ~w20546;
assign w20548 = pi1098 & ~w20547;
assign w20549 = ~pi1098 & w20547;
assign w20550 = ~w20548 & ~w20549;
assign w20551 = ~w20544 & ~w20550;
assign w20552 = w20544 & w20550;
assign w20553 = ~w20551 & ~w20552;
assign w20554 = w20538 & w20553;
assign w20555 = ~w20531 & w20537;
assign w20556 = ~pi4005 & pi9040;
assign w20557 = ~pi4001 & ~pi9040;
assign w20558 = ~w20556 & ~w20557;
assign w20559 = pi1115 & ~w20558;
assign w20560 = ~pi1115 & w20558;
assign w20561 = ~w20559 & ~w20560;
assign w20562 = ~w20555 & ~w20561;
assign w20563 = w20537 & ~w20550;
assign w20564 = ~w20544 & ~w20563;
assign w20565 = w20531 & w20537;
assign w20566 = ~w20531 & ~w20550;
assign w20567 = ~w20565 & ~w20566;
assign w20568 = w20564 & ~w20567;
assign w20569 = ~w20563 & w63741;
assign w20570 = ~w20568 & w63742;
assign w20571 = (~w20554 & w20570) | (~w20554 & w65430) | (w20570 & w65430);
assign w20572 = ~pi3999 & pi9040;
assign w20573 = ~pi3990 & ~pi9040;
assign w20574 = ~w20572 & ~w20573;
assign w20575 = pi1080 & ~w20574;
assign w20576 = ~pi1080 & w20574;
assign w20577 = ~w20575 & ~w20576;
assign w20578 = ~w20571 & w20577;
assign w20579 = ~w20551 & w20561;
assign w20580 = ~w20555 & w20561;
assign w20581 = ~w20579 & ~w20580;
assign w20582 = w20537 & w20552;
assign w20583 = ~w20581 & ~w20582;
assign w20584 = ~w20538 & w20544;
assign w20585 = w20531 & w20550;
assign w20586 = w20584 & ~w20585;
assign w20587 = w20584 & w65431;
assign w20588 = ~w20554 & ~w20587;
assign w20589 = w20583 & ~w20588;
assign w20590 = ~w20561 & w20565;
assign w20591 = w20551 & w20590;
assign w20592 = ~w20537 & ~w20561;
assign w20593 = w20552 & w20592;
assign w20594 = w20538 & w20551;
assign w20595 = ~w20561 & ~w20569;
assign w20596 = ~w20537 & w20550;
assign w20597 = ~w20531 & w20596;
assign w20598 = w20595 & ~w20597;
assign w20599 = ~w20583 & ~w20598;
assign w20600 = ~w20555 & w20586;
assign w20601 = ~w20593 & ~w20594;
assign w20602 = ~w20600 & w20601;
assign w20603 = ~w20599 & w20602;
assign w20604 = ~w20577 & ~w20603;
assign w20605 = ~w20589 & ~w20591;
assign w20606 = ~w20578 & w20605;
assign w20607 = ~w20604 & w20606;
assign w20608 = pi1046 & w20607;
assign w20609 = ~pi1046 & ~w20607;
assign w20610 = ~w20608 & ~w20609;
assign w20611 = w19635 & w19703;
assign w20612 = w19628 & ~w19663;
assign w20613 = ~w20166 & w20612;
assign w20614 = ~w20163 & ~w20259;
assign w20615 = ~w19694 & w20155;
assign w20616 = w20614 & w20615;
assign w20617 = ~w19673 & ~w20613;
assign w20618 = ~w20616 & w20617;
assign w20619 = ~w19628 & ~w20614;
assign w20620 = w19702 & ~w20146;
assign w20621 = ~w19695 & ~w20159;
assign w20622 = w19674 & w20621;
assign w20623 = ~w20620 & w20622;
assign w20624 = ~w20619 & w20623;
assign w20625 = ~w20618 & ~w20624;
assign w20626 = w19691 & ~w20274;
assign w20627 = ~w19664 & ~w20611;
assign w20628 = ~w20626 & w20627;
assign w20629 = ~w20625 & w20628;
assign w20630 = pi1014 & ~w20629;
assign w20631 = ~pi1014 & w20629;
assign w20632 = ~w20630 & ~w20631;
assign w20633 = w20553 & w20555;
assign w20634 = w20551 & w20565;
assign w20635 = ~w20531 & w20544;
assign w20636 = w20596 & ~w20635;
assign w20637 = ~w20563 & w20580;
assign w20638 = ~w20636 & w20637;
assign w20639 = w20579 & ~w20638;
assign w20640 = ~w20538 & ~w20553;
assign w20641 = w20562 & w20640;
assign w20642 = ~w20633 & ~w20634;
assign w20643 = ~w20641 & w20642;
assign w20644 = ~w20639 & w20643;
assign w20645 = w20577 & ~w20644;
assign w20646 = ~w20553 & ~w20555;
assign w20647 = ~w20538 & w20577;
assign w20648 = ~w20561 & ~w20647;
assign w20649 = ~w20633 & w20648;
assign w20650 = ~w20646 & w20649;
assign w20651 = w20563 & w20635;
assign w20652 = ~w20594 & ~w20651;
assign w20653 = w20561 & ~w20652;
assign w20654 = ~w20554 & ~w20577;
assign w20655 = w20638 & w20654;
assign w20656 = ~w20650 & ~w20653;
assign w20657 = ~w20655 & w20656;
assign w20658 = ~w20645 & w20657;
assign w20659 = pi1018 & w20658;
assign w20660 = ~pi1018 & ~w20658;
assign w20661 = ~w20659 & ~w20660;
assign w20662 = w20566 & w20579;
assign w20663 = ~w20563 & w65432;
assign w20664 = (~w20552 & ~w20595) | (~w20552 & w65433) | (~w20595 & w65433);
assign w20665 = ~w20584 & ~w20664;
assign w20666 = ~w20662 & ~w20665;
assign w20667 = ~w20577 & ~w20666;
assign w20668 = ~w20537 & ~w20544;
assign w20669 = ~w20550 & ~w20565;
assign w20670 = ~w20635 & w20669;
assign w20671 = ~w20582 & ~w20668;
assign w20672 = ~w20670 & w20671;
assign w20673 = w20561 & ~w20672;
assign w20674 = ~w20537 & w20635;
assign w20675 = ~w20569 & ~w20674;
assign w20676 = ~w20561 & ~w20675;
assign w20677 = ~w20673 & w63743;
assign w20678 = w20577 & ~w20677;
assign w20679 = ~w20544 & w20590;
assign w20680 = w20552 & w20555;
assign w20681 = ~w20563 & ~w20597;
assign w20682 = w20579 & ~w20681;
assign w20683 = ~w20653 & ~w20682;
assign w20684 = ~w20552 & ~w20662;
assign w20685 = ~w20679 & ~w20680;
assign w20686 = (w20685 & w20683) | (w20685 & w65434) | (w20683 & w65434);
assign w20687 = ~w20678 & w20686;
assign w20688 = w20687 & w65435;
assign w20689 = (pi1019 & ~w20687) | (pi1019 & w65436) | (~w20687 & w65436);
assign w20690 = ~w20688 & ~w20689;
assign w20691 = w20334 & w20481;
assign w20692 = ~w20471 & ~w20691;
assign w20693 = ~w20320 & ~w20327;
assign w20694 = ~w20357 & w20693;
assign w20695 = w20692 & w20694;
assign w20696 = (~w20472 & ~w20694) | (~w20472 & w63744) | (~w20694 & w63744);
assign w20697 = (~w20308 & w20696) | (~w20308 & w65437) | (w20696 & w65437);
assign w20698 = w20325 & ~w20333;
assign w20699 = w20458 & w20698;
assign w20700 = w20308 & ~w20325;
assign w20701 = w20348 & w20700;
assign w20702 = ~w20325 & w20326;
assign w20703 = w20309 & ~w20702;
assign w20704 = ~w20315 & w20321;
assign w20705 = w20308 & ~w20704;
assign w20706 = ~w20459 & w20705;
assign w20707 = ~w20703 & ~w20706;
assign w20708 = ~w20347 & ~w20460;
assign w20709 = w20692 & w20708;
assign w20710 = ~w20707 & w20709;
assign w20711 = w20333 & ~w20710;
assign w20712 = (~w20699 & ~w20695) | (~w20699 & w65438) | (~w20695 & w65438);
assign w20713 = ~w20697 & w20712;
assign w20714 = ~w20711 & w20713;
assign w20715 = pi1010 & ~w20714;
assign w20716 = ~pi1010 & w20714;
assign w20717 = ~w20715 & ~w20716;
assign w20718 = ~w19759 & w19795;
assign w20719 = ~w19795 & w19807;
assign w20720 = w20132 & w20719;
assign w20721 = (~w19742 & w20720) | (~w19742 & w65439) | (w20720 & w65439);
assign w20722 = ~w19754 & w19801;
assign w20723 = (~w19790 & ~w20132) | (~w19790 & w65440) | (~w20132 & w65440);
assign w20724 = ~w20722 & w20723;
assign w20725 = ~w20516 & w20724;
assign w20726 = (w19789 & w20725) | (w19789 & w65441) | (w20725 & w65441);
assign w20727 = w19729 & w19735;
assign w20728 = ~w19755 & w19803;
assign w20729 = (~w19792 & w20727) | (~w19792 & w65442) | (w20727 & w65442);
assign w20730 = w19720 & w19749;
assign w20731 = ~w19807 & w20730;
assign w20732 = (~w19742 & ~w19795) | (~w19742 & w65443) | (~w19795 & w65443);
assign w20733 = ~w20132 & w20732;
assign w20734 = ~w20731 & ~w20733;
assign w20735 = ~w20729 & w20734;
assign w20736 = ~w19789 & ~w20735;
assign w20737 = w19768 & ~w19804;
assign w20738 = ~w19753 & ~w20737;
assign w20739 = ~w20736 & ~w20738;
assign w20740 = ~w20726 & w20739;
assign w20741 = ~pi1011 & w20740;
assign w20742 = pi1011 & ~w20740;
assign w20743 = ~w20741 & ~w20742;
assign w20744 = ~pi4035 & pi9040;
assign w20745 = ~pi4018 & ~pi9040;
assign w20746 = ~w20744 & ~w20745;
assign w20747 = pi1128 & ~w20746;
assign w20748 = ~pi1128 & w20746;
assign w20749 = ~w20747 & ~w20748;
assign w20750 = ~pi3980 & pi9040;
assign w20751 = ~pi4014 & ~pi9040;
assign w20752 = ~w20750 & ~w20751;
assign w20753 = pi1099 & ~w20752;
assign w20754 = ~pi1099 & w20752;
assign w20755 = ~w20753 & ~w20754;
assign w20756 = ~w20749 & ~w20755;
assign w20757 = ~pi3985 & pi9040;
assign w20758 = ~pi3975 & ~pi9040;
assign w20759 = ~w20757 & ~w20758;
assign w20760 = pi1127 & ~w20759;
assign w20761 = ~pi1127 & w20759;
assign w20762 = ~w20760 & ~w20761;
assign w20763 = ~w20756 & ~w20762;
assign w20764 = w20756 & w20762;
assign w20765 = ~w20763 & ~w20764;
assign w20766 = w20749 & w20755;
assign w20767 = ~pi4016 & pi9040;
assign w20768 = ~pi4015 & ~pi9040;
assign w20769 = ~w20767 & ~w20768;
assign w20770 = pi1082 & ~w20769;
assign w20771 = ~pi1082 & w20769;
assign w20772 = ~w20770 & ~w20771;
assign w20773 = ~w20766 & w20772;
assign w20774 = ~w20765 & w20773;
assign w20775 = ~pi3987 & pi9040;
assign w20776 = ~pi3979 & ~pi9040;
assign w20777 = ~w20775 & ~w20776;
assign w20778 = pi1122 & ~w20777;
assign w20779 = ~pi1122 & w20777;
assign w20780 = ~w20778 & ~w20779;
assign w20781 = w20756 & w20780;
assign w20782 = ~w20765 & w65444;
assign w20783 = ~w20762 & ~w20780;
assign w20784 = w20756 & w20783;
assign w20785 = w20749 & ~w20780;
assign w20786 = ~w20755 & ~w20762;
assign w20787 = ~w20756 & ~w20786;
assign w20788 = ~w20785 & ~w20787;
assign w20789 = ~w20749 & w20780;
assign w20790 = w20755 & ~w20785;
assign w20791 = ~w20789 & w20790;
assign w20792 = ~w20788 & ~w20791;
assign w20793 = (~w20784 & ~w20792) | (~w20784 & w20874) | (~w20792 & w20874);
assign w20794 = ~pi4000 & pi9040;
assign w20795 = ~pi4008 & ~pi9040;
assign w20796 = ~w20794 & ~w20795;
assign w20797 = pi1094 & ~w20796;
assign w20798 = ~pi1094 & w20796;
assign w20799 = ~w20797 & ~w20798;
assign w20800 = ~w20793 & w20799;
assign w20801 = w20762 & ~w20780;
assign w20802 = ~w20756 & ~w20766;
assign w20803 = w20801 & ~w20802;
assign w20804 = w20762 & w20780;
assign w20805 = w20749 & w20799;
assign w20806 = w20802 & ~w20805;
assign w20807 = w20804 & w20806;
assign w20808 = ~w20803 & ~w20807;
assign w20809 = ~w20762 & w20780;
assign w20810 = (w20809 & ~w20802) | (w20809 & w65445) | (~w20802 & w65445);
assign w20811 = w20802 & w65446;
assign w20812 = ~w20810 & ~w20811;
assign w20813 = w20808 & w20812;
assign w20814 = ~w20772 & ~w20813;
assign w20815 = w20801 & w20805;
assign w20816 = w20772 & ~w20799;
assign w20817 = ~w20756 & w20816;
assign w20818 = ~w20792 & w20817;
assign w20819 = ~w20782 & ~w20815;
assign w20820 = ~w20818 & w20819;
assign w20821 = ~w20800 & w20820;
assign w20822 = ~w20814 & w20821;
assign w20823 = pi1024 & ~w20822;
assign w20824 = ~pi1024 & w20822;
assign w20825 = ~w20823 & ~w20824;
assign w20826 = ~w20634 & ~w20680;
assign w20827 = w20579 & ~w20585;
assign w20828 = w20681 & w20827;
assign w20829 = ~w20593 & w20826;
assign w20830 = ~w20828 & w20829;
assign w20831 = w20577 & ~w20830;
assign w20832 = w20585 & w20668;
assign w20833 = ~w20581 & ~w20832;
assign w20834 = ~w20561 & ~w20651;
assign w20835 = ~w20568 & w20834;
assign w20836 = ~w20833 & ~w20835;
assign w20837 = ~w20561 & w20681;
assign w20838 = w20826 & w20837;
assign w20839 = ~w20663 & ~w20682;
assign w20840 = ~w20838 & w20839;
assign w20841 = ~w20577 & ~w20840;
assign w20842 = ~w20831 & ~w20836;
assign w20843 = ~w20841 & w20842;
assign w20844 = ~pi1025 & w20843;
assign w20845 = pi1025 & ~w20843;
assign w20846 = ~w20844 & ~w20845;
assign w20847 = ~w20749 & w20809;
assign w20848 = w20799 & ~w20847;
assign w20849 = ~w20766 & w20848;
assign w20850 = ~w20808 & w20849;
assign w20851 = w20755 & w20801;
assign w20852 = ~w20799 & w20851;
assign w20853 = ~w20755 & ~w20780;
assign w20854 = (~w20853 & ~w20790) | (~w20853 & w63745) | (~w20790 & w63745);
assign w20855 = w20763 & ~w20854;
assign w20856 = w20755 & w20762;
assign w20857 = ~w20749 & ~w20799;
assign w20858 = ~w20786 & w20857;
assign w20859 = ~w20856 & w20858;
assign w20860 = ~w20799 & ~w20802;
assign w20861 = (w20809 & w20802) | (w20809 & w65447) | (w20802 & w65447);
assign w20862 = ~w20789 & ~w20853;
assign w20863 = ~w20856 & w20862;
assign w20864 = ~w20861 & ~w20863;
assign w20865 = w20765 & ~w20864;
assign w20866 = w20772 & ~w20859;
assign w20867 = ~w20855 & w20866;
assign w20868 = ~w20865 & w20867;
assign w20869 = w20749 & w20854;
assign w20870 = ~w20799 & ~w20858;
assign w20871 = ~w20869 & w20870;
assign w20872 = ~w20756 & w20799;
assign w20873 = w20854 & w20872;
assign w20874 = ~w20772 & ~w20784;
assign w20875 = ~w20873 & w20874;
assign w20876 = ~w20871 & w20875;
assign w20877 = ~w20868 & ~w20876;
assign w20878 = ~w20850 & ~w20852;
assign w20879 = ~w20877 & w20878;
assign w20880 = pi1035 & ~w20879;
assign w20881 = ~pi1035 & w20879;
assign w20882 = ~w20880 & ~w20881;
assign w20883 = ~w20784 & ~w20787;
assign w20884 = ~w20851 & ~w20883;
assign w20885 = w20884 & w63746;
assign w20886 = ~w20860 & ~w20870;
assign w20887 = ~w20884 & w20886;
assign w20888 = ~w20885 & ~w20887;
assign w20889 = w20772 & ~w20861;
assign w20890 = w20888 & w20889;
assign w20891 = ~w20772 & ~w20888;
assign w20892 = ~w20812 & w20849;
assign w20893 = ~w20869 & w65448;
assign w20894 = ~w20892 & ~w20893;
assign w20895 = ~w20890 & w20894;
assign w20896 = (pi1036 & ~w20895) | (pi1036 & w65449) | (~w20895 & w65449);
assign w20897 = w20895 & w65450;
assign w20898 = ~w20896 & ~w20897;
assign w20899 = ~w20799 & ~w20863;
assign w20900 = ~w20789 & w20856;
assign w20901 = w20848 & ~w20900;
assign w20902 = ~w20899 & ~w20901;
assign w20903 = w20884 & w65451;
assign w20904 = ~w20902 & ~w20903;
assign w20905 = ~w20772 & ~w20904;
assign w20906 = ~w20773 & ~w20857;
assign w20907 = w20804 & ~w20906;
assign w20908 = w20774 & w20848;
assign w20909 = w20801 & w20873;
assign w20910 = ~w20781 & ~w20856;
assign w20911 = w20816 & ~w20910;
assign w20912 = ~w20907 & ~w20911;
assign w20913 = ~w20908 & w20912;
assign w20914 = ~w20909 & w20913;
assign w20915 = ~w20905 & w20914;
assign w20916 = pi1037 & ~w20915;
assign w20917 = ~pi1037 & w20915;
assign w20918 = ~w20916 & ~w20917;
assign w20919 = ~w20340 & ~w20704;
assign w20920 = w20348 & w20919;
assign w20921 = ~w20352 & ~w20484;
assign w20922 = w20920 & w20921;
assign w20923 = w20308 & ~w20464;
assign w20924 = w20333 & ~w20350;
assign w20925 = ~w20923 & w20924;
assign w20926 = ~w20922 & ~w20925;
assign w20927 = w20308 & ~w20351;
assign w20928 = ~w20691 & w20927;
assign w20929 = w20289 & w20316;
assign w20930 = ~w20322 & ~w20929;
assign w20931 = w20333 & ~w20930;
assign w20932 = ~w20308 & ~w20336;
assign w20933 = ~w20931 & w20932;
assign w20934 = ~w20928 & ~w20933;
assign w20935 = ~w20926 & ~w20934;
assign w20936 = ~pi1039 & w20935;
assign w20937 = pi1039 & ~w20935;
assign w20938 = ~w20936 & ~w20937;
assign w20939 = ~pi4210 & pi9040;
assign w20940 = ~pi3947 & ~pi9040;
assign w20941 = ~w20939 & ~w20940;
assign w20942 = pi1182 & ~w20941;
assign w20943 = ~pi1182 & w20941;
assign w20944 = ~w20942 & ~w20943;
assign w20945 = ~pi3937 & pi9040;
assign w20946 = ~pi4277 & ~pi9040;
assign w20947 = ~w20945 & ~w20946;
assign w20948 = pi1146 & ~w20947;
assign w20949 = ~pi1146 & w20947;
assign w20950 = ~w20948 & ~w20949;
assign w20951 = ~pi4025 & pi9040;
assign w20952 = ~pi3954 & ~pi9040;
assign w20953 = ~w20951 & ~w20952;
assign w20954 = pi1175 & ~w20953;
assign w20955 = ~pi1175 & w20953;
assign w20956 = ~w20954 & ~w20955;
assign w20957 = ~pi3934 & pi9040;
assign w20958 = ~pi3971 & ~pi9040;
assign w20959 = ~w20957 & ~w20958;
assign w20960 = pi1131 & ~w20959;
assign w20961 = ~pi1131 & w20959;
assign w20962 = ~w20960 & ~w20961;
assign w20963 = ~w20956 & w20962;
assign w20964 = ~pi3932 & pi9040;
assign w20965 = ~pi3953 & ~pi9040;
assign w20966 = ~w20964 & ~w20965;
assign w20967 = pi1177 & ~w20966;
assign w20968 = ~pi1177 & w20966;
assign w20969 = ~w20967 & ~w20968;
assign w20970 = ~w20962 & ~w20969;
assign w20971 = ~pi3933 & pi9040;
assign w20972 = ~pi4119 & ~pi9040;
assign w20973 = ~w20971 & ~w20972;
assign w20974 = pi1167 & ~w20973;
assign w20975 = ~pi1167 & w20973;
assign w20976 = ~w20974 & ~w20975;
assign w20977 = w20970 & w20976;
assign w20978 = ~w20963 & ~w20977;
assign w20979 = ~w20944 & ~w20969;
assign w20980 = ~w20970 & ~w20976;
assign w20981 = ~w20979 & w20980;
assign w20982 = w20978 & ~w20981;
assign w20983 = w20956 & w20969;
assign w20984 = ~w20944 & w20983;
assign w20985 = w20962 & w20976;
assign w20986 = w20956 & w20985;
assign w20987 = ~w20984 & ~w20986;
assign w20988 = ~w20950 & w20987;
assign w20989 = w20982 & w20988;
assign w20990 = w20956 & ~w20962;
assign w20991 = ~w20976 & w20990;
assign w20992 = w20962 & w20969;
assign w20993 = ~w20970 & ~w20992;
assign w20994 = ~w20956 & ~w20993;
assign w20995 = w20956 & w20993;
assign w20996 = ~w20994 & ~w20995;
assign w20997 = w20985 & w20996;
assign w20998 = ~w20989 & ~w20991;
assign w20999 = ~w20997 & w20998;
assign w21000 = ~w20944 & ~w20999;
assign w21001 = ~w20956 & ~w20976;
assign w21002 = w20944 & w20969;
assign w21003 = w21001 & w21002;
assign w21004 = w20944 & ~w20978;
assign w21005 = w20950 & ~w20984;
assign w21006 = ~w20990 & ~w20992;
assign w21007 = ~w20982 & w21006;
assign w21008 = ~w21004 & w21005;
assign w21009 = ~w21007 & w21008;
assign w21010 = w20944 & ~w20983;
assign w21011 = w20986 & w21010;
assign w21012 = ~w20969 & w20991;
assign w21013 = ~w20950 & ~w21011;
assign w21014 = ~w21012 & w21013;
assign w21015 = ~w20976 & w20992;
assign w21016 = ~w20984 & w21015;
assign w21017 = ~w20963 & ~w20990;
assign w21018 = w20976 & w20993;
assign w21019 = ~w21017 & w21018;
assign w21020 = w21018 & w63747;
assign w21021 = ~w21016 & ~w21020;
assign w21022 = ~w20969 & ~w21001;
assign w21023 = ~w21015 & ~w21022;
assign w21024 = w21010 & ~w21023;
assign w21025 = ~w20994 & ~w21015;
assign w21026 = ~w21001 & ~w21025;
assign w21027 = w21024 & w21026;
assign w21028 = w21014 & w21021;
assign w21029 = ~w21027 & w21028;
assign w21030 = ~w21009 & ~w21029;
assign w21031 = ~w21000 & ~w21003;
assign w21032 = ~w21030 & w21031;
assign w21033 = ~pi4266 & pi9040;
assign w21034 = ~pi4138 & ~pi9040;
assign w21035 = ~w21033 & ~w21034;
assign w21036 = pi1151 & ~w21035;
assign w21037 = ~pi1151 & w21035;
assign w21038 = ~w21036 & ~w21037;
assign w21039 = ~pi4043 & pi9040;
assign w21040 = ~pi3967 & ~pi9040;
assign w21041 = ~w21039 & ~w21040;
assign w21042 = pi1130 & ~w21041;
assign w21043 = ~pi1130 & w21041;
assign w21044 = ~w21042 & ~w21043;
assign w21045 = ~w21038 & ~w21044;
assign w21046 = ~pi3955 & pi9040;
assign w21047 = ~pi4117 & ~pi9040;
assign w21048 = ~w21046 & ~w21047;
assign w21049 = pi1166 & ~w21048;
assign w21050 = ~pi1166 & w21048;
assign w21051 = ~w21049 & ~w21050;
assign w21052 = ~pi3951 & pi9040;
assign w21053 = ~pi3966 & ~pi9040;
assign w21054 = ~w21052 & ~w21053;
assign w21055 = pi1160 & ~w21054;
assign w21056 = ~pi1160 & w21054;
assign w21057 = ~w21055 & ~w21056;
assign w21058 = ~w21051 & w21057;
assign w21059 = w21038 & w21044;
assign w21060 = ~w21045 & ~w21059;
assign w21061 = w21058 & w21060;
assign w21062 = ~w21045 & ~w21061;
assign w21063 = ~pi4132 & pi9040;
assign w21064 = pi4039 & ~pi9040;
assign w21065 = ~w21063 & ~w21064;
assign w21066 = pi1163 & ~w21065;
assign w21067 = ~pi1163 & w21065;
assign w21068 = ~w21066 & ~w21067;
assign w21069 = w21045 & w21058;
assign w21070 = w21044 & ~w21051;
assign w21071 = ~w21044 & w21051;
assign w21072 = ~w21070 & ~w21071;
assign w21073 = ~w21045 & w21072;
assign w21074 = ~w21057 & w21073;
assign w21075 = ~w21068 & ~w21069;
assign w21076 = ~w21074 & w21075;
assign w21077 = ~w21062 & w21076;
assign w21078 = w21038 & w21070;
assign w21079 = ~pi4107 & pi9040;
assign w21080 = pi4022 & ~pi9040;
assign w21081 = ~w21079 & ~w21080;
assign w21082 = pi1161 & ~w21081;
assign w21083 = ~pi1161 & w21081;
assign w21084 = ~w21082 & ~w21083;
assign w21085 = ~w21038 & ~w21057;
assign w21086 = w21073 & w21085;
assign w21087 = w21084 & ~w21086;
assign w21088 = ~w21078 & w21087;
assign w21089 = ~w21069 & ~w21084;
assign w21090 = w21038 & w21051;
assign w21091 = ~w21044 & w21090;
assign w21092 = w21089 & ~w21091;
assign w21093 = ~w21088 & ~w21092;
assign w21094 = ~w21051 & ~w21057;
assign w21095 = w21051 & w21057;
assign w21096 = ~w21094 & ~w21095;
assign w21097 = w21038 & ~w21096;
assign w21098 = ~w21093 & ~w21097;
assign w21099 = w21068 & ~w21098;
assign w21100 = w21051 & ~w21068;
assign w21101 = ~w21071 & ~w21100;
assign w21102 = w21085 & ~w21101;
assign w21103 = ~w21038 & ~w21068;
assign w21104 = w21044 & ~w21103;
assign w21105 = ~w21096 & w21104;
assign w21106 = ~w21084 & ~w21102;
assign w21107 = ~w21105 & w21106;
assign w21108 = w21045 & w21094;
assign w21109 = ~w21038 & w21044;
assign w21110 = w21058 & w21109;
assign w21111 = w21038 & w21057;
assign w21112 = ~w21085 & ~w21111;
assign w21113 = w21060 & ~w21095;
assign w21114 = w21100 & w21112;
assign w21115 = ~w21113 & w21114;
assign w21116 = w21084 & ~w21108;
assign w21117 = ~w21110 & w21116;
assign w21118 = ~w21115 & w21117;
assign w21119 = ~w21107 & ~w21118;
assign w21120 = ~w21077 & ~w21119;
assign w21121 = ~w21099 & w21120;
assign w21122 = ~pi3946 & pi9040;
assign w21123 = ~pi4118 & ~pi9040;
assign w21124 = ~w21122 & ~w21123;
assign w21125 = pi1153 & ~w21124;
assign w21126 = ~pi1153 & w21124;
assign w21127 = ~w21125 & ~w21126;
assign w21128 = ~pi3970 & pi9040;
assign w21129 = ~pi3963 & ~pi9040;
assign w21130 = ~w21128 & ~w21129;
assign w21131 = pi1161 & ~w21130;
assign w21132 = ~pi1161 & w21130;
assign w21133 = ~w21131 & ~w21132;
assign w21134 = ~pi4138 & pi9040;
assign w21135 = ~pi4041 & ~pi9040;
assign w21136 = ~w21134 & ~w21135;
assign w21137 = pi1172 & ~w21136;
assign w21138 = ~pi1172 & w21136;
assign w21139 = ~w21137 & ~w21138;
assign w21140 = w21133 & ~w21139;
assign w21141 = ~pi3949 & pi9040;
assign w21142 = ~pi3950 & ~pi9040;
assign w21143 = ~w21141 & ~w21142;
assign w21144 = pi1130 & ~w21143;
assign w21145 = ~pi1130 & w21143;
assign w21146 = ~w21144 & ~w21145;
assign w21147 = ~pi3968 & pi9040;
assign w21148 = ~pi3969 & ~pi9040;
assign w21149 = ~w21147 & ~w21148;
assign w21150 = pi1175 & ~w21149;
assign w21151 = ~pi1175 & w21149;
assign w21152 = ~w21150 & ~w21151;
assign w21153 = w21146 & ~w21152;
assign w21154 = w21140 & w21153;
assign w21155 = w21127 & ~w21154;
assign w21156 = ~w21140 & ~w21153;
assign w21157 = ~w21146 & w21152;
assign w21158 = ~w21139 & ~w21157;
assign w21159 = w21139 & ~w21152;
assign w21160 = ~w21133 & w21146;
assign w21161 = w21159 & ~w21160;
assign w21162 = ~w21158 & ~w21161;
assign w21163 = ~w21156 & w21162;
assign w21164 = ~w21133 & w21157;
assign w21165 = w21157 & w63748;
assign w21166 = ~w21133 & ~w21139;
assign w21167 = ~w21146 & w21166;
assign w21168 = w21166 & w65452;
assign w21169 = ~w21127 & ~w21165;
assign w21170 = ~w21168 & w21169;
assign w21171 = ~w21163 & w21170;
assign w21172 = ~w21155 & ~w21171;
assign w21173 = w21127 & w21139;
assign w21174 = ~w21133 & ~w21152;
assign w21175 = w21173 & w21174;
assign w21176 = ~w21127 & ~w21154;
assign w21177 = w21140 & ~w21176;
assign w21178 = w21127 & w21146;
assign w21179 = w21133 & w21146;
assign w21180 = w21139 & w21179;
assign w21181 = ~w21178 & ~w21180;
assign w21182 = w21152 & ~w21181;
assign w21183 = ~w21146 & w21159;
assign w21184 = w21133 & w21183;
assign w21185 = ~w21164 & ~w21184;
assign w21186 = ~w21127 & ~w21185;
assign w21187 = ~pi4039 & pi9040;
assign w21188 = pi4130 & ~pi9040;
assign w21189 = ~w21187 & ~w21188;
assign w21190 = pi1177 & ~w21189;
assign w21191 = ~pi1177 & w21189;
assign w21192 = ~w21190 & ~w21191;
assign w21193 = ~w21175 & w21192;
assign w21194 = ~w21177 & w21193;
assign w21195 = ~w21182 & w21194;
assign w21196 = ~w21186 & w21195;
assign w21197 = w21139 & w21160;
assign w21198 = w21160 & w65453;
assign w21199 = w21166 & w65454;
assign w21200 = ~w21198 & ~w21199;
assign w21201 = w21133 & ~w21146;
assign w21202 = w21139 & w21201;
assign w21203 = w21127 & w21202;
assign w21204 = ~w21156 & w21176;
assign w21205 = ~w21192 & ~w21203;
assign w21206 = w21200 & w21205;
assign w21207 = ~w21204 & w21206;
assign w21208 = ~w21196 & ~w21207;
assign w21209 = ~w21172 & ~w21208;
assign w21210 = ~w20983 & w63749;
assign w21211 = w20976 & w20996;
assign w21212 = ~w20976 & w21010;
assign w21213 = w21017 & w21212;
assign w21214 = ~w21211 & ~w21213;
assign w21215 = w21210 & ~w21214;
assign w21216 = w21002 & w21017;
assign w21217 = w20944 & ~w20950;
assign w21218 = ~w20994 & w21014;
assign w21219 = ~w21217 & ~w21218;
assign w21220 = ~w21019 & ~w21216;
assign w21221 = ~w21215 & w21220;
assign w21222 = ~w21219 & w21221;
assign w21223 = w20969 & ~w20976;
assign w21224 = ~w20944 & ~w21223;
assign w21225 = ~w21022 & w21224;
assign w21226 = w20969 & w20991;
assign w21227 = w20950 & ~w20986;
assign w21228 = ~w21225 & w21227;
assign w21229 = ~w21226 & w21228;
assign w21230 = ~w21024 & w21229;
assign w21231 = ~w21222 & ~w21230;
assign w21232 = w21005 & ~w21012;
assign w21233 = (~w20962 & w21210) | (~w20962 & w65455) | (w21210 & w65455);
assign w21234 = ~w20979 & w20985;
assign w21235 = ~w21002 & w21234;
assign w21236 = ~w21233 & ~w21235;
assign w21237 = ~w21232 & ~w21236;
assign w21238 = ~w20950 & ~w20987;
assign w21239 = ~w20944 & ~w20992;
assign w21240 = w20980 & ~w21017;
assign w21241 = w21239 & w21240;
assign w21242 = w21224 & w21236;
assign w21243 = w20996 & ~w21242;
assign w21244 = ~w20996 & ~w21024;
assign w21245 = w21021 & w21244;
assign w21246 = w20950 & ~w21245;
assign w21247 = ~w21243 & w21246;
assign w21248 = ~w21003 & ~w21238;
assign w21249 = ~w21241 & w21248;
assign w21250 = ~w21237 & w21249;
assign w21251 = (~pi1227 & w21247) | (~pi1227 & w65456) | (w21247 & w65456);
assign w21252 = ~w21247 & w65457;
assign w21253 = ~w21251 & ~w21252;
assign w21254 = w21214 & ~w21226;
assign w21255 = w20950 & ~w21254;
assign w21256 = ~w21017 & w21217;
assign w21257 = ~w21226 & w21256;
assign w21258 = w21017 & w21239;
assign w21259 = ~w21257 & ~w21258;
assign w21260 = ~w21026 & w21259;
assign w21261 = ~w20986 & w21005;
assign w21262 = ~w21260 & ~w21261;
assign w21263 = ~w21255 & ~w21262;
assign w21264 = ~pi3969 & pi9040;
assign w21265 = ~pi4107 & ~pi9040;
assign w21266 = ~w21264 & ~w21265;
assign w21267 = pi1166 & ~w21266;
assign w21268 = ~pi1166 & w21266;
assign w21269 = ~w21267 & ~w21268;
assign w21270 = ~pi3966 & pi9040;
assign w21271 = ~pi3948 & ~pi9040;
assign w21272 = ~w21270 & ~w21271;
assign w21273 = pi1169 & ~w21272;
assign w21274 = ~pi1169 & w21272;
assign w21275 = ~w21273 & ~w21274;
assign w21276 = ~pi4117 & pi9040;
assign w21277 = ~pi3970 & ~pi9040;
assign w21278 = ~w21276 & ~w21277;
assign w21279 = pi1181 & ~w21278;
assign w21280 = ~pi1181 & w21278;
assign w21281 = ~w21279 & ~w21280;
assign w21282 = ~w21275 & ~w21281;
assign w21283 = ~pi4130 & pi9040;
assign w21284 = ~pi4023 & ~pi9040;
assign w21285 = ~w21283 & ~w21284;
assign w21286 = pi1155 & ~w21285;
assign w21287 = ~pi1155 & w21285;
assign w21288 = ~w21286 & ~w21287;
assign w21289 = ~pi4131 & pi9040;
assign w21290 = ~pi4266 & ~pi9040;
assign w21291 = ~w21289 & ~w21290;
assign w21292 = pi1151 & ~w21291;
assign w21293 = ~pi1151 & w21291;
assign w21294 = ~w21292 & ~w21293;
assign w21295 = ~w21288 & w21294;
assign w21296 = ~pi4041 & pi9040;
assign w21297 = ~pi3957 & ~pi9040;
assign w21298 = ~w21296 & ~w21297;
assign w21299 = pi1154 & ~w21298;
assign w21300 = ~pi1154 & w21298;
assign w21301 = ~w21299 & ~w21300;
assign w21302 = w21288 & w21301;
assign w21303 = ~w21295 & ~w21302;
assign w21304 = w21282 & ~w21303;
assign w21305 = w21275 & ~w21294;
assign w21306 = ~w21275 & w21294;
assign w21307 = ~w21305 & ~w21306;
assign w21308 = w21288 & w21307;
assign w21309 = (~w21281 & ~w21307) | (~w21281 & w65458) | (~w21307 & w65458);
assign w21310 = w21275 & ~w21288;
assign w21311 = w21301 & w21310;
assign w21312 = w21309 & ~w21311;
assign w21313 = w21275 & w21281;
assign w21314 = w21288 & w21294;
assign w21315 = ~w21310 & ~w21314;
assign w21316 = ~w21301 & ~w21315;
assign w21317 = (w21281 & w21315) | (w21281 & w63750) | (w21315 & w63750);
assign w21318 = w21302 & w21305;
assign w21319 = w21317 & ~w21318;
assign w21320 = (~w21313 & ~w21317) | (~w21313 & w65459) | (~w21317 & w65459);
assign w21321 = w21301 & w21315;
assign w21322 = w21275 & w21294;
assign w21323 = ~w21288 & ~w21301;
assign w21324 = w21322 & w21323;
assign w21325 = ~w21321 & ~w21324;
assign w21326 = ~w21320 & w21325;
assign w21327 = ~w21304 & ~w21312;
assign w21328 = ~w21326 & w21327;
assign w21329 = w21269 & ~w21328;
assign w21330 = ~w21302 & w21313;
assign w21331 = ~w21323 & w21330;
assign w21332 = ~w21301 & w21305;
assign w21333 = ~w21323 & ~w21332;
assign w21334 = w21275 & ~w21301;
assign w21335 = w21288 & w21334;
assign w21336 = ~w21294 & w21335;
assign w21337 = ~w21320 & ~w21336;
assign w21338 = ~w21333 & ~w21337;
assign w21339 = w21302 & w21306;
assign w21340 = w21281 & ~w21301;
assign w21341 = ~w21294 & w21340;
assign w21342 = w21340 & w21353;
assign w21343 = ~w21339 & ~w21342;
assign w21344 = ~w21269 & ~w21304;
assign w21345 = ~w21331 & w21344;
assign w21346 = w21343 & w21345;
assign w21347 = ~w21338 & w21346;
assign w21348 = ~w21329 & ~w21347;
assign w21349 = ~w21288 & w21307;
assign w21350 = ~w21335 & ~w21349;
assign w21351 = w21341 & ~w21350;
assign w21352 = ~w21281 & w21350;
assign w21353 = w21288 & ~w21294;
assign w21354 = w21275 & w21353;
assign w21355 = w21352 & ~w21354;
assign w21356 = w21306 & w21323;
assign w21357 = w21321 & w21349;
assign w21358 = ~w21295 & ~w21353;
assign w21359 = w21317 & w21358;
assign w21360 = ~w21275 & ~w21301;
assign w21361 = ~w21311 & ~w21360;
assign w21362 = ~w21294 & ~w21361;
assign w21363 = w21309 & ~w21362;
assign w21364 = ~w21310 & ~w21318;
assign w21365 = w21363 & ~w21364;
assign w21366 = w21343 & ~w21356;
assign w21367 = ~w21357 & w21366;
assign w21368 = ~w21359 & w21367;
assign w21369 = ~w21365 & w21368;
assign w21370 = ~w21322 & w21369;
assign w21371 = w21355 & ~w21370;
assign w21372 = ~w21348 & ~w21351;
assign w21373 = ~w21371 & w21372;
assign w21374 = ~w21127 & w21167;
assign w21375 = w21174 & w21178;
assign w21376 = ~w21165 & ~w21375;
assign w21377 = w21127 & w21376;
assign w21378 = w21133 & w21153;
assign w21379 = ~w21127 & ~w21378;
assign w21380 = ~w21202 & w21379;
assign w21381 = ~w21377 & ~w21380;
assign w21382 = w21192 & ~w21197;
assign w21383 = ~w21168 & w21382;
assign w21384 = ~w21184 & w21383;
assign w21385 = ~w21381 & w21384;
assign w21386 = w21157 & w21166;
assign w21387 = ~w21139 & w21157;
assign w21388 = ~w21140 & w21146;
assign w21389 = ~w21174 & w21388;
assign w21390 = ~w21387 & ~w21389;
assign w21391 = ~w21127 & ~w21390;
assign w21392 = w21140 & ~w21152;
assign w21393 = w21201 & w65453;
assign w21394 = ~w21392 & ~w21393;
assign w21395 = w21127 & ~w21394;
assign w21396 = w21161 & ~w21201;
assign w21397 = ~w21192 & ~w21386;
assign w21398 = ~w21396 & w21397;
assign w21399 = ~w21391 & w21398;
assign w21400 = ~w21395 & w21399;
assign w21401 = ~w21385 & ~w21400;
assign w21402 = ~w21127 & ~w21146;
assign w21403 = ~w21178 & ~w21192;
assign w21404 = w21140 & w21152;
assign w21405 = ~w21402 & w21404;
assign w21406 = ~w21403 & w21405;
assign w21407 = ~w21374 & ~w21406;
assign w21408 = ~w21401 & w21407;
assign w21409 = w21200 & ~w21387;
assign w21410 = w21171 & ~w21409;
assign w21411 = ~w21139 & w21153;
assign w21412 = ~w21179 & ~w21411;
assign w21413 = (~w21127 & ~w21412) | (~w21127 & w65460) | (~w21412 & w65460);
assign w21414 = ~w21146 & w21392;
assign w21415 = ~w21413 & ~w21414;
assign w21416 = w21192 & ~w21415;
assign w21417 = w21160 & w21159;
assign w21418 = ~w21393 & ~w21417;
assign w21419 = w21412 & w65461;
assign w21420 = ~w21184 & ~w21192;
assign w21421 = w21201 & ~w21420;
assign w21422 = w21418 & ~w21419;
assign w21423 = ~w21421 & w21422;
assign w21424 = w21127 & ~w21423;
assign w21425 = ~w21139 & w21179;
assign w21426 = w21174 & w21402;
assign w21427 = w21157 & w21173;
assign w21428 = ~w21425 & ~w21426;
assign w21429 = ~w21427 & w21428;
assign w21430 = (~w21192 & ~w21429) | (~w21192 & w65462) | (~w21429 & w65462);
assign w21431 = ~w21410 & ~w21430;
assign w21432 = ~w21416 & w21431;
assign w21433 = (~pi1232 & ~w21432) | (~pi1232 & w65463) | (~w21432 & w65463);
assign w21434 = w21432 & w65464;
assign w21435 = ~w21433 & ~w21434;
assign w21436 = ~pi3945 & pi9040;
assign w21437 = ~pi4025 & ~pi9040;
assign w21438 = ~w21436 & ~w21437;
assign w21439 = pi1159 & ~w21438;
assign w21440 = ~pi1159 & w21438;
assign w21441 = ~w21439 & ~w21440;
assign w21442 = ~pi3956 & pi9040;
assign w21443 = ~pi4024 & ~pi9040;
assign w21444 = ~w21442 & ~w21443;
assign w21445 = pi1180 & ~w21444;
assign w21446 = ~pi1180 & w21444;
assign w21447 = ~w21445 & ~w21446;
assign w21448 = w21441 & w21447;
assign w21449 = ~pi4277 & pi9040;
assign w21450 = ~pi3952 & ~pi9040;
assign w21451 = ~w21449 & ~w21450;
assign w21452 = pi1173 & ~w21451;
assign w21453 = ~pi1173 & w21451;
assign w21454 = ~w21452 & ~w21453;
assign w21455 = w21448 & w21454;
assign w21456 = ~w21441 & ~w21454;
assign w21457 = ~pi4040 & pi9040;
assign w21458 = ~pi4021 & ~pi9040;
assign w21459 = ~w21457 & ~w21458;
assign w21460 = pi1174 & ~w21459;
assign w21461 = ~pi1174 & w21459;
assign w21462 = ~w21460 & ~w21461;
assign w21463 = ~w21447 & w21462;
assign w21464 = w21456 & w21463;
assign w21465 = ~w21455 & ~w21464;
assign w21466 = ~pi3964 & pi9040;
assign w21467 = ~pi4133 & ~pi9040;
assign w21468 = ~w21466 & ~w21467;
assign w21469 = pi1176 & ~w21468;
assign w21470 = ~pi1176 & w21468;
assign w21471 = ~w21469 & ~w21470;
assign w21472 = ~w21465 & w21471;
assign w21473 = ~w21454 & ~w21462;
assign w21474 = w21448 & w21473;
assign w21475 = ~w21441 & ~w21447;
assign w21476 = w21454 & ~w21462;
assign w21477 = w21475 & w21476;
assign w21478 = ~w21474 & ~w21477;
assign w21479 = ~w21448 & ~w21475;
assign w21480 = w21462 & ~w21471;
assign w21481 = w21454 & ~w21471;
assign w21482 = w21447 & w21481;
assign w21483 = ~w21480 & ~w21482;
assign w21484 = w21479 & ~w21483;
assign w21485 = ~pi3962 & pi9040;
assign w21486 = ~pi3932 & ~pi9040;
assign w21487 = ~w21485 & ~w21486;
assign w21488 = pi1171 & ~w21487;
assign w21489 = ~pi1171 & w21487;
assign w21490 = ~w21488 & ~w21489;
assign w21491 = w21478 & w21490;
assign w21492 = ~w21472 & w21491;
assign w21493 = ~w21484 & w21492;
assign w21494 = w21447 & w21471;
assign w21495 = ~w21441 & ~w21462;
assign w21496 = w21494 & w21495;
assign w21497 = w21441 & ~w21471;
assign w21498 = ~w21447 & w21497;
assign w21499 = w21454 & w21498;
assign w21500 = ~w21447 & w21456;
assign w21501 = ~w21471 & w21500;
assign w21502 = w21456 & w21494;
assign w21503 = ~w21501 & ~w21502;
assign w21504 = w21447 & w21454;
assign w21505 = w21441 & w21471;
assign w21506 = ~w21454 & ~w21505;
assign w21507 = w21462 & ~w21506;
assign w21508 = ~w21504 & w21507;
assign w21509 = w21503 & ~w21508;
assign w21510 = ~w21455 & ~w21500;
assign w21511 = ~w21462 & ~w21510;
assign w21512 = ~w21490 & ~w21496;
assign w21513 = ~w21499 & w21512;
assign w21514 = ~w21511 & w21513;
assign w21515 = w21509 & w21514;
assign w21516 = ~w21493 & ~w21515;
assign w21517 = ~w21441 & w21482;
assign w21518 = w21462 & w21517;
assign w21519 = w21447 & w21456;
assign w21520 = ~w21479 & w65465;
assign w21521 = ~w21447 & ~w21462;
assign w21522 = ~w21454 & ~w21497;
assign w21523 = w21521 & ~w21522;
assign w21524 = ~w21520 & ~w21523;
assign w21525 = w21473 & ~w21519;
assign w21526 = w21524 & w21525;
assign w21527 = ~w21518 & ~w21526;
assign w21528 = ~w21516 & w21527;
assign w21529 = ~w21281 & ~w21356;
assign w21530 = ~w21337 & ~w21529;
assign w21531 = ~w21282 & w21361;
assign w21532 = w21295 & ~w21531;
assign w21533 = ~w21281 & ~w21334;
assign w21534 = w21288 & ~w21313;
assign w21535 = ~w21533 & w21534;
assign w21536 = w21269 & ~w21332;
assign w21537 = ~w21535 & w21536;
assign w21538 = ~w21357 & w21537;
assign w21539 = ~w21532 & w21538;
assign w21540 = w21352 & ~w21532;
assign w21541 = w21301 & w21322;
assign w21542 = ~w21349 & ~w21541;
assign w21543 = ~w21309 & ~w21542;
assign w21544 = ~w21269 & ~w21543;
assign w21545 = ~w21540 & w21544;
assign w21546 = ~w21539 & ~w21545;
assign w21547 = ~w21530 & ~w21546;
assign w21548 = ~pi4029 & pi9040;
assign w21549 = ~pi3933 & ~pi9040;
assign w21550 = ~w21548 & ~w21549;
assign w21551 = pi1178 & ~w21550;
assign w21552 = ~pi1178 & w21550;
assign w21553 = ~w21551 & ~w21552;
assign w21554 = ~pi4133 & pi9040;
assign w21555 = ~pi3937 & ~pi9040;
assign w21556 = ~w21554 & ~w21555;
assign w21557 = pi1131 & ~w21556;
assign w21558 = ~pi1131 & w21556;
assign w21559 = ~w21557 & ~w21558;
assign w21560 = ~w21553 & ~w21559;
assign w21561 = ~pi3952 & pi9040;
assign w21562 = ~pi4126 & ~pi9040;
assign w21563 = ~w21561 & ~w21562;
assign w21564 = pi1146 & ~w21563;
assign w21565 = ~pi1146 & w21563;
assign w21566 = ~w21564 & ~w21565;
assign w21567 = ~pi3953 & pi9040;
assign w21568 = ~pi3945 & ~pi9040;
assign w21569 = ~w21567 & ~w21568;
assign w21570 = pi1164 & ~w21569;
assign w21571 = ~pi1164 & w21569;
assign w21572 = ~w21570 & ~w21571;
assign w21573 = ~w21566 & w21572;
assign w21574 = w21560 & w21573;
assign w21575 = ~w21553 & w21559;
assign w21576 = w21566 & w21572;
assign w21577 = w21575 & w21576;
assign w21578 = w21553 & ~w21559;
assign w21579 = w21573 & w21578;
assign w21580 = ~w21577 & ~w21579;
assign w21581 = ~w21574 & w21580;
assign w21582 = ~pi3971 & pi9040;
assign w21583 = ~pi3956 & ~pi9040;
assign w21584 = ~w21582 & ~w21583;
assign w21585 = pi1165 & ~w21584;
assign w21586 = ~pi1165 & w21584;
assign w21587 = ~w21585 & ~w21586;
assign w21588 = ~w21581 & ~w21587;
assign w21589 = ~w21578 & ~w21587;
assign w21590 = w21566 & ~w21572;
assign w21591 = ~w21589 & w21590;
assign w21592 = ~pi4021 & pi9040;
assign w21593 = ~pi4192 & ~pi9040;
assign w21594 = ~w21592 & ~w21593;
assign w21595 = pi1158 & ~w21594;
assign w21596 = ~pi1158 & w21594;
assign w21597 = ~w21595 & ~w21596;
assign w21598 = w21572 & ~w21587;
assign w21599 = w21553 & ~w21566;
assign w21600 = w21566 & ~w21578;
assign w21601 = ~w21599 & ~w21600;
assign w21602 = w21598 & w21601;
assign w21603 = ~w21566 & ~w21578;
assign w21604 = ~w21559 & w21572;
assign w21605 = w21589 & ~w21604;
assign w21606 = w21578 & ~w21587;
assign w21607 = ~w21566 & w21606;
assign w21608 = ~w21605 & ~w21607;
assign w21609 = ~w21603 & ~w21608;
assign w21610 = ~w21575 & ~w21578;
assign w21611 = ~w21573 & ~w21610;
assign w21612 = ~w21566 & ~w21575;
assign w21613 = w21587 & ~w21612;
assign w21614 = ~w21611 & w21613;
assign w21615 = ~w21605 & ~w21614;
assign w21616 = ~w21602 & ~w21609;
assign w21617 = ~w21615 & w21616;
assign w21618 = ~w21579 & w21597;
assign w21619 = ~w21591 & w21618;
assign w21620 = ~w21617 & w21619;
assign w21621 = w21603 & w21615;
assign w21622 = w21576 & ~w21610;
assign w21623 = ~w21597 & ~w21622;
assign w21624 = ~w21609 & w21623;
assign w21625 = ~w21621 & w21624;
assign w21626 = ~w21620 & ~w21625;
assign w21627 = ~w21588 & ~w21626;
assign w21628 = ~w21281 & ~w21301;
assign w21629 = w21322 & w21628;
assign w21630 = w21269 & ~w21369;
assign w21631 = ~w21319 & ~w21363;
assign w21632 = w21294 & w21321;
assign w21633 = ~w21631 & ~w21632;
assign w21634 = ~w21269 & ~w21633;
assign w21635 = w21353 & w21360;
assign w21636 = ~w21629 & ~w21635;
assign w21637 = ~w21634 & w21636;
assign w21638 = ~w21630 & w21637;
assign w21639 = w21061 & ~w21103;
assign w21640 = ~w21072 & ~w21111;
assign w21641 = ~w21057 & w21071;
assign w21642 = ~w21109 & ~w21641;
assign w21643 = w21640 & w21642;
assign w21644 = ~w21090 & ~w21108;
assign w21645 = ~w21068 & ~w21644;
assign w21646 = ~w21639 & ~w21643;
assign w21647 = ~w21645 & w21646;
assign w21648 = w21087 & w21647;
assign w21649 = ~w21073 & ~w21085;
assign w21650 = ~w21085 & ~w21090;
assign w21651 = w21072 & ~w21650;
assign w21652 = ~w21649 & ~w21651;
assign w21653 = ~w21068 & ~w21652;
assign w21654 = ~w21058 & w21653;
assign w21655 = ~w21113 & ~w21654;
assign w21656 = ~w21068 & w21109;
assign w21657 = ~w21074 & ~w21656;
assign w21658 = ~w21051 & ~w21657;
assign w21659 = ~w21084 & ~w21658;
assign w21660 = ~w21655 & w21659;
assign w21661 = ~w21648 & ~w21660;
assign w21662 = w21590 & w21610;
assign w21663 = w21580 & ~w21662;
assign w21664 = ~w21566 & w21575;
assign w21665 = w21663 & ~w21664;
assign w21666 = w21587 & ~w21599;
assign w21667 = w21665 & w21666;
assign w21668 = ~w21587 & ~w21665;
assign w21669 = ~w21572 & ~w21606;
assign w21670 = w21599 & w21669;
assign w21671 = ~w21597 & ~w21670;
assign w21672 = ~w21667 & w21671;
assign w21673 = ~w21668 & w21672;
assign w21674 = ~w21572 & w21664;
assign w21675 = w21559 & ~w21663;
assign w21676 = w21560 & ~w21572;
assign w21677 = w21572 & w21599;
assign w21678 = w21587 & ~w21677;
assign w21679 = ~w21676 & w21678;
assign w21680 = w21608 & ~w21679;
assign w21681 = w21559 & w21599;
assign w21682 = w21572 & ~w21681;
assign w21683 = ~w21669 & ~w21682;
assign w21684 = w21597 & ~w21674;
assign w21685 = ~w21683 & w21684;
assign w21686 = ~w21675 & w21685;
assign w21687 = ~w21680 & w21686;
assign w21688 = ~w21673 & ~w21687;
assign w21689 = ~w21051 & ~w21112;
assign w21690 = w21071 & ~w21085;
assign w21691 = w21068 & ~w21078;
assign w21692 = ~w21690 & w21691;
assign w21693 = ~w21689 & w21692;
assign w21694 = ~w21076 & ~w21693;
assign w21695 = w21084 & ~w21694;
assign w21696 = w21068 & w21089;
assign w21697 = ~w21074 & w21696;
assign w21698 = ~w21695 & ~w21697;
assign w21699 = w21057 & ~w21651;
assign w21700 = w21062 & w21699;
assign w21701 = ~w21698 & ~w21700;
assign w21702 = w21044 & w21057;
assign w21703 = ~w21113 & ~w21702;
assign w21704 = w21090 & ~w21703;
assign w21705 = ~w21061 & ~w21704;
assign w21706 = ~w21068 & w21089;
assign w21707 = ~w21640 & w21706;
assign w21708 = w21705 & w21707;
assign w21709 = ~w21701 & ~w21708;
assign w21710 = ~w21068 & w21110;
assign w21711 = w21071 & w21111;
assign w21712 = w21653 & w21703;
assign w21713 = w21068 & w21652;
assign w21714 = ~w21711 & ~w21713;
assign w21715 = ~w21712 & w21714;
assign w21716 = w21084 & ~w21715;
assign w21717 = w21100 & ~w21642;
assign w21718 = w21705 & ~w21717;
assign w21719 = ~w21084 & ~w21718;
assign w21720 = w21038 & ~w21071;
assign w21721 = w21096 & w21720;
assign w21722 = ~w21060 & ~w21084;
assign w21723 = ~w21641 & w21722;
assign w21724 = ~w21721 & ~w21723;
assign w21725 = w21068 & ~w21724;
assign w21726 = ~w21710 & ~w21725;
assign w21727 = ~w21719 & w21726;
assign w21728 = ~w21716 & w21727;
assign w21729 = w21155 & ~w21163;
assign w21730 = ~w21127 & ~w21183;
assign w21731 = ~w21729 & ~w21730;
assign w21732 = ~w21127 & ~w21411;
assign w21733 = ~w21162 & w21732;
assign w21734 = w21133 & w21152;
assign w21735 = w21173 & w21734;
assign w21736 = w21192 & ~w21735;
assign w21737 = w21376 & w21736;
assign w21738 = ~w21733 & w21737;
assign w21739 = w21379 & ~w21412;
assign w21740 = ~w21174 & w21178;
assign w21741 = ~w21734 & w21740;
assign w21742 = w21420 & ~w21741;
assign w21743 = ~w21739 & w21742;
assign w21744 = w21409 & w21743;
assign w21745 = ~w21738 & ~w21744;
assign w21746 = ~w21731 & ~w21745;
assign w21747 = ~pi4193 & pi9040;
assign w21748 = ~pi4132 & ~pi9040;
assign w21749 = ~w21747 & ~w21748;
assign w21750 = pi1169 & ~w21749;
assign w21751 = ~pi1169 & w21749;
assign w21752 = ~w21750 & ~w21751;
assign w21753 = ~pi4023 & pi9040;
assign w21754 = ~pi3968 & ~pi9040;
assign w21755 = ~w21753 & ~w21754;
assign w21756 = pi1183 & ~w21755;
assign w21757 = ~pi1183 & w21755;
assign w21758 = ~w21756 & ~w21757;
assign w21759 = ~w21752 & w21758;
assign w21760 = w21752 & ~w21758;
assign w21761 = ~pi3948 & pi9040;
assign w21762 = ~pi3949 & ~pi9040;
assign w21763 = ~w21761 & ~w21762;
assign w21764 = pi1171 & ~w21763;
assign w21765 = ~pi1171 & w21763;
assign w21766 = ~w21764 & ~w21765;
assign w21767 = w21760 & ~w21766;
assign w21768 = ~w21759 & ~w21767;
assign w21769 = ~pi3957 & pi9040;
assign w21770 = ~pi4043 & ~pi9040;
assign w21771 = ~w21769 & ~w21770;
assign w21772 = pi1173 & ~w21771;
assign w21773 = ~pi1173 & w21771;
assign w21774 = ~w21772 & ~w21773;
assign w21775 = w21766 & w21774;
assign w21776 = ~w21766 & ~w21774;
assign w21777 = ~w21775 & ~w21776;
assign w21778 = ~pi4118 & pi9040;
assign w21779 = ~pi3965 & ~pi9040;
assign w21780 = ~w21778 & ~w21779;
assign w21781 = pi1157 & ~w21780;
assign w21782 = ~pi1157 & w21780;
assign w21783 = ~w21781 & ~w21782;
assign w21784 = ~w21777 & w21783;
assign w21785 = ~w21768 & w21784;
assign w21786 = w21759 & w21766;
assign w21787 = ~w21760 & ~w21786;
assign w21788 = w21774 & ~w21787;
assign w21789 = ~w21752 & ~w21774;
assign w21790 = ~w21758 & w21766;
assign w21791 = w21789 & ~w21790;
assign w21792 = ~w21759 & ~w21776;
assign w21793 = ~w21789 & w21792;
assign w21794 = ~w21791 & ~w21793;
assign w21795 = (w21777 & w21793) | (w21777 & w65466) | (w21793 & w65466);
assign w21796 = ~w21752 & w21766;
assign w21797 = w21774 & w21796;
assign w21798 = w21783 & ~w21797;
assign w21799 = ~w21795 & w21798;
assign w21800 = ~w21775 & ~w21783;
assign w21801 = ~w21758 & w21774;
assign w21802 = w21752 & w21766;
assign w21803 = ~w21801 & ~w21802;
assign w21804 = w21800 & ~w21803;
assign w21805 = ~w21788 & ~w21804;
assign w21806 = ~w21799 & w21805;
assign w21807 = ~pi3963 & pi9040;
assign w21808 = ~pi4131 & ~pi9040;
assign w21809 = ~w21807 & ~w21808;
assign w21810 = pi1155 & ~w21809;
assign w21811 = ~pi1155 & w21809;
assign w21812 = ~w21810 & ~w21811;
assign w21813 = ~w21806 & w21812;
assign w21814 = w21758 & ~w21774;
assign w21815 = ~w21766 & w21814;
assign w21816 = w21800 & ~w21815;
assign w21817 = w21814 & w21816;
assign w21818 = w21760 & w21775;
assign w21819 = ~w21817 & ~w21818;
assign w21820 = w21774 & w21783;
assign w21821 = ~w21816 & ~w21820;
assign w21822 = ~w21812 & ~w21821;
assign w21823 = w21806 & w21822;
assign w21824 = ~w21785 & w21819;
assign w21825 = ~w21813 & w21824;
assign w21826 = ~w21823 & w21825;
assign w21827 = w21559 & w21590;
assign w21828 = ~w21574 & ~w21827;
assign w21829 = w21587 & ~w21828;
assign w21830 = ~w21598 & ~w21607;
assign w21831 = ~w21597 & ~w21601;
assign w21832 = w21682 & ~w21831;
assign w21833 = ~w21830 & ~w21832;
assign w21834 = w21553 & w21572;
assign w21835 = ~w21674 & ~w21834;
assign w21836 = w21678 & ~w21835;
assign w21837 = w21578 & w21836;
assign w21838 = ~w21575 & ~w21599;
assign w21839 = ~w21610 & ~w21838;
assign w21840 = ~w21682 & w21839;
assign w21841 = ~w21597 & ~w21683;
assign w21842 = ~w21840 & w21841;
assign w21843 = ~w21837 & w21842;
assign w21844 = ~w21566 & ~w21587;
assign w21845 = w21560 & w21844;
assign w21846 = w21559 & w21587;
assign w21847 = ~w21573 & w21846;
assign w21848 = w21597 & ~w21845;
assign w21849 = ~w21847 & w21848;
assign w21850 = ~w21662 & w21849;
assign w21851 = ~w21602 & w21850;
assign w21852 = ~w21843 & ~w21851;
assign w21853 = ~w21829 & ~w21833;
assign w21854 = ~w21852 & w21853;
assign w21855 = ~w21447 & ~w21507;
assign w21856 = w21497 & ~w21855;
assign w21857 = w21441 & ~w21481;
assign w21858 = w21521 & w21857;
assign w21859 = w21481 & w21495;
assign w21860 = ~w21464 & ~w21859;
assign w21861 = ~w21858 & w21860;
assign w21862 = w21503 & w21861;
assign w21863 = ~w21856 & w21862;
assign w21864 = ~w21490 & ~w21863;
assign w21865 = ~w21479 & w63751;
assign w21866 = ~w21499 & ~w21519;
assign w21867 = ~w21462 & ~w21866;
assign w21868 = ~w21498 & ~w21517;
assign w21869 = ~w21505 & w21868;
assign w21870 = w21441 & w21454;
assign w21871 = w21462 & ~w21870;
assign w21872 = ~w21869 & w21871;
assign w21873 = ~w21865 & ~w21867;
assign w21874 = ~w21872 & w21873;
assign w21875 = w21490 & ~w21874;
assign w21876 = ~w21501 & ~w21865;
assign w21877 = w21462 & ~w21876;
assign w21878 = ~w21471 & w21474;
assign w21879 = ~w21496 & ~w21878;
assign w21880 = ~w21877 & w21879;
assign w21881 = ~w21864 & w21880;
assign w21882 = ~w21875 & w21881;
assign w21883 = w21281 & ~w21308;
assign w21884 = w21301 & ~w21883;
assign w21885 = ~w21355 & w21884;
assign w21886 = ~w21288 & w21341;
assign w21887 = w21314 & w21340;
assign w21888 = ~w21295 & ~w21887;
assign w21889 = w21316 & w21888;
assign w21890 = w21281 & ~w21333;
assign w21891 = w21269 & ~w21541;
assign w21892 = ~w21889 & w21891;
assign w21893 = ~w21890 & w21892;
assign w21894 = ~w21324 & ~w21339;
assign w21895 = ~w21354 & w21894;
assign w21896 = w21529 & w21895;
assign w21897 = ~w21294 & w21310;
assign w21898 = w21281 & ~w21897;
assign w21899 = ~w21632 & w21898;
assign w21900 = ~w21896 & ~w21899;
assign w21901 = ~w21269 & ~w21635;
assign w21902 = ~w21887 & w21901;
assign w21903 = ~w21900 & w21902;
assign w21904 = ~w21893 & ~w21903;
assign w21905 = ~w21885 & ~w21886;
assign w21906 = ~w21904 & w21905;
assign w21907 = ~w21774 & w21802;
assign w21908 = w21789 & w63752;
assign w21909 = ~w21907 & ~w21908;
assign w21910 = ~w21760 & ~w21909;
assign w21911 = ~w21758 & w21797;
assign w21912 = (~w21783 & w21910) | (~w21783 & w65467) | (w21910 & w65467);
assign w21913 = ~w21790 & ~w21803;
assign w21914 = (w21783 & w21913) | (w21783 & w63753) | (w21913 & w63753);
assign w21915 = ~w21760 & ~w21775;
assign w21916 = ~w21803 & w21915;
assign w21917 = ~w21914 & ~w21916;
assign w21918 = ~w21914 & w65468;
assign w21919 = ~w21912 & ~w21918;
assign w21920 = w21819 & ~w21919;
assign w21921 = w21796 & w21814;
assign w21922 = w21812 & ~w21921;
assign w21923 = ~w21920 & w21922;
assign w21924 = ~w21812 & w21917;
assign w21925 = ~w21923 & ~w21924;
assign w21926 = w21759 & w21776;
assign w21927 = ~w21752 & ~w21775;
assign w21928 = w21812 & ~w21927;
assign w21929 = ~w21913 & w21928;
assign w21930 = ~w21911 & ~w21926;
assign w21931 = ~w21929 & w21930;
assign w21932 = w21783 & ~w21931;
assign w21933 = ~w21794 & ~w21818;
assign w21934 = ~w21760 & ~w21796;
assign w21935 = w21794 & w21934;
assign w21936 = w21812 & ~w21935;
assign w21937 = ~w21783 & ~w21933;
assign w21938 = ~w21936 & w21937;
assign w21939 = ~w21932 & ~w21938;
assign w21940 = ~w21925 & w21939;
assign w21941 = ~pi3959 & pi9040;
assign w21942 = ~pi4210 & ~pi9040;
assign w21943 = ~w21941 & ~w21942;
assign w21944 = pi1158 & ~w21943;
assign w21945 = ~pi1158 & w21943;
assign w21946 = ~w21944 & ~w21945;
assign w21947 = ~pi4119 & pi9040;
assign w21948 = ~pi3962 & ~pi9040;
assign w21949 = ~w21947 & ~w21948;
assign w21950 = pi1168 & ~w21949;
assign w21951 = ~pi1168 & w21949;
assign w21952 = ~w21950 & ~w21951;
assign w21953 = w21946 & w21952;
assign w21954 = ~w21946 & ~w21952;
assign w21955 = ~pi4024 & pi9040;
assign w21956 = ~pi3938 & ~pi9040;
assign w21957 = ~w21955 & ~w21956;
assign w21958 = pi1180 & ~w21957;
assign w21959 = ~pi1180 & w21957;
assign w21960 = ~w21958 & ~w21959;
assign w21961 = ~w21954 & ~w21960;
assign w21962 = ~w21953 & w21961;
assign w21963 = w21946 & w21960;
assign w21964 = ~pi3961 & pi9040;
assign w21965 = ~pi4040 & ~pi9040;
assign w21966 = ~w21964 & ~w21965;
assign w21967 = pi1178 & ~w21966;
assign w21968 = ~pi1178 & w21966;
assign w21969 = ~w21967 & ~w21968;
assign w21970 = w21952 & w21969;
assign w21971 = ~w21963 & w21970;
assign w21972 = ~pi4134 & pi9040;
assign w21973 = ~pi3964 & ~pi9040;
assign w21974 = ~w21972 & ~w21973;
assign w21975 = pi1159 & ~w21974;
assign w21976 = ~pi1159 & w21974;
assign w21977 = ~w21975 & ~w21976;
assign w21978 = w21971 & w21977;
assign w21979 = w21962 & w21978;
assign w21980 = ~pi4126 & pi9040;
assign w21981 = ~pi3934 & ~pi9040;
assign w21982 = ~w21980 & ~w21981;
assign w21983 = pi1145 & ~w21982;
assign w21984 = ~pi1145 & w21982;
assign w21985 = ~w21983 & ~w21984;
assign w21986 = w21960 & ~w21969;
assign w21987 = w21952 & w21986;
assign w21988 = w21946 & ~w21969;
assign w21989 = ~w21954 & ~w21988;
assign w21990 = ~w21946 & ~w21960;
assign w21991 = ~w21963 & ~w21990;
assign w21992 = w21989 & w21991;
assign w21993 = ~w21986 & ~w21992;
assign w21994 = w21977 & ~w21993;
assign w21995 = ~w21952 & ~w21969;
assign w21996 = w21990 & w21995;
assign w21997 = ~w21987 & ~w21996;
assign w21998 = ~w21994 & w21997;
assign w21999 = ~w21985 & ~w21998;
assign w22000 = ~w21970 & ~w21995;
assign w22001 = ~w21991 & w22000;
assign w22002 = w21969 & ~w21985;
assign w22003 = ~w21962 & ~w22002;
assign w22004 = ~w21989 & ~w22003;
assign w22005 = ~w21960 & w21969;
assign w22006 = w21953 & w22005;
assign w22007 = ~w22001 & ~w22006;
assign w22008 = ~w22004 & w22007;
assign w22009 = ~w21946 & w21960;
assign w22010 = w21985 & w22009;
assign w22011 = ~w22000 & w22010;
assign w22012 = w22008 & ~w22011;
assign w22013 = ~w21977 & ~w22012;
assign w22014 = w21977 & w21985;
assign w22015 = ~w21990 & w22014;
assign w22016 = w21993 & w22015;
assign w22017 = ~w21979 & ~w22016;
assign w22018 = ~w21999 & w22017;
assign w22019 = ~w22013 & w22018;
assign w22020 = ~w21796 & w21814;
assign w22021 = ~w21767 & w21798;
assign w22022 = ~w21783 & ~w21907;
assign w22023 = ~w21934 & w22022;
assign w22024 = ~w22021 & ~w22023;
assign w22025 = ~w21812 & ~w22020;
assign w22026 = ~w22024 & w22025;
assign w22027 = w21752 & w21816;
assign w22028 = w21774 & w22027;
assign w22029 = w21752 & ~w21790;
assign w22030 = ~w21789 & ~w22029;
assign w22031 = w21798 & w22030;
assign w22032 = ~w21818 & w21922;
assign w22033 = ~w22031 & w22032;
assign w22034 = ~w22028 & w22033;
assign w22035 = ~w22026 & ~w22034;
assign w22036 = w21768 & w21783;
assign w22037 = w21794 & w22036;
assign w22038 = ~w21912 & ~w22037;
assign w22039 = ~w22035 & w22038;
assign w22040 = w21476 & ~w21868;
assign w22041 = ~w21463 & ~w21877;
assign w22042 = ~w21454 & w21471;
assign w22043 = (w21462 & w21479) | (w21462 & w65469) | (w21479 & w65469);
assign w22044 = ~w21462 & ~w21502;
assign w22045 = ~w21865 & w22044;
assign w22046 = ~w22043 & ~w22045;
assign w22047 = ~w22045 & w65470;
assign w22048 = w21463 & ~w21481;
assign w22049 = ~w21870 & w22048;
assign w22050 = ~w21474 & ~w22049;
assign w22051 = w21868 & w22050;
assign w22052 = ~w22047 & w22051;
assign w22053 = ~w22041 & w22052;
assign w22054 = w21447 & ~w21456;
assign w22055 = ~w21870 & w22054;
assign w22056 = w21478 & ~w22055;
assign w22057 = w21471 & ~w22056;
assign w22058 = w21456 & ~w21463;
assign w22059 = ~w21494 & w22058;
assign w22060 = ~w22057 & ~w22059;
assign w22061 = ~w22053 & w22060;
assign w22062 = w21490 & ~w22061;
assign w22063 = ~w21490 & ~w22052;
assign w22064 = w21480 & ~w22055;
assign w22065 = w21509 & w22064;
assign w22066 = ~w22040 & ~w22065;
assign w22067 = ~w22063 & w22066;
assign w22068 = ~w22062 & w22067;
assign w22069 = ~w21989 & w21991;
assign w22070 = ~w21991 & ~w21995;
assign w22071 = ~w22069 & ~w22070;
assign w22072 = ~w21962 & ~w22009;
assign w22073 = w21977 & ~w21985;
assign w22074 = ~w22071 & w22073;
assign w22075 = ~w22072 & w22074;
assign w22076 = ~w21969 & w22071;
assign w22077 = w21985 & ~w22005;
assign w22078 = w21946 & ~w21952;
assign w22079 = w21969 & w21991;
assign w22080 = ~w22078 & ~w22079;
assign w22081 = w22077 & ~w22080;
assign w22082 = ~w21953 & ~w22005;
assign w22083 = ~w21971 & ~w21985;
assign w22084 = ~w22082 & w22083;
assign w22085 = ~w22076 & ~w22084;
assign w22086 = ~w22081 & w22085;
assign w22087 = (~w21977 & ~w22085) | (~w21977 & w65471) | (~w22085 & w65471);
assign w22088 = w22014 & ~w22078;
assign w22089 = ~w22082 & w22088;
assign w22090 = w21963 & ~w21969;
assign w22091 = ~w21985 & ~w22090;
assign w22092 = w21952 & ~w22077;
assign w22093 = ~w22091 & w22092;
assign w22094 = ~w21978 & ~w22089;
assign w22095 = ~w22093 & w22094;
assign w22096 = ~w22075 & w22095;
assign w22097 = ~w22087 & w22096;
assign w22098 = pi1221 & w22097;
assign w22099 = ~pi1221 & ~w22097;
assign w22100 = ~w22098 & ~w22099;
assign w22101 = ~w22079 & ~w22090;
assign w22102 = ~w21961 & w21985;
assign w22103 = w22101 & w22102;
assign w22104 = w21970 & w22103;
assign w22105 = ~w21960 & w21988;
assign w22106 = w21995 & ~w22009;
assign w22107 = w21952 & ~w21988;
assign w22108 = ~w21990 & w22107;
assign w22109 = ~w21985 & ~w22106;
assign w22110 = ~w22108 & w22109;
assign w22111 = ~w22105 & ~w22110;
assign w22112 = ~w22078 & ~w22111;
assign w22113 = w21985 & ~w22070;
assign w22114 = ~w22069 & w22113;
assign w22115 = ~w22112 & ~w22114;
assign w22116 = ~w21977 & ~w22115;
assign w22117 = w22004 & w22086;
assign w22118 = w21990 & ~w22002;
assign w22119 = ~w21952 & ~w22118;
assign w22120 = w22101 & w22119;
assign w22121 = w22113 & ~w22120;
assign w22122 = w21977 & ~w22110;
assign w22123 = ~w22121 & w22122;
assign w22124 = ~w22104 & ~w22123;
assign w22125 = ~w22116 & w22124;
assign w22126 = ~w22117 & w22125;
assign w22127 = w21985 & w21988;
assign w22128 = ~w22008 & w22091;
assign w22129 = ~w22127 & ~w22128;
assign w22130 = w21952 & ~w22129;
assign w22131 = ~w21985 & ~w22101;
assign w22132 = ~w21977 & ~w21996;
assign w22133 = ~w22103 & w22132;
assign w22134 = ~w22131 & w22133;
assign w22135 = w21962 & w21985;
assign w22136 = w21970 & w22009;
assign w22137 = w21977 & ~w22136;
assign w22138 = ~w22135 & w22137;
assign w22139 = ~w22120 & w22138;
assign w22140 = ~w22134 & ~w22139;
assign w22141 = ~w22130 & ~w22140;
assign w22142 = w21566 & w21597;
assign w22143 = ~w21575 & w22142;
assign w22144 = ~w21834 & w22143;
assign w22145 = ~w21681 & ~w22144;
assign w22146 = ~w21587 & ~w22145;
assign w22147 = w21838 & w21846;
assign w22148 = ~w21560 & w21566;
assign w22149 = w21559 & ~w21598;
assign w22150 = ~w21604 & ~w22148;
assign w22151 = ~w22149 & w22150;
assign w22152 = w21623 & ~w22147;
assign w22153 = ~w22151 & w22152;
assign w22154 = w21587 & w21839;
assign w22155 = ~w21574 & w21597;
assign w22156 = ~w22154 & w22155;
assign w22157 = ~w22153 & ~w22156;
assign w22158 = ~w21836 & ~w22146;
assign w22159 = ~w22157 & w22158;
assign w22160 = pi1213 & w22159;
assign w22161 = ~pi1213 & ~w22159;
assign w22162 = ~w22160 & ~w22161;
assign w22163 = ~w21526 & ~w21867;
assign w22164 = w22052 & ~w22163;
assign w22165 = w21441 & ~w21482;
assign w22166 = ~w21521 & ~w22042;
assign w22167 = w22165 & w22166;
assign w22168 = ~w21517 & ~w22167;
assign w22169 = ~w22164 & w22168;
assign w22170 = ~w21490 & ~w22169;
assign w22171 = w22043 & ~w22165;
assign w22172 = w21509 & w22171;
assign w22173 = w21524 & ~w22172;
assign w22174 = w21490 & ~w22173;
assign w22175 = ~w22046 & ~w22174;
assign w22176 = ~w22170 & w22175;
assign w22177 = ~w21817 & ~w21820;
assign w22178 = ~w21768 & ~w22177;
assign w22179 = w21783 & ~w21909;
assign w22180 = ~w21783 & w21790;
assign w22181 = ~w22179 & ~w22180;
assign w22182 = w21936 & w22181;
assign w22183 = w21766 & ~w21799;
assign w22184 = ~w21803 & ~w22183;
assign w22185 = w21759 & ~w21777;
assign w22186 = ~w21812 & ~w22185;
assign w22187 = ~w22027 & w22186;
assign w22188 = ~w22037 & w22187;
assign w22189 = ~w22184 & w22188;
assign w22190 = ~w22182 & ~w22189;
assign w22191 = ~w22178 & ~w22190;
assign w22192 = ~pi4100 & pi9040;
assign w22193 = ~pi4075 & ~pi9040;
assign w22194 = ~w22192 & ~w22193;
assign w22195 = pi1245 & ~w22194;
assign w22196 = ~pi1245 & w22194;
assign w22197 = ~w22195 & ~w22196;
assign w22198 = ~pi4307 & pi9040;
assign w22199 = ~pi4212 & ~pi9040;
assign w22200 = ~w22198 & ~w22199;
assign w22201 = pi1222 & ~w22200;
assign w22202 = ~pi1222 & w22200;
assign w22203 = ~w22201 & ~w22202;
assign w22204 = w22197 & ~w22203;
assign w22205 = ~pi4125 & pi9040;
assign w22206 = ~pi4307 & ~pi9040;
assign w22207 = ~w22205 & ~w22206;
assign w22208 = pi1239 & ~w22207;
assign w22209 = ~pi1239 & w22207;
assign w22210 = ~w22208 & ~w22209;
assign w22211 = ~pi4110 & pi9040;
assign w22212 = ~pi4125 & ~pi9040;
assign w22213 = ~w22211 & ~w22212;
assign w22214 = pi1240 & ~w22213;
assign w22215 = ~pi1240 & w22213;
assign w22216 = ~w22214 & ~w22215;
assign w22217 = w22210 & w22216;
assign w22218 = w22204 & w22217;
assign w22219 = ~w22203 & ~w22210;
assign w22220 = ~pi4209 & pi9040;
assign w22221 = ~pi4069 & ~pi9040;
assign w22222 = ~w22220 & ~w22221;
assign w22223 = pi1206 & ~w22222;
assign w22224 = ~pi1206 & w22222;
assign w22225 = ~w22223 & ~w22224;
assign w22226 = ~w22197 & w22225;
assign w22227 = w22219 & w22226;
assign w22228 = ~pi4069 & pi9040;
assign w22229 = ~pi4203 & ~pi9040;
assign w22230 = ~w22228 & ~w22229;
assign w22231 = pi1236 & ~w22230;
assign w22232 = ~pi1236 & w22230;
assign w22233 = ~w22231 & ~w22232;
assign w22234 = w22203 & w22210;
assign w22235 = ~w22197 & ~w22225;
assign w22236 = w22234 & w22235;
assign w22237 = w22210 & w22225;
assign w22238 = w22197 & ~w22237;
assign w22239 = w22197 & ~w22225;
assign w22240 = w22203 & w22239;
assign w22241 = w22204 & w22225;
assign w22242 = ~w22240 & ~w22241;
assign w22243 = (w22238 & w22242) | (w22238 & w63754) | (w22242 & w63754);
assign w22244 = ~w22216 & ~w22234;
assign w22245 = (w22244 & w22243) | (w22244 & w65472) | (w22243 & w65472);
assign w22246 = ~w22210 & ~w22225;
assign w22247 = ~w22204 & w22246;
assign w22248 = w22197 & w22237;
assign w22249 = ~w22210 & w22226;
assign w22250 = ~w22248 & ~w22249;
assign w22251 = ~w22247 & w22250;
assign w22252 = ~w22219 & ~w22234;
assign w22253 = w22235 & w22252;
assign w22254 = (w22216 & ~w22252) | (w22216 & w65473) | (~w22252 & w65473);
assign w22255 = ~w22233 & ~w22236;
assign w22256 = (w22255 & w22251) | (w22255 & w65474) | (w22251 & w65474);
assign w22257 = ~w22245 & w22256;
assign w22258 = w22225 & w22234;
assign w22259 = ~w22247 & ~w22258;
assign w22260 = ~w22216 & ~w22259;
assign w22261 = w22216 & w22243;
assign w22262 = ~w22210 & w22225;
assign w22263 = ~w22203 & ~w22216;
assign w22264 = w22262 & w22263;
assign w22265 = w22226 & w22234;
assign w22266 = ~w22264 & ~w22265;
assign w22267 = ~w22253 & w22266;
assign w22268 = (w22233 & w22259) | (w22233 & w65475) | (w22259 & w65475);
assign w22269 = w22267 & w22268;
assign w22270 = ~w22261 & w22269;
assign w22271 = ~w22257 & ~w22270;
assign w22272 = ~w22218 & ~w22227;
assign w22273 = ~w22271 & w22272;
assign w22274 = pi1254 & w22273;
assign w22275 = ~pi1254 & ~w22273;
assign w22276 = ~w22274 & ~w22275;
assign w22277 = ~pi4279 & pi9040;
assign w22278 = ~pi4299 & ~pi9040;
assign w22279 = ~w22277 & ~w22278;
assign w22280 = pi1209 & ~w22279;
assign w22281 = ~pi1209 & w22279;
assign w22282 = ~w22280 & ~w22281;
assign w22283 = ~pi4111 & pi9040;
assign w22284 = ~pi4110 & ~pi9040;
assign w22285 = ~w22283 & ~w22284;
assign w22286 = pi1210 & ~w22285;
assign w22287 = ~pi1210 & w22285;
assign w22288 = ~w22286 & ~w22287;
assign w22289 = ~w22282 & ~w22288;
assign w22290 = ~pi4383 & pi9040;
assign w22291 = ~pi4088 & ~pi9040;
assign w22292 = ~w22290 & ~w22291;
assign w22293 = pi1237 & ~w22292;
assign w22294 = ~pi1237 & w22292;
assign w22295 = ~w22293 & ~w22294;
assign w22296 = ~pi4136 & pi9040;
assign w22297 = ~pi4184 & ~pi9040;
assign w22298 = ~w22296 & ~w22297;
assign w22299 = pi1226 & ~w22298;
assign w22300 = ~pi1226 & w22298;
assign w22301 = ~w22299 & ~w22300;
assign w22302 = w22295 & w22301;
assign w22303 = ~w22295 & ~w22301;
assign w22304 = ~w22302 & ~w22303;
assign w22305 = w22289 & ~w22304;
assign w22306 = ~w22282 & w22288;
assign w22307 = w22295 & w22306;
assign w22308 = ~w22288 & ~w22295;
assign w22309 = w22301 & w22308;
assign w22310 = ~w22307 & ~w22309;
assign w22311 = w22282 & w22301;
assign w22312 = ~w22282 & ~w22301;
assign w22313 = w22288 & ~w22312;
assign w22314 = ~w22282 & w22308;
assign w22315 = ~w22313 & ~w22314;
assign w22316 = ~w22311 & ~w22315;
assign w22317 = ~w22310 & ~w22316;
assign w22318 = (~w22305 & w22316) | (~w22305 & w65476) | (w22316 & w65476);
assign w22319 = ~pi4203 & pi9040;
assign w22320 = ~pi4123 & ~pi9040;
assign w22321 = ~w22319 & ~w22320;
assign w22322 = pi1214 & ~w22321;
assign w22323 = ~pi1214 & w22321;
assign w22324 = ~w22322 & ~w22323;
assign w22325 = ~w22318 & w22324;
assign w22326 = ~pi4216 & pi9040;
assign w22327 = ~pi4136 & ~pi9040;
assign w22328 = ~w22326 & ~w22327;
assign w22329 = pi1246 & ~w22328;
assign w22330 = ~pi1246 & w22328;
assign w22331 = ~w22329 & ~w22330;
assign w22332 = w22282 & ~w22324;
assign w22333 = ~w22288 & w22295;
assign w22334 = w22332 & w22333;
assign w22335 = w22331 & ~w22334;
assign w22336 = w22302 & w22306;
assign w22337 = ~w22324 & ~w22336;
assign w22338 = ~w22314 & w22337;
assign w22339 = w22282 & ~w22295;
assign w22340 = w22288 & ~w22301;
assign w22341 = ~w22339 & ~w22340;
assign w22342 = w22339 & w22340;
assign w22343 = ~w22341 & ~w22342;
assign w22344 = ~w22307 & w22324;
assign w22345 = ~w22343 & w22344;
assign w22346 = ~w22338 & ~w22345;
assign w22347 = w22335 & ~w22346;
assign w22348 = (w22324 & w22304) | (w22324 & w65477) | (w22304 & w65477);
assign w22349 = w22288 & w22311;
assign w22350 = ~w22339 & ~w22349;
assign w22351 = ~w22348 & ~w22350;
assign w22352 = w22288 & w22301;
assign w22353 = ~w22324 & ~w22352;
assign w22354 = w22295 & w22312;
assign w22355 = w22353 & ~w22354;
assign w22356 = w22289 & w22301;
assign w22357 = w22282 & ~w22288;
assign w22358 = w22295 & ~w22301;
assign w22359 = w22357 & w22358;
assign w22360 = w22324 & ~w22356;
assign w22361 = ~w22359 & w22360;
assign w22362 = ~w22355 & ~w22361;
assign w22363 = ~w22331 & ~w22351;
assign w22364 = ~w22362 & w22363;
assign w22365 = ~w22347 & ~w22364;
assign w22366 = ~w22324 & w22342;
assign w22367 = ~w22325 & ~w22366;
assign w22368 = ~w22365 & w22367;
assign w22369 = ~pi1248 & w22368;
assign w22370 = pi1248 & ~w22368;
assign w22371 = ~w22369 & ~w22370;
assign w22372 = ~w22203 & w22260;
assign w22373 = w22204 & w22246;
assign w22374 = ~w22258 & ~w22373;
assign w22375 = w22216 & ~w22374;
assign w22376 = ~w22203 & ~w22225;
assign w22377 = (w22216 & ~w22235) | (w22216 & w63755) | (~w22235 & w63755);
assign w22378 = ~w22376 & w22377;
assign w22379 = ~w22216 & w22242;
assign w22380 = ~w22378 & ~w22379;
assign w22381 = ~w22203 & w22235;
assign w22382 = ~w22219 & ~w22258;
assign w22383 = ~w22381 & w22382;
assign w22384 = (~w22216 & ~w22383) | (~w22216 & w63756) | (~w22383 & w63756);
assign w22385 = w22216 & ~w22248;
assign w22386 = ~w22227 & ~w22240;
assign w22387 = w22385 & w22386;
assign w22388 = ~w22384 & ~w22387;
assign w22389 = (w22233 & ~w22380) | (w22233 & w63757) | (~w22380 & w63757);
assign w22390 = ~w22388 & w22389;
assign w22391 = w22203 & w22216;
assign w22392 = w22226 & w22391;
assign w22393 = ~w22241 & ~w22392;
assign w22394 = ~w22210 & ~w22393;
assign w22395 = ~w22233 & w22266;
assign w22396 = ~w22394 & w22395;
assign w22397 = ~w22380 & w22396;
assign w22398 = ~w22372 & ~w22375;
assign w22399 = (w22398 & w22390) | (w22398 & w65478) | (w22390 & w65478);
assign w22400 = pi1261 & w22399;
assign w22401 = ~pi1261 & ~w22399;
assign w22402 = ~w22400 & ~w22401;
assign w22403 = ~w22203 & w22225;
assign w22404 = ~w22219 & w22250;
assign w22405 = ~w22403 & ~w22404;
assign w22406 = ~w22210 & w22239;
assign w22407 = ~w22236 & ~w22406;
assign w22408 = ~w22233 & ~w22407;
assign w22409 = ~w22405 & ~w22408;
assign w22410 = ~w22216 & ~w22409;
assign w22411 = w22197 & w22262;
assign w22412 = ~w22239 & ~w22246;
assign w22413 = ~w22406 & ~w22412;
assign w22414 = ~w22411 & ~w22413;
assign w22415 = w22391 & ~w22414;
assign w22416 = ~w22226 & ~w22237;
assign w22417 = w22263 & w22416;
assign w22418 = w22197 & w22234;
assign w22419 = w22217 & w22403;
assign w22420 = ~w22373 & ~w22418;
assign w22421 = ~w22419 & w22420;
assign w22422 = (w22233 & ~w22421) | (w22233 & w65479) | (~w22421 & w65479);
assign w22423 = ~w22203 & ~w22217;
assign w22424 = ~w22416 & w22423;
assign w22425 = ~w22265 & ~w22411;
assign w22426 = w22216 & ~w22425;
assign w22427 = w22217 & w22376;
assign w22428 = ~w22424 & ~w22427;
assign w22429 = ~w22426 & w22428;
assign w22430 = ~w22233 & ~w22429;
assign w22431 = ~w22415 & ~w22422;
assign w22432 = ~w22430 & w22431;
assign w22433 = ~w22410 & w22432;
assign w22434 = pi1263 & ~w22433;
assign w22435 = ~pi1263 & w22433;
assign w22436 = ~w22434 & ~w22435;
assign w22437 = ~pi4298 & pi9040;
assign w22438 = ~pi4104 & ~pi9040;
assign w22439 = ~w22437 & ~w22438;
assign w22440 = pi1231 & ~w22439;
assign w22441 = ~pi1231 & w22439;
assign w22442 = ~w22440 & ~w22441;
assign w22443 = ~pi4207 & pi9040;
assign w22444 = ~pi4135 & ~pi9040;
assign w22445 = ~w22443 & ~w22444;
assign w22446 = pi1225 & ~w22445;
assign w22447 = ~pi1225 & w22445;
assign w22448 = ~w22446 & ~w22447;
assign w22449 = w22442 & ~w22448;
assign w22450 = ~pi4038 & pi9040;
assign w22451 = ~pi4100 & ~pi9040;
assign w22452 = ~w22450 & ~w22451;
assign w22453 = pi1220 & ~w22452;
assign w22454 = ~pi1220 & w22452;
assign w22455 = ~w22453 & ~w22454;
assign w22456 = w22449 & ~w22455;
assign w22457 = ~w22442 & w22448;
assign w22458 = ~pi4135 & pi9040;
assign w22459 = ~pi4209 & ~pi9040;
assign w22460 = ~w22458 & ~w22459;
assign w22461 = pi1245 & ~w22460;
assign w22462 = ~pi1245 & w22460;
assign w22463 = ~w22461 & ~w22462;
assign w22464 = w22457 & w22463;
assign w22465 = ~w22456 & ~w22464;
assign w22466 = ~pi4127 & pi9040;
assign w22467 = ~pi4114 & ~pi9040;
assign w22468 = ~w22466 & ~w22467;
assign w22469 = pi1235 & ~w22468;
assign w22470 = ~pi1235 & w22468;
assign w22471 = ~w22469 & ~w22470;
assign w22472 = ~w22465 & w22471;
assign w22473 = ~w22442 & ~w22471;
assign w22474 = w22448 & w22473;
assign w22475 = (w22455 & ~w22473) | (w22455 & w65480) | (~w22473 & w65480);
assign w22476 = w22455 & w22463;
assign w22477 = w22473 & w22476;
assign w22478 = w22442 & w22448;
assign w22479 = ~w22463 & w22471;
assign w22480 = w22478 & w22479;
assign w22481 = ~w22448 & ~w22463;
assign w22482 = w22442 & ~w22471;
assign w22483 = w22481 & w22482;
assign w22484 = ~w22480 & ~w22483;
assign w22485 = ~w22477 & w22484;
assign w22486 = w22475 & ~w22485;
assign w22487 = ~pi4098 & pi9040;
assign w22488 = ~pi4383 & ~pi9040;
assign w22489 = ~w22487 & ~w22488;
assign w22490 = pi1206 & ~w22489;
assign w22491 = ~pi1206 & w22489;
assign w22492 = ~w22490 & ~w22491;
assign w22493 = w22448 & ~w22455;
assign w22494 = w22457 & ~w22463;
assign w22495 = ~w22455 & w22473;
assign w22496 = ~w22494 & ~w22495;
assign w22497 = ~w22493 & ~w22496;
assign w22498 = ~w22478 & ~w22479;
assign w22499 = w22448 & w22471;
assign w22500 = w22463 & ~w22471;
assign w22501 = w22455 & ~w22500;
assign w22502 = ~w22498 & ~w22499;
assign w22503 = ~w22501 & w22502;
assign w22504 = ~w22497 & ~w22503;
assign w22505 = ~w22492 & ~w22504;
assign w22506 = w22463 & w22471;
assign w22507 = ~w22455 & ~w22506;
assign w22508 = ~w22493 & ~w22507;
assign w22509 = ~w22474 & ~w22508;
assign w22510 = ~w22442 & w22471;
assign w22511 = w22481 & w22510;
assign w22512 = (w22455 & ~w22499) | (w22455 & w63758) | (~w22499 & w63758);
assign w22513 = ~w22511 & w22512;
assign w22514 = w22448 & w22463;
assign w22515 = ~w22457 & ~w22471;
assign w22516 = ~w22514 & w22515;
assign w22517 = w22513 & ~w22516;
assign w22518 = ~w22509 & ~w22517;
assign w22519 = ~w22464 & ~w22480;
assign w22520 = ~w22518 & w22519;
assign w22521 = w22492 & ~w22520;
assign w22522 = ~w22472 & ~w22486;
assign w22523 = ~w22505 & w22522;
assign w22524 = ~w22521 & w22523;
assign w22525 = pi1256 & w22524;
assign w22526 = ~pi1256 & ~w22524;
assign w22527 = ~w22525 & ~w22526;
assign w22528 = ~pi4300 & pi9040;
assign w22529 = ~pi4099 & ~pi9040;
assign w22530 = ~w22528 & ~w22529;
assign w22531 = pi1229 & ~w22530;
assign w22532 = ~pi1229 & w22530;
assign w22533 = ~w22531 & ~w22532;
assign w22534 = ~pi4169 & pi9040;
assign w22535 = ~pi4124 & ~pi9040;
assign w22536 = ~w22534 & ~w22535;
assign w22537 = pi1217 & ~w22536;
assign w22538 = ~pi1217 & w22536;
assign w22539 = ~w22537 & ~w22538;
assign w22540 = ~pi4124 & pi9040;
assign w22541 = ~pi4106 & ~pi9040;
assign w22542 = ~w22540 & ~w22541;
assign w22543 = pi1246 & ~w22542;
assign w22544 = ~pi1246 & w22542;
assign w22545 = ~w22543 & ~w22544;
assign w22546 = ~pi4301 & pi9040;
assign w22547 = ~pi4105 & ~pi9040;
assign w22548 = ~w22546 & ~w22547;
assign w22549 = pi1216 & ~w22548;
assign w22550 = ~pi1216 & w22548;
assign w22551 = ~w22549 & ~w22550;
assign w22552 = ~w22545 & ~w22551;
assign w22553 = w22545 & w22551;
assign w22554 = ~w22552 & ~w22553;
assign w22555 = ~pi4121 & pi9040;
assign w22556 = ~pi4295 & ~pi9040;
assign w22557 = ~w22555 & ~w22556;
assign w22558 = pi1247 & ~w22557;
assign w22559 = ~pi1247 & w22557;
assign w22560 = ~w22558 & ~w22559;
assign w22561 = w22545 & w22560;
assign w22562 = ~pi4106 & pi9040;
assign w22563 = ~pi4122 & ~pi9040;
assign w22564 = ~w22562 & ~w22563;
assign w22565 = pi1226 & ~w22564;
assign w22566 = ~pi1226 & w22564;
assign w22567 = ~w22565 & ~w22566;
assign w22568 = w22551 & ~w22567;
assign w22569 = ~w22551 & w22567;
assign w22570 = ~w22568 & ~w22569;
assign w22571 = ~w22561 & w22570;
assign w22572 = ~w22539 & ~w22554;
assign w22573 = ~w22571 & w22572;
assign w22574 = w22554 & w22567;
assign w22575 = ~w22553 & ~w22560;
assign w22576 = ~w22539 & w22545;
assign w22577 = w22567 & w22576;
assign w22578 = ~w22575 & ~w22577;
assign w22579 = w22574 & w22578;
assign w22580 = w22539 & w22579;
assign w22581 = ~w22560 & ~w22576;
assign w22582 = w22539 & w22552;
assign w22583 = ~w22568 & ~w22582;
assign w22584 = w22539 & w22567;
assign w22585 = w22581 & ~w22584;
assign w22586 = w22583 & w22585;
assign w22587 = ~w22573 & ~w22586;
assign w22588 = ~w22580 & w22587;
assign w22589 = ~w22533 & ~w22588;
assign w22590 = w22539 & w22551;
assign w22591 = ~w22545 & w22560;
assign w22592 = ~w22590 & w22591;
assign w22593 = ~w22539 & ~w22567;
assign w22594 = ~w22551 & w22593;
assign w22595 = ~w22592 & ~w22594;
assign w22596 = w22554 & ~w22595;
assign w22597 = w22560 & ~w22583;
assign w22598 = ~w22596 & ~w22597;
assign w22599 = w22533 & ~w22598;
assign w22600 = ~w22560 & w22567;
assign w22601 = w22545 & w22600;
assign w22602 = ~w22539 & ~w22551;
assign w22603 = ~w22545 & ~w22567;
assign w22604 = ~w22602 & w22603;
assign w22605 = ~w22601 & ~w22604;
assign w22606 = ~w22533 & w22560;
assign w22607 = ~w22533 & ~w22590;
assign w22608 = ~w22606 & ~w22607;
assign w22609 = ~w22605 & w22608;
assign w22610 = ~w22554 & ~w22567;
assign w22611 = ~w22554 & w65481;
assign w22612 = w22591 & w22611;
assign w22613 = w22561 & w22593;
assign w22614 = w22600 & w22602;
assign w22615 = ~w22613 & ~w22614;
assign w22616 = ~w22609 & w22615;
assign w22617 = ~w22612 & w22616;
assign w22618 = ~w22599 & w22617;
assign w22619 = ~w22589 & w22618;
assign w22620 = pi1253 & w22619;
assign w22621 = ~pi1253 & ~w22619;
assign w22622 = ~w22620 & ~w22621;
assign w22623 = ~pi4114 & pi9040;
assign w22624 = ~pi4098 & ~pi9040;
assign w22625 = ~w22623 & ~w22624;
assign w22626 = pi1236 & ~w22625;
assign w22627 = ~pi1236 & w22625;
assign w22628 = ~w22626 & ~w22627;
assign w22629 = ~pi4299 & pi9040;
assign w22630 = ~pi4207 & ~pi9040;
assign w22631 = ~w22629 & ~w22630;
assign w22632 = pi1239 & ~w22631;
assign w22633 = ~pi1239 & w22631;
assign w22634 = ~w22632 & ~w22633;
assign w22635 = ~w22628 & ~w22634;
assign w22636 = ~pi4123 & pi9040;
assign w22637 = ~pi4111 & ~pi9040;
assign w22638 = ~w22636 & ~w22637;
assign w22639 = pi1200 & ~w22638;
assign w22640 = ~pi1200 & w22638;
assign w22641 = ~w22639 & ~w22640;
assign w22642 = ~pi4088 & pi9040;
assign w22643 = ~pi4375 & ~pi9040;
assign w22644 = ~w22642 & ~w22643;
assign w22645 = pi1210 & ~w22644;
assign w22646 = ~pi1210 & w22644;
assign w22647 = ~w22645 & ~w22646;
assign w22648 = w22641 & w22647;
assign w22649 = ~w22641 & ~w22647;
assign w22650 = ~w22648 & ~w22649;
assign w22651 = w22635 & ~w22650;
assign w22652 = ~w22628 & ~w22647;
assign w22653 = w22628 & w22647;
assign w22654 = ~w22652 & ~w22653;
assign w22655 = w22634 & w22654;
assign w22656 = ~w22634 & w22653;
assign w22657 = ~pi4375 & pi9040;
assign w22658 = ~pi4298 & ~pi9040;
assign w22659 = ~w22657 & ~w22658;
assign w22660 = pi1241 & ~w22659;
assign w22661 = ~pi1241 & w22659;
assign w22662 = ~w22660 & ~w22661;
assign w22663 = (~w22662 & w22655) | (~w22662 & w65482) | (w22655 & w65482);
assign w22664 = ~w22634 & ~w22647;
assign w22665 = w22634 & w22647;
assign w22666 = ~w22664 & ~w22665;
assign w22667 = ~w22634 & ~w22641;
assign w22668 = w22666 & ~w22667;
assign w22669 = w22663 & ~w22668;
assign w22670 = ~w22651 & ~w22669;
assign w22671 = ~pi4104 & pi9040;
assign w22672 = ~pi4038 & ~pi9040;
assign w22673 = ~w22671 & ~w22672;
assign w22674 = pi1209 & ~w22673;
assign w22675 = ~pi1209 & w22673;
assign w22676 = ~w22674 & ~w22675;
assign w22677 = ~w22670 & w22676;
assign w22678 = w22628 & ~w22641;
assign w22679 = ~w22634 & w22662;
assign w22680 = ~w22664 & ~w22679;
assign w22681 = w22678 & ~w22680;
assign w22682 = ~w22628 & w22641;
assign w22683 = w22664 & w22682;
assign w22684 = w22628 & w22634;
assign w22685 = ~w22647 & w22684;
assign w22686 = ~w22683 & ~w22685;
assign w22687 = ~w22662 & ~w22686;
assign w22688 = (~w22676 & w22687) | (~w22676 & w65483) | (w22687 & w65483);
assign w22689 = w22666 & w22682;
assign w22690 = w22665 & w22678;
assign w22691 = w22628 & w22641;
assign w22692 = ~w22634 & w22691;
assign w22693 = ~w22690 & ~w22692;
assign w22694 = w22676 & ~w22693;
assign w22695 = w22664 & ~w22682;
assign w22696 = ~w22689 & ~w22695;
assign w22697 = ~w22694 & w22696;
assign w22698 = w22662 & ~w22697;
assign w22699 = ~w22678 & ~w22682;
assign w22700 = w22634 & ~w22662;
assign w22701 = w22647 & ~w22676;
assign w22702 = ~w22700 & ~w22701;
assign w22703 = ~w22679 & w22699;
assign w22704 = ~w22702 & w22703;
assign w22705 = ~w22688 & ~w22704;
assign w22706 = ~w22698 & w22705;
assign w22707 = ~w22677 & w22706;
assign w22708 = ~pi1250 & w22707;
assign w22709 = pi1250 & ~w22707;
assign w22710 = ~w22708 & ~w22709;
assign w22711 = ~pi4120 & pi9040;
assign w22712 = ~pi4101 & ~pi9040;
assign w22713 = ~w22711 & ~w22712;
assign w22714 = pi1224 & ~w22713;
assign w22715 = ~pi1224 & w22713;
assign w22716 = ~w22714 & ~w22715;
assign w22717 = ~pi4122 & pi9040;
assign w22718 = ~pi4317 & ~pi9040;
assign w22719 = ~w22717 & ~w22718;
assign w22720 = pi1244 & ~w22719;
assign w22721 = ~pi1244 & w22719;
assign w22722 = ~w22720 & ~w22721;
assign w22723 = ~w22716 & w22722;
assign w22724 = w22716 & ~w22722;
assign w22725 = ~w22723 & ~w22724;
assign w22726 = ~pi4129 & pi9040;
assign w22727 = ~pi4036 & ~pi9040;
assign w22728 = ~w22726 & ~w22727;
assign w22729 = pi1219 & ~w22728;
assign w22730 = ~pi1219 & w22728;
assign w22731 = ~w22729 & ~w22730;
assign w22732 = ~w22725 & w22731;
assign w22733 = ~pi4045 & pi9040;
assign w22734 = ~pi4301 & ~pi9040;
assign w22735 = ~w22733 & ~w22734;
assign w22736 = pi1225 & ~w22735;
assign w22737 = ~pi1225 & w22735;
assign w22738 = ~w22736 & ~w22737;
assign w22739 = w22716 & w22738;
assign w22740 = ~w22716 & ~w22738;
assign w22741 = ~pi4295 & pi9040;
assign w22742 = ~pi4045 & ~pi9040;
assign w22743 = ~w22741 & ~w22742;
assign w22744 = pi1238 & ~w22743;
assign w22745 = ~pi1238 & w22743;
assign w22746 = ~w22744 & ~w22745;
assign w22747 = ~w22740 & ~w22746;
assign w22748 = ~w22740 & w65484;
assign w22749 = ~w22739 & w22748;
assign w22750 = ~w22738 & w22746;
assign w22751 = ~w22740 & ~w22750;
assign w22752 = w22716 & ~w22731;
assign w22753 = w22746 & ~w22752;
assign w22754 = w22722 & ~w22751;
assign w22755 = ~w22753 & w22754;
assign w22756 = ~w22749 & ~w22755;
assign w22757 = ~w22732 & ~w22756;
assign w22758 = ~w22716 & ~w22746;
assign w22759 = ~w22716 & w22731;
assign w22760 = ~w22752 & ~w22759;
assign w22761 = w22738 & w22746;
assign w22762 = w22760 & w22761;
assign w22763 = ~w22758 & ~w22762;
assign w22764 = ~w22722 & ~w22731;
assign w22765 = w22738 & ~w22764;
assign w22766 = ~w22763 & w22765;
assign w22767 = ~w22722 & ~w22746;
assign w22768 = ~w22760 & w22767;
assign w22769 = w22722 & w22731;
assign w22770 = w22716 & ~w22738;
assign w22771 = w22769 & w22770;
assign w22772 = w22740 & w22764;
assign w22773 = w22746 & w22772;
assign w22774 = ~pi4252 & pi9040;
assign w22775 = ~pi4120 & ~pi9040;
assign w22776 = ~w22774 & ~w22775;
assign w22777 = pi1235 & ~w22776;
assign w22778 = ~pi1235 & w22776;
assign w22779 = ~w22777 & ~w22778;
assign w22780 = ~w22771 & w22779;
assign w22781 = ~w22768 & w22780;
assign w22782 = ~w22773 & w22781;
assign w22783 = ~w22766 & w22782;
assign w22784 = w22731 & w22746;
assign w22785 = w22723 & w22784;
assign w22786 = ~w22731 & ~w22738;
assign w22787 = w22723 & w22786;
assign w22788 = w22739 & w22769;
assign w22789 = w22740 & w22784;
assign w22790 = ~w22779 & ~w22789;
assign w22791 = w22724 & w22750;
assign w22792 = ~w22731 & ~w22770;
assign w22793 = ~w22716 & w22738;
assign w22794 = ~w22746 & ~w22793;
assign w22795 = w22792 & w22794;
assign w22796 = w22738 & w22764;
assign w22797 = ~w22785 & ~w22787;
assign w22798 = ~w22788 & ~w22791;
assign w22799 = ~w22796 & w22798;
assign w22800 = w22790 & w22797;
assign w22801 = ~w22795 & w22800;
assign w22802 = w22799 & w22801;
assign w22803 = ~w22783 & ~w22802;
assign w22804 = ~w22757 & ~w22803;
assign w22805 = ~pi1251 & w22804;
assign w22806 = pi1251 & ~w22804;
assign w22807 = ~w22805 & ~w22806;
assign w22808 = w22250 & w22424;
assign w22809 = ~w22241 & w22377;
assign w22810 = ~w22216 & ~w22226;
assign w22811 = ~w22809 & ~w22810;
assign w22812 = w22238 & ~w22252;
assign w22813 = ~w22253 & ~w22812;
assign w22814 = ~w22811 & w22813;
assign w22815 = w22233 & ~w22814;
assign w22816 = ~w22413 & w22809;
assign w22817 = ~w22413 & ~w22418;
assign w22818 = ~w22385 & ~w22817;
assign w22819 = ~w22816 & ~w22818;
assign w22820 = ~w22233 & ~w22819;
assign w22821 = (~w22808 & ~w22380) | (~w22808 & w65485) | (~w22380 & w65485);
assign w22822 = ~w22815 & w22821;
assign w22823 = ~w22820 & w22822;
assign w22824 = pi1285 & ~w22823;
assign w22825 = ~pi1285 & w22823;
assign w22826 = ~w22824 & ~w22825;
assign w22827 = ~w22481 & ~w22514;
assign w22828 = w22482 & w22827;
assign w22829 = ~w22479 & w22501;
assign w22830 = ~w22449 & w22500;
assign w22831 = ~w22508 & ~w22830;
assign w22832 = ~w22513 & ~w22831;
assign w22833 = ~w22474 & w22484;
assign w22834 = ~w22832 & w63759;
assign w22835 = (w22492 & w22834) | (w22492 & w65486) | (w22834 & w65486);
assign w22836 = w22448 & w22455;
assign w22837 = ~w22506 & w22836;
assign w22838 = w22504 & w22837;
assign w22839 = (~w22492 & w22832) | (~w22492 & w65487) | (w22832 & w65487);
assign w22840 = w22449 & w22479;
assign w22841 = w22492 & w22510;
assign w22842 = ~w22840 & ~w22841;
assign w22843 = ~w22455 & ~w22842;
assign w22844 = w22476 & w22828;
assign w22845 = ~w22843 & ~w22844;
assign w22846 = ~w22838 & w22845;
assign w22847 = ~w22839 & w22846;
assign w22848 = (pi1252 & ~w22847) | (pi1252 & w65488) | (~w22847 & w65488);
assign w22849 = w22847 & w65489;
assign w22850 = ~w22848 & ~w22849;
assign w22851 = (w22641 & w22655) | (w22641 & w63760) | (w22655 & w63760);
assign w22852 = ~w22641 & ~w22654;
assign w22853 = ~w22851 & ~w22852;
assign w22854 = ~w22635 & ~w22684;
assign w22855 = w22668 & w22854;
assign w22856 = ~w22853 & w22855;
assign w22857 = w22654 & w22667;
assign w22858 = ~w22682 & ~w22857;
assign w22859 = ~w22680 & ~w22858;
assign w22860 = w22662 & ~w22682;
assign w22861 = w22666 & ~w22691;
assign w22862 = ~w22860 & ~w22861;
assign w22863 = ~w22676 & ~w22862;
assign w22864 = ~w22859 & w22863;
assign w22865 = ~w22856 & w22864;
assign w22866 = w22662 & ~w22854;
assign w22867 = w22858 & w22866;
assign w22868 = w22635 & w22648;
assign w22869 = w22628 & w22649;
assign w22870 = ~w22666 & ~w22869;
assign w22871 = ~w22662 & ~w22870;
assign w22872 = w22868 & w22871;
assign w22873 = w22650 & w22854;
assign w22874 = w22676 & ~w22873;
assign w22875 = ~w22867 & w22874;
assign w22876 = ~w22872 & w22875;
assign w22877 = ~w22865 & ~w22876;
assign w22878 = pi1249 & w22877;
assign w22879 = ~pi1249 & ~w22877;
assign w22880 = ~w22878 & ~w22879;
assign w22881 = ~w22770 & ~w22793;
assign w22882 = ~w22786 & ~w22881;
assign w22883 = w22767 & ~w22882;
assign w22884 = w22723 & w22748;
assign w22885 = ~w22883 & ~w22884;
assign w22886 = ~w22792 & ~w22885;
assign w22887 = w22738 & ~w22746;
assign w22888 = w22722 & w22752;
assign w22889 = w22887 & w22888;
assign w22890 = w22724 & w22761;
assign w22891 = w22746 & ~w22796;
assign w22892 = w22882 & w22891;
assign w22893 = w22758 & ~w22786;
assign w22894 = ~w22765 & w22893;
assign w22895 = w22779 & ~w22787;
assign w22896 = ~w22890 & w22895;
assign w22897 = ~w22894 & w22896;
assign w22898 = ~w22892 & w22897;
assign w22899 = ~w22758 & ~w22793;
assign w22900 = ~w22887 & w22899;
assign w22901 = w22769 & w22900;
assign w22902 = w22747 & ~w22760;
assign w22903 = ~w22739 & w22764;
assign w22904 = ~w22887 & w22903;
assign w22905 = ~w22779 & ~w22902;
assign w22906 = ~w22904 & w22905;
assign w22907 = ~w22901 & w22906;
assign w22908 = ~w22898 & ~w22907;
assign w22909 = ~w22886 & ~w22889;
assign w22910 = ~w22908 & w22909;
assign w22911 = pi1255 & ~w22910;
assign w22912 = ~pi1255 & w22910;
assign w22913 = ~w22911 & ~w22912;
assign w22914 = ~pi4042 & pi9040;
assign w22915 = ~pi4200 & ~pi9040;
assign w22916 = ~w22914 & ~w22915;
assign w22917 = pi1242 & ~w22916;
assign w22918 = ~pi1242 & w22916;
assign w22919 = ~w22917 & ~w22918;
assign w22920 = ~pi4137 & pi9040;
assign w22921 = ~pi4446 & ~pi9040;
assign w22922 = ~w22920 & ~w22921;
assign w22923 = pi1216 & ~w22922;
assign w22924 = ~pi1216 & w22922;
assign w22925 = ~w22923 & ~w22924;
assign w22926 = ~pi4037 & pi9040;
assign w22927 = ~pi4159 & ~pi9040;
assign w22928 = ~w22926 & ~w22927;
assign w22929 = pi1234 & ~w22928;
assign w22930 = ~pi1234 & w22928;
assign w22931 = ~w22929 & ~w22930;
assign w22932 = ~w22925 & w22931;
assign w22933 = ~pi4446 & pi9040;
assign w22934 = ~pi4042 & ~pi9040;
assign w22935 = ~w22933 & ~w22934;
assign w22936 = pi1229 & ~w22935;
assign w22937 = ~pi1229 & w22935;
assign w22938 = ~w22936 & ~w22937;
assign w22939 = w22932 & ~w22938;
assign w22940 = ~pi4036 & pi9040;
assign w22941 = ~pi4252 & ~pi9040;
assign w22942 = ~w22940 & ~w22941;
assign w22943 = pi1230 & ~w22942;
assign w22944 = ~pi1230 & w22942;
assign w22945 = ~w22943 & ~w22944;
assign w22946 = w22931 & ~w22945;
assign w22947 = w22925 & w22938;
assign w22948 = w22946 & w22947;
assign w22949 = ~w22925 & w22945;
assign w22950 = ~w22938 & ~w22949;
assign w22951 = w22938 & w22949;
assign w22952 = ~w22950 & ~w22951;
assign w22953 = ~pi4128 & pi9040;
assign w22954 = ~pi4121 & ~pi9040;
assign w22955 = ~w22953 & ~w22954;
assign w22956 = pi1243 & ~w22955;
assign w22957 = ~pi1243 & w22955;
assign w22958 = ~w22956 & ~w22957;
assign w22959 = ~w22932 & ~w22958;
assign w22960 = w22952 & w22959;
assign w22961 = ~w22939 & ~w22948;
assign w22962 = ~w22960 & w22961;
assign w22963 = ~w22919 & ~w22962;
assign w22964 = w22932 & w23161;
assign w22965 = ~w22931 & w22938;
assign w22966 = ~w22919 & ~w22949;
assign w22967 = w22965 & ~w22966;
assign w22968 = w22938 & w22945;
assign w22969 = w22919 & w22925;
assign w22970 = w22968 & w22969;
assign w22971 = ~w22925 & ~w22945;
assign w22972 = w22938 & w22971;
assign w22973 = w22925 & ~w22945;
assign w22974 = ~w22938 & w22973;
assign w22975 = w22931 & w22974;
assign w22976 = ~w22972 & ~w22975;
assign w22977 = w22919 & ~w22976;
assign w22978 = ~w22946 & w22950;
assign w22979 = ~w22919 & w22978;
assign w22980 = w22958 & ~w22970;
assign w22981 = ~w22964 & w22980;
assign w22982 = ~w22967 & w22981;
assign w22983 = ~w22979 & w22982;
assign w22984 = ~w22977 & w22983;
assign w22985 = w22919 & w22978;
assign w22986 = w22932 & ~w22952;
assign w22987 = ~w22948 & ~w22958;
assign w22988 = ~w22985 & w22987;
assign w22989 = ~w22986 & w22988;
assign w22990 = (~w22963 & w22984) | (~w22963 & w65490) | (w22984 & w65490);
assign w22991 = ~pi1266 & w22990;
assign w22992 = pi1266 & ~w22990;
assign w22993 = ~w22991 & ~w22992;
assign w22994 = ~w22288 & w22324;
assign w22995 = w22358 & w22994;
assign w22996 = ~w22315 & w65491;
assign w22997 = (~w22324 & w22317) | (~w22324 & w65492) | (w22317 & w65492);
assign w22998 = ~w22309 & ~w22336;
assign w22999 = ~w22303 & w22306;
assign w23000 = w22288 & ~w22999;
assign w23001 = w22282 & ~w22352;
assign w23002 = (w22324 & w22352) | (w22324 & w65493) | (w22352 & w65493);
assign w23003 = w23000 & w23002;
assign w23004 = ~w22359 & w22998;
assign w23005 = ~w23003 & w23004;
assign w23006 = w22288 & ~w22324;
assign w23007 = ~w22356 & ~w23006;
assign w23008 = ~w22309 & ~w22313;
assign w23009 = ~w23007 & w23008;
assign w23010 = w22310 & w22348;
assign w23011 = w22302 & w22332;
assign w23012 = ~w23009 & ~w23011;
assign w23013 = ~w23010 & w23012;
assign w23014 = ~w22331 & ~w23013;
assign w23015 = ~w22366 & ~w22995;
assign w23016 = (w23015 & w23005) | (w23015 & w65494) | (w23005 & w65494);
assign w23017 = ~w22997 & w23016;
assign w23018 = ~w23014 & w23017;
assign w23019 = pi1272 & ~w23018;
assign w23020 = ~pi1272 & w23018;
assign w23021 = ~w23019 & ~w23020;
assign w23022 = ~pi4097 & pi9040;
assign w23023 = ~pi4300 & ~pi9040;
assign w23024 = ~w23022 & ~w23023;
assign w23025 = pi1224 & ~w23024;
assign w23026 = ~pi1224 & w23024;
assign w23027 = ~w23025 & ~w23026;
assign w23028 = ~pi4317 & pi9040;
assign w23029 = ~pi4097 & ~pi9040;
assign w23030 = ~w23028 & ~w23029;
assign w23031 = pi1243 & ~w23030;
assign w23032 = ~pi1243 & w23030;
assign w23033 = ~w23031 & ~w23032;
assign w23034 = ~pi4099 & pi9040;
assign w23035 = ~pi4129 & ~pi9040;
assign w23036 = ~w23034 & ~w23035;
assign w23037 = pi1223 & ~w23036;
assign w23038 = ~pi1223 & w23036;
assign w23039 = ~w23037 & ~w23038;
assign w23040 = ~w23033 & w23039;
assign w23041 = ~pi4105 & pi9040;
assign w23042 = ~pi4169 & ~pi9040;
assign w23043 = ~w23041 & ~w23042;
assign w23044 = pi1219 & ~w23043;
assign w23045 = ~pi1219 & w23043;
assign w23046 = ~w23044 & ~w23045;
assign w23047 = ~w23033 & w23046;
assign w23048 = w23033 & ~w23046;
assign w23049 = ~w23047 & ~w23048;
assign w23050 = ~w23040 & ~w23049;
assign w23051 = ~pi4101 & pi9040;
assign w23052 = ~pi4190 & ~pi9040;
assign w23053 = ~w23051 & ~w23052;
assign w23054 = pi1230 & ~w23053;
assign w23055 = ~pi1230 & w23053;
assign w23056 = ~w23054 & ~w23055;
assign w23057 = ~pi4044 & pi9040;
assign w23058 = ~pi4037 & ~pi9040;
assign w23059 = ~w23057 & ~w23058;
assign w23060 = pi1208 & ~w23059;
assign w23061 = ~pi1208 & w23059;
assign w23062 = ~w23060 & ~w23061;
assign w23063 = w23056 & w23062;
assign w23064 = ~w23033 & ~w23046;
assign w23065 = w23033 & w23046;
assign w23066 = w23056 & w23065;
assign w23067 = ~w23056 & ~w23065;
assign w23068 = ~w23066 & ~w23067;
assign w23069 = ~w23064 & w23068;
assign w23070 = ~w23062 & ~w23064;
assign w23071 = w23056 & ~w23062;
assign w23072 = w23039 & w23071;
assign w23073 = ~w23070 & ~w23072;
assign w23074 = ~w23069 & ~w23073;
assign w23075 = (~w23063 & w23069) | (~w23063 & w63761) | (w23069 & w63761);
assign w23076 = w23050 & ~w23075;
assign w23077 = ~w23056 & ~w23062;
assign w23078 = w23049 & ~w23077;
assign w23079 = ~w23063 & w23078;
assign w23080 = w23040 & w23071;
assign w23081 = ~w23079 & ~w23080;
assign w23082 = (~w23027 & w23076) | (~w23027 & w65495) | (w23076 & w65495);
assign w23083 = w23064 & w23077;
assign w23084 = w23047 & w23062;
assign w23085 = ~w23046 & w23056;
assign w23086 = w23033 & w23085;
assign w23087 = ~w23084 & ~w23086;
assign w23088 = w23046 & ~w23056;
assign w23089 = (~w23088 & w23087) | (~w23088 & w63762) | (w23087 & w63762);
assign w23090 = ~w23027 & ~w23062;
assign w23091 = (~w23087 & w65496) | (~w23087 & w65497) | (w65496 & w65497);
assign w23092 = ~w23083 & ~w23091;
assign w23093 = w23039 & ~w23092;
assign w23094 = w23039 & ~w23064;
assign w23095 = ~w23063 & w23064;
assign w23096 = w23027 & ~w23094;
assign w23097 = ~w23095 & w23096;
assign w23098 = w23089 & w23097;
assign w23099 = ~w23093 & ~w23098;
assign w23100 = ~w23082 & w23099;
assign w23101 = pi1273 & ~w23100;
assign w23102 = ~pi1273 & w23100;
assign w23103 = ~w23101 & ~w23102;
assign w23104 = w22652 & w22679;
assign w23105 = ~w22663 & ~w23104;
assign w23106 = w22641 & ~w23105;
assign w23107 = ~w22654 & w65498;
assign w23108 = w22662 & ~w23107;
assign w23109 = w22634 & w22682;
assign w23110 = ~w22662 & ~w23109;
assign w23111 = ~w22665 & w22699;
assign w23112 = ~w22855 & w23111;
assign w23113 = ~w22655 & w23110;
assign w23114 = ~w23112 & w23113;
assign w23115 = (~w22655 & w65499) | (~w22655 & w65500) | (w65499 & w65500);
assign w23116 = (w23115 & w23114) | (w23115 & w63763) | (w23114 & w63763);
assign w23117 = ~w22851 & w65501;
assign w23118 = ~w22662 & w23107;
assign w23119 = ~w22676 & ~w22683;
assign w23120 = ~w23118 & w23119;
assign w23121 = ~w23117 & w23120;
assign w23122 = (~w23106 & w23116) | (~w23106 & w65502) | (w23116 & w65502);
assign w23123 = pi1260 & w23122;
assign w23124 = ~pi1260 & ~w23122;
assign w23125 = ~w23123 & ~w23124;
assign w23126 = w23046 & w23080;
assign w23127 = w23033 & w23062;
assign w23128 = ~w23085 & ~w23127;
assign w23129 = ~w23039 & ~w23128;
assign w23130 = ~w23046 & w23063;
assign w23131 = ~w23129 & ~w23130;
assign w23132 = w23066 & ~w23131;
assign w23133 = ~w23033 & ~w23056;
assign w23134 = ~w23039 & ~w23133;
assign w23135 = w23128 & ~w23134;
assign w23136 = w23048 & w23135;
assign w23137 = ~w23046 & w23062;
assign w23138 = (w23040 & w23070) | (w23040 & w63764) | (w23070 & w63764);
assign w23139 = ~w23048 & ~w23137;
assign w23140 = ~w23039 & w23139;
assign w23141 = ~w23056 & w23127;
assign w23142 = ~w23140 & w23141;
assign w23143 = ~w23138 & ~w23142;
assign w23144 = (~w23039 & ~w23049) | (~w23039 & w63765) | (~w23049 & w63765);
assign w23145 = ~w23069 & w65503;
assign w23146 = (w23027 & ~w23143) | (w23027 & w63766) | (~w23143 & w63766);
assign w23147 = ~w23145 & w23146;
assign w23148 = w23049 & w23077;
assign w23149 = w23087 & ~w23148;
assign w23150 = ~w23039 & ~w23149;
assign w23151 = ~w23027 & ~w23080;
assign w23152 = ~w23142 & w65504;
assign w23153 = ~w23150 & w23152;
assign w23154 = ~w23126 & ~w23136;
assign w23155 = ~w23132 & w23154;
assign w23156 = (w23155 & w23147) | (w23155 & w65505) | (w23147 & w65505);
assign w23157 = pi1267 & ~w23156;
assign w23158 = ~pi1267 & w23156;
assign w23159 = ~w23157 & ~w23158;
assign w23160 = ~w22919 & ~w22925;
assign w23161 = ~w22938 & w22945;
assign w23162 = ~w22925 & ~w22931;
assign w23163 = ~w23161 & ~w23162;
assign w23164 = ~w23160 & w23163;
assign w23165 = w22931 & ~w22938;
assign w23166 = w22971 & w23165;
assign w23167 = ~w22967 & ~w23166;
assign w23168 = w23164 & ~w23167;
assign w23169 = ~w22949 & ~w22973;
assign w23170 = w22965 & w23169;
assign w23171 = ~w22931 & w22945;
assign w23172 = w23160 & w23171;
assign w23173 = w22925 & w23161;
assign w23174 = w23161 & w63767;
assign w23175 = ~w23172 & ~w23174;
assign w23176 = ~w22938 & ~w22969;
assign w23177 = ~w23175 & w23176;
assign w23178 = (~w22919 & w22986) | (~w22919 & w65506) | (w22986 & w65506);
assign w23179 = w22969 & ~w23165;
assign w23180 = w22950 & w23160;
assign w23181 = w22958 & ~w23179;
assign w23182 = ~w23170 & w23181;
assign w23183 = ~w23180 & w23182;
assign w23184 = ~w23177 & w23183;
assign w23185 = ~w23178 & w23184;
assign w23186 = w22919 & ~w22951;
assign w23187 = w22919 & ~w23171;
assign w23188 = (~w23187 & ~w22952) | (~w23187 & w63768) | (~w22952 & w63768);
assign w23189 = (~w22958 & w23188) | (~w22958 & w65507) | (w23188 & w65507);
assign w23190 = ~w22931 & ~w22968;
assign w23191 = ~w23169 & w23190;
assign w23192 = w23175 & ~w23191;
assign w23193 = w23189 & w23192;
assign w23194 = (~w23168 & w23185) | (~w23168 & w65508) | (w23185 & w65508);
assign w23195 = pi1262 & w23194;
assign w23196 = ~pi1262 & ~w23194;
assign w23197 = ~w23195 & ~w23196;
assign w23198 = ~w22746 & w22771;
assign w23199 = w22760 & w22794;
assign w23200 = ~w22725 & w22887;
assign w23201 = ~w22887 & w22888;
assign w23202 = ~w22772 & w22790;
assign w23203 = ~w23199 & ~w23200;
assign w23204 = ~w23201 & w23203;
assign w23205 = w23202 & w23204;
assign w23206 = ~w22722 & w22750;
assign w23207 = ~w22768 & ~w23206;
assign w23208 = ~w22881 & ~w23207;
assign w23209 = w22740 & w22769;
assign w23210 = w22779 & ~w23209;
assign w23211 = ~w22762 & w23210;
assign w23212 = ~w22889 & w23211;
assign w23213 = ~w23208 & w23212;
assign w23214 = ~w23205 & ~w23213;
assign w23215 = ~w22722 & ~w22893;
assign w23216 = ~w22763 & w23215;
assign w23217 = ~w22785 & ~w23198;
assign w23218 = ~w23216 & w23217;
assign w23219 = ~w23214 & w23218;
assign w23220 = ~pi1265 & ~w23219;
assign w23221 = pi1265 & w23219;
assign w23222 = ~w23220 & ~w23221;
assign w23223 = w22288 & w22339;
assign w23224 = w22331 & ~w23223;
assign w23225 = ~w23008 & w23224;
assign w23226 = ~w22314 & ~w23225;
assign w23227 = w22324 & ~w23226;
assign w23228 = w22301 & w22339;
assign w23229 = w23006 & w23228;
assign w23230 = w22331 & ~w23229;
assign w23231 = ~w22324 & w23009;
assign w23232 = ~w22994 & w23228;
assign w23233 = ~w22308 & w22324;
assign w23234 = w23001 & w23233;
assign w23235 = w22308 & w22312;
assign w23236 = ~w22307 & ~w22359;
assign w23237 = ~w23235 & w23236;
assign w23238 = ~w23232 & ~w23234;
assign w23239 = w23237 & w23238;
assign w23240 = ~w23231 & w23239;
assign w23241 = ~w23230 & ~w23240;
assign w23242 = ~w22306 & ~w22357;
assign w23243 = w22304 & ~w23242;
assign w23244 = ~w22304 & ~w22332;
assign w23245 = w22331 & ~w22352;
assign w23246 = ~w23243 & w23245;
assign w23247 = ~w23244 & w23246;
assign w23248 = ~w23227 & ~w23247;
assign w23249 = ~w23241 & w23248;
assign w23250 = ~pi1258 & w23249;
assign w23251 = pi1258 & ~w23249;
assign w23252 = ~w23250 & ~w23251;
assign w23253 = w23068 & w23094;
assign w23254 = ~w23069 & w23140;
assign w23255 = ~w23027 & ~w23083;
assign w23256 = ~w23253 & w23255;
assign w23257 = ~w23254 & w23256;
assign w23258 = w23047 & w23063;
assign w23259 = ~w23039 & ~w23127;
assign w23260 = ~w23139 & w23259;
assign w23261 = w23027 & ~w23258;
assign w23262 = ~w23260 & w23261;
assign w23263 = ~w23074 & w23262;
assign w23264 = ~w23257 & ~w23263;
assign w23265 = ~w23056 & ~w23094;
assign w23266 = w23039 & w23086;
assign w23267 = ~w23265 & ~w23266;
assign w23268 = w23062 & ~w23259;
assign w23269 = ~w23267 & w23268;
assign w23270 = ~w23264 & ~w23269;
assign w23271 = ~pi1284 & w23270;
assign w23272 = pi1284 & ~w23270;
assign w23273 = ~w23271 & ~w23272;
assign w23274 = ~w23039 & w23130;
assign w23275 = w23131 & ~w23135;
assign w23276 = ~w23056 & ~w23149;
assign w23277 = ~w23275 & ~w23276;
assign w23278 = ~w23027 & ~w23277;
assign w23279 = w23027 & w23063;
assign w23280 = (~w23279 & w23140) | (~w23279 & w65509) | (w23140 & w65509);
assign w23281 = w23068 & ~w23280;
assign w23282 = ~w23070 & w23129;
assign w23283 = ~w23136 & ~w23138;
assign w23284 = ~w23282 & w23283;
assign w23285 = w23027 & ~w23284;
assign w23286 = ~w23274 & ~w23281;
assign w23287 = ~w23278 & w23286;
assign w23288 = (pi1274 & ~w23287) | (pi1274 & w65510) | (~w23287 & w65510);
assign w23289 = w23287 & w65511;
assign w23290 = ~w23288 & ~w23289;
assign w23291 = w22567 & ~w22602;
assign w23292 = w22592 & w23291;
assign w23293 = w22576 & w22569;
assign w23294 = ~w22545 & ~w22593;
assign w23295 = w22553 & w22593;
assign w23296 = ~w23294 & ~w23295;
assign w23297 = w22560 & ~w23296;
assign w23298 = w22581 & ~w23294;
assign w23299 = w22567 & w22590;
assign w23300 = ~w23293 & ~w23299;
assign w23301 = ~w23298 & w23300;
assign w23302 = ~w23297 & w23301;
assign w23303 = w22533 & ~w23302;
assign w23304 = w22539 & w22554;
assign w23305 = ~w22570 & ~w23304;
assign w23306 = ~w22571 & ~w23305;
assign w23307 = ~w22554 & ~w22560;
assign w23308 = ~w23291 & w23307;
assign w23309 = ~w23306 & ~w23308;
assign w23310 = ~w22533 & ~w23309;
assign w23311 = ~w23292 & ~w23303;
assign w23312 = ~w23310 & w23311;
assign w23313 = ~pi1276 & w23312;
assign w23314 = pi1276 & ~w23312;
assign w23315 = ~w23313 & ~w23314;
assign w23316 = (~w22331 & w23000) | (~w22331 & w65512) | (w23000 & w65512);
assign w23317 = w22316 & ~w22998;
assign w23318 = (w22324 & w23317) | (w22324 & w65513) | (w23317 & w65513);
assign w23319 = ~w22999 & ~w23235;
assign w23320 = w22337 & ~w23319;
assign w23321 = ~w22303 & w22324;
assign w23322 = w22357 & ~w23321;
assign w23323 = ~w22335 & w23322;
assign w23324 = ~w22353 & ~w22357;
assign w23325 = w22302 & ~w23324;
assign w23326 = ~w22307 & ~w22994;
assign w23327 = w22312 & ~w23326;
assign w23328 = ~w23223 & ~w23325;
assign w23329 = ~w23327 & w23328;
assign w23330 = w22331 & ~w23329;
assign w23331 = ~w23320 & ~w23323;
assign w23332 = ~w23318 & w23331;
assign w23333 = ~w23330 & w23332;
assign w23334 = pi1270 & ~w23333;
assign w23335 = ~pi1270 & w23333;
assign w23336 = ~w23334 & ~w23335;
assign w23337 = ~w22779 & ~w23206;
assign w23338 = ~w22739 & w22746;
assign w23339 = w22760 & w23338;
assign w23340 = ~w22722 & w22731;
assign w23341 = (w23340 & ~w22899) | (w23340 & w65514) | (~w22899 & w65514);
assign w23342 = ~w23339 & ~w23341;
assign w23343 = ~w23337 & ~w23342;
assign w23344 = ~w22731 & w22779;
assign w23345 = w22751 & w23344;
assign w23346 = ~w22762 & ~w22789;
assign w23347 = ~w23345 & w23346;
assign w23348 = w22722 & ~w23347;
assign w23349 = w22739 & w22784;
assign w23350 = w22724 & ~w22891;
assign w23351 = w23342 & w23350;
assign w23352 = ~w22755 & w65515;
assign w23353 = ~w23351 & w23352;
assign w23354 = ~w22779 & ~w23353;
assign w23355 = ~w23343 & ~w23348;
assign w23356 = ~w23354 & w23355;
assign w23357 = pi1264 & ~w23356;
assign w23358 = ~pi1264 & w23356;
assign w23359 = ~w23357 & ~w23358;
assign w23360 = ~w22471 & w22481;
assign w23361 = w22442 & w22506;
assign w23362 = ~w23360 & ~w23361;
assign w23363 = w22475 & w23362;
assign w23364 = ~w22476 & ~w22499;
assign w23365 = w23362 & w65516;
assign w23366 = w22493 & w23361;
assign w23367 = ~w22510 & w22827;
assign w23368 = ~w22495 & ~w22827;
assign w23369 = ~w23367 & ~w23368;
assign w23370 = ~w22840 & ~w23366;
assign w23371 = ~w23369 & w23370;
assign w23372 = (w22492 & ~w23371) | (w22492 & w65517) | (~w23371 & w65517);
assign w23373 = ~w22457 & ~w22506;
assign w23374 = w22827 & w23373;
assign w23375 = ~w22455 & ~w22511;
assign w23376 = ~w23374 & w23375;
assign w23377 = ~w22499 & ~w22500;
assign w23378 = ~w22442 & ~w23377;
assign w23379 = ~w22455 & ~w22479;
assign w23380 = ~w23378 & w23379;
assign w23381 = w22457 & w22479;
assign w23382 = ~w22483 & ~w23381;
assign w23383 = ~w23380 & w23382;
assign w23384 = ~w23376 & ~w23383;
assign w23385 = (w23376 & ~w23371) | (w23376 & w65518) | (~w23371 & w65518);
assign w23386 = ~w22492 & ~w23363;
assign w23387 = ~w23385 & w23386;
assign w23388 = ~w23372 & ~w23384;
assign w23389 = ~w23387 & w23388;
assign w23390 = ~pi1269 & w23389;
assign w23391 = pi1269 & ~w23389;
assign w23392 = ~w23390 & ~w23391;
assign w23393 = (~w22662 & w22855) | (~w22662 & w65519) | (w22855 & w65519);
assign w23394 = w22641 & w22685;
assign w23395 = w22650 & ~w22667;
assign w23396 = w22860 & w23395;
assign w23397 = ~w23104 & ~w23394;
assign w23398 = ~w23396 & w23397;
assign w23399 = ~w23393 & w23398;
assign w23400 = w22676 & ~w23399;
assign w23401 = ~w22690 & w23110;
assign w23402 = w22662 & ~w22868;
assign w23403 = ~w23401 & ~w23402;
assign w23404 = (w22662 & ~w22653) | (w22662 & w65520) | (~w22653 & w65520);
assign w23405 = ~w22869 & w23404;
assign w23406 = ~w22871 & ~w23405;
assign w23407 = ~w22650 & w22684;
assign w23408 = ~w22689 & ~w23407;
assign w23409 = (~w22676 & w23406) | (~w22676 & w65521) | (w23406 & w65521);
assign w23410 = ~w23403 & ~w23409;
assign w23411 = ~w23400 & w23410;
assign w23412 = ~pi1257 & w23411;
assign w23413 = pi1257 & ~w23411;
assign w23414 = ~w23412 & ~w23413;
assign w23415 = w22570 & ~w22578;
assign w23416 = ~w22611 & ~w23415;
assign w23417 = ~w22601 & ~w23299;
assign w23418 = w22533 & w23417;
assign w23419 = ~w23416 & ~w23418;
assign w23420 = ~w22570 & ~w22577;
assign w23421 = w22606 & w23420;
assign w23422 = w22533 & w22539;
assign w23423 = ~w22574 & ~w22610;
assign w23424 = w23422 & w23423;
assign w23425 = w22533 & ~w22539;
assign w23426 = ~w23420 & w23425;
assign w23427 = ~w23415 & w23426;
assign w23428 = ~w23421 & ~w23424;
assign w23429 = ~w23427 & w23428;
assign w23430 = ~w23419 & w23429;
assign w23431 = pi1283 & ~w23430;
assign w23432 = ~pi1283 & w23430;
assign w23433 = ~w23431 & ~w23432;
assign w23434 = ~w22946 & ~w23171;
assign w23435 = w22947 & ~w23434;
assign w23436 = w22965 & w22971;
assign w23437 = ~w22974 & ~w23436;
assign w23438 = (~w22958 & ~w23437) | (~w22958 & w65522) | (~w23437 & w65522);
assign w23439 = ~w23435 & ~w23438;
assign w23440 = w22919 & ~w22958;
assign w23441 = ~w23439 & ~w23440;
assign w23442 = ~w23161 & w23440;
assign w23443 = ~w23163 & ~w23187;
assign w23444 = ~w23164 & ~w23443;
assign w23445 = w22973 & w65523;
assign w23446 = w23175 & ~w23445;
assign w23447 = ~w23444 & w23446;
assign w23448 = (~w23442 & w23447) | (~w23442 & w65524) | (w23447 & w65524);
assign w23449 = w23439 & ~w23448;
assign w23450 = ~w22938 & w23171;
assign w23451 = w23189 & w23450;
assign w23452 = ~w23441 & ~w23451;
assign w23453 = ~w23449 & w23452;
assign w23454 = pi1278 & ~w23453;
assign w23455 = ~pi1278 & w23453;
assign w23456 = ~w23454 & ~w23455;
assign w23457 = w22590 & w22601;
assign w23458 = w22575 & ~w22576;
assign w23459 = w23423 & w23458;
assign w23460 = w22533 & ~w23295;
assign w23461 = ~w22579 & w23460;
assign w23462 = ~w22612 & w23461;
assign w23463 = ~w23459 & w23462;
assign w23464 = ~w22591 & ~w23307;
assign w23465 = w22590 & ~w23464;
assign w23466 = ~w22533 & ~w22594;
assign w23467 = w23417 & w23466;
assign w23468 = ~w23465 & w23467;
assign w23469 = ~w22560 & ~w22605;
assign w23470 = w23305 & w23469;
assign w23471 = w22569 & w22591;
assign w23472 = ~w23422 & w23471;
assign w23473 = ~w22613 & ~w23457;
assign w23474 = ~w23472 & w23473;
assign w23475 = ~w23470 & w23474;
assign w23476 = (w23475 & w23463) | (w23475 & w65525) | (w23463 & w65525);
assign w23477 = pi1286 & w23476;
assign w23478 = ~pi1286 & ~w23476;
assign w23479 = ~w23477 & ~w23478;
assign w23480 = w22831 & w23369;
assign w23481 = ~w22449 & ~w22479;
assign w23482 = w22479 & ~w22836;
assign w23483 = ~w22492 & ~w23482;
assign w23484 = (~w23483 & w22831) | (~w23483 & w65526) | (w22831 & w65526);
assign w23485 = ~w23481 & ~w23484;
assign w23486 = w22514 & ~w23361;
assign w23487 = ~w22512 & w23486;
assign w23488 = w22829 & w23362;
assign w23489 = w22492 & ~w22840;
assign w23490 = ~w23487 & w23489;
assign w23491 = ~w23488 & w23490;
assign w23492 = ~w22477 & ~w22492;
assign w23493 = ~w23380 & w23492;
assign w23494 = ~w23491 & ~w23493;
assign w23495 = ~w22844 & ~w23480;
assign w23496 = ~w23485 & w23495;
assign w23497 = ~w23494 & w23496;
assign w23498 = pi1282 & ~w23497;
assign w23499 = ~pi1282 & w23497;
assign w23500 = ~w23498 & ~w23499;
assign w23501 = ~w22968 & ~w23445;
assign w23502 = w23187 & ~w23501;
assign w23503 = ~w22971 & ~w23171;
assign w23504 = w22938 & w22958;
assign w23505 = ~w23503 & w23504;
assign w23506 = ~w23173 & ~w23505;
assign w23507 = ~w22919 & ~w23506;
assign w23508 = ~w23169 & w23186;
assign w23509 = w22958 & ~w23166;
assign w23510 = ~w23508 & w23509;
assign w23511 = w22925 & ~w22931;
assign w23512 = ~w22932 & w23176;
assign w23513 = ~w22925 & ~w23165;
assign w23514 = w23434 & w23513;
assign w23515 = ~w23512 & ~w23514;
assign w23516 = ~w23511 & ~w23515;
assign w23517 = ~w22970 & w22987;
assign w23518 = ~w23516 & w23517;
assign w23519 = ~w23510 & ~w23518;
assign w23520 = ~w23502 & ~w23507;
assign w23521 = ~w23519 & w23520;
assign w23522 = pi1292 & w23521;
assign w23523 = ~pi1292 & ~w23521;
assign w23524 = ~w23522 & ~w23523;
assign w23525 = ~pi4379 & pi9040;
assign w23526 = ~pi4306 & ~pi9040;
assign w23527 = ~w23525 & ~w23526;
assign w23528 = pi1310 & ~w23527;
assign w23529 = ~pi1310 & w23527;
assign w23530 = ~w23528 & ~w23529;
assign w23531 = ~pi4303 & pi9040;
assign w23532 = ~pi4309 & ~pi9040;
assign w23533 = ~w23531 & ~w23532;
assign w23534 = pi1271 & ~w23533;
assign w23535 = ~pi1271 & w23533;
assign w23536 = ~w23534 & ~w23535;
assign w23537 = ~pi4505 & pi9040;
assign w23538 = ~pi4214 & ~pi9040;
assign w23539 = ~w23537 & ~w23538;
assign w23540 = pi1307 & ~w23539;
assign w23541 = ~pi1307 & w23539;
assign w23542 = ~w23540 & ~w23541;
assign w23543 = w23536 & ~w23542;
assign w23544 = ~pi4491 & pi9040;
assign w23545 = ~pi4292 & ~pi9040;
assign w23546 = ~w23544 & ~w23545;
assign w23547 = pi1302 & ~w23546;
assign w23548 = ~pi1302 & w23546;
assign w23549 = ~w23547 & ~w23548;
assign w23550 = w23543 & ~w23549;
assign w23551 = ~pi4306 & pi9040;
assign w23552 = ~pi4491 & ~pi9040;
assign w23553 = ~w23551 & ~w23552;
assign w23554 = pi1288 & ~w23553;
assign w23555 = ~pi1288 & w23553;
assign w23556 = ~w23554 & ~w23555;
assign w23557 = w23542 & w23556;
assign w23558 = ~pi4302 & pi9040;
assign w23559 = ~pi4308 & ~pi9040;
assign w23560 = ~w23558 & ~w23559;
assign w23561 = pi1306 & ~w23560;
assign w23562 = ~pi1306 & w23560;
assign w23563 = ~w23561 & ~w23562;
assign w23564 = w23536 & ~w23563;
assign w23565 = ~w23549 & ~w23564;
assign w23566 = ~w23536 & w23563;
assign w23567 = ~w23565 & ~w23566;
assign w23568 = ~w23565 & w65527;
assign w23569 = ~w23542 & ~w23556;
assign w23570 = ~w23536 & w23549;
assign w23571 = w23563 & ~w23570;
assign w23572 = w23569 & ~w23571;
assign w23573 = w23542 & ~w23549;
assign w23574 = w23566 & w23573;
assign w23575 = ~w23550 & ~w23574;
assign w23576 = ~w23572 & w23575;
assign w23577 = (~w23530 & ~w23576) | (~w23530 & w65528) | (~w23576 & w65528);
assign w23578 = ~w23556 & ~w23574;
assign w23579 = ~w23536 & ~w23563;
assign w23580 = ~w23542 & w23579;
assign w23581 = w23542 & w23564;
assign w23582 = ~w23580 & ~w23581;
assign w23583 = w23563 & w23569;
assign w23584 = w23542 & ~w23556;
assign w23585 = w23536 & w23563;
assign w23586 = ~w23542 & w23549;
assign w23587 = w23585 & ~w23586;
assign w23588 = ~w23584 & w23587;
assign w23589 = ~w23583 & ~w23588;
assign w23590 = ~w23549 & w23578;
assign w23591 = w23582 & w23590;
assign w23592 = w23589 & w23591;
assign w23593 = ~w23536 & w23573;
assign w23594 = ~w23550 & ~w23593;
assign w23595 = w23556 & w23563;
assign w23596 = ~w23594 & w23595;
assign w23597 = w23530 & ~w23574;
assign w23598 = w23579 & w63769;
assign w23599 = ~w23556 & ~w23598;
assign w23600 = (~w23542 & w23564) | (~w23542 & w23586) | (w23564 & w23586);
assign w23601 = ~w23599 & w23600;
assign w23602 = (~w23542 & ~w23569) | (~w23542 & w65529) | (~w23569 & w65529);
assign w23603 = ~w23549 & ~w23602;
assign w23604 = (w23536 & w23601) | (w23536 & w65530) | (w23601 & w65530);
assign w23605 = ~w23549 & w23556;
assign w23606 = w23566 & w23605;
assign w23607 = w23542 & w23549;
assign w23608 = w23579 & w23607;
assign w23609 = ~w23606 & ~w23608;
assign w23610 = ~w23572 & w23609;
assign w23611 = ~w23588 & w23597;
assign w23612 = w23610 & w23611;
assign w23613 = ~w23604 & w23612;
assign w23614 = ~w23577 & ~w23596;
assign w23615 = ~w23592 & w23614;
assign w23616 = ~w23613 & w23615;
assign w23617 = pi1318 & ~w23616;
assign w23618 = ~pi1318 & w23616;
assign w23619 = ~w23617 & ~w23618;
assign w23620 = ~w23549 & w23581;
assign w23621 = w23556 & ~w23620;
assign w23622 = w23564 & w23586;
assign w23623 = ~w23598 & ~w23622;
assign w23624 = w23621 & w23623;
assign w23625 = ~w23578 & ~w23624;
assign w23626 = w23549 & ~w23556;
assign w23627 = w23564 & w23626;
assign w23628 = ~w23530 & ~w23608;
assign w23629 = w23557 & w23570;
assign w23630 = w23580 & ~w23626;
assign w23631 = ~w23627 & ~w23629;
assign w23632 = w23628 & w23631;
assign w23633 = ~w23630 & w23632;
assign w23634 = w23589 & w23633;
assign w23635 = w23549 & ~w23582;
assign w23636 = ~w23582 & w65531;
assign w23637 = ~w23556 & w23594;
assign w23638 = ~w23542 & w23566;
assign w23639 = w23556 & ~w23581;
assign w23640 = ~w23638 & w23639;
assign w23641 = ~w23637 & ~w23640;
assign w23642 = w23585 & w23607;
assign w23643 = w23597 & ~w23642;
assign w23644 = ~w23636 & w23643;
assign w23645 = ~w23641 & w23644;
assign w23646 = ~w23634 & ~w23645;
assign w23647 = ~w23625 & ~w23646;
assign w23648 = ~pi1317 & w23647;
assign w23649 = pi1317 & ~w23647;
assign w23650 = ~w23648 & ~w23649;
assign w23651 = w23566 & w23586;
assign w23652 = ~w23642 & ~w23651;
assign w23653 = w23599 & w23652;
assign w23654 = ~w23621 & ~w23653;
assign w23655 = w23530 & ~w23651;
assign w23656 = w23557 & w23579;
assign w23657 = w23564 & ~w23573;
assign w23658 = ~w23574 & ~w23657;
assign w23659 = ~w23556 & ~w23658;
assign w23660 = w23587 & ~w23603;
assign w23661 = w23655 & ~w23656;
assign w23662 = ~w23659 & w23661;
assign w23663 = ~w23660 & w23662;
assign w23664 = ~w23598 & ~w23606;
assign w23665 = w23628 & w23664;
assign w23666 = ~w23636 & w23665;
assign w23667 = ~w23604 & w23666;
assign w23668 = ~w23663 & ~w23667;
assign w23669 = ~w23629 & ~w23654;
assign w23670 = ~w23668 & w23669;
assign w23671 = ~pi1320 & ~w23670;
assign w23672 = pi1320 & w23670;
assign w23673 = ~w23671 & ~w23672;
assign w23674 = ~pi4211 & pi9040;
assign w23675 = ~pi4246 & ~pi9040;
assign w23676 = ~w23674 & ~w23675;
assign w23677 = pi1291 & ~w23676;
assign w23678 = ~pi1291 & w23676;
assign w23679 = ~w23677 & ~w23678;
assign w23680 = ~pi4246 & pi9040;
assign w23681 = ~pi4505 & ~pi9040;
assign w23682 = ~w23680 & ~w23681;
assign w23683 = pi1259 & ~w23682;
assign w23684 = ~pi1259 & w23682;
assign w23685 = ~w23683 & ~w23684;
assign w23686 = ~pi4249 & pi9040;
assign w23687 = ~pi4215 & ~pi9040;
assign w23688 = ~w23686 & ~w23687;
assign w23689 = pi1309 & ~w23688;
assign w23690 = ~pi1309 & w23688;
assign w23691 = ~w23689 & ~w23690;
assign w23692 = ~w23685 & w23691;
assign w23693 = ~pi4404 & pi9040;
assign w23694 = ~pi4297 & ~pi9040;
assign w23695 = ~w23693 & ~w23694;
assign w23696 = pi1304 & ~w23695;
assign w23697 = ~pi1304 & w23695;
assign w23698 = ~w23696 & ~w23697;
assign w23699 = ~w23691 & w23698;
assign w23700 = ~w23692 & ~w23699;
assign w23701 = ~pi4292 & pi9040;
assign w23702 = ~pi4379 & ~pi9040;
assign w23703 = ~w23701 & ~w23702;
assign w23704 = pi1294 & ~w23703;
assign w23705 = ~pi1294 & w23703;
assign w23706 = ~w23704 & ~w23705;
assign w23707 = ~pi4493 & pi9040;
assign w23708 = ~pi4249 & ~pi9040;
assign w23709 = ~w23707 & ~w23708;
assign w23710 = pi1296 & ~w23709;
assign w23711 = ~pi1296 & w23709;
assign w23712 = ~w23710 & ~w23711;
assign w23713 = ~w23706 & ~w23712;
assign w23714 = w23700 & w23713;
assign w23715 = w23685 & ~w23691;
assign w23716 = w23706 & w23712;
assign w23717 = ~w23715 & ~w23716;
assign w23718 = w23706 & ~w23717;
assign w23719 = w23706 & ~w23712;
assign w23720 = w23700 & w23719;
assign w23721 = w23698 & w23712;
assign w23722 = w23715 & w23721;
assign w23723 = ~w23685 & w23698;
assign w23724 = ~w23692 & w23712;
assign w23725 = w23692 & ~w23712;
assign w23726 = ~w23724 & ~w23725;
assign w23727 = w23723 & w23726;
assign w23728 = ~w23720 & ~w23722;
assign w23729 = ~w23727 & w23728;
assign w23730 = w23685 & ~w23698;
assign w23731 = ~w23712 & w23723;
assign w23732 = ~w23730 & ~w23731;
assign w23733 = ~w23698 & ~w23712;
assign w23734 = ~w23713 & ~w23733;
assign w23735 = w23692 & w23721;
assign w23736 = (~w23735 & ~w23732) | (~w23735 & w65532) | (~w23732 & w65532);
assign w23737 = w23692 & w23736;
assign w23738 = (~w23714 & ~w23729) | (~w23714 & w63770) | (~w23729 & w63770);
assign w23739 = (w23679 & ~w23738) | (w23679 & w65533) | (~w23738 & w65533);
assign w23740 = ~w23722 & ~w23731;
assign w23741 = ~w23706 & ~w23740;
assign w23742 = ~w23706 & ~w23723;
assign w23743 = ~w23726 & w23742;
assign w23744 = (~w23679 & ~w23729) | (~w23679 & w65534) | (~w23729 & w65534);
assign w23745 = ~w23741 & ~w23744;
assign w23746 = ~w23739 & w23745;
assign w23747 = ~pi1319 & ~w23746;
assign w23748 = pi1319 & w23746;
assign w23749 = ~w23747 & ~w23748;
assign w23750 = ~pi4391 & pi9040;
assign w23751 = ~pi4311 & ~pi9040;
assign w23752 = ~w23750 & ~w23751;
assign w23753 = pi1300 & ~w23752;
assign w23754 = ~pi1300 & w23752;
assign w23755 = ~w23753 & ~w23754;
assign w23756 = ~pi4311 & pi9040;
assign w23757 = ~pi4284 & ~pi9040;
assign w23758 = ~w23756 & ~w23757;
assign w23759 = pi1289 & ~w23758;
assign w23760 = ~pi1289 & w23758;
assign w23761 = ~w23759 & ~w23760;
assign w23762 = ~pi4484 & pi9040;
assign w23763 = ~pi4293 & ~pi9040;
assign w23764 = ~w23762 & ~w23763;
assign w23765 = pi1280 & ~w23764;
assign w23766 = ~pi1280 & w23764;
assign w23767 = ~w23765 & ~w23766;
assign w23768 = ~w23761 & ~w23767;
assign w23769 = ~pi4497 & pi9040;
assign w23770 = ~pi4588 & ~pi9040;
assign w23771 = ~w23769 & ~w23770;
assign w23772 = pi1268 & ~w23771;
assign w23773 = ~pi1268 & w23771;
assign w23774 = ~w23772 & ~w23773;
assign w23775 = ~pi4588 & pi9040;
assign w23776 = ~pi4316 & ~pi9040;
assign w23777 = ~w23775 & ~w23776;
assign w23778 = pi1279 & ~w23777;
assign w23779 = ~pi1279 & w23777;
assign w23780 = ~w23778 & ~w23779;
assign w23781 = w23774 & ~w23780;
assign w23782 = w23768 & w23781;
assign w23783 = w23761 & ~w23774;
assign w23784 = ~w23767 & ~w23780;
assign w23785 = ~w23783 & w23784;
assign w23786 = w23767 & w23774;
assign w23787 = w23780 & w23786;
assign w23788 = ~w23785 & ~w23787;
assign w23789 = ~pi4285 & pi9040;
assign w23790 = ~pi4593 & ~pi9040;
assign w23791 = ~w23789 & ~w23790;
assign w23792 = pi1303 & ~w23791;
assign w23793 = ~pi1303 & w23791;
assign w23794 = ~w23792 & ~w23793;
assign w23795 = w23761 & w23767;
assign w23796 = w23767 & w23780;
assign w23797 = ~w23795 & ~w23796;
assign w23798 = ~w23774 & w23797;
assign w23799 = w23797 & w65535;
assign w23800 = ~w23774 & ~w23794;
assign w23801 = ~w23796 & w23800;
assign w23802 = ~w23761 & w23786;
assign w23803 = ~w23801 & ~w23802;
assign w23804 = w23780 & ~w23803;
assign w23805 = ~w23799 & ~w23804;
assign w23806 = ~w23768 & ~w23795;
assign w23807 = w23780 & ~w23806;
assign w23808 = ~w23785 & ~w23807;
assign w23809 = ~w23774 & w23780;
assign w23810 = w23794 & ~w23809;
assign w23811 = w23761 & w23810;
assign w23812 = w23808 & w23811;
assign w23813 = (~w23782 & w23788) | (~w23782 & w65536) | (w23788 & w65536);
assign w23814 = w23805 & w23813;
assign w23815 = (w23755 & ~w23814) | (w23755 & w65537) | (~w23814 & w65537);
assign w23816 = ~w23755 & w23794;
assign w23817 = ~w23782 & w23816;
assign w23818 = ~w23808 & w23817;
assign w23819 = ~w23755 & ~w23794;
assign w23820 = ~w23761 & w23780;
assign w23821 = w23774 & ~w23820;
assign w23822 = ~w23781 & ~w23796;
assign w23823 = w23821 & w23822;
assign w23824 = w23767 & w23809;
assign w23825 = ~w23823 & ~w23824;
assign w23826 = w23819 & ~w23825;
assign w23827 = w23768 & w23809;
assign w23828 = w23767 & w23794;
assign w23829 = ~w23780 & w23819;
assign w23830 = ~w23828 & ~w23829;
assign w23831 = w23783 & ~w23830;
assign w23832 = w23780 & ~w23783;
assign w23833 = ~w23755 & ~w23832;
assign w23834 = w23802 & w23833;
assign w23835 = ~w23827 & ~w23831;
assign w23836 = ~w23834 & w23835;
assign w23837 = ~w23818 & ~w23826;
assign w23838 = w23836 & w23837;
assign w23839 = ~w23815 & w23838;
assign w23840 = pi1316 & w23839;
assign w23841 = ~pi1316 & ~w23839;
assign w23842 = ~w23840 & ~w23841;
assign w23843 = ~pi4214 & pi9040;
assign w23844 = ~pi4211 & ~pi9040;
assign w23845 = ~w23843 & ~w23844;
assign w23846 = pi1299 & ~w23845;
assign w23847 = ~pi1299 & w23845;
assign w23848 = ~w23846 & ~w23847;
assign w23849 = ~pi4698 & pi9040;
assign w23850 = ~pi4213 & ~pi9040;
assign w23851 = ~w23849 & ~w23850;
assign w23852 = pi1259 & ~w23851;
assign w23853 = ~pi1259 & w23851;
assign w23854 = ~w23852 & ~w23853;
assign w23855 = w23848 & w23854;
assign w23856 = ~pi4310 & pi9040;
assign w23857 = ~pi4286 & ~pi9040;
assign w23858 = ~w23856 & ~w23857;
assign w23859 = pi1295 & ~w23858;
assign w23860 = ~pi1295 & w23858;
assign w23861 = ~w23859 & ~w23860;
assign w23862 = w23848 & ~w23861;
assign w23863 = ~w23848 & w23861;
assign w23864 = ~w23862 & ~w23863;
assign w23865 = ~w23855 & ~w23864;
assign w23866 = ~pi4373 & pi9040;
assign w23867 = ~pi4493 & ~pi9040;
assign w23868 = ~w23866 & ~w23867;
assign w23869 = pi1308 & ~w23868;
assign w23870 = ~pi1308 & w23868;
assign w23871 = ~w23869 & ~w23870;
assign w23872 = w23848 & ~w23871;
assign w23873 = w23854 & ~w23872;
assign w23874 = ~pi4215 & pi9040;
assign w23875 = ~pi4373 & ~pi9040;
assign w23876 = ~w23874 & ~w23875;
assign w23877 = pi1298 & ~w23876;
assign w23878 = ~pi1298 & w23876;
assign w23879 = ~w23877 & ~w23878;
assign w23880 = (~w23879 & w23865) | (~w23879 & w65538) | (w23865 & w65538);
assign w23881 = ~w23848 & w23871;
assign w23882 = ~w23854 & ~w23861;
assign w23883 = w23854 & w23861;
assign w23884 = ~w23882 & ~w23883;
assign w23885 = w23881 & w23884;
assign w23886 = ~pi4398 & pi9040;
assign w23887 = ~pi4205 & ~pi9040;
assign w23888 = ~w23886 & ~w23887;
assign w23889 = pi1296 & ~w23888;
assign w23890 = ~pi1296 & w23888;
assign w23891 = ~w23889 & ~w23890;
assign w23892 = w23848 & w23879;
assign w23893 = ~w23871 & w23892;
assign w23894 = w23891 & ~w23893;
assign w23895 = ~w23885 & w23894;
assign w23896 = ~w23880 & w23895;
assign w23897 = ~w23861 & ~w23879;
assign w23898 = ~w23861 & w23871;
assign w23899 = ~w23897 & ~w23898;
assign w23900 = w23855 & ~w23899;
assign w23901 = w23861 & w23879;
assign w23902 = ~w23848 & ~w23854;
assign w23903 = ~w23855 & ~w23902;
assign w23904 = w23871 & w23901;
assign w23905 = w23903 & w23904;
assign w23906 = ~w23900 & ~w23905;
assign w23907 = w23879 & w23902;
assign w23908 = ~w23861 & w23907;
assign w23909 = ~w23891 & ~w23908;
assign w23910 = w23906 & w23909;
assign w23911 = ~w23896 & ~w23910;
assign w23912 = w23848 & w23871;
assign w23913 = w23897 & w23912;
assign w23914 = ~w23901 & ~w23903;
assign w23915 = ~w23861 & ~w23892;
assign w23916 = w23914 & ~w23915;
assign w23917 = w23881 & w23916;
assign w23918 = w23879 & ~w23903;
assign w23919 = ~w23854 & w23879;
assign w23920 = w23854 & ~w23879;
assign w23921 = ~w23919 & ~w23920;
assign w23922 = w23903 & ~w23921;
assign w23923 = ~w23918 & ~w23922;
assign w23924 = ~w23884 & ~w23923;
assign w23925 = ~w23891 & ~w23892;
assign w23926 = ~w23920 & w23925;
assign w23927 = ~w23865 & w23926;
assign w23928 = ~w23924 & ~w23927;
assign w23929 = ~w23871 & ~w23928;
assign w23930 = ~w23913 & ~w23917;
assign w23931 = ~w23911 & w23930;
assign w23932 = ~w23929 & w23931;
assign w23933 = pi1312 & ~w23932;
assign w23934 = ~pi1312 & w23932;
assign w23935 = ~w23933 & ~w23934;
assign w23936 = ~pi4247 & pi9040;
assign w23937 = ~pi4280 & ~pi9040;
assign w23938 = ~w23936 & ~w23937;
assign w23939 = pi1287 & ~w23938;
assign w23940 = ~pi1287 & w23938;
assign w23941 = ~w23939 & ~w23940;
assign w23942 = ~pi4380 & pi9040;
assign w23943 = ~pi4208 & ~pi9040;
assign w23944 = ~w23942 & ~w23943;
assign w23945 = pi1298 & ~w23944;
assign w23946 = ~pi1298 & w23944;
assign w23947 = ~w23945 & ~w23946;
assign w23948 = w23941 & w23947;
assign w23949 = ~pi4254 & pi9040;
assign w23950 = ~pi4495 & ~pi9040;
assign w23951 = ~w23949 & ~w23950;
assign w23952 = pi1290 & ~w23951;
assign w23953 = ~pi1290 & w23951;
assign w23954 = ~w23952 & ~w23953;
assign w23955 = ~pi4294 & pi9040;
assign w23956 = ~pi4281 & ~pi9040;
assign w23957 = ~w23955 & ~w23956;
assign w23958 = pi1305 & ~w23957;
assign w23959 = ~pi1305 & w23957;
assign w23960 = ~w23958 & ~w23959;
assign w23961 = w23954 & ~w23960;
assign w23962 = ~w23954 & w23960;
assign w23963 = ~w23947 & w23962;
assign w23964 = ~w23961 & ~w23963;
assign w23965 = ~w23963 & w65539;
assign w23966 = ~pi4204 & pi9040;
assign w23967 = ~pi4296 & ~pi9040;
assign w23968 = ~w23966 & ~w23967;
assign w23969 = pi1275 & ~w23968;
assign w23970 = ~pi1275 & w23968;
assign w23971 = ~w23969 & ~w23970;
assign w23972 = ~w23965 & ~w23971;
assign w23973 = ~pi4281 & pi9040;
assign w23974 = ~pi4204 & ~pi9040;
assign w23975 = ~w23973 & ~w23974;
assign w23976 = pi1299 & ~w23975;
assign w23977 = ~pi1299 & w23975;
assign w23978 = ~w23976 & ~w23977;
assign w23979 = ~w23947 & w23954;
assign w23980 = w23941 & ~w23960;
assign w23981 = w23979 & w23980;
assign w23982 = ~w23971 & ~w23981;
assign w23983 = ~w23941 & ~w23954;
assign w23984 = ~w23947 & ~w23960;
assign w23985 = w23983 & w23984;
assign w23986 = ~w23941 & w23960;
assign w23987 = w23947 & w23986;
assign w23988 = w23986 & w63771;
assign w23989 = w23941 & ~w23947;
assign w23990 = ~w23961 & ~w23989;
assign w23991 = ~w23979 & ~w23980;
assign w23992 = ~w23990 & w23991;
assign w23993 = w23971 & ~w23985;
assign w23994 = ~w23988 & w23993;
assign w23995 = ~w23941 & w23954;
assign w23996 = w23960 & w23995;
assign w23997 = w23995 & w65540;
assign w23998 = w23994 & w63772;
assign w23999 = ~w23982 & ~w23998;
assign w24000 = w23947 & w23971;
assign w24001 = w23983 & w24000;
assign w24002 = ~w23981 & ~w23990;
assign w24003 = w23947 & ~w23980;
assign w24004 = ~w23990 & ~w24003;
assign w24005 = w23954 & w23960;
assign w24006 = ~w23986 & ~w24005;
assign w24007 = ~w24004 & w24006;
assign w24008 = ~w24007 & w63327;
assign w24009 = ~w24002 & w24008;
assign w24010 = ~w23978 & ~w24001;
assign w24011 = ~w23972 & w24010;
assign w24012 = ~w23999 & w24011;
assign w24013 = ~w24009 & w24012;
assign w24014 = w23948 & w23962;
assign w24015 = w23994 & w65541;
assign w24016 = ~w23960 & w23983;
assign w24017 = ~w23996 & ~w24016;
assign w24018 = w23982 & w24017;
assign w24019 = ~w24015 & ~w24018;
assign w24020 = w23978 & ~w24014;
assign w24021 = ~w24019 & w24020;
assign w24022 = (pi1314 & w24013) | (pi1314 & w65542) | (w24013 & w65542);
assign w24023 = ~w24013 & w65543;
assign w24024 = ~w24022 & ~w24023;
assign w24025 = ~w23715 & ~w23725;
assign w24026 = (~w23698 & w23725) | (~w23698 & w63773) | (w23725 & w63773);
assign w24027 = ~w23679 & ~w24026;
assign w24028 = ~w23698 & w23712;
assign w24029 = ~w23726 & ~w24028;
assign w24030 = w24027 & ~w24029;
assign w24031 = ~w23685 & ~w23691;
assign w24032 = ~w23713 & ~w24028;
assign w24033 = w24031 & ~w24032;
assign w24034 = w23685 & w23691;
assign w24035 = w24028 & w24034;
assign w24036 = w23679 & ~w24035;
assign w24037 = ~w24033 & w24036;
assign w24038 = w23698 & ~w23712;
assign w24039 = ~w24031 & ~w24038;
assign w24040 = ~w23717 & ~w24039;
assign w24041 = ~w23727 & ~w24040;
assign w24042 = w24037 & w24041;
assign w24043 = (~w23706 & w24042) | (~w23706 & w63774) | (w24042 & w63774);
assign w24044 = ~w23699 & ~w24028;
assign w24045 = ~w23732 & ~w24044;
assign w24046 = ~w24026 & w65544;
assign w24047 = w23685 & ~w24038;
assign w24048 = w24037 & ~w24047;
assign w24049 = ~w24046 & ~w24048;
assign w24050 = w23706 & ~w24045;
assign w24051 = ~w24049 & w24050;
assign w24052 = ~w24043 & ~w24051;
assign w24053 = w23679 & w23734;
assign w24054 = ~w23685 & ~w23706;
assign w24055 = (~w24054 & w24039) | (~w24054 & w65545) | (w24039 & w65545);
assign w24056 = w23691 & ~w23723;
assign w24057 = ~w24053 & w24056;
assign w24058 = ~w24055 & w24057;
assign w24059 = ~w24052 & w65546;
assign w24060 = (pi1322 & w24052) | (pi1322 & w65547) | (w24052 & w65547);
assign w24061 = ~w24059 & ~w24060;
assign w24062 = w23691 & ~w23712;
assign w24063 = (~w23712 & w24056) | (~w23712 & w63775) | (w24056 & w63775);
assign w24064 = ~w23698 & w24031;
assign w24065 = (w23712 & ~w24031) | (w23712 & w23721) | (~w24031 & w23721);
assign w24066 = ~w23679 & ~w24065;
assign w24067 = ~w24063 & w24066;
assign w24068 = ~w23722 & ~w24035;
assign w24069 = ~w24067 & w24068;
assign w24070 = ~w24067 & w65548;
assign w24071 = ~w24062 & ~w24070;
assign w24072 = ~w24055 & w24062;
assign w24073 = ~w23679 & ~w24072;
assign w24074 = ~w24071 & w24073;
assign w24075 = ~w23706 & ~w24069;
assign w24076 = ~w24028 & ~w24038;
assign w24077 = w24034 & ~w24076;
assign w24078 = ~w24039 & w65549;
assign w24079 = ~w24055 & ~w24078;
assign w24080 = w23715 & w24076;
assign w24081 = ~w24077 & ~w24080;
assign w24082 = ~w24079 & w24081;
assign w24083 = w23679 & ~w24082;
assign w24084 = ~w24075 & ~w24083;
assign w24085 = ~w24074 & w24084;
assign w24086 = ~pi1340 & w24085;
assign w24087 = pi1340 & ~w24085;
assign w24088 = ~w24086 & ~w24087;
assign w24089 = ~w23806 & w23829;
assign w24090 = ~w23761 & ~w23794;
assign w24091 = w23824 & w24090;
assign w24092 = ~w23783 & ~w23828;
assign w24093 = w23797 & ~w24092;
assign w24094 = (w24093 & w23804) | (w24093 & w65550) | (w23804 & w65550);
assign w24095 = w23761 & w23784;
assign w24096 = w23833 & ~w24095;
assign w24097 = ~w23795 & w23819;
assign w24098 = ~w24096 & ~w24097;
assign w24099 = ~w24094 & ~w24098;
assign w24100 = w23783 & w23794;
assign w24101 = ~w24090 & ~w24100;
assign w24102 = w23780 & ~w24101;
assign w24103 = w23781 & ~w23806;
assign w24104 = w23755 & ~w24093;
assign w24105 = ~w24103 & w24104;
assign w24106 = ~w23799 & ~w24102;
assign w24107 = w24105 & w24106;
assign w24108 = ~w24099 & ~w24107;
assign w24109 = ~w24089 & ~w24091;
assign w24110 = ~w24108 & w24109;
assign w24111 = pi1329 & ~w24110;
assign w24112 = ~pi1329 & w24110;
assign w24113 = ~w24111 & ~w24112;
assign w24114 = ~pi4382 & pi9040;
assign w24115 = ~pi4220 & ~pi9040;
assign w24116 = ~w24114 & ~w24115;
assign w24117 = pi1293 & ~w24116;
assign w24118 = ~pi1293 & w24116;
assign w24119 = ~w24117 & ~w24118;
assign w24120 = ~pi4280 & pi9040;
assign w24121 = ~pi4382 & ~pi9040;
assign w24122 = ~w24120 & ~w24121;
assign w24123 = pi1280 & ~w24122;
assign w24124 = ~pi1280 & w24122;
assign w24125 = ~w24123 & ~w24124;
assign w24126 = ~pi4495 & pi9040;
assign w24127 = ~pi4380 & ~pi9040;
assign w24128 = ~w24126 & ~w24127;
assign w24129 = pi1287 & ~w24128;
assign w24130 = ~pi1287 & w24128;
assign w24131 = ~w24129 & ~w24130;
assign w24132 = w24125 & w24131;
assign w24133 = ~pi4288 & pi9040;
assign w24134 = ~pi4497 & ~pi9040;
assign w24135 = ~w24133 & ~w24134;
assign w24136 = pi1300 & ~w24135;
assign w24137 = ~pi1300 & w24135;
assign w24138 = ~w24136 & ~w24137;
assign w24139 = ~pi4208 & pi9040;
assign w24140 = ~pi4254 & ~pi9040;
assign w24141 = ~w24139 & ~w24140;
assign w24142 = pi1281 & ~w24141;
assign w24143 = ~pi1281 & w24141;
assign w24144 = ~w24142 & ~w24143;
assign w24145 = ~w24138 & w24144;
assign w24146 = ~w24125 & ~w24131;
assign w24147 = ~w24145 & ~w24146;
assign w24148 = w24145 & w24146;
assign w24149 = ~w24132 & ~w24147;
assign w24150 = ~w24148 & w24149;
assign w24151 = w24119 & w24150;
assign w24152 = w24131 & ~w24138;
assign w24153 = ~w24131 & w24138;
assign w24154 = ~w24152 & ~w24153;
assign w24155 = w24125 & ~w24154;
assign w24156 = w24119 & w24138;
assign w24157 = ~w24119 & ~w24144;
assign w24158 = w24152 & w24157;
assign w24159 = w24138 & w24144;
assign w24160 = ~w24138 & ~w24144;
assign w24161 = ~w24159 & ~w24160;
assign w24162 = w24132 & ~w24161;
assign w24163 = ~w24125 & ~w24144;
assign w24164 = ~w24153 & ~w24156;
assign w24165 = w24163 & ~w24164;
assign w24166 = ~w24158 & ~w24162;
assign w24167 = ~w24165 & w24166;
assign w24168 = w24166 & w65551;
assign w24169 = ~w24144 & w24154;
assign w24170 = ~w24125 & ~w24138;
assign w24171 = w24154 & w63776;
assign w24172 = ~w24119 & w24171;
assign w24173 = w24131 & w24144;
assign w24174 = ~w24131 & ~w24144;
assign w24175 = ~w24173 & ~w24174;
assign w24176 = ~w24138 & ~w24175;
assign w24177 = (~w24125 & w24172) | (~w24125 & w65552) | (w24172 & w65552);
assign w24178 = ~w24168 & ~w24177;
assign w24179 = ~pi4282 & pi9040;
assign w24180 = ~pi4221 & ~pi9040;
assign w24181 = ~w24179 & ~w24180;
assign w24182 = pi1290 & ~w24181;
assign w24183 = ~pi1290 & w24181;
assign w24184 = ~w24182 & ~w24183;
assign w24185 = ~w24155 & w24184;
assign w24186 = ~w24178 & w24185;
assign w24187 = ~w24119 & ~w24152;
assign w24188 = (w24187 & ~w24149) | (w24187 & w63777) | (~w24149 & w63777);
assign w24189 = ~w24171 & w24188;
assign w24190 = w24167 & ~w24189;
assign w24191 = ~w24184 & ~w24190;
assign w24192 = ~w24119 & w24125;
assign w24193 = w24152 & w24184;
assign w24194 = w24161 & ~w24193;
assign w24195 = w24192 & ~w24194;
assign w24196 = ~w24151 & ~w24195;
assign w24197 = ~w24191 & w24196;
assign w24198 = (pi1313 & ~w24197) | (pi1313 & w65553) | (~w24197 & w65553);
assign w24199 = w24197 & w65554;
assign w24200 = ~w24198 & ~w24199;
assign w24201 = w23784 & w23800;
assign w24202 = ~w23761 & w24201;
assign w24203 = w23761 & ~w23822;
assign w24204 = (w23794 & w24203) | (w23794 & w65555) | (w24203 & w65555);
assign w24205 = ~w23781 & ~w23809;
assign w24206 = w23761 & ~w24205;
assign w24207 = (~w23794 & ~w23786) | (~w23794 & w65556) | (~w23786 & w65556);
assign w24208 = ~w23798 & w24207;
assign w24209 = ~w24206 & w24208;
assign w24210 = (w23755 & w24209) | (w23755 & w65557) | (w24209 & w65557);
assign w24211 = ~w23784 & w24093;
assign w24212 = w23810 & ~w23821;
assign w24213 = ~w23804 & ~w24212;
assign w24214 = ~w24211 & w24213;
assign w24215 = ~w23755 & ~w24214;
assign w24216 = w23784 & w23783;
assign w24217 = ~w23787 & ~w24216;
assign w24218 = w23794 & ~w24217;
assign w24219 = ~w24205 & w65558;
assign w24220 = ~w24202 & ~w24219;
assign w24221 = ~w24218 & w24220;
assign w24222 = ~w24094 & w24221;
assign w24223 = ~w24210 & w24222;
assign w24224 = ~w24215 & w24223;
assign w24225 = pi1327 & ~w24224;
assign w24226 = ~pi1327 & w24224;
assign w24227 = ~w24225 & ~w24226;
assign w24228 = w24125 & w24138;
assign w24229 = ~w24170 & ~w24228;
assign w24230 = ~w24119 & w24159;
assign w24231 = ~w24131 & w24161;
assign w24232 = (~w24231 & w63778) | (~w24231 & w63779) | (w63778 & w63779);
assign w24233 = (~w24229 & ~w24232) | (~w24229 & w65559) | (~w24232 & w65559);
assign w24234 = ~w24175 & w24229;
assign w24235 = ~w24233 & ~w24234;
assign w24236 = w24184 & ~w24235;
assign w24237 = ~w24132 & ~w24146;
assign w24238 = ~w24119 & ~w24237;
assign w24239 = w24232 & ~w24238;
assign w24240 = ~w24184 & ~w24234;
assign w24241 = w24239 & w24240;
assign w24242 = ~w24236 & ~w24241;
assign w24243 = pi1315 & ~w24242;
assign w24244 = ~pi1315 & w24242;
assign w24245 = ~w24243 & ~w24244;
assign w24246 = ~w23871 & w23925;
assign w24247 = w23914 & w24246;
assign w24248 = w23884 & w65560;
assign w24249 = w23882 & w23892;
assign w24250 = w23891 & ~w24249;
assign w24251 = w23879 & w23883;
assign w24252 = ~w23848 & ~w23897;
assign w24253 = w23855 & w23897;
assign w24254 = ~w24252 & ~w24253;
assign w24255 = w23871 & ~w24254;
assign w24256 = ~w23862 & ~w23871;
assign w24257 = ~w24252 & w24256;
assign w24258 = w24250 & ~w24251;
assign w24259 = ~w24257 & w24258;
assign w24260 = ~w24255 & w24259;
assign w24261 = w23861 & w23922;
assign w24262 = w23912 & w23921;
assign w24263 = ~w23891 & ~w24262;
assign w24264 = ~w24261 & w24263;
assign w24265 = ~w24260 & ~w24264;
assign w24266 = ~w24247 & ~w24248;
assign w24267 = ~w24265 & w24266;
assign w24268 = ~pi1321 & w24267;
assign w24269 = pi1321 & ~w24267;
assign w24270 = ~w24268 & ~w24269;
assign w24271 = ~w23556 & ~w23635;
assign w24272 = w23543 & ~w23622;
assign w24273 = ~w23638 & ~w24272;
assign w24274 = w23530 & ~w24273;
assign w24275 = w23556 & ~w23608;
assign w24276 = w23652 & w24275;
assign w24277 = ~w24274 & w24276;
assign w24278 = ~w24271 & ~w24277;
assign w24279 = ~w23556 & w24272;
assign w24280 = w23623 & ~w23656;
assign w24281 = w24275 & ~w24280;
assign w24282 = ~w23530 & ~w23574;
assign w24283 = ~w23642 & w24282;
assign w24284 = ~w23620 & w24283;
assign w24285 = ~w24279 & w24284;
assign w24286 = ~w24281 & w24285;
assign w24287 = ~w23567 & w23584;
assign w24288 = ~w23635 & w23655;
assign w24289 = ~w24287 & w24288;
assign w24290 = ~w24286 & ~w24289;
assign w24291 = ~w24290 & w65561;
assign w24292 = (pi1337 & w24290) | (pi1337 & w65562) | (w24290 & w65562);
assign w24293 = ~w24291 & ~w24292;
assign w24294 = ~w23755 & w23827;
assign w24295 = ~w23824 & ~w24095;
assign w24296 = ~w23755 & ~w24295;
assign w24297 = ~w23825 & ~w24296;
assign w24298 = (w23794 & w24297) | (w23794 & w65563) | (w24297 & w65563);
assign w24299 = w23774 & w23807;
assign w24300 = ~w23834 & ~w24296;
assign w24301 = ~w24299 & w24300;
assign w24302 = ~w23794 & ~w24301;
assign w24303 = w23801 & ~w23820;
assign w24304 = w23774 & w23795;
assign w24305 = ~w24216 & ~w24304;
assign w24306 = ~w24303 & w24305;
assign w24307 = w23755 & ~w24306;
assign w24308 = w23786 & ~w23820;
assign w24309 = ~w23768 & w23816;
assign w24310 = ~w24308 & w24309;
assign w24311 = w24295 & w24310;
assign w24312 = ~w24201 & ~w24294;
assign w24313 = ~w24311 & w24312;
assign w24314 = ~w24307 & w24313;
assign w24315 = ~w24298 & w24314;
assign w24316 = ~w24302 & w24315;
assign w24317 = pi1323 & ~w24316;
assign w24318 = ~pi1323 & w24316;
assign w24319 = ~w24317 & ~w24318;
assign w24320 = ~w23879 & w23903;
assign w24321 = ~w23918 & ~w24320;
assign w24322 = ~w23879 & w23882;
assign w24323 = ~w24248 & ~w24322;
assign w24324 = w23898 & ~w24323;
assign w24325 = (w24250 & w24321) | (w24250 & w65564) | (w24321 & w65564);
assign w24326 = ~w24324 & w24325;
assign w24327 = (~w23920 & ~w23922) | (~w23920 & w65565) | (~w23922 & w65565);
assign w24328 = w23871 & ~w24327;
assign w24329 = w23871 & w23907;
assign w24330 = ~w23891 & ~w24329;
assign w24331 = ~w23916 & w24330;
assign w24332 = ~w24328 & w24331;
assign w24333 = ~w24326 & ~w24332;
assign w24334 = ~w23883 & ~w23891;
assign w24335 = ~w23864 & w23879;
assign w24336 = ~w24334 & ~w24335;
assign w24337 = ~w23871 & w23921;
assign w24338 = ~w24336 & w24337;
assign w24339 = ~w24333 & ~w24338;
assign w24340 = ~pi1333 & w24339;
assign w24341 = pi1333 & ~w24339;
assign w24342 = ~w24340 & ~w24341;
assign w24343 = w23718 & w24044;
assign w24344 = w23706 & ~w24025;
assign w24345 = w23717 & ~w24044;
assign w24346 = ~w24344 & ~w24345;
assign w24347 = w23679 & ~w24346;
assign w24348 = ~w23679 & w23716;
assign w24349 = ~w23713 & ~w24348;
assign w24350 = w24034 & ~w24349;
assign w24351 = ~w23722 & ~w24064;
assign w24352 = w23736 & w24351;
assign w24353 = ~w23679 & ~w24352;
assign w24354 = ~w24343 & ~w24350;
assign w24355 = ~w24347 & w24354;
assign w24356 = ~w24353 & w24355;
assign w24357 = pi1348 & ~w24356;
assign w24358 = ~pi1348 & w24356;
assign w24359 = ~w24357 & ~w24358;
assign w24360 = ~pi4228 & pi9040;
assign w24361 = ~pi4698 & ~pi9040;
assign w24362 = ~w24360 & ~w24361;
assign w24363 = pi1271 & ~w24362;
assign w24364 = ~pi1271 & w24362;
assign w24365 = ~w24363 & ~w24364;
assign w24366 = ~pi4287 & pi9040;
assign w24367 = ~pi4228 & ~pi9040;
assign w24368 = ~w24366 & ~w24367;
assign w24369 = pi1309 & ~w24368;
assign w24370 = ~pi1309 & w24368;
assign w24371 = ~w24369 & ~w24370;
assign w24372 = ~pi4205 & pi9040;
assign w24373 = ~pi4404 & ~pi9040;
assign w24374 = ~w24372 & ~w24373;
assign w24375 = pi1307 & ~w24374;
assign w24376 = ~pi1307 & w24374;
assign w24377 = ~w24375 & ~w24376;
assign w24378 = ~w24371 & w24377;
assign w24379 = ~pi4309 & pi9040;
assign w24380 = ~pi4302 & ~pi9040;
assign w24381 = ~w24379 & ~w24380;
assign w24382 = pi1291 & ~w24381;
assign w24383 = ~pi1291 & w24381;
assign w24384 = ~w24382 & ~w24383;
assign w24385 = ~w24371 & w24384;
assign w24386 = ~w24377 & ~w24384;
assign w24387 = w24377 & w24384;
assign w24388 = ~w24386 & ~w24387;
assign w24389 = ~pi4213 & pi9040;
assign w24390 = ~pi4287 & ~pi9040;
assign w24391 = ~w24389 & ~w24390;
assign w24392 = pi1297 & ~w24391;
assign w24393 = ~pi1297 & w24391;
assign w24394 = ~w24392 & ~w24393;
assign w24395 = ~w24384 & ~w24394;
assign w24396 = ~w24385 & ~w24395;
assign w24397 = w24388 & w24396;
assign w24398 = ~pi4206 & pi9040;
assign w24399 = ~pi4310 & ~pi9040;
assign w24400 = ~w24398 & ~w24399;
assign w24401 = pi1277 & ~w24400;
assign w24402 = ~pi1277 & w24400;
assign w24403 = ~w24401 & ~w24402;
assign w24404 = (w24403 & w24397) | (w24403 & w63780) | (w24397 & w63780);
assign w24405 = w24371 & w24394;
assign w24406 = w24386 & w24405;
assign w24407 = ~w24386 & ~w24403;
assign w24408 = ~w24397 & w65566;
assign w24409 = ~w24404 & ~w24406;
assign w24410 = (w24365 & ~w24409) | (w24365 & w65567) | (~w24409 & w65567);
assign w24411 = ~w24384 & w24403;
assign w24412 = (w24371 & ~w24388) | (w24371 & w63781) | (~w24388 & w63781);
assign w24413 = ~w24394 & w24412;
assign w24414 = ~w24371 & ~w24394;
assign w24415 = w24388 & w63782;
assign w24416 = ~w24413 & ~w24415;
assign w24417 = ~w24371 & w24388;
assign w24418 = ~w24412 & ~w24417;
assign w24419 = w24394 & w24418;
assign w24420 = w24416 & ~w24419;
assign w24421 = ~w24365 & ~w24420;
assign w24422 = ~w24386 & ~w24394;
assign w24423 = ~w24377 & w24394;
assign w24424 = ~w24422 & ~w24423;
assign w24425 = ~w24371 & w24403;
assign w24426 = w24424 & w24425;
assign w24427 = ~w24410 & ~w24426;
assign w24428 = ~w24421 & w24427;
assign w24429 = pi1330 & ~w24428;
assign w24430 = ~pi1330 & w24428;
assign w24431 = ~w24429 & ~w24430;
assign w24432 = ~w24385 & w24403;
assign w24433 = w24419 & w24432;
assign w24434 = ~w24377 & w24403;
assign w24435 = ~w24387 & ~w24434;
assign w24436 = w24384 & w24394;
assign w24437 = ~w24378 & ~w24395;
assign w24438 = ~w24436 & w24437;
assign w24439 = w24435 & w24438;
assign w24440 = (~w24394 & w24417) | (~w24394 & w65568) | (w24417 & w65568);
assign w24441 = ~w24418 & w24440;
assign w24442 = w24365 & ~w24439;
assign w24443 = ~w24441 & w24442;
assign w24444 = w24386 & w24414;
assign w24445 = (~w24385 & ~w24388) | (~w24385 & w65569) | (~w24388 & w65569);
assign w24446 = ~w24403 & ~w24423;
assign w24447 = w24445 & w24446;
assign w24448 = w24403 & ~w24445;
assign w24449 = ~w24417 & w24448;
assign w24450 = ~w24365 & ~w24444;
assign w24451 = ~w24447 & w24450;
assign w24452 = ~w24449 & w24451;
assign w24453 = ~w24443 & ~w24452;
assign w24454 = w24394 & ~w24403;
assign w24455 = w24385 & w24454;
assign w24456 = ~w24433 & ~w24455;
assign w24457 = ~w24453 & w24456;
assign w24458 = pi1326 & ~w24457;
assign w24459 = ~pi1326 & w24457;
assign w24460 = ~w24458 & ~w24459;
assign w24461 = ~w24388 & w24414;
assign w24462 = ~w24397 & ~w24461;
assign w24463 = ~w24403 & ~w24462;
assign w24464 = w24403 & ~w24414;
assign w24465 = ~w24388 & ~w24464;
assign w24466 = (w24465 & w24462) | (w24465 & w63389) | (w24462 & w63389);
assign w24467 = ~w24386 & w24394;
assign w24468 = w24432 & w24467;
assign w24469 = ~w24415 & ~w24468;
assign w24470 = w24385 & w24394;
assign w24471 = ~w24411 & ~w24470;
assign w24472 = ~w24466 & w63783;
assign w24473 = (~w24365 & w24472) | (~w24365 & w65570) | (w24472 & w65570);
assign w24474 = w24436 & w24447;
assign w24475 = (w24365 & w24466) | (w24365 & w65571) | (w24466 & w65571);
assign w24476 = ~w24416 & w24448;
assign w24477 = ~w24474 & ~w24476;
assign w24478 = ~w24475 & w24477;
assign w24479 = w24478 & w65572;
assign w24480 = (~pi1332 & ~w24478) | (~pi1332 & w65573) | (~w24478 & w65573);
assign w24481 = ~w24479 & ~w24480;
assign w24482 = w24387 & w24472;
assign w24483 = ~w24371 & ~w24462;
assign w24484 = w24371 & ~w24377;
assign w24485 = ~w24436 & ~w24484;
assign w24486 = ~w24403 & ~w24485;
assign w24487 = ~w24371 & ~w24384;
assign w24488 = ~w24403 & ~w24487;
assign w24489 = ~w24387 & w24405;
assign w24490 = ~w24485 & ~w24489;
assign w24491 = ~w24488 & ~w24490;
assign w24492 = ~w24486 & ~w24491;
assign w24493 = ~w24483 & ~w24492;
assign w24494 = w24454 & w24484;
assign w24495 = (w24411 & w24422) | (w24411 & w65574) | (w24422 & w65574);
assign w24496 = ~w24422 & w24486;
assign w24497 = ~w24489 & ~w24495;
assign w24498 = ~w24496 & w24497;
assign w24499 = (w24365 & w24476) | (w24365 & w65575) | (w24476 & w65575);
assign w24500 = (~w24494 & w24493) | (~w24494 & w63784) | (w24493 & w63784);
assign w24501 = ~w24482 & w24500;
assign w24502 = (~pi1342 & ~w24501) | (~pi1342 & w65576) | (~w24501 & w65576);
assign w24503 = w24501 & w65577;
assign w24504 = ~w24502 & ~w24503;
assign w24505 = ~pi4316 & pi9040;
assign w24506 = ~pi4288 & ~pi9040;
assign w24507 = ~w24505 & ~w24506;
assign w24508 = pi1301 & ~w24507;
assign w24509 = ~pi1301 & w24507;
assign w24510 = ~w24508 & ~w24509;
assign w24511 = ~pi4293 & pi9040;
assign w24512 = ~pi4282 & ~pi9040;
assign w24513 = ~w24511 & ~w24512;
assign w24514 = pi1289 & ~w24513;
assign w24515 = ~pi1289 & w24513;
assign w24516 = ~w24514 & ~w24515;
assign w24517 = ~pi4593 & pi9040;
assign w24518 = ~pi4384 & ~pi9040;
assign w24519 = ~w24517 & ~w24518;
assign w24520 = pi1306 & ~w24519;
assign w24521 = ~pi1306 & w24519;
assign w24522 = ~w24520 & ~w24521;
assign w24523 = ~w24516 & ~w24522;
assign w24524 = w24516 & w24522;
assign w24525 = ~pi4221 & pi9040;
assign w24526 = ~pi4484 & ~pi9040;
assign w24527 = ~w24525 & ~w24526;
assign w24528 = pi1310 & ~w24527;
assign w24529 = ~pi1310 & w24527;
assign w24530 = ~w24528 & ~w24529;
assign w24531 = ~pi4384 & pi9040;
assign w24532 = ~pi4374 & ~pi9040;
assign w24533 = ~w24531 & ~w24532;
assign w24534 = pi1311 & ~w24533;
assign w24535 = ~pi1311 & w24533;
assign w24536 = ~w24534 & ~w24535;
assign w24537 = ~w24530 & w24536;
assign w24538 = ~w24524 & w24537;
assign w24539 = ~w24523 & w24538;
assign w24540 = ~w24510 & w24539;
assign w24541 = ~w24523 & ~w24524;
assign w24542 = ~w24530 & ~w24536;
assign w24543 = ~w24522 & w24536;
assign w24544 = ~w24542 & ~w24543;
assign w24545 = w24541 & ~w24544;
assign w24546 = ~w24510 & ~w24545;
assign w24547 = w24530 & ~w24536;
assign w24548 = ~w24516 & w24522;
assign w24549 = ~w24547 & ~w24548;
assign w24550 = ~w24536 & w24541;
assign w24551 = ~w24549 & ~w24550;
assign w24552 = w24546 & ~w24551;
assign w24553 = w24523 & ~w24530;
assign w24554 = w24522 & w24542;
assign w24555 = w24516 & w24530;
assign w24556 = w24536 & w24555;
assign w24557 = (w24510 & ~w24542) | (w24510 & w64404) | (~w24542 & w64404);
assign w24558 = ~w24556 & w24557;
assign w24559 = ~w24553 & w24558;
assign w24560 = ~pi4284 & pi9040;
assign w24561 = ~pi4304 & ~pi9040;
assign w24562 = ~w24560 & ~w24561;
assign w24563 = pi1279 & ~w24562;
assign w24564 = ~pi1279 & w24562;
assign w24565 = ~w24563 & ~w24564;
assign w24566 = ~w24552 & w65578;
assign w24567 = w24522 & w24530;
assign w24568 = ~w24516 & ~w24567;
assign w24569 = w24558 & ~w24568;
assign w24570 = ~w24542 & ~w24556;
assign w24571 = w24546 & ~w24570;
assign w24572 = ~w24516 & w24530;
assign w24573 = ~w24547 & ~w24572;
assign w24574 = ~w24551 & ~w24573;
assign w24575 = ~w24569 & ~w24571;
assign w24576 = (w24565 & ~w24575) | (w24565 & w65579) | (~w24575 & w65579);
assign w24577 = w24547 & w24548;
assign w24578 = w24523 & w24537;
assign w24579 = ~w24577 & ~w24578;
assign w24580 = w24510 & ~w24579;
assign w24581 = ~w24540 & ~w24580;
assign w24582 = ~w24566 & w24581;
assign w24583 = ~w24576 & w24582;
assign w24584 = pi1336 & ~w24583;
assign w24585 = ~pi1336 & w24583;
assign w24586 = ~w24584 & ~w24585;
assign w24587 = w24542 & w24559;
assign w24588 = ~w24522 & ~w24536;
assign w24589 = ~w24555 & ~w24588;
assign w24590 = ~w24538 & w24589;
assign w24591 = w24551 & w24590;
assign w24592 = (~w24578 & ~w24551) | (~w24578 & w65580) | (~w24551 & w65580);
assign w24593 = ~w24522 & w24555;
assign w24594 = w24565 & ~w24593;
assign w24595 = ~w24590 & w24594;
assign w24596 = w24592 & ~w24595;
assign w24597 = w24510 & ~w24596;
assign w24598 = w24516 & ~w24536;
assign w24599 = w24522 & w24598;
assign w24600 = ~w24554 & ~w24593;
assign w24601 = (~w24599 & w24600) | (~w24599 & w63785) | (w24600 & w63785);
assign w24602 = (w24565 & w24591) | (w24565 & w65581) | (w24591 & w65581);
assign w24603 = ~w24522 & ~w24530;
assign w24604 = ~w24510 & ~w24603;
assign w24605 = ~w24523 & ~w24537;
assign w24606 = (~w24543 & w24605) | (~w24543 & w63786) | (w24605 & w63786);
assign w24607 = w24604 & ~w24606;
assign w24608 = w24522 & w24555;
assign w24609 = ~w24536 & w24608;
assign w24610 = w24510 & ~w24548;
assign w24611 = ~w24604 & ~w24610;
assign w24612 = ~w24536 & ~w24611;
assign w24613 = w24524 & ~w24530;
assign w24614 = (w24536 & ~w24524) | (w24536 & w65582) | (~w24524 & w65582);
assign w24615 = ~w24565 & ~w24614;
assign w24616 = ~w24612 & w24615;
assign w24617 = ~w24607 & ~w24609;
assign w24618 = ~w24616 & w24617;
assign w24619 = ~w24587 & w24618;
assign w24620 = ~w24602 & w24619;
assign w24621 = (pi1328 & ~w24620) | (pi1328 & w65583) | (~w24620 & w65583);
assign w24622 = w24620 & w65584;
assign w24623 = ~w24621 & ~w24622;
assign w24624 = w23883 & w23893;
assign w24625 = ~w23871 & w23922;
assign w24626 = ~w24329 & ~w24625;
assign w24627 = ~w23861 & ~w24626;
assign w24628 = (w24256 & w24320) | (w24256 & w65585) | (w24320 & w65585);
assign w24629 = w23906 & ~w24255;
assign w24630 = w24321 & ~w24629;
assign w24631 = w23891 & ~w24628;
assign w24632 = ~w24630 & w24631;
assign w24633 = ~w23872 & ~w23881;
assign w24634 = w23883 & ~w24633;
assign w24635 = ~w23893 & ~w24251;
assign w24636 = ~w24322 & w24635;
assign w24637 = ~w24634 & w24636;
assign w24638 = w24330 & w24637;
assign w24639 = ~w24632 & ~w24638;
assign w24640 = ~w23913 & ~w24624;
assign w24641 = ~w24627 & w24640;
assign w24642 = (pi1344 & w24639) | (pi1344 & w65586) | (w24639 & w65586);
assign w24643 = ~w24639 & w65587;
assign w24644 = ~w24642 & ~w24643;
assign w24645 = w23941 & w23979;
assign w24646 = ~w23996 & ~w24645;
assign w24647 = w23971 & ~w24646;
assign w24648 = (w24008 & w63787) | (w24008 & w63788) | (w63787 & w63788);
assign w24649 = w23971 & ~w24003;
assign w24650 = (~w23997 & ~w24007) | (~w23997 & w65588) | (~w24007 & w65588);
assign w24651 = (w23978 & w24648) | (w23978 & w65589) | (w24648 & w65589);
assign w24652 = ~w23954 & ~w23971;
assign w24653 = w23989 & w24652;
assign w24654 = w23989 & ~w24005;
assign w24655 = w24649 & ~w24654;
assign w24656 = w23947 & ~w23971;
assign w24657 = w24005 & w24656;
assign w24658 = ~w24653 & ~w24657;
assign w24659 = ~w23988 & w24658;
assign w24660 = ~w24655 & w24659;
assign w24661 = ~w23978 & ~w24660;
assign w24662 = w23982 & ~w23992;
assign w24663 = w23971 & ~w23986;
assign w24664 = ~w24000 & ~w24663;
assign w24665 = ~w24662 & w24664;
assign w24666 = ~w24661 & ~w24665;
assign w24667 = ~w24651 & w24666;
assign w24668 = ~pi1354 & w24667;
assign w24669 = pi1354 & ~w24667;
assign w24670 = ~w24668 & ~w24669;
assign w24671 = w24119 & w24171;
assign w24672 = ~w24153 & ~w24170;
assign w24673 = ~w24161 & ~w24672;
assign w24674 = ~w24155 & ~w24673;
assign w24675 = ~w24119 & ~w24674;
assign w24676 = w24173 & w24229;
assign w24677 = ~w24154 & w63789;
assign w24678 = ~w24676 & ~w24677;
assign w24679 = w24145 & w24192;
assign w24680 = ~w24675 & w24678;
assign w24681 = (w24184 & ~w24680) | (w24184 & w63790) | (~w24680 & w63790);
assign w24682 = ~w24153 & w24237;
assign w24683 = (w24119 & w24175) | (w24119 & w63791) | (w24175 & w63791);
assign w24684 = ~w24682 & w24683;
assign w24685 = ~w24677 & ~w24684;
assign w24686 = ~w24684 & w24678;
assign w24687 = ~w24239 & ~w24686;
assign w24688 = w24119 & ~w24169;
assign w24689 = w24678 & w24688;
assign w24690 = ~w24148 & ~w24172;
assign w24691 = ~w24689 & w24690;
assign w24692 = ~w24184 & ~w24691;
assign w24693 = ~w24681 & ~w24687;
assign w24694 = w24693 & w65590;
assign w24695 = (~pi1331 & ~w24693) | (~pi1331 & w65591) | (~w24693 & w65591);
assign w24696 = ~w24694 & ~w24695;
assign w24697 = w24523 & w24547;
assign w24698 = w24510 & ~w24697;
assign w24699 = ~w24608 & w24698;
assign w24700 = ~w24591 & w63792;
assign w24701 = w24543 & w24572;
assign w24702 = w24547 & w24565;
assign w24703 = ~w24701 & ~w24702;
assign w24704 = ~w24510 & ~w24703;
assign w24705 = ~w24510 & w24613;
assign w24706 = w24516 & w24542;
assign w24707 = (~w24510 & ~w24555) | (~w24510 & w65592) | (~w24555 & w65592);
assign w24708 = ~w24706 & w24707;
assign w24709 = ~w24699 & ~w24708;
assign w24710 = ~w24554 & ~w24565;
assign w24711 = ~w24705 & w24710;
assign w24712 = ~w24709 & w24711;
assign w24713 = w24592 & w24712;
assign w24714 = ~w24536 & w24553;
assign w24715 = ~w24593 & ~w24714;
assign w24716 = w24510 & ~w24715;
assign w24717 = ~w24539 & w24565;
assign w24718 = ~w24716 & w24717;
assign w24719 = ~w24713 & ~w24718;
assign w24720 = (~w24704 & w24700) | (~w24704 & w65593) | (w24700 & w65593);
assign w24721 = ~w24719 & w65594;
assign w24722 = (~pi1325 & w24719) | (~pi1325 & w65595) | (w24719 & w65595);
assign w24723 = ~w24721 & ~w24722;
assign w24724 = w23941 & ~w23964;
assign w24725 = w23978 & ~w24724;
assign w24726 = (~w24008 & w63793) | (~w24008 & w63794) | (w63793 & w63794);
assign w24727 = w24725 & ~w24726;
assign w24728 = w23984 & w23995;
assign w24729 = ~w23978 & ~w24728;
assign w24730 = (~w24008 & w65596) | (~w24008 & w65597) | (w65596 & w65597);
assign w24731 = ~w24727 & ~w24730;
assign w24732 = w23983 & w65598;
assign w24733 = ~w23947 & w23978;
assign w24734 = w23983 & w24733;
assign w24735 = w23971 & ~w24014;
assign w24736 = ~w24734 & w24735;
assign w24737 = ~w24732 & w24736;
assign w24738 = (~w24003 & w24007) | (~w24003 & w65599) | (w24007 & w65599);
assign w24739 = ~w23960 & w23978;
assign w24740 = w23995 & ~w24739;
assign w24741 = ~w23971 & ~w24740;
assign w24742 = ~w24738 & w24741;
assign w24743 = ~w24737 & ~w24742;
assign w24744 = ~w24731 & w65600;
assign w24745 = (pi1349 & w24731) | (pi1349 & w65601) | (w24731 & w65601);
assign w24746 = ~w24744 & ~w24745;
assign w24747 = w23971 & w24016;
assign w24748 = w23948 & ~w23978;
assign w24749 = ~w24656 & ~w24748;
assign w24750 = w23961 & ~w24749;
assign w24751 = ~w24725 & w24750;
assign w24752 = ~w23984 & w24663;
assign w24753 = ~w24724 & w24752;
assign w24754 = ~w23984 & ~w23987;
assign w24755 = w23954 & ~w23971;
assign w24756 = ~w24754 & w24755;
assign w24757 = ~w23947 & ~w23995;
assign w24758 = ~w24006 & w24757;
assign w24759 = w23978 & ~w24732;
assign w24760 = ~w24758 & w24759;
assign w24761 = ~w24756 & w24760;
assign w24762 = ~w24753 & w24761;
assign w24763 = ~w23941 & ~w24656;
assign w24764 = w23962 & ~w24763;
assign w24765 = ~w23978 & ~w23985;
assign w24766 = ~w24653 & w24765;
assign w24767 = ~w23997 & ~w24764;
assign w24768 = w24766 & w24767;
assign w24769 = ~w24647 & w24768;
assign w24770 = ~w24762 & ~w24769;
assign w24771 = ~w24747 & ~w24751;
assign w24772 = ~w24770 & w24771;
assign w24773 = pi1338 & ~w24772;
assign w24774 = ~pi1338 & w24772;
assign w24775 = ~w24773 & ~w24774;
assign w24776 = ~w24154 & w24163;
assign w24777 = w24238 & ~w24776;
assign w24778 = w24173 & w24228;
assign w24779 = ~w24163 & w24237;
assign w24780 = w24161 & w24779;
assign w24781 = ~w24132 & w24156;
assign w24782 = ~w24673 & w24781;
assign w24783 = ~w24184 & ~w24778;
assign w24784 = ~w24777 & w24783;
assign w24785 = ~w24780 & ~w24782;
assign w24786 = w24784 & w24785;
assign w24787 = w24229 & w24779;
assign w24788 = (~w24119 & w24787) | (~w24119 & w65602) | (w24787 & w65602);
assign w24789 = w24184 & w24685;
assign w24790 = ~w24788 & w24789;
assign w24791 = ~w24786 & ~w24790;
assign w24792 = w24239 & ~w24788;
assign w24793 = ~w24146 & w24161;
assign w24794 = ~w24792 & w24793;
assign w24795 = (pi1324 & w24791) | (pi1324 & w65603) | (w24791 & w65603);
assign w24796 = ~w24791 & w65604;
assign w24797 = ~w24795 & ~w24796;
assign w24798 = ~w24572 & ~w24598;
assign w24799 = ~w24593 & ~w24798;
assign w24800 = ~w24510 & ~w24799;
assign w24801 = ~w24567 & ~w24706;
assign w24802 = w24699 & ~w24801;
assign w24803 = w24543 & ~w24572;
assign w24804 = ~w24565 & ~w24803;
assign w24805 = ~w24800 & w24804;
assign w24806 = ~w24802 & w24805;
assign w24807 = w24510 & ~w24572;
assign w24808 = ~w24549 & w24807;
assign w24809 = w24565 & ~w24701;
assign w24810 = ~w24609 & w24809;
assign w24811 = ~w24705 & ~w24808;
assign w24812 = w24810 & w24811;
assign w24813 = w24543 & w24569;
assign w24814 = ~w24715 & w24798;
assign w24815 = ~w24510 & ~w24577;
assign w24816 = ~w24814 & w24815;
assign w24817 = ~w24698 & ~w24816;
assign w24818 = (~w24813 & w24806) | (~w24813 & w65605) | (w24806 & w65605);
assign w24819 = ~w24817 & w24818;
assign w24820 = pi1347 & ~w24819;
assign w24821 = ~pi1347 & w24819;
assign w24822 = ~w24820 & ~w24821;
assign w24823 = ~pi4805 & pi9040;
assign w24824 = ~pi4490 & ~pi9040;
assign w24825 = ~w24823 & ~w24824;
assign w24826 = pi1367 & ~w24825;
assign w24827 = ~pi1367 & w24825;
assign w24828 = ~w24826 & ~w24827;
assign w24829 = ~pi4521 & pi9040;
assign w24830 = ~pi4735 & ~pi9040;
assign w24831 = ~w24829 & ~w24830;
assign w24832 = pi1341 & ~w24831;
assign w24833 = ~pi1341 & w24831;
assign w24834 = ~w24832 & ~w24833;
assign w24835 = ~w24828 & w24834;
assign w24836 = ~pi4477 & pi9040;
assign w24837 = ~pi4482 & ~pi9040;
assign w24838 = ~w24836 & ~w24837;
assign w24839 = pi1346 & ~w24838;
assign w24840 = ~pi1346 & w24838;
assign w24841 = ~w24839 & ~w24840;
assign w24842 = w24835 & w24841;
assign w24843 = w24828 & w24834;
assign w24844 = ~pi4409 & pi9040;
assign w24845 = ~pi4402 & ~pi9040;
assign w24846 = ~w24844 & ~w24845;
assign w24847 = pi1335 & ~w24846;
assign w24848 = ~pi1335 & w24846;
assign w24849 = ~w24847 & ~w24848;
assign w24850 = ~w24843 & ~w24849;
assign w24851 = ~pi4678 & pi9040;
assign w24852 = ~pi4553 & ~pi9040;
assign w24853 = ~w24851 & ~w24852;
assign w24854 = pi1373 & ~w24853;
assign w24855 = ~pi1373 & w24853;
assign w24856 = ~w24854 & ~w24855;
assign w24857 = w24828 & w24856;
assign w24858 = ~w24828 & ~w24856;
assign w24859 = ~w24857 & ~w24858;
assign w24860 = w24850 & ~w24859;
assign w24861 = w24842 & w24860;
assign w24862 = ~pi4482 & pi9040;
assign w24863 = ~pi4578 & ~pi9040;
assign w24864 = ~w24862 & ~w24863;
assign w24865 = pi1371 & ~w24864;
assign w24866 = ~pi1371 & w24864;
assign w24867 = ~w24865 & ~w24866;
assign w24868 = ~w24834 & w24849;
assign w24869 = ~w24841 & w24868;
assign w24870 = w24868 & w63795;
assign w24871 = w24849 & ~w24870;
assign w24872 = ~w24834 & w24841;
assign w24873 = w24856 & w24872;
assign w24874 = w24872 & w24876;
assign w24875 = w24871 & ~w24874;
assign w24876 = ~w24828 & w24856;
assign w24877 = ~w24841 & w24876;
assign w24878 = w24850 & ~w24877;
assign w24879 = ~w24875 & ~w24878;
assign w24880 = ~w24834 & ~w24856;
assign w24881 = (w24849 & w24859) | (w24849 & w65606) | (w24859 & w65606);
assign w24882 = ~w24843 & w24856;
assign w24883 = w24841 & ~w24882;
assign w24884 = ~w24881 & w24883;
assign w24885 = ~w24879 & ~w24884;
assign w24886 = ~w24867 & ~w24885;
assign w24887 = w24841 & ~w24856;
assign w24888 = ~w24835 & ~w24887;
assign w24889 = w24834 & ~w24841;
assign w24890 = w24856 & w24889;
assign w24891 = w24828 & w24880;
assign w24892 = ~w24890 & ~w24891;
assign w24893 = ~w24888 & ~w24892;
assign w24894 = ~w24834 & ~w24841;
assign w24895 = ~w24859 & w24894;
assign w24896 = (w24849 & w24893) | (w24849 & w65607) | (w24893 & w65607);
assign w24897 = w24857 & w24889;
assign w24898 = ~w24849 & ~w24897;
assign w24899 = ~w24841 & w24880;
assign w24900 = ~w24873 & ~w24899;
assign w24901 = w24898 & w24900;
assign w24902 = ~w24842 & ~w24888;
assign w24903 = w24849 & ~w24902;
assign w24904 = ~w24841 & w24843;
assign w24905 = ~w24842 & ~w24904;
assign w24906 = w24856 & ~w24905;
assign w24907 = w24903 & ~w24906;
assign w24908 = w24867 & ~w24901;
assign w24909 = ~w24907 & w24908;
assign w24910 = ~w24861 & ~w24896;
assign w24911 = ~w24909 & w24910;
assign w24912 = ~w24886 & w24911;
assign w24913 = pi1384 & w24912;
assign w24914 = ~pi1384 & ~w24912;
assign w24915 = ~w24913 & ~w24914;
assign w24916 = ~pi4603 & pi9040;
assign w24917 = ~pi4479 & ~pi9040;
assign w24918 = ~w24916 & ~w24917;
assign w24919 = pi1346 & ~w24918;
assign w24920 = ~pi1346 & w24918;
assign w24921 = ~w24919 & ~w24920;
assign w24922 = ~pi4561 & pi9040;
assign w24923 = ~pi4678 & ~pi9040;
assign w24924 = ~w24922 & ~w24923;
assign w24925 = pi1345 & ~w24924;
assign w24926 = ~pi1345 & w24924;
assign w24927 = ~w24925 & ~w24926;
assign w24928 = ~pi4735 & pi9040;
assign w24929 = ~pi4409 & ~pi9040;
assign w24930 = ~w24928 & ~w24929;
assign w24931 = pi1341 & ~w24930;
assign w24932 = ~pi1341 & w24930;
assign w24933 = ~w24931 & ~w24932;
assign w24934 = ~pi4483 & pi9040;
assign w24935 = ~pi4805 & ~pi9040;
assign w24936 = ~w24934 & ~w24935;
assign w24937 = pi1358 & ~w24936;
assign w24938 = ~pi1358 & w24936;
assign w24939 = ~w24937 & ~w24938;
assign w24940 = ~w24933 & ~w24939;
assign w24941 = ~pi4401 & pi9040;
assign w24942 = ~pi4730 & ~pi9040;
assign w24943 = ~w24941 & ~w24942;
assign w24944 = pi1363 & ~w24943;
assign w24945 = ~pi1363 & w24943;
assign w24946 = ~w24944 & ~w24945;
assign w24947 = w24940 & w24946;
assign w24948 = ~w24927 & w24947;
assign w24949 = ~w24921 & ~w24948;
assign w24950 = ~w24927 & w24946;
assign w24951 = w24927 & ~w24946;
assign w24952 = ~w24950 & ~w24951;
assign w24953 = ~pi4507 & pi9040;
assign w24954 = ~pi4561 & ~pi9040;
assign w24955 = ~w24953 & ~w24954;
assign w24956 = pi1370 & ~w24955;
assign w24957 = ~pi1370 & w24955;
assign w24958 = ~w24956 & ~w24957;
assign w24959 = ~w24939 & w24958;
assign w24960 = w24933 & ~w24959;
assign w24961 = w24952 & w24960;
assign w24962 = w24940 & w24951;
assign w24963 = ~w24933 & w24946;
assign w24964 = w24939 & w24963;
assign w24965 = ~w24962 & ~w24964;
assign w24966 = ~w24958 & ~w24965;
assign w24967 = w24933 & ~w24939;
assign w24968 = w24950 & w24967;
assign w24969 = w24958 & w24968;
assign w24970 = ~w24961 & ~w24969;
assign w24971 = w24949 & w24970;
assign w24972 = ~w24966 & w24971;
assign w24973 = w24946 & w24958;
assign w24974 = w24927 & w24939;
assign w24975 = w24933 & w24939;
assign w24976 = ~w24927 & ~w24975;
assign w24977 = ~w24974 & ~w24976;
assign w24978 = ~w24976 & w65608;
assign w24979 = w24927 & ~w24967;
assign w24980 = w24933 & ~w24946;
assign w24981 = ~w24963 & ~w24980;
assign w24982 = ~w24979 & w24981;
assign w24983 = w24940 & w24982;
assign w24984 = w24951 & w24967;
assign w24985 = ~w24983 & ~w24984;
assign w24986 = ~w24946 & w24975;
assign w24987 = ~w24968 & ~w24986;
assign w24988 = ~w24958 & ~w24987;
assign w24989 = w24921 & ~w24978;
assign w24990 = ~w24988 & w24989;
assign w24991 = w24985 & w24990;
assign w24992 = ~w24972 & ~w24991;
assign w24993 = ~w24940 & ~w24975;
assign w24994 = w24951 & w24993;
assign w24995 = ~w24947 & ~w24994;
assign w24996 = ~w24983 & w24995;
assign w24997 = w24958 & ~w24996;
assign w24998 = w24939 & ~w24958;
assign w24999 = w24952 & w24998;
assign w25000 = ~w24997 & ~w24999;
assign w25001 = ~w24992 & w25000;
assign w25002 = ~pi1377 & w25001;
assign w25003 = pi1377 & ~w25001;
assign w25004 = ~w25002 & ~w25003;
assign w25005 = ~w24927 & ~w24940;
assign w25006 = w24981 & w25005;
assign w25007 = ~w24962 & ~w25006;
assign w25008 = ~w24946 & ~w25007;
assign w25009 = ~w24958 & ~w24993;
assign w25010 = ~w24959 & ~w24974;
assign w25011 = w24980 & ~w25010;
assign w25012 = ~w25009 & ~w25011;
assign w25013 = w24958 & ~w24967;
assign w25014 = w24927 & w24946;
assign w25015 = ~w25013 & w25014;
assign w25016 = w24949 & ~w25015;
assign w25017 = w25012 & w25016;
assign w25018 = ~w25008 & w25017;
assign w25019 = w24939 & w24973;
assign w25020 = ~w24985 & w25012;
assign w25021 = w24979 & ~w24995;
assign w25022 = ~w24927 & ~w24987;
assign w25023 = w24921 & ~w25019;
assign w25024 = ~w25022 & w25023;
assign w25025 = ~w25021 & w25024;
assign w25026 = ~w25020 & w25025;
assign w25027 = ~w25018 & ~w25026;
assign w25028 = ~pi1380 & w25027;
assign w25029 = pi1380 & ~w25027;
assign w25030 = ~w25028 & ~w25029;
assign w25031 = ~pi4485 & pi9040;
assign w25032 = ~pi4852 & ~pi9040;
assign w25033 = ~w25031 & ~w25032;
assign w25034 = pi1374 & ~w25033;
assign w25035 = ~pi1374 & w25033;
assign w25036 = ~w25034 & ~w25035;
assign w25037 = ~pi4393 & pi9040;
assign w25038 = ~pi4509 & ~pi9040;
assign w25039 = ~w25037 & ~w25038;
assign w25040 = pi1371 & ~w25039;
assign w25041 = ~pi1371 & w25039;
assign w25042 = ~w25040 & ~w25041;
assign w25043 = w25036 & w25042;
assign w25044 = ~pi4492 & pi9040;
assign w25045 = ~pi4510 & ~pi9040;
assign w25046 = ~w25044 & ~w25045;
assign w25047 = pi1355 & ~w25046;
assign w25048 = ~pi1355 & w25046;
assign w25049 = ~w25047 & ~w25048;
assign w25050 = ~w25043 & w25049;
assign w25051 = ~pi4650 & pi9040;
assign w25052 = ~pi4403 & ~pi9040;
assign w25053 = ~w25051 & ~w25052;
assign w25054 = pi1367 & ~w25053;
assign w25055 = ~pi1367 & w25053;
assign w25056 = ~w25054 & ~w25055;
assign w25057 = ~pi4718 & pi9040;
assign w25058 = ~pi4394 & ~pi9040;
assign w25059 = ~w25057 & ~w25058;
assign w25060 = pi1339 & ~w25059;
assign w25061 = ~pi1339 & w25059;
assign w25062 = ~w25060 & ~w25061;
assign w25063 = w25056 & ~w25062;
assign w25064 = w25042 & ~w25049;
assign w25065 = w25063 & ~w25064;
assign w25066 = ~w25050 & w25065;
assign w25067 = ~w25049 & ~w25056;
assign w25068 = w25042 & w25062;
assign w25069 = w25067 & w25068;
assign w25070 = ~w25066 & ~w25069;
assign w25071 = ~w25049 & ~w25062;
assign w25072 = w25056 & ~w25071;
assign w25073 = w25064 & w25072;
assign w25074 = w25049 & w25062;
assign w25075 = w25056 & w25074;
assign w25076 = w25074 & w65609;
assign w25077 = ~w25073 & ~w25076;
assign w25078 = (w25036 & w25073) | (w25036 & w65610) | (w25073 & w65610);
assign w25079 = w25070 & ~w25078;
assign w25080 = ~pi4591 & pi9040;
assign w25081 = ~pi4396 & ~pi9040;
assign w25082 = ~w25080 & ~w25081;
assign w25083 = pi1356 & ~w25082;
assign w25084 = ~pi1356 & w25082;
assign w25085 = ~w25083 & ~w25084;
assign w25086 = ~w25079 & ~w25085;
assign w25087 = ~w25042 & ~w25062;
assign w25088 = ~w25068 & ~w25087;
assign w25089 = ~w25072 & ~w25088;
assign w25090 = ~w25085 & ~w25089;
assign w25091 = w25036 & ~w25042;
assign w25092 = ~w25074 & w25091;
assign w25093 = ~w25071 & w25092;
assign w25094 = w25043 & w25067;
assign w25095 = ~w25036 & w25042;
assign w25096 = w25056 & w25095;
assign w25097 = ~w25056 & w25062;
assign w25098 = ~w25095 & w25097;
assign w25099 = w25049 & ~w25056;
assign w25100 = w25042 & ~w25099;
assign w25101 = ~w25042 & w25049;
assign w25102 = ~w25100 & ~w25101;
assign w25103 = ~w25056 & ~w25068;
assign w25104 = ~w25102 & w25103;
assign w25105 = ~w25096 & ~w25098;
assign w25106 = (w25085 & w25104) | (w25085 & w65611) | (w25104 & w65611);
assign w25107 = ~w25049 & w25063;
assign w25108 = ~w25063 & ~w25097;
assign w25109 = w25042 & w25108;
assign w25110 = ~w25042 & ~w25108;
assign w25111 = ~w25109 & ~w25110;
assign w25112 = w25074 & ~w25111;
assign w25113 = ~w25085 & ~w25097;
assign w25114 = w25102 & w25113;
assign w25115 = ~w25107 & ~w25114;
assign w25116 = ~w25112 & w25115;
assign w25117 = ~w25036 & ~w25116;
assign w25118 = (~w25094 & w25090) | (~w25094 & w65612) | (w25090 & w65612);
assign w25119 = ~w25106 & w25118;
assign w25120 = ~w25086 & w25119;
assign w25121 = ~w25117 & w25120;
assign w25122 = ~pi1382 & ~w25121;
assign w25123 = pi1382 & w25121;
assign w25124 = ~w25122 & ~w25123;
assign w25125 = ~pi4615 & pi9040;
assign w25126 = ~pi4400 & ~pi9040;
assign w25127 = ~w25125 & ~w25126;
assign w25128 = pi1350 & ~w25127;
assign w25129 = ~pi1350 & w25127;
assign w25130 = ~w25128 & ~w25129;
assign w25131 = ~pi4578 & pi9040;
assign w25132 = ~pi4475 & ~pi9040;
assign w25133 = ~w25131 & ~w25132;
assign w25134 = pi1368 & ~w25133;
assign w25135 = ~pi1368 & w25133;
assign w25136 = ~w25134 & ~w25135;
assign w25137 = ~w25130 & ~w25136;
assign w25138 = ~pi4479 & pi9040;
assign w25139 = ~pi4507 & ~pi9040;
assign w25140 = ~w25138 & ~w25139;
assign w25141 = pi1361 & ~w25140;
assign w25142 = ~pi1361 & w25140;
assign w25143 = ~w25141 & ~w25142;
assign w25144 = ~pi4475 & pi9040;
assign w25145 = ~pi4603 & ~pi9040;
assign w25146 = ~w25144 & ~w25145;
assign w25147 = pi1334 & ~w25146;
assign w25148 = ~pi1334 & w25146;
assign w25149 = ~w25147 & ~w25148;
assign w25150 = ~w25143 & ~w25149;
assign w25151 = ~pi4473 & pi9040;
assign w25152 = ~pi4413 & ~pi9040;
assign w25153 = ~w25151 & ~w25152;
assign w25154 = pi1358 & ~w25153;
assign w25155 = ~pi1358 & w25153;
assign w25156 = ~w25154 & ~w25155;
assign w25157 = w25150 & ~w25156;
assign w25158 = w25137 & w25157;
assign w25159 = ~pi4553 & pi9040;
assign w25160 = ~pi4401 & ~pi9040;
assign w25161 = ~w25159 & ~w25160;
assign w25162 = pi1363 & ~w25161;
assign w25163 = ~pi1363 & w25161;
assign w25164 = ~w25162 & ~w25163;
assign w25165 = w25130 & w25136;
assign w25166 = (w25143 & ~w25165) | (w25143 & w63796) | (~w25165 & w63796);
assign w25167 = ~w25130 & w25136;
assign w25168 = w25156 & w25167;
assign w25169 = w25137 & ~w25156;
assign w25170 = ~w25168 & ~w25169;
assign w25171 = w25170 & w63797;
assign w25172 = ~w25149 & w25165;
assign w25173 = w25149 & ~w25167;
assign w25174 = w25130 & ~w25136;
assign w25175 = ~w25156 & w25174;
assign w25176 = (~w25149 & ~w25174) | (~w25149 & w25198) | (~w25174 & w25198);
assign w25177 = ~w25173 & ~w25176;
assign w25178 = ~w25172 & ~w25177;
assign w25179 = ~w25166 & ~w25178;
assign w25180 = w25149 & w25174;
assign w25181 = w25174 & w25189;
assign w25182 = ~w25171 & ~w25181;
assign w25183 = ~w25179 & w25182;
assign w25184 = ~w25164 & ~w25183;
assign w25185 = ~w25149 & ~w25156;
assign w25186 = w25136 & w25185;
assign w25187 = ~w25171 & ~w25186;
assign w25188 = w25150 & w65613;
assign w25189 = w25149 & w25156;
assign w25190 = w25137 & ~w25185;
assign w25191 = ~w25189 & w25190;
assign w25192 = ~w25181 & ~w25188;
assign w25193 = ~w25191 & w25192;
assign w25194 = ~w25187 & ~w25193;
assign w25195 = w25156 & w25165;
assign w25196 = (w25143 & ~w25165) | (w25143 & w65614) | (~w25165 & w65614);
assign w25197 = ~w25177 & w25196;
assign w25198 = ~w25149 & w25156;
assign w25199 = ~w25137 & w25198;
assign w25200 = ~w25165 & w25199;
assign w25201 = w25130 & w25156;
assign w25202 = w25173 & ~w25201;
assign w25203 = ~w25143 & ~w25200;
assign w25204 = ~w25202 & w25203;
assign w25205 = w25164 & ~w25197;
assign w25206 = ~w25204 & w25205;
assign w25207 = w25149 & w25201;
assign w25208 = w25185 & w25167;
assign w25209 = ~w25207 & ~w25208;
assign w25210 = w25143 & ~w25209;
assign w25211 = w25143 & ~w25164;
assign w25212 = ~w25130 & ~w25149;
assign w25213 = ~w25180 & ~w25212;
assign w25214 = (w25211 & w25180) | (w25211 & w65615) | (w25180 & w65615);
assign w25215 = ~w25158 & ~w25214;
assign w25216 = ~w25210 & w25215;
assign w25217 = ~w25194 & w25216;
assign w25218 = ~w25206 & w25217;
assign w25219 = (pi1376 & ~w25218) | (pi1376 & w65616) | (~w25218 & w65616);
assign w25220 = w25218 & w65617;
assign w25221 = ~w25219 & ~w25220;
assign w25222 = ~pi4481 & pi9040;
assign w25223 = ~pi4579 & ~pi9040;
assign w25224 = ~w25222 & ~w25223;
assign w25225 = pi1353 & ~w25224;
assign w25226 = ~pi1353 & w25224;
assign w25227 = ~w25225 & ~w25226;
assign w25228 = ~pi4852 & pi9040;
assign w25229 = ~pi4511 & ~pi9040;
assign w25230 = ~w25228 & ~w25229;
assign w25231 = pi1369 & ~w25230;
assign w25232 = ~pi1369 & w25230;
assign w25233 = ~w25231 & ~w25232;
assign w25234 = w25227 & ~w25233;
assign w25235 = ~pi4394 & pi9040;
assign w25236 = ~pi4711 & ~pi9040;
assign w25237 = ~w25235 & ~w25236;
assign w25238 = pi1352 & ~w25237;
assign w25239 = ~pi1352 & w25237;
assign w25240 = ~w25238 & ~w25239;
assign w25241 = ~w25233 & w25240;
assign w25242 = ~pi4711 & pi9040;
assign w25243 = ~pi4397 & ~pi9040;
assign w25244 = ~w25242 & ~w25243;
assign w25245 = pi1365 & ~w25244;
assign w25246 = ~pi1365 & w25244;
assign w25247 = ~w25245 & ~w25246;
assign w25248 = w25241 & ~w25247;
assign w25249 = ~pi4480 & pi9040;
assign w25250 = ~pi4602 & ~pi9040;
assign w25251 = ~w25249 & ~w25250;
assign w25252 = pi1366 & ~w25251;
assign w25253 = ~pi1366 & w25251;
assign w25254 = ~w25252 & ~w25253;
assign w25255 = (w25254 & w25248) | (w25254 & w65618) | (w25248 & w65618);
assign w25256 = ~w25241 & w25254;
assign w25257 = ~w25227 & ~w25240;
assign w25258 = ~w25247 & w25257;
assign w25259 = w25256 & ~w25258;
assign w25260 = ~w25255 & ~w25259;
assign w25261 = w25233 & w25254;
assign w25262 = w25227 & ~w25240;
assign w25263 = w25233 & ~w25247;
assign w25264 = w25262 & w25263;
assign w25265 = ~w25254 & ~w25264;
assign w25266 = ~w25261 & ~w25265;
assign w25267 = w25260 & w25266;
assign w25268 = ~w25227 & w25240;
assign w25269 = ~w25234 & ~w25268;
assign w25270 = ~w25247 & w25268;
assign w25271 = ~w25254 & ~w25270;
assign w25272 = ~w25269 & w25271;
assign w25273 = w25233 & w25247;
assign w25274 = w25257 & w25273;
assign w25275 = ~pi4579 & pi9040;
assign w25276 = ~pi4485 & ~pi9040;
assign w25277 = ~w25275 & ~w25276;
assign w25278 = pi1372 & ~w25277;
assign w25279 = ~pi1372 & w25277;
assign w25280 = ~w25278 & ~w25279;
assign w25281 = ~w25274 & ~w25280;
assign w25282 = w25233 & ~w25240;
assign w25283 = w25247 & w25254;
assign w25284 = w25282 & w25283;
assign w25285 = w25227 & w25240;
assign w25286 = ~w25248 & ~w25261;
assign w25287 = w25285 & ~w25286;
assign w25288 = w25247 & ~w25254;
assign w25289 = ~w25233 & w25257;
assign w25290 = ~w25288 & w25289;
assign w25291 = w25281 & ~w25284;
assign w25292 = ~w25290 & w25291;
assign w25293 = w25292 & w65619;
assign w25294 = w25288 & w25289;
assign w25295 = w25256 & ~w25269;
assign w25296 = w25273 & w25285;
assign w25297 = ~w25264 & ~w25296;
assign w25298 = ~w25241 & ~w25282;
assign w25299 = ~w25247 & ~w25254;
assign w25300 = ~w25298 & w25299;
assign w25301 = w25280 & ~w25294;
assign w25302 = ~w25295 & w25297;
assign w25303 = ~w25300 & w25302;
assign w25304 = w25301 & w25303;
assign w25305 = ~w25293 & ~w25304;
assign w25306 = w25263 & w25268;
assign w25307 = w25254 & w25306;
assign w25308 = ~w25267 & ~w25307;
assign w25309 = ~w25305 & w25308;
assign w25310 = pi1383 & w25309;
assign w25311 = ~pi1383 & ~w25309;
assign w25312 = ~w25310 & ~w25311;
assign w25313 = ~pi4413 & pi9040;
assign w25314 = ~pi4521 & ~pi9040;
assign w25315 = ~w25313 & ~w25314;
assign w25316 = pi1375 & ~w25315;
assign w25317 = ~pi1375 & w25315;
assign w25318 = ~w25316 & ~w25317;
assign w25319 = ~pi4730 & pi9040;
assign w25320 = ~pi4381 & ~pi9040;
assign w25321 = ~w25319 & ~w25320;
assign w25322 = pi1368 & ~w25321;
assign w25323 = ~pi1368 & w25321;
assign w25324 = ~w25322 & ~w25323;
assign w25325 = ~w25318 & w25324;
assign w25326 = w25318 & ~w25324;
assign w25327 = ~w25325 & ~w25326;
assign w25328 = ~pi4400 & pi9040;
assign w25329 = ~pi4506 & ~pi9040;
assign w25330 = ~w25328 & ~w25329;
assign w25331 = pi1372 & ~w25330;
assign w25332 = ~pi1372 & w25330;
assign w25333 = ~w25331 & ~w25332;
assign w25334 = w25318 & ~w25333;
assign w25335 = ~pi4506 & pi9040;
assign w25336 = ~pi4512 & ~pi9040;
assign w25337 = ~w25335 & ~w25336;
assign w25338 = pi1353 & ~w25337;
assign w25339 = ~pi1353 & w25337;
assign w25340 = ~w25338 & ~w25339;
assign w25341 = ~w25334 & w25340;
assign w25342 = ~w25327 & w25341;
assign w25343 = w25324 & ~w25340;
assign w25344 = ~w25324 & w25340;
assign w25345 = ~w25343 & ~w25344;
assign w25346 = w25334 & ~w25345;
assign w25347 = ~w25318 & w25333;
assign w25348 = w25345 & w25347;
assign w25349 = ~w25346 & ~w25348;
assign w25350 = w25333 & w25340;
assign w25351 = ~w25333 & ~w25340;
assign w25352 = ~w25350 & ~w25351;
assign w25353 = ~w25324 & w25333;
assign w25354 = ~w25352 & ~w25353;
assign w25355 = ~pi4408 & pi9040;
assign w25356 = ~pi4473 & ~pi9040;
assign w25357 = ~w25355 & ~w25356;
assign w25358 = pi1360 & ~w25357;
assign w25359 = ~pi1360 & w25357;
assign w25360 = ~w25358 & ~w25359;
assign w25361 = w25349 & w63798;
assign w25362 = ~w25318 & w25340;
assign w25363 = ~w25333 & w25362;
assign w25364 = w25333 & w25343;
assign w25365 = ~w25360 & ~w25364;
assign w25366 = ~w25363 & w25365;
assign w25367 = (~w25342 & w25361) | (~w25342 & w65620) | (w25361 & w65620);
assign w25368 = ~pi4402 & pi9040;
assign w25369 = ~pi4615 & ~pi9040;
assign w25370 = ~w25368 & ~w25369;
assign w25371 = pi1350 & ~w25370;
assign w25372 = ~pi1350 & w25370;
assign w25373 = ~w25371 & ~w25372;
assign w25374 = ~w25367 & w25373;
assign w25375 = ~w25343 & ~w25351;
assign w25376 = ~w25341 & w25375;
assign w25377 = ~w25324 & w25360;
assign w25378 = w25362 & w25377;
assign w25379 = ~w25347 & ~w25360;
assign w25380 = ~w25347 & w65621;
assign w25381 = ~w25340 & ~w25380;
assign w25382 = ~w25341 & ~w25344;
assign w25383 = ~w25381 & w25382;
assign w25384 = (~w25378 & ~w25376) | (~w25378 & w65622) | (~w25376 & w65622);
assign w25385 = ~w25383 & w25384;
assign w25386 = ~w25373 & ~w25385;
assign w25387 = w25325 & w25350;
assign w25388 = w25333 & ~w25340;
assign w25389 = w25379 & w25388;
assign w25390 = w25326 & ~w25352;
assign w25391 = w25340 & w25360;
assign w25392 = (w25360 & ~w25325) | (w25360 & w65623) | (~w25325 & w65623);
assign w25393 = w25326 & w25388;
assign w25394 = ~w25391 & ~w25393;
assign w25395 = ~w25392 & w25394;
assign w25396 = ~w25390 & ~w25395;
assign w25397 = ~w25325 & ~w25334;
assign w25398 = ~w25375 & w25397;
assign w25399 = w25360 & ~w25364;
assign w25400 = ~w25398 & w25399;
assign w25401 = ~w25387 & ~w25389;
assign w25402 = (w25401 & w25396) | (w25401 & w65624) | (w25396 & w65624);
assign w25403 = ~w25386 & w25402;
assign w25404 = ~w25374 & w25403;
assign w25405 = pi1381 & ~w25404;
assign w25406 = ~pi1381 & w25404;
assign w25407 = ~w25405 & ~w25406;
assign w25408 = ~w25233 & ~w25254;
assign w25409 = w25227 & w25247;
assign w25410 = ~w25240 & ~w25408;
assign w25411 = w25409 & w25410;
assign w25412 = w25247 & ~w25285;
assign w25413 = w25298 & w25412;
assign w25414 = ~w25227 & w25413;
assign w25415 = (~w25258 & ~w25413) | (~w25258 & w65625) | (~w25413 & w65625);
assign w25416 = ~w25408 & ~w25415;
assign w25417 = w25262 & w25408;
assign w25418 = ~w25288 & ~w25417;
assign w25419 = ~w25412 & ~w25418;
assign w25420 = ~w25411 & ~w25419;
assign w25421 = ~w25416 & w25420;
assign w25422 = w25280 & ~w25421;
assign w25423 = ~w25268 & w25299;
assign w25424 = ~w25280 & w25283;
assign w25425 = ~w25423 & ~w25424;
assign w25426 = w25233 & ~w25262;
assign w25427 = ~w25425 & w25426;
assign w25428 = w25227 & ~w25247;
assign w25429 = ~w25280 & ~w25285;
assign w25430 = ~w25428 & w25429;
assign w25431 = ~w25270 & ~w25430;
assign w25432 = w25408 & ~w25431;
assign w25433 = w25254 & w25428;
assign w25434 = w25282 & w25433;
assign w25435 = w25280 & ~w25434;
assign w25436 = w25261 & w25268;
assign w25437 = ~w25248 & ~w25264;
assign w25438 = ~w25436 & w25437;
assign w25439 = ~w25435 & ~w25438;
assign w25440 = w25241 & w25433;
assign w25441 = ~w25427 & ~w25440;
assign w25442 = ~w25432 & w25441;
assign w25443 = ~w25439 & w25442;
assign w25444 = ~w25422 & w25443;
assign w25445 = pi1386 & ~w25444;
assign w25446 = ~pi1386 & w25444;
assign w25447 = ~w25445 & ~w25446;
assign w25448 = ~w25164 & w25189;
assign w25449 = w25137 & w25448;
assign w25450 = w25165 & w65626;
assign w25451 = ~w25208 & ~w25450;
assign w25452 = w25143 & ~w25168;
assign w25453 = w25451 & w25452;
assign w25454 = ~w25130 & ~w25156;
assign w25455 = ~w25186 & w25454;
assign w25456 = ~w25143 & ~w25207;
assign w25457 = ~w25455 & w25456;
assign w25458 = ~w25453 & ~w25457;
assign w25459 = w25193 & ~w25458;
assign w25460 = w25164 & ~w25459;
assign w25461 = w25174 & w25185;
assign w25462 = ~w25143 & ~w25164;
assign w25463 = ~w25199 & w25451;
assign w25464 = w25462 & ~w25463;
assign w25465 = w25149 & w25169;
assign w25466 = ~w25175 & ~w25195;
assign w25467 = ~w25455 & w25466;
assign w25468 = w25211 & ~w25465;
assign w25469 = ~w25467 & w25468;
assign w25470 = w25136 & w25143;
assign w25471 = w25198 & w25470;
assign w25472 = ~w25461 & ~w25471;
assign w25473 = ~w25449 & w25472;
assign w25474 = ~w25469 & w25473;
assign w25475 = ~w25464 & w25474;
assign w25476 = ~w25460 & w25475;
assign w25477 = pi1378 & ~w25476;
assign w25478 = ~pi1378 & w25476;
assign w25479 = ~w25477 & ~w25478;
assign w25480 = ~w24834 & ~w24857;
assign w25481 = (w24834 & ~w24876) | (w24834 & w63799) | (~w24876 & w63799);
assign w25482 = ~w24887 & w25481;
assign w25483 = (~w24869 & w25482) | (~w24869 & w65627) | (w25482 & w65627);
assign w25484 = ~w24870 & ~w25483;
assign w25485 = w24867 & ~w25484;
assign w25486 = (w24849 & ~w24843) | (w24849 & w65628) | (~w24843 & w65628);
assign w25487 = w25481 & w25486;
assign w25488 = ~w24870 & ~w25487;
assign w25489 = w24849 & ~w24858;
assign w25490 = w24872 & ~w25489;
assign w25491 = ~w24867 & ~w25490;
assign w25492 = w25488 & w25491;
assign w25493 = ~w25485 & ~w25492;
assign w25494 = ~w24891 & ~w24897;
assign w25495 = w24903 & ~w25494;
assign w25496 = (~w24890 & w24900) | (~w24890 & w65629) | (w24900 & w65629);
assign w25497 = ~w24873 & ~w24904;
assign w25498 = w25496 & w25497;
assign w25499 = w24898 & ~w25498;
assign w25500 = ~w25495 & ~w25499;
assign w25501 = ~w25493 & w25500;
assign w25502 = pi1417 & ~w25501;
assign w25503 = ~pi1417 & w25501;
assign w25504 = ~w25502 & ~w25503;
assign w25505 = w24828 & ~w24867;
assign w25506 = ~w24868 & w25505;
assign w25507 = (~w25506 & w24875) | (~w25506 & w65630) | (w24875 & w65630);
assign w25508 = w24887 & ~w25507;
assign w25509 = ~w24842 & ~w24873;
assign w25510 = w24849 & ~w25509;
assign w25511 = ~w24835 & ~w24857;
assign w25512 = ~w24841 & ~w24849;
assign w25513 = ~w25511 & w25512;
assign w25514 = ~w24867 & ~w25513;
assign w25515 = ~w25510 & w25514;
assign w25516 = w25496 & w25515;
assign w25517 = ~w24891 & ~w25482;
assign w25518 = w25489 & ~w25517;
assign w25519 = ~w24842 & ~w24894;
assign w25520 = w24859 & ~w25519;
assign w25521 = (w24867 & ~w24860) | (w24867 & w65631) | (~w24860 & w65631);
assign w25522 = ~w25520 & w25521;
assign w25523 = ~w25518 & w25522;
assign w25524 = ~w25516 & ~w25523;
assign w25525 = ~w24856 & w24869;
assign w25526 = ~w25508 & ~w25525;
assign w25527 = ~w25524 & w25526;
assign w25528 = pi1403 & ~w25527;
assign w25529 = ~pi1403 & w25527;
assign w25530 = ~w25528 & ~w25529;
assign w25531 = ~pi4385 & pi9040;
assign w25532 = ~pi4650 & ~pi9040;
assign w25533 = ~w25531 & ~w25532;
assign w25534 = pi1362 & ~w25533;
assign w25535 = ~pi1362 & w25533;
assign w25536 = ~w25534 & ~w25535;
assign w25537 = ~pi4602 & pi9040;
assign w25538 = ~pi4393 & ~pi9040;
assign w25539 = ~w25537 & ~w25538;
assign w25540 = pi1356 & ~w25539;
assign w25541 = ~pi1356 & w25539;
assign w25542 = ~w25540 & ~w25541;
assign w25543 = ~w25536 & ~w25542;
assign w25544 = ~pi4397 & pi9040;
assign w25545 = ~pi4425 & ~pi9040;
assign w25546 = ~w25544 & ~w25545;
assign w25547 = pi1364 & ~w25546;
assign w25548 = ~pi1364 & w25546;
assign w25549 = ~w25547 & ~w25548;
assign w25550 = ~pi4403 & pi9040;
assign w25551 = ~pi4492 & ~pi9040;
assign w25552 = ~w25550 & ~w25551;
assign w25553 = pi1339 & ~w25552;
assign w25554 = ~pi1339 & w25552;
assign w25555 = ~w25553 & ~w25554;
assign w25556 = ~w25549 & ~w25555;
assign w25557 = ~pi4583 & pi9040;
assign w25558 = ~pi4508 & ~pi9040;
assign w25559 = ~w25557 & ~w25558;
assign w25560 = pi1359 & ~w25559;
assign w25561 = ~pi1359 & w25559;
assign w25562 = ~w25560 & ~w25561;
assign w25563 = w25549 & ~w25562;
assign w25564 = ~w25536 & ~w25563;
assign w25565 = (~w25543 & ~w25564) | (~w25543 & w65632) | (~w25564 & w65632);
assign w25566 = ~w25542 & w25562;
assign w25567 = w25556 & w25566;
assign w25568 = w25542 & ~w25562;
assign w25569 = w25556 & w25568;
assign w25570 = w25549 & ~w25555;
assign w25571 = w25566 & w25570;
assign w25572 = ~w25549 & w25562;
assign w25573 = ~w25556 & ~w25566;
assign w25574 = w25572 & w25573;
assign w25575 = ~w25569 & ~w25571;
assign w25576 = ~w25574 & w25575;
assign w25577 = ~w25567 & w25576;
assign w25578 = ~w25565 & ~w25577;
assign w25579 = ~pi4425 & pi9040;
assign w25580 = ~pi4494 & ~pi9040;
assign w25581 = ~w25579 & ~w25580;
assign w25582 = pi1357 & ~w25581;
assign w25583 = ~pi1357 & w25581;
assign w25584 = ~w25582 & ~w25583;
assign w25585 = w25549 & w25555;
assign w25586 = w25573 & ~w25585;
assign w25587 = w25573 & w65633;
assign w25588 = ~w25542 & ~w25570;
assign w25589 = w25542 & w25570;
assign w25590 = ~w25588 & ~w25589;
assign w25591 = ~w25536 & w25590;
assign w25592 = ~w25555 & w25572;
assign w25593 = w25590 & w63800;
assign w25594 = ~w25542 & ~w25556;
assign w25595 = ~w25556 & w63801;
assign w25596 = ~w25542 & ~w25595;
assign w25597 = ~w25586 & ~w25596;
assign w25598 = ~w25536 & ~w25572;
assign w25599 = w25588 & ~w25598;
assign w25600 = ~w25597 & w25599;
assign w25601 = ~w25587 & ~w25593;
assign w25602 = ~w25600 & w25601;
assign w25603 = ~w25584 & ~w25602;
assign w25604 = (w25568 & ~w25590) | (w25568 & w65634) | (~w25590 & w65634);
assign w25605 = w25536 & w25597;
assign w25606 = w25588 & w25598;
assign w25607 = ~w25571 & ~w25606;
assign w25608 = ~w25604 & w25607;
assign w25609 = ~w25605 & w25608;
assign w25610 = w25584 & ~w25609;
assign w25611 = ~w25578 & ~w25603;
assign w25612 = w25611 & w65635;
assign w25613 = (~pi1394 & ~w25611) | (~pi1394 & w65636) | (~w25611 & w65636);
assign w25614 = ~w25612 & ~w25613;
assign w25615 = ~w25362 & ~w25388;
assign w25616 = ~w25345 & w25615;
assign w25617 = w25392 & ~w25616;
assign w25618 = ~w25395 & ~w25617;
assign w25619 = w25348 & w25377;
assign w25620 = (~w25360 & w25345) | (~w25360 & w65637) | (w25345 & w65637);
assign w25621 = ~w25350 & ~w25620;
assign w25622 = w25350 & ~w25360;
assign w25623 = w25324 & ~w25622;
assign w25624 = ~w25621 & w25623;
assign w25625 = ~w25363 & ~w25373;
assign w25626 = ~w25390 & w25625;
assign w25627 = ~w25619 & w25626;
assign w25628 = ~w25624 & w25627;
assign w25629 = ~w25379 & ~w25400;
assign w25630 = ~w25346 & w25373;
assign w25631 = ~w25629 & w25630;
assign w25632 = ~w25628 & ~w25631;
assign w25633 = ~w25618 & ~w25632;
assign w25634 = ~pi1379 & w25633;
assign w25635 = pi1379 & ~w25633;
assign w25636 = ~w25634 & ~w25635;
assign w25637 = ~w24899 & w24905;
assign w25638 = ~w24871 & ~w25511;
assign w25639 = w25637 & w25638;
assign w25640 = w24881 & w24892;
assign w25641 = ~w24867 & ~w25640;
assign w25642 = ~w25639 & w25641;
assign w25643 = ~w25488 & w25519;
assign w25644 = w24867 & ~w24874;
assign w25645 = w25494 & w25644;
assign w25646 = ~w25643 & w25645;
assign w25647 = ~w25642 & ~w25646;
assign w25648 = w24868 & w24876;
assign w25649 = (w24867 & ~w24905) | (w24867 & w65638) | (~w24905 & w65638);
assign w25650 = ~w24893 & ~w25649;
assign w25651 = ~w24849 & ~w25650;
assign w25652 = ~w24861 & ~w25648;
assign w25653 = ~w25651 & w25652;
assign w25654 = ~w25647 & w25653;
assign w25655 = pi1425 & w25654;
assign w25656 = ~pi1425 & ~w25654;
assign w25657 = ~w25655 & ~w25656;
assign w25658 = w24967 & w25014;
assign w25659 = w24974 & ~w24981;
assign w25660 = ~w25658 & ~w25659;
assign w25661 = w24958 & ~w25006;
assign w25662 = (~w24958 & ~w24951) | (~w24958 & w65639) | (~w24951 & w65639);
assign w25663 = w24939 & ~w24981;
assign w25664 = ~w24927 & ~w24939;
assign w25665 = ~w24963 & ~w25664;
assign w25666 = ~w24950 & ~w25665;
assign w25667 = w25662 & ~w25663;
assign w25668 = ~w25666 & w25667;
assign w25669 = (w25660 & w25668) | (w25660 & w65640) | (w25668 & w65640);
assign w25670 = w24921 & ~w25669;
assign w25671 = ~w24921 & ~w24982;
assign w25672 = ~w25659 & w25671;
assign w25673 = w24958 & ~w24962;
assign w25674 = ~w25672 & w25673;
assign w25675 = ~w24921 & ~w25007;
assign w25676 = ~w24958 & w25660;
assign w25677 = ~w25675 & w25676;
assign w25678 = ~w25674 & ~w25677;
assign w25679 = ~w25670 & ~w25678;
assign w25680 = ~pi1387 & w25679;
assign w25681 = pi1387 & ~w25679;
assign w25682 = ~w25680 & ~w25681;
assign w25683 = w25536 & w25562;
assign w25684 = w25555 & ~w25562;
assign w25685 = ~w25683 & ~w25684;
assign w25686 = ~w25567 & ~w25604;
assign w25687 = ~w25685 & ~w25686;
assign w25688 = w25536 & w25555;
assign w25689 = ~w25566 & w25688;
assign w25690 = w25589 & w25683;
assign w25691 = ~w25556 & ~w25585;
assign w25692 = w25542 & w25549;
assign w25693 = w25691 & w65641;
assign w25694 = w25566 & w25585;
assign w25695 = ~w25536 & ~w25555;
assign w25696 = w25563 & w25695;
assign w25697 = ~w25694 & ~w25696;
assign w25698 = ~w25690 & w25697;
assign w25699 = ~w25693 & w25698;
assign w25700 = w25564 & ~w25590;
assign w25701 = w25699 & w25700;
assign w25702 = w25543 & ~w25697;
assign w25703 = w25568 & ~w25691;
assign w25704 = w25584 & ~w25689;
assign w25705 = ~w25703 & w25704;
assign w25706 = ~w25702 & w25705;
assign w25707 = ~w25701 & w25706;
assign w25708 = ~w25568 & w25591;
assign w25709 = w25698 & w65642;
assign w25710 = ~w25708 & w25709;
assign w25711 = (~w25687 & w25707) | (~w25687 & w65643) | (w25707 & w65643);
assign w25712 = pi1390 & w25711;
assign w25713 = ~pi1390 & ~w25711;
assign w25714 = ~w25712 & ~w25713;
assign w25715 = w25150 & w25201;
assign w25716 = ~w25461 & ~w25715;
assign w25717 = w25165 & w65614;
assign w25718 = (~w25164 & ~w25716) | (~w25164 & w65644) | (~w25716 & w65644);
assign w25719 = ~w25143 & w25466;
assign w25720 = (w25149 & ~w25170) | (w25149 & w65645) | (~w25170 & w65645);
assign w25721 = ~w25719 & w25720;
assign w25722 = w25156 & w25214;
assign w25723 = ~w25198 & w25462;
assign w25724 = w25170 & w25723;
assign w25725 = ~w25157 & ~w25724;
assign w25726 = ~w25130 & ~w25725;
assign w25727 = w25150 & w25716;
assign w25728 = ~w25150 & w25156;
assign w25729 = ~w25137 & w25728;
assign w25730 = w25213 & w25729;
assign w25731 = ~w25208 & ~w25727;
assign w25732 = ~w25730 & w25731;
assign w25733 = w25164 & ~w25732;
assign w25734 = ~w25718 & ~w25722;
assign w25735 = ~w25721 & w25734;
assign w25736 = ~w25726 & w25735;
assign w25737 = ~w25733 & w25736;
assign w25738 = ~pi1385 & w25737;
assign w25739 = pi1385 & ~w25737;
assign w25740 = ~w25738 & ~w25739;
assign w25741 = w25298 & w25409;
assign w25742 = ~w25290 & ~w25741;
assign w25743 = ~w25254 & ~w25742;
assign w25744 = w25241 & w25254;
assign w25745 = w25292 & w65646;
assign w25746 = ~w25283 & w25289;
assign w25747 = ~w25240 & ~w25433;
assign w25748 = w25240 & ~w25263;
assign w25749 = ~w25423 & w25748;
assign w25750 = ~w25747 & ~w25749;
assign w25751 = w25281 & ~w25746;
assign w25752 = ~w25750 & w25751;
assign w25753 = ~w25263 & w25268;
assign w25754 = ~w25264 & ~w25753;
assign w25755 = ~w25254 & ~w25754;
assign w25756 = w25257 & w25261;
assign w25757 = ~w25440 & ~w25756;
assign w25758 = ~w25741 & w25757;
assign w25759 = w25280 & ~w25755;
assign w25760 = w25758 & w25759;
assign w25761 = ~w25752 & ~w25760;
assign w25762 = ~w25284 & ~w25307;
assign w25763 = ~w25743 & w25762;
assign w25764 = ~w25745 & w25763;
assign w25765 = ~w25761 & w25764;
assign w25766 = pi1393 & ~w25765;
assign w25767 = ~pi1393 & w25765;
assign w25768 = ~w25766 & ~w25767;
assign w25769 = w25288 & w25414;
assign w25770 = (~w25263 & ~w25410) | (~w25263 & w65647) | (~w25410 & w65647);
assign w25771 = w25271 & ~w25770;
assign w25772 = ~w25255 & ~w25413;
assign w25773 = ~w25771 & w25772;
assign w25774 = w25280 & ~w25773;
assign w25775 = (w25283 & ~w25757) | (w25283 & w65648) | (~w25757 & w65648);
assign w25776 = w25234 & w25240;
assign w25777 = w25271 & ~w25776;
assign w25778 = w25260 & ~w25777;
assign w25779 = w25297 & ~w25306;
assign w25780 = ~w25778 & w25779;
assign w25781 = ~w25280 & ~w25780;
assign w25782 = ~w25769 & ~w25775;
assign w25783 = ~w25774 & w25782;
assign w25784 = ~w25781 & w25783;
assign w25785 = pi1402 & ~w25784;
assign w25786 = ~pi1402 & w25784;
assign w25787 = ~w25785 & ~w25786;
assign w25788 = w24958 & ~w24984;
assign w25789 = w24950 & w24975;
assign w25790 = w25662 & ~w25789;
assign w25791 = ~w25788 & ~w25790;
assign w25792 = w24927 & w24964;
assign w25793 = ~w24981 & w25664;
assign w25794 = w24981 & ~w25664;
assign w25795 = w24993 & w25794;
assign w25796 = (~w24958 & w25795) | (~w24958 & w65649) | (w25795 & w65649);
assign w25797 = ~w24977 & ~w25666;
assign w25798 = w25013 & ~w25797;
assign w25799 = w24921 & ~w25792;
assign w25800 = ~w25798 & w25799;
assign w25801 = ~w25796 & w25800;
assign w25802 = ~w24964 & ~w24974;
assign w25803 = ~w25659 & ~w25802;
assign w25804 = w24973 & ~w24975;
assign w25805 = ~w24951 & ~w25804;
assign w25806 = ~w24979 & ~w25805;
assign w25807 = w25009 & ~w25793;
assign w25808 = ~w24921 & ~w25803;
assign w25809 = ~w25806 & ~w25807;
assign w25810 = w25808 & w25809;
assign w25811 = (~w25791 & w25801) | (~w25791 & w65650) | (w25801 & w65650);
assign w25812 = ~pi1397 & w25811;
assign w25813 = pi1397 & ~w25811;
assign w25814 = ~w25812 & ~w25813;
assign w25815 = ~pi4508 & pi9040;
assign w25816 = ~pi4609 & ~pi9040;
assign w25817 = ~w25815 & ~w25816;
assign w25818 = pi1352 & ~w25817;
assign w25819 = ~pi1352 & w25817;
assign w25820 = ~w25818 & ~w25819;
assign w25821 = ~pi4399 & pi9040;
assign w25822 = ~pi4385 & ~pi9040;
assign w25823 = ~w25821 & ~w25822;
assign w25824 = pi1357 & ~w25823;
assign w25825 = ~pi1357 & w25823;
assign w25826 = ~w25824 & ~w25825;
assign w25827 = ~pi4419 & pi9040;
assign w25828 = ~pi4392 & ~pi9040;
assign w25829 = ~w25827 & ~w25828;
assign w25830 = pi1369 & ~w25829;
assign w25831 = ~pi1369 & w25829;
assign w25832 = ~w25830 & ~w25831;
assign w25833 = ~w25826 & ~w25832;
assign w25834 = w25826 & w25832;
assign w25835 = ~w25833 & ~w25834;
assign w25836 = ~pi4392 & pi9040;
assign w25837 = ~pi4481 & ~pi9040;
assign w25838 = ~w25836 & ~w25837;
assign w25839 = pi1364 & ~w25838;
assign w25840 = ~pi1364 & w25838;
assign w25841 = ~w25839 & ~w25840;
assign w25842 = ~pi4396 & pi9040;
assign w25843 = ~pi4399 & ~pi9040;
assign w25844 = ~w25842 & ~w25843;
assign w25845 = pi1351 & ~w25844;
assign w25846 = ~pi1351 & w25844;
assign w25847 = ~w25845 & ~w25846;
assign w25848 = ~w25841 & ~w25847;
assign w25849 = ~w25835 & ~w25848;
assign w25850 = ~pi4494 & pi9040;
assign w25851 = ~pi4583 & ~pi9040;
assign w25852 = ~w25850 & ~w25851;
assign w25853 = pi1343 & ~w25852;
assign w25854 = ~pi1343 & w25852;
assign w25855 = ~w25853 & ~w25854;
assign w25856 = w25849 & ~w25855;
assign w25857 = w25835 & ~w25841;
assign w25858 = w25841 & w25847;
assign w25859 = ~w25848 & ~w25858;
assign w25860 = w25826 & ~w25832;
assign w25861 = ~w25859 & w25860;
assign w25862 = ~w25826 & ~w25847;
assign w25863 = w25841 & w25855;
assign w25864 = w25862 & w25863;
assign w25865 = ~w25861 & ~w25864;
assign w25866 = w25832 & ~w25855;
assign w25867 = ~w25826 & w25866;
assign w25868 = ~w25859 & w25867;
assign w25869 = w25865 & ~w25868;
assign w25870 = (w25857 & ~w25865) | (w25857 & w63802) | (~w25865 & w63802);
assign w25871 = w25832 & w25862;
assign w25872 = w25833 & w25847;
assign w25873 = ~w25871 & ~w25872;
assign w25874 = ~w25826 & ~w25841;
assign w25875 = w25859 & ~w25874;
assign w25876 = w25855 & w25873;
assign w25877 = ~w25875 & w25876;
assign w25878 = ~w25856 & ~w25877;
assign w25879 = (w25820 & ~w25878) | (w25820 & w63803) | (~w25878 & w63803);
assign w25880 = ~w25835 & w25848;
assign w25881 = w25826 & w25847;
assign w25882 = ~w25841 & w25881;
assign w25883 = w25833 & w25841;
assign w25884 = ~w25882 & ~w25883;
assign w25885 = w25873 & w25884;
assign w25886 = ~w25834 & ~w25848;
assign w25887 = (~w25880 & ~w25885) | (~w25880 & w63804) | (~w25885 & w63804);
assign w25888 = ~w25855 & ~w25887;
assign w25889 = (~w25855 & ~w25881) | (~w25855 & w65651) | (~w25881 & w65651);
assign w25890 = ~w25866 & ~w25889;
assign w25891 = ~w25885 & w25890;
assign w25892 = (~w25820 & w25888) | (~w25820 & w65652) | (w25888 & w65652);
assign w25893 = ~w25832 & ~w25855;
assign w25894 = ~w25862 & ~w25881;
assign w25895 = w25893 & w25894;
assign w25896 = w25832 & ~w25841;
assign w25897 = ~w25835 & ~w25896;
assign w25898 = ~w25857 & ~w25897;
assign w25899 = w25889 & ~w25895;
assign w25900 = ~w25898 & w25899;
assign w25901 = w25858 & w25900;
assign w25902 = ~w25832 & w25841;
assign w25903 = ~w25881 & ~w25902;
assign w25904 = w25855 & w25903;
assign w25905 = ~w25865 & w25904;
assign w25906 = ~w25901 & ~w25905;
assign w25907 = ~w25879 & w25906;
assign w25908 = (pi1398 & ~w25907) | (pi1398 & w65653) | (~w25907 & w65653);
assign w25909 = w25907 & w65654;
assign w25910 = ~w25908 & ~w25909;
assign w25911 = (~w25728 & w25177) | (~w25728 & w65655) | (w25177 & w65655);
assign w25912 = ~w25178 & ~w25911;
assign w25913 = ~w25143 & w25174;
assign w25914 = ~w25191 & ~w25913;
assign w25915 = w25187 & w25914;
assign w25916 = (w25164 & ~w25915) | (w25164 & w65656) | (~w25915 & w65656);
assign w25917 = ~w25170 & w25462;
assign w25918 = ~w25136 & w25715;
assign w25919 = w25165 & w25448;
assign w25920 = ~w25137 & ~w25164;
assign w25921 = ~w25172 & w25920;
assign w25922 = w25452 & w25921;
assign w25923 = ~w25918 & ~w25919;
assign w25924 = ~w25917 & w25923;
assign w25925 = ~w25922 & w25924;
assign w25926 = ~w25194 & w25925;
assign w25927 = ~w25916 & w25926;
assign w25928 = pi1392 & w25927;
assign w25929 = ~pi1392 & ~w25927;
assign w25930 = ~w25928 & ~w25929;
assign w25931 = ~w25324 & w25350;
assign w25932 = (w25324 & ~w25362) | (w25324 & w63392) | (~w25362 & w63392);
assign w25933 = ~w25397 & w25932;
assign w25934 = ~w25931 & ~w25933;
assign w25935 = (w25360 & w25933) | (w25360 & w65657) | (w25933 & w65657);
assign w25936 = ~w25348 & ~w25616;
assign w25937 = ~w25325 & ~w25353;
assign w25938 = ~w25615 & w25937;
assign w25939 = w25360 & ~w25376;
assign w25940 = w25934 & w25939;
assign w25941 = (~w25938 & w25936) | (~w25938 & w63393) | (w25936 & w63393);
assign w25942 = ~w25940 & w25941;
assign w25943 = ~w25334 & w25936;
assign w25944 = (~w25935 & ~w25942) | (~w25935 & w63805) | (~w25942 & w63805);
assign w25945 = w25373 & ~w25944;
assign w25946 = w25326 & w25351;
assign w25947 = w25344 & w25347;
assign w25948 = w25360 & ~w25946;
assign w25949 = ~w25947 & w25948;
assign w25950 = ~w25620 & ~w25949;
assign w25951 = (~w25950 & w25942) | (~w25950 & w65658) | (w25942 & w65658);
assign w25952 = ~w25945 & w65659;
assign w25953 = (pi1391 & w25945) | (pi1391 & w65660) | (w25945 & w65660);
assign w25954 = ~w25952 & ~w25953;
assign w25955 = w25075 & w25095;
assign w25956 = ~w25042 & ~w25067;
assign w25957 = ~w25069 & ~w25956;
assign w25958 = w25036 & ~w25957;
assign w25959 = ~w25076 & ~w25110;
assign w25960 = w25958 & ~w25959;
assign w25961 = w25088 & ~w25108;
assign w25962 = ~w25036 & w25961;
assign w25963 = (~w25049 & w25960) | (~w25049 & w65661) | (w25960 & w65661);
assign w25964 = w25074 & ~w25098;
assign w25965 = ~w25056 & w25071;
assign w25966 = ~w25096 & ~w25965;
assign w25967 = ~w25964 & w25966;
assign w25968 = (~w25085 & w25960) | (~w25085 & w65662) | (w25960 & w65662);
assign w25969 = ~w25036 & ~w25100;
assign w25970 = w25070 & w25111;
assign w25971 = ~w25958 & w25970;
assign w25972 = (w25085 & w25111) | (w25085 & w65663) | (w25111 & w65663);
assign w25973 = ~w25971 & w25972;
assign w25974 = ~w25094 & ~w25955;
assign w25975 = ~w25963 & w25974;
assign w25976 = ~w25968 & ~w25973;
assign w25977 = (pi1396 & ~w25976) | (pi1396 & w65664) | (~w25976 & w65664);
assign w25978 = w25976 & w65665;
assign w25979 = ~w25977 & ~w25978;
assign w25980 = w25847 & w25896;
assign w25981 = (~w25896 & ~w25885) | (~w25896 & w63806) | (~w25885 & w63806);
assign w25982 = (w25885 & w65666) | (w25885 & w65667) | (w65666 & w65667);
assign w25983 = w25833 & w25848;
assign w25984 = ~w25980 & ~w25983;
assign w25985 = ~w25982 & w25984;
assign w25986 = w25855 & ~w25985;
assign w25987 = (~w25820 & ~w25869) | (~w25820 & w63807) | (~w25869 & w63807);
assign w25988 = w25848 & w25860;
assign w25989 = (w25820 & ~w25873) | (w25820 & w65668) | (~w25873 & w65668);
assign w25990 = w25858 & w25989;
assign w25991 = w25820 & ~w25855;
assign w25992 = ~w25833 & w25991;
assign w25993 = w25981 & w25992;
assign w25994 = ~w25987 & ~w25990;
assign w25995 = ~w25993 & w25994;
assign w25996 = (pi1408 & ~w25995) | (pi1408 & w65669) | (~w25995 & w65669);
assign w25997 = w25995 & w65670;
assign w25998 = ~w25996 & ~w25997;
assign w25999 = ~w25841 & ~w25887;
assign w26000 = ~w25874 & w25903;
assign w26001 = ~w25832 & w25858;
assign w26002 = w25855 & ~w26001;
assign w26003 = ~w26000 & ~w26002;
assign w26004 = ~w25904 & ~w26003;
assign w26005 = (~w25820 & w25999) | (~w25820 & w65671) | (w25999 & w65671);
assign w26006 = w25832 & w25882;
assign w26007 = ~w25989 & ~w26006;
assign w26008 = w25855 & ~w26007;
assign w26009 = ~w25820 & ~w25893;
assign w26010 = ~w25834 & w25858;
assign w26011 = ~w26009 & w26010;
assign w26012 = ~w25881 & ~w25883;
assign w26013 = w25991 & ~w26012;
assign w26014 = ~w26011 & ~w26013;
assign w26015 = ~w26008 & w26014;
assign w26016 = ~w26005 & w26015;
assign w26017 = pi1399 & ~w26016;
assign w26018 = ~pi1399 & w26016;
assign w26019 = ~w26017 & ~w26018;
assign w26020 = w25036 & w25109;
assign w26021 = ~w25036 & w25089;
assign w26022 = w25049 & w25961;
assign w26023 = ~w25085 & ~w26020;
assign w26024 = ~w26021 & ~w26022;
assign w26025 = w26023 & w26024;
assign w26026 = w25042 & w25107;
assign w26027 = w25085 & ~w26026;
assign w26028 = ~w25036 & ~w25064;
assign w26029 = ~w25956 & w26028;
assign w26030 = ~w25075 & ~w26029;
assign w26031 = ~w25958 & w26030;
assign w26032 = w26027 & w26031;
assign w26033 = ~w26025 & ~w26032;
assign w26034 = w25072 & w25092;
assign w26035 = ~w26033 & ~w26034;
assign w26036 = ~pi1389 & w26035;
assign w26037 = pi1389 & ~w26035;
assign w26038 = ~w26036 & ~w26037;
assign w26039 = ~w25542 & w25563;
assign w26040 = w25697 & w26039;
assign w26041 = w25568 & w25585;
assign w26042 = ~w25595 & ~w26041;
assign w26043 = w25576 & w26042;
assign w26044 = (~w25536 & ~w25576) | (~w25536 & w65672) | (~w25576 & w65672);
assign w26045 = w25536 & ~w25594;
assign w26046 = w26043 & w26045;
assign w26047 = ~w25584 & ~w26040;
assign w26048 = ~w26044 & w26047;
assign w26049 = ~w26046 & w26048;
assign w26050 = w25536 & ~w25572;
assign w26051 = ~w25573 & w26050;
assign w26052 = ~w25589 & ~w25592;
assign w26053 = ~w26041 & w26052;
assign w26054 = ~w25536 & ~w26053;
assign w26055 = ~w25562 & ~w26042;
assign w26056 = ~w25574 & w25584;
assign w26057 = w25697 & ~w26051;
assign w26058 = w26056 & w26057;
assign w26059 = ~w26054 & w26058;
assign w26060 = ~w26055 & w26059;
assign w26061 = ~w26049 & ~w26060;
assign w26062 = pi1401 & w26061;
assign w26063 = ~pi1401 & ~w26061;
assign w26064 = ~w26062 & ~w26063;
assign w26065 = ~w25398 & ~w25947;
assign w26066 = ~w25360 & ~w26065;
assign w26067 = w25345 & ~w25391;
assign w26068 = w25349 & w65673;
assign w26069 = w25392 & ~w25931;
assign w26070 = ~w25325 & ~w25344;
assign w26071 = w26069 & ~w26070;
assign w26072 = w25373 & ~w25387;
assign w26073 = ~w26071 & w26072;
assign w26074 = ~w26068 & w26073;
assign w26075 = w25318 & ~w25375;
assign w26076 = w25365 & ~w25937;
assign w26077 = ~w26069 & ~w26076;
assign w26078 = ~w25373 & ~w26075;
assign w26079 = ~w26077 & w26078;
assign w26080 = ~w26074 & ~w26079;
assign w26081 = ~w25340 & w25360;
assign w26082 = ~w25349 & w26081;
assign w26083 = ~w26066 & ~w26082;
assign w26084 = ~w26080 & w26083;
assign w26085 = pi1407 & ~w26084;
assign w26086 = ~pi1407 & w26084;
assign w26087 = ~w26085 & ~w26086;
assign w26088 = ~w25036 & ~w25077;
assign w26089 = ~w25088 & w25099;
assign w26090 = ~w25065 & ~w25097;
assign w26091 = w25036 & ~w26090;
assign w26092 = ~w25068 & w25108;
assign w26093 = ~w25036 & w26092;
assign w26094 = ~w25073 & ~w25085;
assign w26095 = ~w26089 & w26094;
assign w26096 = ~w26091 & ~w26093;
assign w26097 = w26095 & w26096;
assign w26098 = w25036 & ~w25049;
assign w26099 = w26092 & w26098;
assign w26100 = w25049 & ~w25111;
assign w26101 = w26027 & ~w26099;
assign w26102 = ~w26100 & w26101;
assign w26103 = ~w26097 & ~w26102;
assign w26104 = ~w26088 & ~w26103;
assign w26105 = ~pi1388 & w26104;
assign w26106 = pi1388 & ~w26104;
assign w26107 = ~w26105 & ~w26106;
assign w26108 = w25832 & w26010;
assign w26109 = w25833 & ~w25863;
assign w26110 = ~w25847 & ~w26109;
assign w26111 = ~w25898 & w26110;
assign w26112 = ~w25895 & ~w26108;
assign w26113 = (w25820 & w26111) | (w25820 & w65674) | (w26111 & w65674);
assign w26114 = w25855 & ~w25884;
assign w26115 = ~w25872 & w26002;
assign w26116 = ~w25889 & ~w26114;
assign w26117 = ~w26115 & w26116;
assign w26118 = w25855 & w25898;
assign w26119 = ~w25900 & ~w25983;
assign w26120 = (~w25820 & ~w26119) | (~w25820 & w65675) | (~w26119 & w65675);
assign w26121 = ~w26113 & ~w26117;
assign w26122 = ~w26120 & w26121;
assign w26123 = pi1409 & w26122;
assign w26124 = ~pi1409 & ~w26122;
assign w26125 = ~w26123 & ~w26124;
assign w26126 = w25543 & w25585;
assign w26127 = (w25536 & ~w25691) | (w25536 & w65676) | (~w25691 & w65676);
assign w26128 = w25565 & ~w26127;
assign w26129 = ~w25567 & ~w26128;
assign w26130 = w25584 & ~w26129;
assign w26131 = ~w25555 & w25562;
assign w26132 = ~w25542 & w25685;
assign w26133 = ~w25556 & ~w26132;
assign w26134 = ~w26131 & ~w26133;
assign w26135 = w25688 & w25692;
assign w26136 = ~w25587 & ~w26135;
assign w26137 = ~w26134 & w26136;
assign w26138 = ~w25584 & ~w26137;
assign w26139 = ~w25568 & w26050;
assign w26140 = ~w25596 & w26139;
assign w26141 = ~w26126 & ~w26140;
assign w26142 = ~w26130 & w26141;
assign w26143 = ~w26138 & w26142;
assign w26144 = pi1437 & ~w26143;
assign w26145 = ~pi1437 & w26143;
assign w26146 = ~w26144 & ~w26145;
assign w26147 = ~pi4958 & pi9040;
assign w26148 = ~pi4616 & ~pi9040;
assign w26149 = ~w26147 & ~w26148;
assign w26150 = pi1438 & ~w26149;
assign w26151 = ~pi1438 & w26149;
assign w26152 = ~w26150 & ~w26151;
assign w26153 = ~pi4604 & pi9040;
assign w26154 = ~pi4816 & ~pi9040;
assign w26155 = ~w26153 & ~w26154;
assign w26156 = pi1406 & ~w26155;
assign w26157 = ~pi1406 & w26155;
assign w26158 = ~w26156 & ~w26157;
assign w26159 = ~pi4689 & pi9040;
assign w26160 = ~pi4590 & ~pi9040;
assign w26161 = ~w26159 & ~w26160;
assign w26162 = pi1404 & ~w26161;
assign w26163 = ~pi1404 & w26161;
assign w26164 = ~w26162 & ~w26163;
assign w26165 = ~w26158 & ~w26164;
assign w26166 = ~pi4754 & pi9040;
assign w26167 = ~pi4710 & ~pi9040;
assign w26168 = ~w26166 & ~w26167;
assign w26169 = pi1427 & ~w26168;
assign w26170 = ~pi1427 & w26168;
assign w26171 = ~w26169 & ~w26170;
assign w26172 = w26165 & ~w26171;
assign w26173 = ~pi4695 & pi9040;
assign w26174 = ~pi4715 & ~pi9040;
assign w26175 = ~w26173 & ~w26174;
assign w26176 = pi1414 & ~w26175;
assign w26177 = ~pi1414 & w26175;
assign w26178 = ~w26176 & ~w26177;
assign w26179 = w26172 & w26178;
assign w26180 = w26152 & ~w26179;
assign w26181 = ~w26171 & w26178;
assign w26182 = w26158 & ~w26164;
assign w26183 = ~w26158 & w26164;
assign w26184 = ~w26182 & ~w26183;
assign w26185 = w26181 & ~w26184;
assign w26186 = ~w26165 & ~w26185;
assign w26187 = w26180 & ~w26186;
assign w26188 = ~w26152 & w26164;
assign w26189 = ~w26164 & w26171;
assign w26190 = w26164 & ~w26171;
assign w26191 = ~w26189 & ~w26190;
assign w26192 = w26158 & ~w26191;
assign w26193 = w26171 & ~w26178;
assign w26194 = w26183 & w26193;
assign w26195 = ~w26192 & ~w26194;
assign w26196 = (w26188 & w26192) | (w26188 & w65677) | (w26192 & w65677);
assign w26197 = ~pi4937 & pi9040;
assign w26198 = ~pi4604 & ~pi9040;
assign w26199 = ~w26197 & ~w26198;
assign w26200 = pi1423 & ~w26199;
assign w26201 = ~pi1423 & w26199;
assign w26202 = ~w26200 & ~w26201;
assign w26203 = w26181 & w26183;
assign w26204 = w26172 & ~w26178;
assign w26205 = w26152 & w26171;
assign w26206 = ~w26181 & ~w26193;
assign w26207 = w26152 & ~w26158;
assign w26208 = w26164 & ~w26207;
assign w26209 = w26206 & w26208;
assign w26210 = ~w26158 & ~w26178;
assign w26211 = w26171 & ~w26188;
assign w26212 = w26210 & w26211;
assign w26213 = ~w26209 & ~w26212;
assign w26214 = ~w26182 & w26205;
assign w26215 = w26213 & w26214;
assign w26216 = w26202 & ~w26203;
assign w26217 = ~w26204 & w26216;
assign w26218 = ~w26196 & w26217;
assign w26219 = ~w26215 & w26218;
assign w26220 = ~w26179 & ~w26182;
assign w26221 = w26171 & w26178;
assign w26222 = w26183 & w26221;
assign w26223 = ~w26171 & w26182;
assign w26224 = ~w26152 & ~w26222;
assign w26225 = ~w26223 & w26224;
assign w26226 = ~w26220 & w26225;
assign w26227 = ~w26202 & w26213;
assign w26228 = ~w26226 & w26227;
assign w26229 = ~w26219 & ~w26228;
assign w26230 = ~w26152 & w26158;
assign w26231 = w26206 & w26230;
assign w26232 = ~w26187 & ~w26231;
assign w26233 = ~w26229 & w26232;
assign w26234 = ~pi1442 & ~w26233;
assign w26235 = pi1442 & w26233;
assign w26236 = ~w26234 & ~w26235;
assign w26237 = ~pi4772 & pi9040;
assign w26238 = ~pi4623 & ~pi9040;
assign w26239 = ~w26237 & ~w26238;
assign w26240 = pi1431 & ~w26239;
assign w26241 = ~pi1431 & w26239;
assign w26242 = ~w26240 & ~w26241;
assign w26243 = ~pi4815 & pi9040;
assign w26244 = ~pi4737 & ~pi9040;
assign w26245 = ~w26243 & ~w26244;
assign w26246 = pi1413 & ~w26245;
assign w26247 = ~pi1413 & w26245;
assign w26248 = ~w26246 & ~w26247;
assign w26249 = ~w26242 & w26248;
assign w26250 = w26242 & ~w26248;
assign w26251 = ~w26249 & ~w26250;
assign w26252 = ~pi4817 & pi9040;
assign w26253 = ~pi4618 & ~pi9040;
assign w26254 = ~w26252 & ~w26253;
assign w26255 = pi1419 & ~w26254;
assign w26256 = ~pi1419 & w26254;
assign w26257 = ~w26255 & ~w26256;
assign w26258 = ~w26242 & ~w26257;
assign w26259 = ~pi4617 & pi9040;
assign w26260 = ~pi4850 & ~pi9040;
assign w26261 = ~w26259 & ~w26260;
assign w26262 = pi1433 & ~w26261;
assign w26263 = ~pi1433 & w26261;
assign w26264 = ~w26262 & ~w26263;
assign w26265 = ~w26258 & ~w26264;
assign w26266 = w26248 & w26264;
assign w26267 = w26258 & w26266;
assign w26268 = ~w26265 & ~w26267;
assign w26269 = ~pi4738 & pi9040;
assign w26270 = ~pi4817 & ~pi9040;
assign w26271 = ~w26269 & ~w26270;
assign w26272 = pi1434 & ~w26271;
assign w26273 = ~pi1434 & w26271;
assign w26274 = ~w26272 & ~w26273;
assign w26275 = ~w26268 & w26274;
assign w26276 = ~w26268 & w65678;
assign w26277 = ~w26242 & w26276;
assign w26278 = ~pi4850 & pi9040;
assign w26279 = ~pi4619 & ~pi9040;
assign w26280 = ~w26278 & ~w26279;
assign w26281 = pi1412 & ~w26280;
assign w26282 = ~pi1412 & w26280;
assign w26283 = ~w26281 & ~w26282;
assign w26284 = ~w26248 & ~w26257;
assign w26285 = ~w26242 & ~w26264;
assign w26286 = ~w26284 & w26285;
assign w26287 = w26264 & ~w26274;
assign w26288 = w26242 & w26287;
assign w26289 = ~w26248 & ~w26264;
assign w26290 = ~w26264 & w26274;
assign w26291 = w26248 & ~w26290;
assign w26292 = ~w26250 & ~w26257;
assign w26293 = ~w26289 & w26292;
assign w26294 = ~w26291 & w26293;
assign w26295 = ~w26249 & ~w26257;
assign w26296 = ~w26249 & ~w26289;
assign w26297 = w26274 & ~w26295;
assign w26298 = ~w26296 & w26297;
assign w26299 = ~w26286 & ~w26288;
assign w26300 = ~w26294 & w26299;
assign w26301 = ~w26298 & w26300;
assign w26302 = (w26283 & ~w26300) | (w26283 & w65679) | (~w26300 & w65679);
assign w26303 = w26264 & w26274;
assign w26304 = ~w26257 & w26264;
assign w26305 = w26250 & ~w26304;
assign w26306 = w26303 & w26305;
assign w26307 = ~w26267 & ~w26306;
assign w26308 = ~w26274 & ~w26304;
assign w26309 = ~w26242 & w26257;
assign w26310 = w26296 & w26309;
assign w26311 = ~w26295 & ~w26310;
assign w26312 = w26308 & ~w26311;
assign w26313 = w26248 & w26257;
assign w26314 = ~w26284 & ~w26313;
assign w26315 = w26242 & ~w26264;
assign w26316 = ~w26291 & w26315;
assign w26317 = ~w26314 & w26316;
assign w26318 = w26307 & ~w26317;
assign w26319 = ~w26312 & w26318;
assign w26320 = ~w26283 & ~w26319;
assign w26321 = w26242 & ~w26284;
assign w26322 = w26304 & w26321;
assign w26323 = w26274 & ~w26283;
assign w26324 = w26321 & w65680;
assign w26325 = w26258 & w26303;
assign w26326 = ~w26266 & ~w26289;
assign w26327 = w26309 & ~w26326;
assign w26328 = ~w26266 & ~w26274;
assign w26329 = w26251 & w26328;
assign w26330 = ~w26327 & ~w26329;
assign w26331 = ~w26274 & ~w26314;
assign w26332 = w26330 & w26331;
assign w26333 = ~w26324 & ~w26325;
assign w26334 = ~w26332 & w26333;
assign w26335 = ~w26277 & w26334;
assign w26336 = ~w26302 & w26335;
assign w26337 = (pi1441 & ~w26336) | (pi1441 & w65681) | (~w26336 & w65681);
assign w26338 = w26336 & w65682;
assign w26339 = ~w26337 & ~w26338;
assign w26340 = ~pi4774 & pi9040;
assign w26341 = ~pi4959 & ~pi9040;
assign w26342 = ~w26340 & ~w26341;
assign w26343 = pi1404 & ~w26342;
assign w26344 = ~pi1404 & w26342;
assign w26345 = ~w26343 & ~w26344;
assign w26346 = ~pi4654 & pi9040;
assign w26347 = ~pi4736 & ~pi9040;
assign w26348 = ~w26346 & ~w26347;
assign w26349 = pi1428 & ~w26348;
assign w26350 = ~pi1428 & w26348;
assign w26351 = ~w26349 & ~w26350;
assign w26352 = w26345 & ~w26351;
assign w26353 = ~pi4831 & pi9040;
assign w26354 = ~pi4608 & ~pi9040;
assign w26355 = ~w26353 & ~w26354;
assign w26356 = pi1431 & ~w26355;
assign w26357 = ~pi1431 & w26355;
assign w26358 = ~w26356 & ~w26357;
assign w26359 = ~pi4692 & pi9040;
assign w26360 = ~pi4612 & ~pi9040;
assign w26361 = ~w26359 & ~w26360;
assign w26362 = pi1423 & ~w26361;
assign w26363 = ~pi1423 & w26361;
assign w26364 = ~w26362 & ~w26363;
assign w26365 = ~w26358 & ~w26364;
assign w26366 = w26345 & w26365;
assign w26367 = (~w26358 & ~w26365) | (~w26358 & w65683) | (~w26365 & w65683);
assign w26368 = ~w26352 & ~w26367;
assign w26369 = w26358 & w26364;
assign w26370 = ~w26345 & w26364;
assign w26371 = ~w26369 & ~w26370;
assign w26372 = ~w26351 & ~w26371;
assign w26373 = ~w26366 & ~w26372;
assign w26374 = w26368 & ~w26373;
assign w26375 = ~w26345 & ~w26364;
assign w26376 = w26351 & ~w26358;
assign w26377 = ~w26345 & ~w26351;
assign w26378 = w26358 & w26377;
assign w26379 = ~w26376 & ~w26378;
assign w26380 = w26375 & w26379;
assign w26381 = ~pi4816 & pi9040;
assign w26382 = ~pi4709 & ~pi9040;
assign w26383 = ~w26381 & ~w26382;
assign w26384 = pi1410 & ~w26383;
assign w26385 = ~pi1410 & w26383;
assign w26386 = ~w26384 & ~w26385;
assign w26387 = (w26386 & w26374) | (w26386 & w65684) | (w26374 & w65684);
assign w26388 = w26345 & w26358;
assign w26389 = ~w26386 & ~w26388;
assign w26390 = ~w26351 & w26364;
assign w26391 = ~w26358 & w26390;
assign w26392 = w26351 & ~w26364;
assign w26393 = ~w26390 & ~w26392;
assign w26394 = ~w26386 & w26393;
assign w26395 = w26393 & w63808;
assign w26396 = (w26389 & w26395) | (w26389 & w65685) | (w26395 & w65685);
assign w26397 = w26345 & w26396;
assign w26398 = ~pi4959 & pi9040;
assign w26399 = ~pi4754 & ~pi9040;
assign w26400 = ~w26398 & ~w26399;
assign w26401 = pi1433 & ~w26400;
assign w26402 = ~pi1433 & w26400;
assign w26403 = ~w26401 & ~w26402;
assign w26404 = ~w26345 & w26393;
assign w26405 = w26388 & w26392;
assign w26406 = ~w26404 & ~w26405;
assign w26407 = (~w26386 & w26404) | (~w26386 & w65686) | (w26404 & w65686);
assign w26408 = w26345 & w26351;
assign w26409 = ~w26369 & w26408;
assign w26410 = ~w26372 & w65687;
assign w26411 = w26386 & ~w26410;
assign w26412 = w26403 & ~w26407;
assign w26413 = ~w26411 & w26412;
assign w26414 = w26369 & w26408;
assign w26415 = w26352 & ~w26358;
assign w26416 = w26386 & ~w26415;
assign w26417 = w26390 & ~w26416;
assign w26418 = w26351 & w26365;
assign w26419 = w26389 & ~w26418;
assign w26420 = w26370 & w26376;
assign w26421 = w26358 & w26375;
assign w26422 = w26386 & ~w26420;
assign w26423 = ~w26421 & w26422;
assign w26424 = ~w26419 & ~w26423;
assign w26425 = ~w26403 & ~w26414;
assign w26426 = ~w26417 & w26425;
assign w26427 = ~w26424 & w26426;
assign w26428 = ~w26413 & ~w26427;
assign w26429 = ~w26387 & ~w26397;
assign w26430 = ~w26428 & w26429;
assign w26431 = pi1443 & ~w26430;
assign w26432 = ~pi1443 & w26430;
assign w26433 = ~w26431 & ~w26432;
assign w26434 = ~pi4733 & pi9040;
assign w26435 = ~pi4675 & ~pi9040;
assign w26436 = ~w26434 & ~w26435;
assign w26437 = pi1411 & ~w26436;
assign w26438 = ~pi1411 & w26436;
assign w26439 = ~w26437 & ~w26438;
assign w26440 = ~pi4675 & pi9040;
assign w26441 = ~pi4831 & ~pi9040;
assign w26442 = ~w26440 & ~w26441;
assign w26443 = pi1424 & ~w26442;
assign w26444 = ~pi1424 & w26442;
assign w26445 = ~w26443 & ~w26444;
assign w26446 = w26439 & w26445;
assign w26447 = ~w26439 & ~w26445;
assign w26448 = ~w26446 & ~w26447;
assign w26449 = ~pi4606 & pi9040;
assign w26450 = ~pi4780 & ~pi9040;
assign w26451 = ~w26449 & ~w26450;
assign w26452 = pi1406 & ~w26451;
assign w26453 = ~pi1406 & w26451;
assign w26454 = ~w26452 & ~w26453;
assign w26455 = ~pi4590 & pi9040;
assign w26456 = ~pi4949 & ~pi9040;
assign w26457 = ~w26455 & ~w26456;
assign w26458 = pi1432 & ~w26457;
assign w26459 = ~pi1432 & w26457;
assign w26460 = ~w26458 & ~w26459;
assign w26461 = ~w26454 & w26460;
assign w26462 = w26454 & ~w26460;
assign w26463 = ~w26461 & ~w26462;
assign w26464 = ~w26448 & ~w26463;
assign w26465 = ~w26439 & ~w26460;
assign w26466 = ~pi4709 & pi9040;
assign w26467 = ~pi4691 & ~pi9040;
assign w26468 = ~w26466 & ~w26467;
assign w26469 = pi1400 & ~w26468;
assign w26470 = ~pi1400 & w26468;
assign w26471 = ~w26469 & ~w26470;
assign w26472 = w26454 & ~w26471;
assign w26473 = ~w26465 & w26472;
assign w26474 = w26439 & w26471;
assign w26475 = w26461 & w26474;
assign w26476 = ~w26439 & ~w26454;
assign w26477 = w26460 & ~w26471;
assign w26478 = w26476 & w26477;
assign w26479 = ~w26475 & ~w26478;
assign w26480 = ~w26439 & w26454;
assign w26481 = ~pi4612 & pi9040;
assign w26482 = ~pi4606 & ~pi9040;
assign w26483 = ~w26481 & ~w26482;
assign w26484 = pi1427 & ~w26483;
assign w26485 = ~pi1427 & w26483;
assign w26486 = ~w26484 & ~w26485;
assign w26487 = (~w26473 & ~w26479) | (~w26473 & w65688) | (~w26479 & w65688);
assign w26488 = ~w26439 & w26471;
assign w26489 = w26463 & w26488;
assign w26490 = (w26445 & ~w26463) | (w26445 & w63810) | (~w26463 & w63810);
assign w26491 = ~w26487 & w26490;
assign w26492 = w26454 & w26474;
assign w26493 = ~w26476 & ~w26492;
assign w26494 = (w26471 & ~w26474) | (w26471 & w63811) | (~w26474 & w63811);
assign w26495 = ~w26473 & ~w26494;
assign w26496 = w26463 & w26493;
assign w26497 = w26495 & w26496;
assign w26498 = ~w26491 & ~w26497;
assign w26499 = ~w26464 & ~w26498;
assign w26500 = ~w26439 & ~w26471;
assign w26501 = w26462 & w26500;
assign w26502 = ~w26489 & ~w26501;
assign w26503 = (~w26460 & w26489) | (~w26460 & w63812) | (w26489 & w63812);
assign w26504 = w26445 & ~w26465;
assign w26505 = (w26504 & ~w26479) | (w26504 & w63813) | (~w26479 & w63813);
assign w26506 = ~w26460 & w26471;
assign w26507 = w26454 & ~w26506;
assign w26508 = w26448 & ~w26476;
assign w26509 = w26448 & w63814;
assign w26510 = (~w26507 & w26509) | (~w26507 & w65689) | (w26509 & w65689);
assign w26511 = ~w26446 & w26454;
assign w26512 = w26477 & ~w26511;
assign w26513 = (~w26445 & w26492) | (~w26445 & w63815) | (w26492 & w63815);
assign w26514 = ~w26512 & w26513;
assign w26515 = w26486 & ~w26503;
assign w26516 = ~w26505 & ~w26514;
assign w26517 = w26515 & w26516;
assign w26518 = ~w26510 & w26517;
assign w26519 = ~w26473 & w26479;
assign w26520 = ~w26445 & ~w26519;
assign w26521 = w26462 & w26488;
assign w26522 = ~w26486 & ~w26521;
assign w26523 = ~w26520 & w26522;
assign w26524 = ~w26518 & ~w26523;
assign w26525 = ~w26524 & w65690;
assign w26526 = (pi1452 & w26524) | (pi1452 & w65691) | (w26524 & w65691);
assign w26527 = ~w26525 & ~w26526;
assign w26528 = ~w26463 & w26509;
assign w26529 = w26486 & ~w26528;
assign w26530 = w26439 & w26477;
assign w26531 = ~w26454 & w26530;
assign w26532 = ~w26500 & ~w26506;
assign w26533 = w26490 & ~w26532;
assign w26534 = ~w26531 & ~w26533;
assign w26535 = ~w26510 & w26534;
assign w26536 = ~w26529 & ~w26535;
assign w26537 = w26447 & w26463;
assign w26538 = ~w26480 & w26504;
assign w26539 = ~w26530 & w26538;
assign w26540 = ~w26537 & ~w26539;
assign w26541 = ~w26493 & ~w26494;
assign w26542 = ~w26540 & w26541;
assign w26543 = w26460 & ~w26474;
assign w26544 = ~w26500 & w26543;
assign w26545 = (~w26486 & ~w26543) | (~w26486 & w65692) | (~w26543 & w65692);
assign w26546 = ~w26495 & ~w26544;
assign w26547 = w26486 & ~w26546;
assign w26548 = ~w26445 & ~w26545;
assign w26549 = ~w26547 & w26548;
assign w26550 = (~w26488 & ~w26534) | (~w26488 & w65693) | (~w26534 & w65693);
assign w26551 = w26445 & w26547;
assign w26552 = ~w26550 & w26551;
assign w26553 = ~w26542 & ~w26549;
assign w26554 = ~w26536 & w26553;
assign w26555 = w26554 & w65694;
assign w26556 = (pi1449 & ~w26554) | (pi1449 & w65695) | (~w26554 & w65695);
assign w26557 = ~w26555 & ~w26556;
assign w26558 = ~pi4734 & pi9040;
assign w26559 = ~pi4617 & ~pi9040;
assign w26560 = ~w26558 & ~w26559;
assign w26561 = pi1421 & ~w26560;
assign w26562 = ~pi1421 & w26560;
assign w26563 = ~w26561 & ~w26562;
assign w26564 = ~pi4619 & pi9040;
assign w26565 = ~pi4839 & ~pi9040;
assign w26566 = ~w26564 & ~w26565;
assign w26567 = pi1420 & ~w26566;
assign w26568 = ~pi1420 & w26566;
assign w26569 = ~w26567 & ~w26568;
assign w26570 = ~w26563 & ~w26569;
assign w26571 = ~pi4947 & pi9040;
assign w26572 = ~pi4652 & ~pi9040;
assign w26573 = ~w26571 & ~w26572;
assign w26574 = pi1429 & ~w26573;
assign w26575 = ~pi1429 & w26573;
assign w26576 = ~w26574 & ~w26575;
assign w26577 = ~pi4690 & pi9040;
assign w26578 = ~pi4772 & ~pi9040;
assign w26579 = ~w26577 & ~w26578;
assign w26580 = pi1418 & ~w26579;
assign w26581 = ~pi1418 & w26579;
assign w26582 = ~w26580 & ~w26581;
assign w26583 = ~w26576 & w26582;
assign w26584 = ~pi4737 & pi9040;
assign w26585 = ~pi4947 & ~pi9040;
assign w26586 = ~w26584 & ~w26585;
assign w26587 = pi1430 & ~w26586;
assign w26588 = ~pi1430 & w26586;
assign w26589 = ~w26587 & ~w26588;
assign w26590 = ~w26563 & ~w26576;
assign w26591 = w26569 & w26590;
assign w26592 = w26590 & w63394;
assign w26593 = w26589 & ~w26592;
assign w26594 = (w26583 & w26592) | (w26583 & w65696) | (w26592 & w65696);
assign w26595 = ~w26569 & ~w26582;
assign w26596 = w26576 & w26595;
assign w26597 = ~w26594 & ~w26596;
assign w26598 = w26570 & ~w26597;
assign w26599 = w26563 & ~w26569;
assign w26600 = w26582 & ~w26599;
assign w26601 = (~w26589 & w26599) | (~w26589 & w63816) | (w26599 & w63816);
assign w26602 = w26563 & ~w26589;
assign w26603 = ~w26569 & ~w26576;
assign w26604 = ~w26582 & w26603;
assign w26605 = ~w26602 & ~w26604;
assign w26606 = ~w26601 & ~w26605;
assign w26607 = w26569 & ~w26582;
assign w26608 = ~w26569 & w26582;
assign w26609 = ~w26607 & ~w26608;
assign w26610 = w26582 & w26589;
assign w26611 = ~w26576 & ~w26610;
assign w26612 = w26563 & ~w26609;
assign w26613 = ~w26611 & w26612;
assign w26614 = ~w26606 & ~w26613;
assign w26615 = ~w26598 & w26614;
assign w26616 = ~pi4610 & pi9040;
assign w26617 = ~pi4707 & ~pi9040;
assign w26618 = ~w26616 & ~w26617;
assign w26619 = pi1436 & ~w26618;
assign w26620 = ~pi1436 & w26618;
assign w26621 = ~w26619 & ~w26620;
assign w26622 = ~w26615 & w26621;
assign w26623 = ~w26563 & w26576;
assign w26624 = w26608 & w26623;
assign w26625 = w26576 & w26589;
assign w26626 = w26607 & w26625;
assign w26627 = ~w26624 & ~w26626;
assign w26628 = ~w26591 & w26627;
assign w26629 = ~w26610 & w26621;
assign w26630 = ~w26628 & ~w26629;
assign w26631 = ~w26576 & w26601;
assign w26632 = w26563 & ~w26608;
assign w26633 = w26625 & w26632;
assign w26634 = ~w26631 & ~w26633;
assign w26635 = ~w26621 & ~w26634;
assign w26636 = ~w26589 & ~w26624;
assign w26637 = ~w26563 & w26607;
assign w26638 = ~w26623 & ~w26637;
assign w26639 = w26576 & w26607;
assign w26640 = w26636 & ~w26639;
assign w26641 = ~w26638 & w26640;
assign w26642 = ~w26630 & ~w26641;
assign w26643 = ~w26635 & w26642;
assign w26644 = ~w26622 & w26643;
assign w26645 = pi1444 & ~w26644;
assign w26646 = ~pi1444 & w26644;
assign w26647 = ~w26645 & ~w26646;
assign w26648 = ~pi4707 & pi9040;
assign w26649 = ~pi4794 & ~pi9040;
assign w26650 = ~w26648 & ~w26649;
assign w26651 = pi1413 & ~w26650;
assign w26652 = ~pi1413 & w26650;
assign w26653 = ~w26651 & ~w26652;
assign w26654 = ~pi4839 & pi9040;
assign w26655 = ~pi4605 & ~pi9040;
assign w26656 = ~w26654 & ~w26655;
assign w26657 = pi1412 & ~w26656;
assign w26658 = ~pi1412 & w26656;
assign w26659 = ~w26657 & ~w26658;
assign w26660 = w26653 & ~w26659;
assign w26661 = ~pi4716 & pi9040;
assign w26662 = ~pi4613 & ~pi9040;
assign w26663 = ~w26661 & ~w26662;
assign w26664 = pi1416 & ~w26663;
assign w26665 = ~pi1416 & w26663;
assign w26666 = ~w26664 & ~w26665;
assign w26667 = ~w26660 & ~w26666;
assign w26668 = ~pi4699 & pi9040;
assign w26669 = ~pi4620 & ~pi9040;
assign w26670 = ~w26668 & ~w26669;
assign w26671 = pi1426 & ~w26670;
assign w26672 = ~pi1426 & w26670;
assign w26673 = ~w26671 & ~w26672;
assign w26674 = w26653 & ~w26673;
assign w26675 = w26659 & ~w26674;
assign w26676 = ~pi4794 & pi9040;
assign w26677 = ~pi4690 & ~pi9040;
assign w26678 = ~w26676 & ~w26677;
assign w26679 = pi1435 & ~w26678;
assign w26680 = ~pi1435 & w26678;
assign w26681 = ~w26679 & ~w26680;
assign w26682 = ~w26675 & w26681;
assign w26683 = ~w26653 & w26673;
assign w26684 = w26659 & w26683;
assign w26685 = ~w26659 & ~w26673;
assign w26686 = ~w26684 & ~w26685;
assign w26687 = ~w26653 & ~w26673;
assign w26688 = w26681 & w26687;
assign w26689 = ~pi4613 & pi9040;
assign w26690 = ~pi4607 & ~pi9040;
assign w26691 = ~w26689 & ~w26690;
assign w26692 = pi1415 & ~w26691;
assign w26693 = ~pi1415 & w26691;
assign w26694 = ~w26692 & ~w26693;
assign w26695 = ~w26688 & ~w26694;
assign w26696 = w26686 & w26695;
assign w26697 = ~w26682 & ~w26696;
assign w26698 = w26667 & ~w26697;
assign w26699 = ~w26666 & ~w26683;
assign w26700 = ~w26659 & ~w26681;
assign w26701 = w26673 & w26681;
assign w26702 = ~w26659 & w26701;
assign w26703 = ~w26700 & ~w26702;
assign w26704 = w26699 & ~w26703;
assign w26705 = ~w26674 & ~w26683;
assign w26706 = w26659 & w26681;
assign w26707 = ~w26705 & w26706;
assign w26708 = ~w26659 & w26705;
assign w26709 = ~w26699 & ~w26700;
assign w26710 = ~w26707 & w26709;
assign w26711 = ~w26708 & w26710;
assign w26712 = w26694 & ~w26704;
assign w26713 = ~w26711 & w26712;
assign w26714 = ~w26694 & ~w26707;
assign w26715 = ~w26659 & w26681;
assign w26716 = w26687 & w26715;
assign w26717 = w26666 & ~w26683;
assign w26718 = ~w26703 & w26717;
assign w26719 = w26714 & ~w26716;
assign w26720 = ~w26718 & w26719;
assign w26721 = ~w26713 & ~w26720;
assign w26722 = ~w26698 & ~w26721;
assign w26723 = ~pi1447 & w26722;
assign w26724 = pi1447 & ~w26722;
assign w26725 = ~w26723 & ~w26724;
assign w26726 = ~w26604 & ~w26639;
assign w26727 = ~w26563 & ~w26726;
assign w26728 = w26627 & w63328;
assign w26729 = w26589 & ~w26728;
assign w26730 = ~w26727 & w26729;
assign w26731 = ~w26636 & ~w26730;
assign w26732 = w26563 & w26576;
assign w26733 = w26595 & w26732;
assign w26734 = ~w26621 & ~w26733;
assign w26735 = ~w26570 & ~w26607;
assign w26736 = w26625 & w26735;
assign w26737 = w26602 & ~w26607;
assign w26738 = ~w26605 & ~w26737;
assign w26739 = ~w26736 & ~w26738;
assign w26740 = ~w26738 & w65697;
assign w26741 = w26734 & w26740;
assign w26742 = w26600 & w26732;
assign w26743 = w26739 & w63817;
assign w26744 = ~w26570 & ~w26590;
assign w26745 = ~w26589 & ~w26603;
assign w26746 = ~w26744 & w26745;
assign w26747 = w26621 & w26627;
assign w26748 = ~w26742 & ~w26746;
assign w26749 = w26747 & w26748;
assign w26750 = ~w26743 & w26749;
assign w26751 = ~w26741 & ~w26750;
assign w26752 = ~w26751 & w65698;
assign w26753 = (pi1446 & w26751) | (pi1446 & w65699) | (w26751 & w65699);
assign w26754 = ~w26752 & ~w26753;
assign w26755 = w26583 & w26599;
assign w26756 = ~w26742 & ~w26755;
assign w26757 = w26607 & ~w26623;
assign w26758 = w26636 & ~w26757;
assign w26759 = w26593 & ~w26596;
assign w26760 = ~w26758 & ~w26759;
assign w26761 = w26756 & ~w26760;
assign w26762 = ~w26760 & w65700;
assign w26763 = w26570 & w26610;
assign w26764 = w26569 & w26614;
assign w26765 = w26761 & w26764;
assign w26766 = w26734 & ~w26763;
assign w26767 = (w26729 & w63818) | (w26729 & w63819) | (w63818 & w63819);
assign w26768 = ~w26765 & w26767;
assign w26769 = ~w26589 & ~w26637;
assign w26770 = ~w26727 & w26756;
assign w26771 = ~w26599 & ~w26637;
assign w26772 = w26625 & ~w26771;
assign w26773 = (~w26772 & w26770) | (~w26772 & w65701) | (w26770 & w65701);
assign w26774 = (~w26768 & w65702) | (~w26768 & w65703) | (w65702 & w65703);
assign w26775 = (w26768 & w65704) | (w26768 & w65705) | (w65704 & w65705);
assign w26776 = ~w26774 & ~w26775;
assign w26777 = w26164 & ~w26178;
assign w26778 = ~w26195 & w26777;
assign w26779 = w26165 & w26171;
assign w26780 = ~w26223 & ~w26779;
assign w26781 = w26178 & ~w26780;
assign w26782 = ~w26152 & w26203;
assign w26783 = w26158 & w26171;
assign w26784 = ~w26204 & ~w26783;
assign w26785 = w26152 & ~w26784;
assign w26786 = w26202 & ~w26782;
assign w26787 = ~w26781 & w26786;
assign w26788 = ~w26778 & w26787;
assign w26789 = ~w26785 & w26788;
assign w26790 = ~w26202 & ~w26222;
assign w26791 = ~w26178 & ~w26780;
assign w26792 = w26152 & ~w26181;
assign w26793 = ~w26184 & ~w26221;
assign w26794 = ~w26792 & ~w26793;
assign w26795 = w26190 & w26207;
assign w26796 = w26790 & ~w26795;
assign w26797 = ~w26791 & w26796;
assign w26798 = ~w26794 & w26797;
assign w26799 = ~w26789 & ~w26798;
assign w26800 = ~pi1440 & w26799;
assign w26801 = pi1440 & ~w26799;
assign w26802 = ~w26800 & ~w26801;
assign w26803 = ~w26301 & w26315;
assign w26804 = w26242 & w26313;
assign w26805 = w26283 & ~w26804;
assign w26806 = w26250 & w26304;
assign w26807 = ~w26265 & w26308;
assign w26808 = w26805 & ~w26806;
assign w26809 = ~w26807 & w26808;
assign w26810 = ~w26275 & w26809;
assign w26811 = w26251 & w26264;
assign w26812 = w26274 & w26811;
assign w26813 = ~w26274 & ~w26321;
assign w26814 = ~w26326 & w26813;
assign w26815 = ~w26251 & w26326;
assign w26816 = w26257 & w26815;
assign w26817 = ~w26283 & ~w26812;
assign w26818 = ~w26814 & ~w26816;
assign w26819 = w26817 & w26818;
assign w26820 = ~w26810 & ~w26819;
assign w26821 = ~w26803 & ~w26820;
assign w26822 = ~pi1451 & w26821;
assign w26823 = pi1451 & ~w26821;
assign w26824 = ~w26822 & ~w26823;
assign w26825 = ~w26681 & w26687;
assign w26826 = (w26666 & ~w26687) | (w26666 & w65706) | (~w26687 & w65706);
assign w26827 = ~w26683 & ~w26706;
assign w26828 = ~w26660 & w26827;
assign w26829 = w26826 & w26828;
assign w26830 = ~w26666 & w26681;
assign w26831 = (w26830 & w26684) | (w26830 & w65707) | (w26684 & w65707);
assign w26832 = w26653 & w26666;
assign w26833 = ~w26715 & w26832;
assign w26834 = w26667 & w26685;
assign w26835 = ~w26674 & w63821;
assign w26836 = ~w26683 & w26835;
assign w26837 = ~w26660 & ~w26700;
assign w26838 = w26653 & ~w26830;
assign w26839 = ~w26837 & ~w26838;
assign w26840 = ~w26666 & ~w26701;
assign w26841 = w26683 & w26840;
assign w26842 = w26701 & w26660;
assign w26843 = ~w26841 & ~w26842;
assign w26844 = w26839 & ~w26843;
assign w26845 = w26694 & ~w26833;
assign w26846 = ~w26834 & w26845;
assign w26847 = w26846 & w65708;
assign w26848 = ~w26844 & w26847;
assign w26849 = ~w26675 & ~w26705;
assign w26850 = ~w26681 & w26849;
assign w26851 = (~w26666 & ~w26683) | (~w26666 & w65709) | (~w26683 & w65709);
assign w26852 = ~w26827 & w26851;
assign w26853 = ~w26702 & w26826;
assign w26854 = w26674 & w26700;
assign w26855 = ~w26701 & ~w26854;
assign w26856 = w26853 & ~w26855;
assign w26857 = w26683 & w26856;
assign w26858 = ~w26841 & w65710;
assign w26859 = ~w26850 & ~w26852;
assign w26860 = w26858 & w26859;
assign w26861 = ~w26857 & w26860;
assign w26862 = (~w26829 & w26861) | (~w26829 & w65711) | (w26861 & w65711);
assign w26863 = pi1458 & ~w26862;
assign w26864 = ~pi1458 & w26862;
assign w26865 = ~w26863 & ~w26864;
assign w26866 = ~w26461 & w26509;
assign w26867 = ~w26497 & ~w26866;
assign w26868 = w26464 & ~w26472;
assign w26869 = ~w26497 & w65712;
assign w26870 = ~w26486 & ~w26869;
assign w26871 = ~w26475 & w26490;
assign w26872 = ~w26454 & w26500;
assign w26873 = w26463 & w26474;
assign w26874 = ~w26445 & ~w26872;
assign w26875 = ~w26873 & w26874;
assign w26876 = ~w26871 & ~w26875;
assign w26877 = ~w26445 & ~w26471;
assign w26878 = ~w26478 & ~w26877;
assign w26879 = ~w26507 & w26878;
assign w26880 = w26486 & ~w26879;
assign w26881 = (~w26876 & ~w26867) | (~w26876 & w65713) | (~w26867 & w65713);
assign w26882 = ~w26870 & w26881;
assign w26883 = pi1466 & w26882;
assign w26884 = ~pi1466 & ~w26882;
assign w26885 = ~w26883 & ~w26884;
assign w26886 = ~pi4608 & pi9040;
assign w26887 = ~pi4937 & ~pi9040;
assign w26888 = ~w26886 & ~w26887;
assign w26889 = pi1411 & ~w26888;
assign w26890 = ~pi1411 & w26888;
assign w26891 = ~w26889 & ~w26890;
assign w26892 = ~pi4781 & pi9040;
assign w26893 = ~pi4958 & ~pi9040;
assign w26894 = ~w26892 & ~w26893;
assign w26895 = pi1436 & ~w26894;
assign w26896 = ~pi1436 & w26894;
assign w26897 = ~w26895 & ~w26896;
assign w26898 = ~pi4949 & pi9040;
assign w26899 = ~pi4774 & ~pi9040;
assign w26900 = ~w26898 & ~w26899;
assign w26901 = pi1432 & ~w26900;
assign w26902 = ~pi1432 & w26900;
assign w26903 = ~w26901 & ~w26902;
assign w26904 = w26897 & ~w26903;
assign w26905 = ~pi4883 & pi9040;
assign w26906 = ~pi4695 & ~pi9040;
assign w26907 = ~w26905 & ~w26906;
assign w26908 = pi1418 & ~w26907;
assign w26909 = ~pi1418 & w26907;
assign w26910 = ~w26908 & ~w26909;
assign w26911 = w26904 & w26910;
assign w26912 = ~w26897 & ~w26910;
assign w26913 = ~w26903 & w26912;
assign w26914 = ~w26911 & ~w26913;
assign w26915 = ~pi4710 & pi9040;
assign w26916 = ~pi4692 & ~pi9040;
assign w26917 = ~w26915 & ~w26916;
assign w26918 = pi1439 & ~w26917;
assign w26919 = ~pi1439 & w26917;
assign w26920 = ~w26918 & ~w26919;
assign w26921 = ~w26914 & w26920;
assign w26922 = ~w26897 & ~w26920;
assign w26923 = w26910 & w26922;
assign w26924 = ~w26897 & w26920;
assign w26925 = w26910 & ~w26924;
assign w26926 = w26897 & w26920;
assign w26927 = ~w26903 & ~w26926;
assign w26928 = ~w26925 & w26927;
assign w26929 = ~pi4736 & pi9040;
assign w26930 = ~pi4883 & ~pi9040;
assign w26931 = ~w26929 & ~w26930;
assign w26932 = pi1405 & ~w26931;
assign w26933 = ~pi1405 & w26931;
assign w26934 = ~w26932 & ~w26933;
assign w26935 = w26897 & w26903;
assign w26936 = w26910 & w26935;
assign w26937 = ~w26928 & w65714;
assign w26938 = (~w26934 & ~w26935) | (~w26934 & w65715) | (~w26935 & w65715);
assign w26939 = w26903 & w26910;
assign w26940 = w26903 & ~w26920;
assign w26941 = ~w26939 & ~w26940;
assign w26942 = ~w26897 & ~w26941;
assign w26943 = ~w26897 & w26934;
assign w26944 = (~w26943 & w26942) | (~w26943 & w65716) | (w26942 & w65716);
assign w26945 = ~w26937 & w26944;
assign w26946 = ~w26921 & ~w26923;
assign w26947 = ~w26945 & w26946;
assign w26948 = ~w26891 & ~w26947;
assign w26949 = ~w26910 & w26926;
assign w26950 = ~w26934 & w26949;
assign w26951 = ~w26920 & w26943;
assign w26952 = ~w26950 & ~w26951;
assign w26953 = ~w26903 & w26934;
assign w26954 = ~w26904 & ~w26910;
assign w26955 = w26922 & ~w26934;
assign w26956 = w26954 & ~w26955;
assign w26957 = ~w26953 & ~w26956;
assign w26958 = ~w26952 & w26957;
assign w26959 = ~w26903 & ~w26910;
assign w26960 = ~w26939 & ~w26959;
assign w26961 = w26920 & ~w26935;
assign w26962 = w26934 & w26961;
assign w26963 = w26891 & w26924;
assign w26964 = ~w26962 & ~w26963;
assign w26965 = w26960 & ~w26964;
assign w26966 = (w26934 & ~w26922) | (w26934 & w26953) | (~w26922 & w26953);
assign w26967 = w26891 & ~w26924;
assign w26968 = w26954 & w26967;
assign w26969 = w26966 & w26968;
assign w26970 = w26897 & ~w26920;
assign w26971 = w26891 & ~w26934;
assign w26972 = w26970 & w26971;
assign w26973 = ~w26969 & ~w26972;
assign w26974 = ~w26958 & w26973;
assign w26975 = ~w26965 & w26974;
assign w26976 = ~w26948 & w26975;
assign w26977 = pi1448 & ~w26976;
assign w26978 = ~pi1448 & w26976;
assign w26979 = ~w26977 & ~w26978;
assign w26980 = w26921 & w26934;
assign w26981 = ~w26923 & w26938;
assign w26982 = ~w26912 & w26937;
assign w26983 = w26891 & ~w26981;
assign w26984 = ~w26982 & w26983;
assign w26985 = w26953 & w26970;
assign w26986 = ~w26951 & ~w26985;
assign w26987 = w26891 & w26910;
assign w26988 = w26960 & ~w26987;
assign w26989 = ~w26986 & w26988;
assign w26990 = ~w26920 & w26936;
assign w26991 = ~w26904 & ~w26940;
assign w26992 = ~w26922 & w26927;
assign w26993 = w26987 & ~w26991;
assign w26994 = ~w26992 & w26993;
assign w26995 = ~w26891 & ~w26925;
assign w26996 = w26957 & w26995;
assign w26997 = ~w26950 & ~w26990;
assign w26998 = ~w26989 & w26997;
assign w26999 = ~w26994 & w26998;
assign w27000 = ~w26980 & ~w26996;
assign w27001 = w26999 & w27000;
assign w27002 = ~w26984 & w27001;
assign w27003 = ~pi1445 & w27002;
assign w27004 = pi1445 & ~w27002;
assign w27005 = ~w27003 & ~w27004;
assign w27006 = ~pi4685 & pi9040;
assign w27007 = ~pi4699 & ~pi9040;
assign w27008 = ~w27006 & ~w27007;
assign w27009 = pi1415 & ~w27008;
assign w27010 = ~pi1415 & w27008;
assign w27011 = ~w27009 & ~w27010;
assign w27012 = ~pi4607 & pi9040;
assign w27013 = ~pi4685 & ~pi9040;
assign w27014 = ~w27012 & ~w27013;
assign w27015 = pi1429 & ~w27014;
assign w27016 = ~pi1429 & w27014;
assign w27017 = ~w27015 & ~w27016;
assign w27018 = ~w27011 & ~w27017;
assign w27019 = ~pi4611 & pi9040;
assign w27020 = ~pi4734 & ~pi9040;
assign w27021 = ~w27019 & ~w27020;
assign w27022 = pi1422 & ~w27021;
assign w27023 = ~pi1422 & w27021;
assign w27024 = ~w27022 & ~w27023;
assign w27025 = ~pi4891 & pi9040;
assign w27026 = ~pi4716 & ~pi9040;
assign w27027 = ~w27025 & ~w27026;
assign w27028 = pi1426 & ~w27027;
assign w27029 = ~pi1426 & w27027;
assign w27030 = ~w27028 & ~w27029;
assign w27031 = w27024 & w27030;
assign w27032 = ~pi4618 & pi9040;
assign w27033 = ~pi4610 & ~pi9040;
assign w27034 = ~w27032 & ~w27033;
assign w27035 = pi1420 & ~w27034;
assign w27036 = ~pi1420 & w27034;
assign w27037 = ~w27035 & ~w27036;
assign w27038 = w27031 & w27037;
assign w27039 = w27018 & w27038;
assign w27040 = ~w27011 & w27017;
assign w27041 = w27011 & ~w27017;
assign w27042 = ~w27040 & ~w27041;
assign w27043 = ~w27030 & w27042;
assign w27044 = w27030 & w27041;
assign w27045 = ~w27043 & ~w27044;
assign w27046 = w27024 & ~w27045;
assign w27047 = ~w27024 & w27030;
assign w27048 = ~pi4623 & pi9040;
assign w27049 = ~pi4891 & ~pi9040;
assign w27050 = ~w27048 & ~w27049;
assign w27051 = pi1395 & ~w27050;
assign w27052 = ~pi1395 & w27050;
assign w27053 = ~w27051 & ~w27052;
assign w27054 = w27017 & w27053;
assign w27055 = (w27047 & w27042) | (w27047 & w63822) | (w27042 & w63822);
assign w27056 = ~w27024 & ~w27030;
assign w27057 = ~w27042 & w63823;
assign w27058 = w27024 & w27040;
assign w27059 = ~w27017 & w27030;
assign w27060 = w27011 & w27024;
assign w27061 = ~w27059 & ~w27060;
assign w27062 = ~w27011 & ~w27030;
assign w27063 = ~w27053 & ~w27062;
assign w27064 = w27061 & w27063;
assign w27065 = w27058 & w27064;
assign w27066 = ~w27055 & ~w27057;
assign w27067 = ~w27065 & w27066;
assign w27068 = ~w27046 & w27067;
assign w27069 = ~w27037 & ~w27068;
assign w27070 = w27017 & ~w27030;
assign w27071 = w27024 & w27070;
assign w27072 = w27053 & ~w27071;
assign w27073 = w27018 & w27056;
assign w27074 = w27072 & ~w27073;
assign w27075 = ~w27044 & ~w27058;
assign w27076 = ~w27070 & w27075;
assign w27077 = ~w27018 & w27037;
assign w27078 = w27075 & w65717;
assign w27079 = ~w27053 & ~w27078;
assign w27080 = ~w27074 & ~w27079;
assign w27081 = w27037 & w27053;
assign w27082 = ~w27076 & w27081;
assign w27083 = ~w27039 & ~w27082;
assign w27084 = ~w27080 & w27083;
assign w27085 = ~w27069 & w27084;
assign w27086 = ~pi1461 & w27085;
assign w27087 = pi1461 & ~w27085;
assign w27088 = ~w27086 & ~w27087;
assign w27089 = ~w26460 & w26508;
assign w27090 = w26486 & ~w26512;
assign w27091 = w26502 & w27090;
assign w27092 = ~w27089 & w27091;
assign w27093 = w26460 & w26492;
assign w27094 = ~w26486 & ~w27093;
assign w27095 = w26540 & w27094;
assign w27096 = ~w27092 & ~w27095;
assign w27097 = ~w26528 & ~w27096;
assign w27098 = ~pi1468 & w27097;
assign w27099 = pi1468 & ~w27097;
assign w27100 = ~w27098 & ~w27099;
assign w27101 = w26288 & w26313;
assign w27102 = w26250 & w26290;
assign w27103 = ~w26274 & w26815;
assign w27104 = ~w27102 & ~w27103;
assign w27105 = ~w26257 & ~w27104;
assign w27106 = ~w26287 & ~w26290;
assign w27107 = w26313 & ~w27106;
assign w27108 = w26251 & ~w26314;
assign w27109 = ~w26283 & ~w26288;
assign w27110 = ~w27102 & w27109;
assign w27111 = ~w27107 & ~w27108;
assign w27112 = w27110 & w27111;
assign w27113 = ~w26251 & ~w26264;
assign w27114 = ~w26310 & ~w27113;
assign w27115 = ~w26274 & ~w27114;
assign w27116 = ~w26306 & w65718;
assign w27117 = ~w26276 & w27116;
assign w27118 = ~w27115 & w27117;
assign w27119 = ~w27112 & ~w27118;
assign w27120 = ~w26325 & ~w27101;
assign w27121 = ~w27105 & w27120;
assign w27122 = ~w27119 & w27121;
assign w27123 = pi1459 & ~w27122;
assign w27124 = ~pi1459 & w27122;
assign w27125 = ~w27123 & ~w27124;
assign w27126 = ~w26191 & w65719;
assign w27127 = ~w26222 & ~w27126;
assign w27128 = ~w26178 & w26191;
assign w27129 = w26191 & w65720;
assign w27130 = w26152 & ~w27129;
assign w27131 = (~w26152 & ~w26181) | (~w26152 & w65721) | (~w26181 & w65721);
assign w27132 = ~w26189 & ~w26210;
assign w27133 = ~w26193 & ~w27132;
assign w27134 = ~w26192 & w27131;
assign w27135 = ~w27133 & w27134;
assign w27136 = (w27127 & w27135) | (w27127 & w65722) | (w27135 & w65722);
assign w27137 = w26202 & ~w27136;
assign w27138 = w26790 & ~w27128;
assign w27139 = ~w27126 & w27138;
assign w27140 = w26180 & ~w27139;
assign w27141 = ~w26179 & ~w27129;
assign w27142 = ~w26202 & ~w27141;
assign w27143 = ~w26152 & w27127;
assign w27144 = ~w27142 & w27143;
assign w27145 = ~w27140 & ~w27144;
assign w27146 = ~w27137 & ~w27145;
assign w27147 = ~pi1462 & w27146;
assign w27148 = pi1462 & ~w27146;
assign w27149 = ~w27147 & ~w27148;
assign w27150 = w27042 & w27056;
assign w27151 = w27075 & ~w27150;
assign w27152 = ~w27053 & ~w27151;
assign w27153 = ~w27017 & ~w27024;
assign w27154 = w27011 & w27017;
assign w27155 = w27030 & w27154;
assign w27156 = ~w27153 & ~w27155;
assign w27157 = w27011 & ~w27156;
assign w27158 = ~w27041 & ~w27053;
assign w27159 = w27151 & ~w27158;
assign w27160 = ~w27157 & w27159;
assign w27161 = (~w27037 & w27160) | (~w27037 & w65723) | (w27160 & w65723);
assign w27162 = ~w27018 & w27053;
assign w27163 = ~w27155 & w27162;
assign w27164 = ~w27067 & w27163;
assign w27165 = ~w27031 & ~w27037;
assign w27166 = ~w27040 & ~w27056;
assign w27167 = w27158 & w27166;
assign w27168 = ~w27057 & ~w27167;
assign w27169 = w27017 & w27062;
assign w27170 = (w27158 & ~w27156) | (w27158 & w63824) | (~w27156 & w63824);
assign w27171 = ~w27037 & ~w27170;
assign w27172 = ~w27165 & ~w27168;
assign w27173 = ~w27171 & w27172;
assign w27174 = ~w27047 & w27081;
assign w27175 = (w27174 & ~w27159) | (w27174 & w65724) | (~w27159 & w65724);
assign w27176 = ~w27164 & ~w27173;
assign w27177 = ~w27175 & w27176;
assign w27178 = (pi1454 & ~w27177) | (pi1454 & w65725) | (~w27177 & w65725);
assign w27179 = w27177 & w65726;
assign w27180 = ~w27178 & ~w27179;
assign w27181 = ~w26811 & ~w27113;
assign w27182 = w26257 & ~w27181;
assign w27183 = ~w26322 & w26330;
assign w27184 = w26295 & w27114;
assign w27185 = w27183 & w27184;
assign w27186 = (w26283 & w27185) | (w26283 & w65727) | (w27185 & w65727);
assign w27187 = ~w26288 & w26805;
assign w27188 = ~w26249 & ~w26305;
assign w27189 = w26323 & ~w27188;
assign w27190 = w27183 & ~w27189;
assign w27191 = ~w27187 & ~w27190;
assign w27192 = ~w27186 & ~w27191;
assign w27193 = ~pi1471 & w27192;
assign w27194 = pi1471 & ~w27192;
assign w27195 = ~w27193 & ~w27194;
assign w27196 = ~w26949 & ~w26955;
assign w27197 = ~w26960 & ~w27196;
assign w27198 = w26920 & w26935;
assign w27199 = w26938 & w27198;
assign w27200 = w26960 & w26970;
assign w27201 = ~w26913 & ~w26923;
assign w27202 = ~w27198 & w27201;
assign w27203 = ~w26928 & w65728;
assign w27204 = w27202 & w27203;
assign w27205 = ~w27197 & w65729;
assign w27206 = ~w27204 & w27205;
assign w27207 = w26891 & ~w27206;
assign w27208 = (~w26891 & ~w27201) | (~w26891 & w65730) | (~w27201 & w65730);
assign w27209 = ~w26914 & w26992;
assign w27210 = ~w27208 & ~w27209;
assign w27211 = w26934 & ~w27210;
assign w27212 = ~w26960 & ~w26970;
assign w27213 = ~w26934 & ~w26967;
assign w27214 = ~w27200 & w27213;
assign w27215 = ~w27212 & w27214;
assign w27216 = ~w27211 & ~w27215;
assign w27217 = ~w27207 & w27216;
assign w27218 = pi1456 & w27217;
assign w27219 = ~pi1456 & ~w27217;
assign w27220 = ~w27218 & ~w27219;
assign w27221 = ~w26345 & w26351;
assign w27222 = w26358 & ~w26386;
assign w27223 = ~w26369 & ~w27222;
assign w27224 = w27221 & ~w27223;
assign w27225 = ~w26345 & w26386;
assign w27226 = ~w26408 & ~w27225;
assign w27227 = w26365 & ~w27226;
assign w27228 = w26352 & w26364;
assign w27229 = ~w27227 & ~w27228;
assign w27230 = w26403 & ~w27224;
assign w27231 = w27229 & w27230;
assign w27232 = ~w26389 & ~w26391;
assign w27233 = w26345 & w26364;
assign w27234 = ~w26415 & ~w27233;
assign w27235 = ~w26421 & w27234;
assign w27236 = (w26386 & ~w27234) | (w26386 & w65731) | (~w27234 & w65731);
assign w27237 = (~w26403 & w27232) | (~w26403 & w65732) | (w27232 & w65732);
assign w27238 = ~w27236 & w27237;
assign w27239 = ~w27231 & ~w27238;
assign w27240 = ~w26388 & ~w26408;
assign w27241 = ~w26372 & w63825;
assign w27242 = (w26386 & w27241) | (w26386 & w65733) | (w27241 & w65733);
assign w27243 = ~w26406 & w27242;
assign w27244 = w26366 & ~w26386;
assign w27245 = ~w26394 & ~w27244;
assign w27246 = w27235 & ~w27245;
assign w27247 = ~w27239 & ~w27246;
assign w27248 = ~w27243 & w27247;
assign w27249 = pi1492 & ~w27248;
assign w27250 = ~pi1492 & w27248;
assign w27251 = ~w27249 & ~w27250;
assign w27252 = w26602 & ~w26726;
assign w27253 = w26569 & w26583;
assign w27254 = w26769 & ~w27253;
assign w27255 = w26570 & ~w26582;
assign w27256 = ~w26728 & w63826;
assign w27257 = ~w26609 & w26623;
assign w27258 = ~w26742 & ~w27257;
assign w27259 = (w27258 & w27256) | (w27258 & w65734) | (w27256 & w65734);
assign w27260 = ~w26621 & ~w27259;
assign w27261 = (w26589 & w26591) | (w26589 & w65735) | (w26591 & w65735);
assign w27262 = (w26563 & w26639) | (w26563 & w65736) | (w26639 & w65736);
assign w27263 = w26576 & ~w26632;
assign w27264 = w26769 & w27263;
assign w27265 = ~w27261 & ~w27262;
assign w27266 = ~w27264 & w27265;
assign w27267 = w26621 & ~w27266;
assign w27268 = ~w26742 & w65737;
assign w27269 = w26589 & ~w27268;
assign w27270 = ~w27252 & ~w27269;
assign w27271 = ~w27267 & w27270;
assign w27272 = ~w27260 & w27271;
assign w27273 = pi1457 & w27272;
assign w27274 = ~pi1457 & ~w27272;
assign w27275 = ~w27273 & ~w27274;
assign w27276 = ~w26404 & ~w27222;
assign w27277 = w27229 & ~w27242;
assign w27278 = ~w27276 & ~w27277;
assign w27279 = w26364 & w26386;
assign w27280 = ~w26377 & w27279;
assign w27281 = ~w26388 & w27280;
assign w27282 = ~w26403 & ~w27244;
assign w27283 = ~w26358 & w26404;
assign w27284 = ~w27222 & w27240;
assign w27285 = ~w26393 & ~w27284;
assign w27286 = ~w27281 & w27282;
assign w27287 = ~w27283 & ~w27285;
assign w27288 = w27286 & w27287;
assign w27289 = ~w26366 & w26371;
assign w27290 = ~w26379 & w27289;
assign w27291 = w26403 & ~w27290;
assign w27292 = ~w26396 & w27291;
assign w27293 = ~w27242 & w27292;
assign w27294 = ~w27288 & ~w27293;
assign w27295 = ~w27294 & w65738;
assign w27296 = (pi1465 & w27294) | (pi1465 & w65739) | (w27294 & w65739);
assign w27297 = ~w27295 & ~w27296;
assign w27298 = w26673 & w26700;
assign w27299 = w26843 & w27298;
assign w27300 = ~w26675 & ~w26828;
assign w27301 = (w26666 & w27300) | (w26666 & w65740) | (w27300 & w65740);
assign w27302 = w26683 & w26715;
assign w27303 = ~w26666 & w26673;
assign w27304 = (~w27303 & w26836) | (~w27303 & w65741) | (w26836 & w65741);
assign w27305 = (w26653 & w26707) | (w26653 & w63827) | (w26707 & w63827);
assign w27306 = ~w27302 & ~w27305;
assign w27307 = ~w27304 & w27306;
assign w27308 = ~w27301 & ~w27307;
assign w27309 = ~w26694 & ~w27299;
assign w27310 = ~w27308 & w27309;
assign w27311 = ~w26688 & w26851;
assign w27312 = ~w26853 & ~w27311;
assign w27313 = w26694 & ~w26854;
assign w27314 = w26843 & w27313;
assign w27315 = ~w27305 & w27314;
assign w27316 = ~w27312 & w27315;
assign w27317 = ~w27310 & w65742;
assign w27318 = (~pi1472 & w27310) | (~pi1472 & w65743) | (w27310 & w65743);
assign w27319 = ~w27317 & ~w27318;
assign w27320 = w26376 & w27225;
assign w27321 = ~w26386 & ~w27221;
assign w27322 = ~w26373 & w65744;
assign w27323 = w26351 & w26421;
assign w27324 = ~w26368 & w26416;
assign w27325 = ~w26395 & ~w27323;
assign w27326 = w27282 & w27325;
assign w27327 = ~w27324 & w27326;
assign w27328 = w27236 & ~w27289;
assign w27329 = w27289 & w27321;
assign w27330 = ~w26378 & w26403;
assign w27331 = ~w26405 & ~w26420;
assign w27332 = w27330 & w27331;
assign w27333 = ~w27329 & w27332;
assign w27334 = ~w27328 & w27333;
assign w27335 = ~w27327 & ~w27334;
assign w27336 = ~w27320 & ~w27322;
assign w27337 = ~w26397 & w27336;
assign w27338 = ~w27335 & w27337;
assign w27339 = pi1479 & w27338;
assign w27340 = ~pi1479 & ~w27338;
assign w27341 = ~w27339 & ~w27340;
assign w27342 = w26182 & w26221;
assign w27343 = ~w26191 & w26210;
assign w27344 = w26225 & ~w27343;
assign w27345 = (~w26777 & w27132) | (~w26777 & w65745) | (w27132 & w65745);
assign w27346 = ~w26210 & ~w27345;
assign w27347 = w26152 & ~w26172;
assign w27348 = ~w27346 & w27347;
assign w27349 = ~w27344 & ~w27348;
assign w27350 = w26152 & ~w26203;
assign w27351 = w26777 & w26783;
assign w27352 = w27131 & ~w27351;
assign w27353 = ~w27350 & ~w27352;
assign w27354 = w26202 & ~w27342;
assign w27355 = ~w27353 & w27354;
assign w27356 = ~w27349 & w27355;
assign w27357 = w26225 & w65746;
assign w27358 = ~w26205 & ~w26783;
assign w27359 = ~w27346 & ~w27358;
assign w27360 = ~w26185 & ~w26202;
assign w27361 = ~w27357 & w27360;
assign w27362 = ~w27359 & w27361;
assign w27363 = ~w27356 & ~w27362;
assign w27364 = ~pi1460 & w27363;
assign w27365 = pi1460 & ~w27363;
assign w27366 = ~w27364 & ~w27365;
assign w27367 = w27046 & w27072;
assign w27368 = ~w27011 & ~w27024;
assign w27369 = ~w27070 & ~w27166;
assign w27370 = ~w27017 & ~w27053;
assign w27371 = ~w27060 & w27370;
assign w27372 = ~w27369 & ~w27371;
assign w27373 = (~w27368 & w27369) | (~w27368 & w65747) | (w27369 & w65747);
assign w27374 = ~w27055 & ~w27368;
assign w27375 = w27372 & ~w27374;
assign w27376 = w27037 & ~w27373;
assign w27377 = ~w27375 & w27376;
assign w27378 = ~w27030 & ~w27154;
assign w27379 = w27163 & ~w27378;
assign w27380 = ~w27073 & ~w27379;
assign w27381 = w27171 & w27380;
assign w27382 = ~w27377 & ~w27381;
assign w27383 = ~w27030 & ~w27053;
assign w27384 = w27060 & w27383;
assign w27385 = ~w27367 & ~w27384;
assign w27386 = ~w27382 & w27385;
assign w27387 = pi1453 & ~w27386;
assign w27388 = ~pi1453 & w27386;
assign w27389 = ~w27387 & ~w27388;
assign w27390 = ~w27060 & ~w27368;
assign w27391 = ~w27017 & ~w27390;
assign w27392 = w27075 & w27081;
assign w27393 = (~w27038 & ~w27392) | (~w27038 & w65748) | (~w27392 & w65748);
assign w27394 = ~w27154 & ~w27393;
assign w27395 = ~w27030 & ~w27151;
assign w27396 = ~w27064 & ~w27395;
assign w27397 = ~w27037 & ~w27396;
assign w27398 = ~w27018 & ~w27060;
assign w27399 = w27024 & w27059;
assign w27400 = ~w27037 & ~w27399;
assign w27401 = w27063 & ~w27398;
assign w27402 = ~w27400 & w27401;
assign w27403 = ~w27070 & ~w27400;
assign w27404 = w27053 & ~w27061;
assign w27405 = ~w27403 & w27404;
assign w27406 = ~w27402 & ~w27405;
assign w27407 = ~w27394 & w27406;
assign w27408 = ~w27397 & w27407;
assign w27409 = pi1455 & ~w27408;
assign w27410 = ~pi1455 & w27408;
assign w27411 = ~w27409 & ~w27410;
assign w27412 = ~w26911 & w26966;
assign w27413 = w26940 & w27412;
assign w27414 = (~w26949 & ~w27412) | (~w26949 & w65749) | (~w27412 & w65749);
assign w27415 = ~w26903 & ~w27414;
assign w27416 = ~w26926 & w26939;
assign w27417 = ~w26943 & w27416;
assign w27418 = ~w27413 & ~w27417;
assign w27419 = ~w27415 & w27418;
assign w27420 = w26891 & ~w27419;
assign w27421 = w26938 & ~w26991;
assign w27422 = w26920 & w26954;
assign w27423 = w27412 & ~w27422;
assign w27424 = ~w26891 & ~w27421;
assign w27425 = ~w27423 & w27424;
assign w27426 = w26903 & w26962;
assign w27427 = ~w26985 & ~w27426;
assign w27428 = ~w26910 & ~w27427;
assign w27429 = w26914 & ~w26949;
assign w27430 = ~w26934 & ~w26961;
assign w27431 = ~w27429 & w27430;
assign w27432 = ~w27425 & ~w27431;
assign w27433 = ~w27428 & w27432;
assign w27434 = ~w27420 & w27433;
assign w27435 = pi1474 & w27434;
assign w27436 = ~pi1474 & ~w27434;
assign w27437 = ~w27435 & ~w27436;
assign w27438 = w26675 & w26832;
assign w27439 = ~w26825 & ~w26839;
assign w27440 = ~w27438 & w27439;
assign w27441 = w26714 & w27440;
assign w27442 = ~w26840 & ~w26849;
assign w27443 = ~w26666 & ~w26675;
assign w27444 = ~w27442 & ~w27443;
assign w27445 = w26694 & ~w26716;
assign w27446 = ~w27444 & w27445;
assign w27447 = ~w27441 & ~w27446;
assign w27448 = w26660 & w27303;
assign w27449 = ~w26856 & ~w27448;
assign w27450 = ~w27447 & w27449;
assign w27451 = pi1498 & w27450;
assign w27452 = ~pi1498 & ~w27450;
assign w27453 = ~w27451 & ~w27452;
assign w27454 = ~pi4906 & pi9040;
assign w27455 = ~pi4967 & ~pi9040;
assign w27456 = ~w27454 & ~w27455;
assign w27457 = pi1469 & ~w27456;
assign w27458 = ~pi1469 & w27456;
assign w27459 = ~w27457 & ~w27458;
assign w27460 = ~pi4841 & pi9040;
assign w27461 = ~pi4821 & ~pi9040;
assign w27462 = ~w27460 & ~w27461;
assign w27463 = pi1463 & ~w27462;
assign w27464 = ~pi1463 & w27462;
assign w27465 = ~w27463 & ~w27464;
assign w27466 = w27459 & ~w27465;
assign w27467 = ~w27459 & w27465;
assign w27468 = ~w27466 & ~w27467;
assign w27469 = ~pi5187 & pi9040;
assign w27470 = ~pi4843 & ~pi9040;
assign w27471 = ~w27469 & ~w27470;
assign w27472 = pi1476 & ~w27471;
assign w27473 = ~pi1476 & w27471;
assign w27474 = ~w27472 & ~w27473;
assign w27475 = ~w27465 & w27474;
assign w27476 = w27468 & ~w27475;
assign w27477 = ~pi4874 & pi9040;
assign w27478 = ~pi5184 & ~pi9040;
assign w27479 = ~w27477 & ~w27478;
assign w27480 = pi1493 & ~w27479;
assign w27481 = ~pi1493 & w27479;
assign w27482 = ~w27480 & ~w27481;
assign w27483 = ~w27465 & w27482;
assign w27484 = w27474 & ~w27483;
assign w27485 = ~w27459 & w27482;
assign w27486 = ~w27474 & w27485;
assign w27487 = ~w27484 & ~w27486;
assign w27488 = ~pi4845 & pi9040;
assign w27489 = ~pi5150 & ~pi9040;
assign w27490 = ~w27488 & ~w27489;
assign w27491 = pi1489 & ~w27490;
assign w27492 = ~pi1489 & w27490;
assign w27493 = ~w27491 & ~w27492;
assign w27494 = ~w27487 & w27493;
assign w27495 = w27476 & w27494;
assign w27496 = ~w27465 & ~w27493;
assign w27497 = ~w27459 & w27474;
assign w27498 = w27496 & w27497;
assign w27499 = ~w27474 & ~w27482;
assign w27500 = ~w27468 & w27499;
assign w27501 = w27459 & ~w27482;
assign w27502 = w27465 & w27474;
assign w27503 = w27501 & w27502;
assign w27504 = ~w27498 & ~w27503;
assign w27505 = ~w27500 & w27504;
assign w27506 = w27459 & w27493;
assign w27507 = w27499 & w27506;
assign w27508 = ~w27459 & ~w27465;
assign w27509 = w27482 & w27508;
assign w27510 = ~w27507 & ~w27509;
assign w27511 = ~w27505 & ~w27510;
assign w27512 = ~w27483 & ~w27493;
assign w27513 = ~w27474 & w27508;
assign w27514 = w27512 & w27513;
assign w27515 = ~w27474 & w27482;
assign w27516 = w27459 & w27474;
assign w27517 = w27465 & ~w27515;
assign w27518 = ~w27516 & w27517;
assign w27519 = w27496 & w27516;
assign w27520 = ~w27482 & w27519;
assign w27521 = w27466 & w27515;
assign w27522 = ~w27518 & ~w27521;
assign w27523 = (~w27493 & ~w27522) | (~w27493 & w65750) | (~w27522 & w65750);
assign w27524 = w27465 & w27482;
assign w27525 = ~w27475 & ~w27524;
assign w27526 = w27474 & w27485;
assign w27527 = w27493 & ~w27501;
assign w27528 = ~w27526 & w27527;
assign w27529 = ~w27525 & w27528;
assign w27530 = ~pi4832 & pi9040;
assign w27531 = ~pi4836 & ~pi9040;
assign w27532 = ~w27530 & ~w27531;
assign w27533 = pi1484 & ~w27532;
assign w27534 = ~pi1484 & w27532;
assign w27535 = ~w27533 & ~w27534;
assign w27536 = ~w27529 & w27535;
assign w27537 = ~w27523 & w27536;
assign w27538 = ~w27503 & ~w27526;
assign w27539 = ~w27518 & ~w27538;
assign w27540 = w27465 & ~w27474;
assign w27541 = w27493 & ~w27540;
assign w27542 = ~w27484 & ~w27525;
assign w27543 = ~w27541 & ~w27542;
assign w27544 = w27493 & ~w27525;
assign w27545 = ~w27543 & ~w27544;
assign w27546 = ~w27498 & ~w27535;
assign w27547 = ~w27507 & w27546;
assign w27548 = ~w27539 & w27547;
assign w27549 = ~w27545 & w27548;
assign w27550 = ~w27537 & ~w27549;
assign w27551 = ~w27495 & ~w27514;
assign w27552 = ~w27511 & w27551;
assign w27553 = ~w27550 & w27552;
assign w27554 = pi1504 & ~w27553;
assign w27555 = ~pi1504 & w27553;
assign w27556 = ~w27554 & ~w27555;
assign w27557 = ~pi4987 & pi9040;
assign w27558 = ~pi4842 & ~pi9040;
assign w27559 = ~w27557 & ~w27558;
assign w27560 = pi1484 & ~w27559;
assign w27561 = ~pi1484 & w27559;
assign w27562 = ~w27560 & ~w27561;
assign w27563 = ~pi4967 & pi9040;
assign w27564 = ~pi5187 & ~pi9040;
assign w27565 = ~w27563 & ~w27564;
assign w27566 = pi1470 & ~w27565;
assign w27567 = ~pi1470 & w27565;
assign w27568 = ~w27566 & ~w27567;
assign w27569 = ~w27562 & w27568;
assign w27570 = w27562 & ~w27568;
assign w27571 = ~w27569 & ~w27570;
assign w27572 = ~pi4843 & pi9040;
assign w27573 = ~pi4874 & ~pi9040;
assign w27574 = ~w27572 & ~w27573;
assign w27575 = pi1469 & ~w27574;
assign w27576 = ~pi1469 & w27574;
assign w27577 = ~w27575 & ~w27576;
assign w27578 = w27571 & w27577;
assign w27579 = ~pi4964 & pi9040;
assign w27580 = ~pi4890 & ~pi9040;
assign w27581 = ~w27579 & ~w27580;
assign w27582 = pi1496 & ~w27581;
assign w27583 = ~pi1496 & w27581;
assign w27584 = ~w27582 & ~w27583;
assign w27585 = ~pi4876 & pi9040;
assign w27586 = ~pi4987 & ~pi9040;
assign w27587 = ~w27585 & ~w27586;
assign w27588 = pi1481 & ~w27587;
assign w27589 = ~pi1481 & w27587;
assign w27590 = ~w27588 & ~w27589;
assign w27591 = ~w27577 & ~w27590;
assign w27592 = w27562 & ~w27590;
assign w27593 = ~w27591 & ~w27592;
assign w27594 = ~w27569 & w27591;
assign w27595 = ~pi4965 & pi9040;
assign w27596 = ~pi4876 & ~pi9040;
assign w27597 = ~w27595 & ~w27596;
assign w27598 = pi1480 & ~w27597;
assign w27599 = ~pi1480 & w27597;
assign w27600 = ~w27598 & ~w27599;
assign w27601 = ~w27593 & ~w27600;
assign w27602 = ~w27594 & w27601;
assign w27603 = ~w27578 & ~w27584;
assign w27604 = ~w27602 & w27603;
assign w27605 = w27577 & w27590;
assign w27606 = ~w27591 & ~w27605;
assign w27607 = w27569 & w27606;
assign w27608 = w27584 & ~w27594;
assign w27609 = ~w27607 & w27608;
assign w27610 = ~w27604 & ~w27609;
assign w27611 = ~w27568 & ~w27577;
assign w27612 = ~w27584 & w27590;
assign w27613 = w27562 & w27611;
assign w27614 = ~w27612 & w27613;
assign w27615 = ~w27605 & ~w27612;
assign w27616 = w27571 & ~w27615;
assign w27617 = ~w27600 & ~w27614;
assign w27618 = ~w27616 & w27617;
assign w27619 = ~w27562 & ~w27577;
assign w27620 = w27568 & w27590;
assign w27621 = ~w27568 & ~w27590;
assign w27622 = ~w27620 & ~w27621;
assign w27623 = w27619 & ~w27622;
assign w27624 = w27562 & w27584;
assign w27625 = w27568 & ~w27577;
assign w27626 = ~w27568 & w27605;
assign w27627 = ~w27625 & ~w27626;
assign w27628 = w27624 & ~w27627;
assign w27629 = w27562 & w27577;
assign w27630 = ~w27619 & ~w27629;
assign w27631 = w27612 & ~w27625;
assign w27632 = w27630 & w27631;
assign w27633 = w27600 & ~w27623;
assign w27634 = ~w27632 & w27633;
assign w27635 = ~w27628 & w27634;
assign w27636 = ~w27618 & ~w27635;
assign w27637 = ~w27610 & ~w27636;
assign w27638 = pi1509 & w27637;
assign w27639 = ~pi1509 & ~w27637;
assign w27640 = ~w27638 & ~w27639;
assign w27641 = w27501 & w27540;
assign w27642 = w27485 & w27502;
assign w27643 = ~w27496 & ~w27642;
assign w27644 = ~w27467 & w27515;
assign w27645 = ~w27642 & ~w27644;
assign w27646 = w27493 & ~w27645;
assign w27647 = w27459 & ~w27502;
assign w27648 = ~w27497 & w27512;
assign w27649 = ~w27647 & w27648;
assign w27650 = w27505 & ~w27646;
assign w27651 = w27650 & w63828;
assign w27652 = ~w27500 & w27645;
assign w27653 = (~w27641 & ~w27652) | (~w27641 & w65751) | (~w27652 & w65751);
assign w27654 = (~w27535 & w27651) | (~w27535 & w65752) | (w27651 & w65752);
assign w27655 = w27483 & w27506;
assign w27656 = (w27535 & ~w27650) | (w27535 & w65753) | (~w27650 & w65753);
assign w27657 = w27474 & ~w27482;
assign w27658 = w27508 & w27657;
assign w27659 = ~w27655 & ~w27658;
assign w27660 = ~w27656 & w27659;
assign w27661 = ~w27654 & w27660;
assign w27662 = pi1505 & ~w27661;
assign w27663 = ~pi1505 & w27661;
assign w27664 = ~w27662 & ~w27663;
assign w27665 = ~w27493 & w27657;
assign w27666 = ~w27496 & ~w27525;
assign w27667 = w27487 & w27666;
assign w27668 = w27535 & ~w27665;
assign w27669 = ~w27500 & w27668;
assign w27670 = w27510 & w27669;
assign w27671 = ~w27667 & w27670;
assign w27672 = w27516 & w27524;
assign w27673 = ~w27485 & ~w27501;
assign w27674 = ~w27474 & ~w27493;
assign w27675 = w27673 & w27674;
assign w27676 = ~w27535 & ~w27672;
assign w27677 = ~w27675 & w27676;
assign w27678 = ~w27494 & w27677;
assign w27679 = ~w27511 & w27678;
assign w27680 = ~w27671 & ~w27679;
assign w27681 = ~w27520 & ~w27680;
assign w27682 = ~pi1511 & w27681;
assign w27683 = pi1511 & ~w27681;
assign w27684 = ~w27682 & ~w27683;
assign w27685 = ~pi4890 & pi9040;
assign w27686 = ~pi4960 & ~pi9040;
assign w27687 = ~w27685 & ~w27686;
assign w27688 = pi1476 & ~w27687;
assign w27689 = ~pi1476 & w27687;
assign w27690 = ~w27688 & ~w27689;
assign w27691 = ~pi4836 & pi9040;
assign w27692 = ~pi4988 & ~pi9040;
assign w27693 = ~w27691 & ~w27692;
assign w27694 = pi1478 & ~w27693;
assign w27695 = ~pi1478 & w27693;
assign w27696 = ~w27694 & ~w27695;
assign w27697 = ~pi5184 & pi9040;
assign w27698 = ~pi4818 & ~pi9040;
assign w27699 = ~w27697 & ~w27698;
assign w27700 = pi1503 & ~w27699;
assign w27701 = ~pi1503 & w27699;
assign w27702 = ~w27700 & ~w27701;
assign w27703 = w27696 & ~w27702;
assign w27704 = ~pi4990 & pi9040;
assign w27705 = ~pi4964 & ~pi9040;
assign w27706 = ~w27704 & ~w27705;
assign w27707 = pi1495 & ~w27706;
assign w27708 = ~pi1495 & w27706;
assign w27709 = ~w27707 & ~w27708;
assign w27710 = ~pi4911 & pi9040;
assign w27711 = ~pi4957 & ~pi9040;
assign w27712 = ~w27710 & ~w27711;
assign w27713 = pi1483 & ~w27712;
assign w27714 = ~pi1483 & w27712;
assign w27715 = ~w27713 & ~w27714;
assign w27716 = ~w27709 & w27715;
assign w27717 = ~w27703 & ~w27716;
assign w27718 = ~w27696 & w27702;
assign w27719 = ~w27709 & ~w27718;
assign w27720 = w27717 & w27719;
assign w27721 = ~pi4881 & pi9040;
assign w27722 = ~pi5038 & ~pi9040;
assign w27723 = ~w27721 & ~w27722;
assign w27724 = pi1493 & ~w27723;
assign w27725 = ~pi1493 & w27723;
assign w27726 = ~w27724 & ~w27725;
assign w27727 = w27696 & w27726;
assign w27728 = w27702 & ~w27715;
assign w27729 = w27727 & w27728;
assign w27730 = w27696 & ~w27709;
assign w27731 = ~w27726 & ~w27730;
assign w27732 = ~w27717 & w27731;
assign w27733 = ~w27720 & ~w27729;
assign w27734 = (~w27690 & ~w27733) | (~w27690 & w65754) | (~w27733 & w65754);
assign w27735 = ~w27702 & w27715;
assign w27736 = w27727 & w27735;
assign w27737 = w27703 & ~w27715;
assign w27738 = (w27709 & ~w27703) | (w27709 & w64412) | (~w27703 & w64412);
assign w27739 = ~w27715 & w27726;
assign w27740 = ~w27702 & w27739;
assign w27741 = w27715 & ~w27726;
assign w27742 = w27696 & w27741;
assign w27743 = w27741 & w63829;
assign w27744 = ~w27696 & ~w27726;
assign w27745 = w27728 & w27744;
assign w27746 = ~w27743 & ~w27745;
assign w27747 = ~w27740 & w27746;
assign w27748 = w27738 & ~w27747;
assign w27749 = w27716 & w27718;
assign w27750 = w27703 & w27739;
assign w27751 = ~w27743 & ~w27750;
assign w27752 = ~w27696 & w27726;
assign w27753 = w27715 & w27752;
assign w27754 = ~w27737 & ~w27753;
assign w27755 = ~w27709 & ~w27754;
assign w27756 = (w27709 & ~w27741) | (w27709 & w65755) | (~w27741 & w65755);
assign w27757 = w27702 & w27715;
assign w27758 = w27744 & w27757;
assign w27759 = ~w27729 & ~w27758;
assign w27760 = w27754 & w27759;
assign w27761 = w27756 & w27760;
assign w27762 = w27751 & ~w27755;
assign w27763 = ~w27761 & w27762;
assign w27764 = w27690 & ~w27763;
assign w27765 = ~w27736 & ~w27749;
assign w27766 = ~w27734 & w27765;
assign w27767 = ~w27748 & w27766;
assign w27768 = ~w27764 & w27767;
assign w27769 = pi1512 & ~w27768;
assign w27770 = ~pi1512 & w27768;
assign w27771 = ~w27769 & ~w27770;
assign w27772 = ~pi4962 & pi9040;
assign w27773 = ~pi4844 & ~pi9040;
assign w27774 = ~w27772 & ~w27773;
assign w27775 = pi1494 & ~w27774;
assign w27776 = ~pi1494 & w27774;
assign w27777 = ~w27775 & ~w27776;
assign w27778 = ~pi5278 & pi9040;
assign w27779 = ~pi4898 & ~pi9040;
assign w27780 = ~w27778 & ~w27779;
assign w27781 = pi1488 & ~w27780;
assign w27782 = ~pi1488 & w27780;
assign w27783 = ~w27781 & ~w27782;
assign w27784 = ~pi4833 & pi9040;
assign w27785 = ~pi5063 & ~pi9040;
assign w27786 = ~w27784 & ~w27785;
assign w27787 = pi1497 & ~w27786;
assign w27788 = ~pi1497 & w27786;
assign w27789 = ~w27787 & ~w27788;
assign w27790 = ~pi5063 & pi9040;
assign w27791 = ~pi4854 & ~pi9040;
assign w27792 = ~w27790 & ~w27791;
assign w27793 = pi1467 & ~w27792;
assign w27794 = ~pi1467 & w27792;
assign w27795 = ~w27793 & ~w27794;
assign w27796 = ~w27789 & ~w27795;
assign w27797 = w27789 & w27795;
assign w27798 = ~w27796 & ~w27797;
assign w27799 = ~pi5039 & pi9040;
assign w27800 = ~pi4961 & ~pi9040;
assign w27801 = ~w27799 & ~w27800;
assign w27802 = pi1487 & ~w27801;
assign w27803 = ~pi1487 & w27801;
assign w27804 = ~w27802 & ~w27803;
assign w27805 = w27795 & w27804;
assign w27806 = w27783 & w27805;
assign w27807 = ~pi4854 & pi9040;
assign w27808 = ~pi4840 & ~pi9040;
assign w27809 = ~w27807 & ~w27808;
assign w27810 = pi1501 & ~w27809;
assign w27811 = ~pi1501 & w27809;
assign w27812 = ~w27810 & ~w27811;
assign w27813 = w27804 & ~w27812;
assign w27814 = w27789 & w27813;
assign w27815 = ~w27806 & ~w27814;
assign w27816 = ~w27783 & ~w27804;
assign w27817 = ~w27795 & w27816;
assign w27818 = w27815 & ~w27817;
assign w27819 = w27815 & w63396;
assign w27820 = ~w27783 & ~w27819;
assign w27821 = w27789 & w27804;
assign w27822 = ~w27783 & ~w27795;
assign w27823 = w27821 & w27822;
assign w27824 = w27812 & ~w27823;
assign w27825 = w27798 & w27824;
assign w27826 = w27824 & w63397;
assign w27827 = w27783 & ~w27826;
assign w27828 = ~w27820 & ~w27827;
assign w27829 = w27783 & ~w27789;
assign w27830 = w27795 & ~w27804;
assign w27831 = ~w27829 & ~w27830;
assign w27832 = ~w27789 & ~w27812;
assign w27833 = w27783 & ~w27812;
assign w27834 = ~w27832 & ~w27833;
assign w27835 = ~w27821 & w27831;
assign w27836 = ~w27834 & w27835;
assign w27837 = (~w27777 & w27828) | (~w27777 & w63830) | (w27828 & w63830);
assign w27838 = ~w27789 & ~w27804;
assign w27839 = ~w27821 & ~w27838;
assign w27840 = w27795 & ~w27839;
assign w27841 = w27833 & w27840;
assign w27842 = w27789 & w27812;
assign w27843 = w27816 & w27842;
assign w27844 = ~w27832 & ~w27842;
assign w27845 = ~w27795 & ~w27804;
assign w27846 = w27783 & w27845;
assign w27847 = w27844 & w27846;
assign w27848 = w27812 & w27847;
assign w27849 = w27813 & w27822;
assign w27850 = ~w27795 & w27839;
assign w27851 = ~w27825 & ~w27850;
assign w27852 = w27820 & ~w27851;
assign w27853 = ~w27805 & w27812;
assign w27854 = ~w27831 & w27853;
assign w27855 = ~w27822 & w27838;
assign w27856 = ~w27814 & ~w27855;
assign w27857 = (w27777 & w27852) | (w27777 & w65756) | (w27852 & w65756);
assign w27858 = ~w27843 & ~w27849;
assign w27859 = ~w27841 & w27858;
assign w27860 = ~w27848 & w27859;
assign w27861 = ~w27837 & w27860;
assign w27862 = w27861 & w65757;
assign w27863 = (pi1508 & ~w27861) | (pi1508 & w65758) | (~w27861 & w65758);
assign w27864 = ~w27862 & ~w27863;
assign w27865 = ~pi5060 & pi9040;
assign w27866 = ~pi4909 & ~pi9040;
assign w27867 = ~w27865 & ~w27866;
assign w27868 = pi1500 & ~w27867;
assign w27869 = ~pi1500 & w27867;
assign w27870 = ~w27868 & ~w27869;
assign w27871 = ~pi4898 & pi9040;
assign w27872 = ~pi5116 & ~pi9040;
assign w27873 = ~w27871 & ~w27872;
assign w27874 = pi1478 & ~w27873;
assign w27875 = ~pi1478 & w27873;
assign w27876 = ~w27874 & ~w27875;
assign w27877 = ~pi4844 & pi9040;
assign w27878 = ~pi5278 & ~pi9040;
assign w27879 = ~w27877 & ~w27878;
assign w27880 = pi1502 & ~w27879;
assign w27881 = ~pi1502 & w27879;
assign w27882 = ~w27880 & ~w27881;
assign w27883 = ~w27876 & w27882;
assign w27884 = ~pi4849 & pi9040;
assign w27885 = ~pi5060 & ~pi9040;
assign w27886 = ~w27884 & ~w27885;
assign w27887 = pi1473 & ~w27886;
assign w27888 = ~pi1473 & w27886;
assign w27889 = ~w27887 & ~w27888;
assign w27890 = ~w27870 & ~w27889;
assign w27891 = w27870 & w27889;
assign w27892 = ~w27890 & ~w27891;
assign w27893 = ~pi4835 & pi9040;
assign w27894 = ~pi4847 & ~pi9040;
assign w27895 = ~w27893 & ~w27894;
assign w27896 = pi1486 & ~w27895;
assign w27897 = ~pi1486 & w27895;
assign w27898 = ~w27896 & ~w27897;
assign w27899 = ~w27892 & w27898;
assign w27900 = ~w27870 & ~w27882;
assign w27901 = w27876 & w27889;
assign w27902 = w27876 & ~w27898;
assign w27903 = w27900 & ~w27901;
assign w27904 = ~w27902 & w27903;
assign w27905 = w27892 & ~w27898;
assign w27906 = ~w27876 & ~w27889;
assign w27907 = w27892 & w63832;
assign w27908 = w27870 & w27882;
assign w27909 = w27876 & ~w27889;
assign w27910 = ~w27889 & ~w27898;
assign w27911 = ~w27902 & ~w27910;
assign w27912 = w27911 & w65759;
assign w27913 = ~w27904 & ~w27907;
assign w27914 = ~w27912 & w27913;
assign w27915 = w27883 & ~w27899;
assign w27916 = w27914 & w27915;
assign w27917 = ~w27870 & w27916;
assign w27918 = w27876 & w27900;
assign w27919 = ~w27901 & ~w27906;
assign w27920 = w27889 & w27908;
assign w27921 = w27870 & w27898;
assign w27922 = ~w27870 & w27882;
assign w27923 = ~w27921 & ~w27922;
assign w27924 = ~w27889 & ~w27923;
assign w27925 = ~w27870 & ~w27898;
assign w27926 = ~w27920 & ~w27925;
assign w27927 = ~w27924 & w27926;
assign w27928 = ~w27919 & ~w27927;
assign w27929 = w27892 & w65760;
assign w27930 = w27909 & w27929;
assign w27931 = ~pi4966 & pi9040;
assign w27932 = ~pi4837 & ~pi9040;
assign w27933 = ~w27931 & ~w27932;
assign w27934 = pi1483 & ~w27933;
assign w27935 = ~pi1483 & w27933;
assign w27936 = ~w27934 & ~w27935;
assign w27937 = ~w27923 & w65761;
assign w27938 = w27883 & w27891;
assign w27939 = ~w27898 & w27938;
assign w27940 = ~w27937 & ~w27939;
assign w27941 = ~w27876 & ~w27882;
assign w27942 = w27898 & w27941;
assign w27943 = w27889 & w27942;
assign w27944 = ~w27918 & ~w27936;
assign w27945 = ~w27943 & w27944;
assign w27946 = ~w27928 & w27945;
assign w27947 = ~w27930 & w27940;
assign w27948 = w27946 & w27947;
assign w27949 = w27901 & w27921;
assign w27950 = w27936 & ~w27949;
assign w27951 = w27890 & w27942;
assign w27952 = ~w27900 & ~w27921;
assign w27953 = w27909 & w27952;
assign w27954 = ~w27938 & w27950;
assign w27955 = ~w27951 & ~w27953;
assign w27956 = w27954 & w27955;
assign w27957 = ~w27929 & w27956;
assign w27958 = ~w27948 & ~w27957;
assign w27959 = ~w27958 & w65762;
assign w27960 = (~pi1514 & w27958) | (~pi1514 & w65763) | (w27958 & w65763);
assign w27961 = ~w27959 & ~w27960;
assign w27962 = (w27493 & ~w27538) | (w27493 & w63833) | (~w27538 & w63833);
assign w27963 = ~w27519 & ~w27658;
assign w27964 = ~w27962 & w27963;
assign w27965 = ~w27535 & ~w27964;
assign w27966 = w27476 & w27482;
assign w27967 = ~w27475 & ~w27496;
assign w27968 = ~w27962 & w65764;
assign w27969 = ~w27966 & ~w27968;
assign w27970 = w27535 & ~w27969;
assign w27971 = (w27493 & w27652) | (w27493 & w65765) | (w27652 & w65765);
assign w27972 = ~w27486 & ~w27641;
assign w27973 = ~w27535 & ~w27972;
assign w27974 = w27502 & w27673;
assign w27975 = ~w27493 & ~w27513;
assign w27976 = ~w27974 & w27975;
assign w27977 = ~w27973 & w27976;
assign w27978 = ~w27971 & ~w27977;
assign w27979 = ~w27965 & ~w27978;
assign w27980 = ~w27970 & w27979;
assign w27981 = ~pi1515 & w27980;
assign w27982 = pi1515 & ~w27980;
assign w27983 = ~w27981 & ~w27982;
assign w27984 = ~pi5150 & pi9040;
assign w27985 = ~pi4881 & ~pi9040;
assign w27986 = ~w27984 & ~w27985;
assign w27987 = pi1464 & ~w27986;
assign w27988 = ~pi1464 & w27986;
assign w27989 = ~w27987 & ~w27988;
assign w27990 = ~pi5038 & pi9040;
assign w27991 = ~pi4990 & ~pi9040;
assign w27992 = ~w27990 & ~w27991;
assign w27993 = pi1480 & ~w27992;
assign w27994 = ~pi1480 & w27992;
assign w27995 = ~w27993 & ~w27994;
assign w27996 = ~pi4821 & pi9040;
assign w27997 = ~pi4832 & ~pi9040;
assign w27998 = ~w27996 & ~w27997;
assign w27999 = pi1481 & ~w27998;
assign w28000 = ~pi1481 & w27998;
assign w28001 = ~w27999 & ~w28000;
assign w28002 = ~w27995 & ~w28001;
assign w28003 = ~pi4818 & pi9040;
assign w28004 = ~pi4911 & ~pi9040;
assign w28005 = ~w28003 & ~w28004;
assign w28006 = pi1485 & ~w28005;
assign w28007 = ~pi1485 & w28005;
assign w28008 = ~w28006 & ~w28007;
assign w28009 = ~pi4957 & pi9040;
assign w28010 = ~pi4841 & ~pi9040;
assign w28011 = ~w28009 & ~w28010;
assign w28012 = pi1487 & ~w28011;
assign w28013 = ~pi1487 & w28011;
assign w28014 = ~w28012 & ~w28013;
assign w28015 = w28008 & ~w28014;
assign w28016 = ~w28008 & w28014;
assign w28017 = ~w28015 & ~w28016;
assign w28018 = w28002 & w28017;
assign w28019 = w27995 & ~w28008;
assign w28020 = w28001 & ~w28014;
assign w28021 = ~w28019 & ~w28020;
assign w28022 = w28001 & ~w28008;
assign w28023 = ~w27995 & w28001;
assign w28024 = ~w28014 & ~w28023;
assign w28025 = ~w28022 & ~w28024;
assign w28026 = ~w28021 & w28025;
assign w28027 = w28002 & w28014;
assign w28028 = w27995 & ~w28001;
assign w28029 = w28008 & w28028;
assign w28030 = w28028 & w28015;
assign w28031 = ~w28027 & ~w28030;
assign w28032 = ~pi5185 & pi9040;
assign w28033 = ~pi4906 & ~pi9040;
assign w28034 = ~w28032 & ~w28033;
assign w28035 = pi1497 & ~w28034;
assign w28036 = ~pi1497 & w28034;
assign w28037 = ~w28035 & ~w28036;
assign w28038 = ~w28031 & ~w28037;
assign w28039 = ~w28018 & ~w28026;
assign w28040 = (w27989 & ~w28039) | (w27989 & w65766) | (~w28039 & w65766);
assign w28041 = ~w27989 & w27995;
assign w28042 = ~w28014 & w28022;
assign w28043 = w28041 & w28042;
assign w28044 = w28001 & w28014;
assign w28045 = w27995 & w28001;
assign w28046 = w28008 & w28045;
assign w28047 = w27989 & ~w28046;
assign w28048 = w28044 & ~w28047;
assign w28049 = ~w27989 & ~w27995;
assign w28050 = w28015 & w28049;
assign w28051 = w27989 & ~w28042;
assign w28052 = w28019 & ~w28051;
assign w28053 = ~w28037 & ~w28050;
assign w28054 = ~w28048 & w28053;
assign w28055 = ~w28052 & w28054;
assign w28056 = ~w27995 & w28044;
assign w28057 = w28008 & w28056;
assign w28058 = w28002 & ~w28008;
assign w28059 = ~w28029 & ~w28058;
assign w28060 = ~w27989 & ~w28059;
assign w28061 = w27989 & ~w27995;
assign w28062 = ~w28051 & ~w28061;
assign w28063 = ~w28021 & ~w28062;
assign w28064 = w28037 & ~w28057;
assign w28065 = ~w28060 & w28064;
assign w28066 = ~w28063 & w28065;
assign w28067 = ~w28055 & ~w28066;
assign w28068 = ~w28040 & ~w28043;
assign w28069 = ~w28067 & w28068;
assign w28070 = pi1506 & ~w28069;
assign w28071 = ~pi1506 & w28069;
assign w28072 = ~w28070 & ~w28071;
assign w28073 = ~w27914 & ~w27936;
assign w28074 = w27882 & w27902;
assign w28075 = ~w27941 & ~w28074;
assign w28076 = w27905 & ~w28075;
assign w28077 = w27870 & ~w27882;
assign w28078 = (w28077 & ~w27911) | (w28077 & w65767) | (~w27911 & w65767);
assign w28079 = w27889 & w28078;
assign w28080 = w27898 & ~w27901;
assign w28081 = w27876 & w27890;
assign w28082 = ~w27898 & ~w28081;
assign w28083 = ~w27882 & ~w28080;
assign w28084 = ~w28082 & w28083;
assign w28085 = w27906 & w27952;
assign w28086 = ~w27902 & ~w27922;
assign w28087 = (~w27889 & ~w27902) | (~w27889 & w65768) | (~w27902 & w65768);
assign w28088 = w27902 & w65769;
assign w28089 = ~w28086 & ~w28087;
assign w28090 = ~w28088 & w28089;
assign w28091 = w27919 & ~w27923;
assign w28092 = ~w28090 & w28091;
assign w28093 = ~w28084 & ~w28085;
assign w28094 = ~w28092 & w28093;
assign w28095 = w27936 & ~w28094;
assign w28096 = ~w28076 & ~w28079;
assign w28097 = ~w28073 & w28096;
assign w28098 = ~w28095 & w28097;
assign w28099 = pi1518 & ~w28098;
assign w28100 = ~pi1518 & w28098;
assign w28101 = ~w28099 & ~w28100;
assign w28102 = ~w27727 & ~w27744;
assign w28103 = w27728 & w28102;
assign w28104 = ~w27744 & ~w27757;
assign w28105 = ~w27741 & ~w28104;
assign w28106 = ~w28104 & w63834;
assign w28107 = ~w27753 & ~w28106;
assign w28108 = (w27690 & w28106) | (w27690 & w65770) | (w28106 & w65770);
assign w28109 = w27751 & ~w28103;
assign w28110 = ~w28108 & w28109;
assign w28111 = w27709 & ~w28110;
assign w28112 = (~w27735 & ~w28102) | (~w27735 & w65771) | (~w28102 & w65771);
assign w28113 = w27690 & ~w27709;
assign w28114 = ~w28112 & w28113;
assign w28115 = (w27749 & w27763) | (w27749 & w63835) | (w27763 & w63835);
assign w28116 = w27730 & w27739;
assign w28117 = w27760 & w63836;
assign w28118 = w27719 & w27752;
assign w28119 = ~w27737 & ~w28116;
assign w28120 = ~w28118 & w28119;
assign w28121 = w27746 & w28120;
assign w28122 = ~w28117 & w28121;
assign w28123 = ~w27690 & ~w28122;
assign w28124 = ~w28111 & ~w28114;
assign w28125 = ~w28115 & ~w28123;
assign w28126 = w28125 & w65772;
assign w28127 = (~pi1513 & ~w28125) | (~pi1513 & w65773) | (~w28125 & w65773);
assign w28128 = ~w28126 & ~w28127;
assign w28129 = ~w27562 & w27590;
assign w28130 = ~w27592 & ~w28129;
assign w28131 = ~w27619 & w28130;
assign w28132 = w28130 & w63837;
assign w28133 = w27568 & w27577;
assign w28134 = ~w28130 & w28133;
assign w28135 = ~w28132 & ~w28134;
assign w28136 = ~w27571 & ~w27577;
assign w28137 = ~w28131 & ~w28136;
assign w28138 = (~w27584 & ~w27569) | (~w27584 & w65774) | (~w27569 & w65774);
assign w28139 = ~w28137 & w28138;
assign w28140 = ~w27568 & w28130;
assign w28141 = w28130 & w65775;
assign w28142 = w27584 & ~w28141;
assign w28143 = (w28135 & w28139) | (w28135 & w65776) | (w28139 & w65776);
assign w28144 = w27600 & ~w28143;
assign w28145 = w27569 & w27591;
assign w28146 = ~w27600 & ~w28140;
assign w28147 = w28135 & w28146;
assign w28148 = w27584 & ~w28145;
assign w28149 = ~w28147 & w28148;
assign w28150 = ~w28141 & ~w28145;
assign w28151 = ~w27600 & ~w28150;
assign w28152 = ~w27584 & w28135;
assign w28153 = ~w28151 & w28152;
assign w28154 = ~w28149 & ~w28153;
assign w28155 = ~w28144 & ~w28154;
assign w28156 = ~pi1522 & w28155;
assign w28157 = pi1522 & ~w28155;
assign w28158 = ~w28156 & ~w28157;
assign w28159 = ~w27789 & ~w27816;
assign w28160 = w27797 & w27816;
assign w28161 = ~w28159 & ~w28160;
assign w28162 = ~w27834 & ~w28159;
assign w28163 = ~w27823 & ~w28162;
assign w28164 = (~w27806 & w28161) | (~w27806 & w65777) | (w28161 & w65777);
assign w28165 = w28163 & w28164;
assign w28166 = w27777 & ~w28165;
assign w28167 = ~w27789 & w27804;
assign w28168 = (w28167 & w27852) | (w28167 & w63838) | (w27852 & w63838);
assign w28169 = ~w27805 & ~w27845;
assign w28170 = w27842 & ~w28169;
assign w28171 = ~w27812 & ~w27821;
assign w28172 = ~w27840 & ~w27850;
assign w28173 = (w28172 & w65778) | (w28172 & w65779) | (w65778 & w65779);
assign w28174 = w27783 & ~w27839;
assign w28175 = w28169 & w28174;
assign w28176 = ~w28170 & ~w28175;
assign w28177 = ~w28173 & w28176;
assign w28178 = ~w27777 & ~w28177;
assign w28179 = ~w28166 & ~w28168;
assign w28180 = w28179 & w65780;
assign w28181 = (pi1510 & ~w28179) | (pi1510 & w65781) | (~w28179 & w65781);
assign w28182 = ~w28180 & ~w28181;
assign w28183 = ~pi5059 & pi9040;
assign w28184 = ~pi4963 & ~pi9040;
assign w28185 = ~w28183 & ~w28184;
assign w28186 = pi1494 & ~w28185;
assign w28187 = ~pi1494 & w28185;
assign w28188 = ~w28186 & ~w28187;
assign w28189 = ~pi4840 & pi9040;
assign w28190 = ~pi4923 & ~pi9040;
assign w28191 = ~w28189 & ~w28190;
assign w28192 = pi1490 & ~w28191;
assign w28193 = ~pi1490 & w28191;
assign w28194 = ~w28192 & ~w28193;
assign w28195 = w28188 & w28194;
assign w28196 = ~pi4846 & pi9040;
assign w28197 = ~pi4962 & ~pi9040;
assign w28198 = ~w28196 & ~w28197;
assign w28199 = pi1499 & ~w28198;
assign w28200 = ~pi1499 & w28198;
assign w28201 = ~w28199 & ~w28200;
assign w28202 = ~pi4838 & pi9040;
assign w28203 = ~pi4984 & ~pi9040;
assign w28204 = ~w28202 & ~w28203;
assign w28205 = pi1467 & ~w28204;
assign w28206 = ~pi1467 & w28204;
assign w28207 = ~w28205 & ~w28206;
assign w28208 = w28201 & ~w28207;
assign w28209 = ~pi4923 & pi9040;
assign w28210 = ~pi4943 & ~pi9040;
assign w28211 = ~w28209 & ~w28210;
assign w28212 = pi1491 & ~w28211;
assign w28213 = ~pi1491 & w28211;
assign w28214 = ~w28212 & ~w28213;
assign w28215 = w28208 & ~w28214;
assign w28216 = ~w28195 & ~w28215;
assign w28217 = w28208 & w28214;
assign w28218 = (~w28214 & ~w28208) | (~w28214 & w63840) | (~w28208 & w63840);
assign w28219 = ~w28217 & ~w28218;
assign w28220 = ~w28216 & ~w28219;
assign w28221 = ~w28201 & w28207;
assign w28222 = ~w28208 & ~w28221;
assign w28223 = w28188 & w28201;
assign w28224 = ~w28222 & ~w28223;
assign w28225 = ~w28194 & w28224;
assign w28226 = ~w28220 & ~w28225;
assign w28227 = ~pi5116 & pi9040;
assign w28228 = ~pi4882 & ~pi9040;
assign w28229 = ~w28227 & ~w28228;
assign w28230 = pi1482 & ~w28229;
assign w28231 = ~pi1482 & w28229;
assign w28232 = ~w28230 & ~w28231;
assign w28233 = ~w28226 & ~w28232;
assign w28234 = ~w28188 & w28201;
assign w28235 = w28207 & w28234;
assign w28236 = (w28194 & ~w28234) | (w28194 & w28241) | (~w28234 & w28241);
assign w28237 = (~w28194 & ~w28208) | (~w28194 & w65782) | (~w28208 & w65782);
assign w28238 = ~w28236 & ~w28237;
assign w28239 = w28207 & w28214;
assign w28240 = ~w28194 & w28207;
assign w28241 = w28194 & ~w28207;
assign w28242 = ~w28188 & ~w28241;
assign w28243 = ~w28239 & ~w28240;
assign w28244 = w28242 & w28243;
assign w28245 = w28232 & ~w28244;
assign w28246 = w28238 & ~w28245;
assign w28247 = ~w28188 & ~w28201;
assign w28248 = ~w28240 & ~w28247;
assign w28249 = w28214 & ~w28242;
assign w28250 = ~w28248 & w28249;
assign w28251 = ~w28188 & w28194;
assign w28252 = w28239 & ~w28251;
assign w28253 = ~w28201 & ~w28207;
assign w28254 = ~w28194 & w28253;
assign w28255 = w28188 & w28254;
assign w28256 = w28223 & w28240;
assign w28257 = w28195 & ~w28222;
assign w28258 = (~w28247 & w28222) | (~w28247 & w63398) | (w28222 & w63398);
assign w28259 = w28195 & w28221;
assign w28260 = ~w28256 & ~w28259;
assign w28261 = ~w28188 & w28221;
assign w28262 = w28221 & w65783;
assign w28263 = w28260 & ~w28262;
assign w28264 = ~w28214 & ~w28258;
assign w28265 = w28263 & w28264;
assign w28266 = ~w28252 & ~w28256;
assign w28267 = ~w28255 & w28266;
assign w28268 = ~w28265 & w28267;
assign w28269 = w28232 & ~w28268;
assign w28270 = ~w28246 & ~w28250;
assign w28271 = ~w28233 & w28270;
assign w28272 = ~w28269 & w28271;
assign w28273 = ~pi1519 & ~w28272;
assign w28274 = pi1519 & w28272;
assign w28275 = ~w28273 & ~w28274;
assign w28276 = w27577 & w27624;
assign w28277 = w27622 & w27630;
assign w28278 = ~w27584 & ~w27606;
assign w28279 = w28129 & ~w28138;
assign w28280 = ~w28277 & w28279;
assign w28281 = ~w28132 & ~w28278;
assign w28282 = ~w28280 & w28281;
assign w28283 = w27623 & w28282;
assign w28284 = w27600 & ~w28276;
assign w28285 = ~w28277 & w28284;
assign w28286 = ~w28283 & w28285;
assign w28287 = ~w27611 & ~w27624;
assign w28288 = ~w28129 & w28287;
assign w28289 = w27571 & w28288;
assign w28290 = ~w27590 & w28136;
assign w28291 = ~w27600 & ~w28289;
assign w28292 = ~w28290 & w28291;
assign w28293 = w28282 & w28292;
assign w28294 = ~w28286 & ~w28293;
assign w28295 = pi1521 & w28294;
assign w28296 = ~pi1521 & ~w28294;
assign w28297 = ~w28295 & ~w28296;
assign w28298 = w27738 & ~w28105;
assign w28299 = ~w27726 & ~w27742;
assign w28300 = w28298 & ~w28299;
assign w28301 = (w27719 & w28105) | (w27719 & w63841) | (w28105 & w63841);
assign w28302 = w27735 & w28102;
assign w28303 = ~w27758 & ~w28302;
assign w28304 = ~w28301 & w28303;
assign w28305 = ~w28300 & w28304;
assign w28306 = ~w27709 & ~w28103;
assign w28307 = ~w27702 & w27742;
assign w28308 = w27709 & ~w27745;
assign w28309 = ~w28307 & w28308;
assign w28310 = ~w28306 & ~w28309;
assign w28311 = (w28306 & ~w28304) | (w28306 & w65784) | (~w28304 & w65784);
assign w28312 = ~w27690 & ~w28298;
assign w28313 = ~w28311 & w28312;
assign w28314 = (~w28310 & w28305) | (~w28310 & w65785) | (w28305 & w65785);
assign w28315 = ~w28313 & w28314;
assign w28316 = pi1520 & w28315;
assign w28317 = ~pi1520 & ~w28315;
assign w28318 = ~w28316 & ~w28317;
assign w28319 = ~w27892 & w65786;
assign w28320 = w27906 & w27925;
assign w28321 = ~w28319 & ~w28320;
assign w28322 = ~w27882 & ~w28321;
assign w28323 = w27906 & w27908;
assign w28324 = ~w28319 & ~w28323;
assign w28325 = ~w27870 & w28088;
assign w28326 = ~w27929 & ~w27942;
assign w28327 = w27919 & ~w28326;
assign w28328 = w27936 & ~w28325;
assign w28329 = w28324 & w28328;
assign w28330 = ~w28327 & w28329;
assign w28331 = ~w27892 & w28082;
assign w28332 = w27906 & w27921;
assign w28333 = ~w27936 & ~w28332;
assign w28334 = ~w27951 & w28333;
assign w28335 = ~w28331 & w28334;
assign w28336 = ~w28090 & w28335;
assign w28337 = ~w28330 & ~w28336;
assign w28338 = w27940 & ~w28322;
assign w28339 = ~w28337 & w28338;
assign w28340 = ~pi1526 & w28339;
assign w28341 = pi1526 & ~w28339;
assign w28342 = ~w28340 & ~w28341;
assign w28343 = ~w28188 & ~w28208;
assign w28344 = ~w28236 & w28343;
assign w28345 = ~w28214 & w28344;
assign w28346 = w28223 & w28239;
assign w28347 = ~w28254 & ~w28346;
assign w28348 = ~w28244 & w28347;
assign w28349 = ~w28257 & w28348;
assign w28350 = w28348 & w63842;
assign w28351 = w28214 & w28344;
assign w28352 = ~w28242 & ~w28258;
assign w28353 = ~w28201 & w28241;
assign w28354 = w28218 & ~w28353;
assign w28355 = ~w28343 & w28354;
assign w28356 = ~w28351 & ~w28352;
assign w28357 = w28214 & ~w28234;
assign w28358 = w28356 & w63843;
assign w28359 = ~w28345 & ~w28350;
assign w28360 = ~w28358 & w28359;
assign w28361 = w28232 & ~w28360;
assign w28362 = (~w28232 & ~w28356) | (~w28232 & w65787) | (~w28356 & w65787);
assign w28363 = w28234 & w28241;
assign w28364 = ~w28352 & ~w28363;
assign w28365 = w28218 & ~w28364;
assign w28366 = ~w28362 & ~w28365;
assign w28367 = ~w28361 & w65788;
assign w28368 = (pi1517 & w28361) | (pi1517 & w65789) | (w28361 & w65789);
assign w28369 = ~w28367 & ~w28368;
assign w28370 = ~w27777 & w27783;
assign w28371 = ~w27822 & ~w28370;
assign w28372 = ~w27795 & ~w28167;
assign w28373 = w27844 & ~w28371;
assign w28374 = ~w28372 & w28373;
assign w28375 = ~w27840 & ~w27849;
assign w28376 = ~w28163 & ~w28375;
assign w28377 = ~w27777 & w27818;
assign w28378 = w27832 & w28169;
assign w28379 = w27777 & ~w28160;
assign w28380 = ~w27847 & w28379;
assign w28381 = ~w28378 & w28380;
assign w28382 = ~w27826 & w28381;
assign w28383 = ~w28377 & ~w28382;
assign w28384 = ~w27843 & ~w28374;
assign w28385 = ~w28376 & w28384;
assign w28386 = ~w28383 & w28385;
assign w28387 = ~pi1516 & w28386;
assign w28388 = pi1516 & ~w28386;
assign w28389 = ~w28387 & ~w28388;
assign w28390 = ~w28169 & w28171;
assign w28391 = ~w27840 & ~w28390;
assign w28392 = w27820 & w28391;
assign w28393 = w27777 & w27815;
assign w28394 = ~w27783 & ~w27805;
assign w28395 = (w28172 & w65790) | (w28172 & w65791) | (w65790 & w65791);
assign w28396 = ~w28390 & ~w28395;
assign w28397 = ~w28393 & ~w28396;
assign w28398 = ~w27777 & w28169;
assign w28399 = w27824 & w28398;
assign w28400 = (~w28392 & w65792) | (~w28392 & w65793) | (w65792 & w65793);
assign w28401 = ~w28397 & w28400;
assign w28402 = pi1507 & w28401;
assign w28403 = ~pi1507 & ~w28401;
assign w28404 = ~w28402 & ~w28403;
assign w28405 = ~pi4909 & pi9040;
assign w28406 = ~pi5039 & ~pi9040;
assign w28407 = ~w28405 & ~w28406;
assign w28408 = pi1473 & ~w28407;
assign w28409 = ~pi1473 & w28407;
assign w28410 = ~w28408 & ~w28409;
assign w28411 = ~pi4837 & pi9040;
assign w28412 = ~pi4834 & ~pi9040;
assign w28413 = ~w28411 & ~w28412;
assign w28414 = pi1475 & ~w28413;
assign w28415 = ~pi1475 & w28413;
assign w28416 = ~w28414 & ~w28415;
assign w28417 = ~pi4834 & pi9040;
assign w28418 = ~pi4833 & ~pi9040;
assign w28419 = ~w28417 & ~w28418;
assign w28420 = pi1482 & ~w28419;
assign w28421 = ~pi1482 & w28419;
assign w28422 = ~w28420 & ~w28421;
assign w28423 = ~pi4961 & pi9040;
assign w28424 = ~pi4835 & ~pi9040;
assign w28425 = ~w28423 & ~w28424;
assign w28426 = pi1500 & ~w28425;
assign w28427 = ~pi1500 & w28425;
assign w28428 = ~w28426 & ~w28427;
assign w28429 = ~w28422 & ~w28428;
assign w28430 = w28422 & w28428;
assign w28431 = ~w28429 & ~w28430;
assign w28432 = ~pi4882 & pi9040;
assign w28433 = ~pi5059 & ~pi9040;
assign w28434 = ~w28432 & ~w28433;
assign w28435 = pi1477 & ~w28434;
assign w28436 = ~pi1477 & w28434;
assign w28437 = ~w28435 & ~w28436;
assign w28438 = ~pi4984 & pi9040;
assign w28439 = ~pi4846 & ~pi9040;
assign w28440 = ~w28438 & ~w28439;
assign w28441 = pi1499 & ~w28440;
assign w28442 = ~pi1499 & w28440;
assign w28443 = ~w28441 & ~w28442;
assign w28444 = ~w28437 & ~w28443;
assign w28445 = (~w28444 & w28431) | (~w28444 & w65794) | (w28431 & w65794);
assign w28446 = ~w28422 & w28428;
assign w28447 = ~w28416 & w28446;
assign w28448 = w28422 & ~w28428;
assign w28449 = ~w28447 & ~w28448;
assign w28450 = ~w28447 & w65795;
assign w28451 = ~w28445 & ~w28450;
assign w28452 = w28410 & w28451;
assign w28453 = w28422 & w28437;
assign w28454 = ~w28443 & w28447;
assign w28455 = w28428 & ~w28443;
assign w28456 = w28429 & w28437;
assign w28457 = ~w28437 & w28448;
assign w28458 = ~w28456 & ~w28457;
assign w28459 = ~w28431 & w65796;
assign w28460 = w28458 & w28459;
assign w28461 = ~w28454 & ~w28460;
assign w28462 = w28453 & ~w28461;
assign w28463 = ~w28437 & w28446;
assign w28464 = ~w28443 & w28453;
assign w28465 = w28429 & w28443;
assign w28466 = ~w28464 & ~w28465;
assign w28467 = ~w28463 & w28466;
assign w28468 = w28466 & w65797;
assign w28469 = ~w28428 & w28443;
assign w28470 = ~w28455 & ~w28469;
assign w28471 = w28422 & w28470;
assign w28472 = ~w28410 & ~w28416;
assign w28473 = (w28472 & ~w28470) | (w28472 & w65798) | (~w28470 & w65798);
assign w28474 = ~w28437 & w28443;
assign w28475 = w28410 & w28416;
assign w28476 = ~w28474 & w28475;
assign w28477 = ~w28473 & ~w28476;
assign w28478 = w28468 & ~w28477;
assign w28479 = ~w28458 & ~w28474;
assign w28480 = ~w28463 & ~w28479;
assign w28481 = ~w28422 & ~w28443;
assign w28482 = w28416 & ~w28429;
assign w28483 = ~w28481 & w28482;
assign w28484 = ~w28480 & w28483;
assign w28485 = ~w28410 & ~w28447;
assign w28486 = ~w28451 & w28485;
assign w28487 = ~w28468 & w28486;
assign w28488 = ~w28452 & ~w28478;
assign w28489 = ~w28484 & w28488;
assign w28490 = ~w28462 & ~w28487;
assign w28491 = w28489 & w28490;
assign w28492 = pi1533 & ~w28491;
assign w28493 = ~pi1533 & w28491;
assign w28494 = ~w28492 & ~w28493;
assign w28495 = w28429 & w28444;
assign w28496 = ~w28455 & ~w28495;
assign w28497 = w28467 & ~w28496;
assign w28498 = ~w28453 & ~w28469;
assign w28499 = w28437 & w28469;
assign w28500 = w28416 & ~w28498;
assign w28501 = ~w28499 & w28500;
assign w28502 = ~w28497 & ~w28501;
assign w28503 = ~w28410 & ~w28502;
assign w28504 = w28437 & w28443;
assign w28505 = w28410 & w28504;
assign w28506 = w28469 & w65799;
assign w28507 = ~w28505 & ~w28506;
assign w28508 = ~w28430 & ~w28507;
assign w28509 = w28475 & ~w28480;
assign w28510 = w28472 & w28498;
assign w28511 = w28416 & w28437;
assign w28512 = w28455 & w28511;
assign w28513 = ~w28510 & ~w28512;
assign w28514 = ~w28481 & ~w28513;
assign w28515 = w28410 & ~w28416;
assign w28516 = ~w28453 & ~w28465;
assign w28517 = w28515 & ~w28516;
assign w28518 = ~w28508 & ~w28517;
assign w28519 = ~w28514 & w28518;
assign w28520 = ~w28509 & w28519;
assign w28521 = ~w28503 & w28520;
assign w28522 = pi1532 & ~w28521;
assign w28523 = ~pi1532 & w28521;
assign w28524 = ~w28522 & ~w28523;
assign w28525 = ~w28238 & w28263;
assign w28526 = w28194 & w28234;
assign w28527 = (w28214 & ~w28253) | (w28214 & w65800) | (~w28253 & w65800);
assign w28528 = ~w28526 & w28527;
assign w28529 = ~w28354 & ~w28528;
assign w28530 = (w28232 & ~w28525) | (w28232 & w65801) | (~w28525 & w65801);
assign w28531 = ~w28261 & ~w28363;
assign w28532 = ~w28255 & w28531;
assign w28533 = ~w28232 & ~w28532;
assign w28534 = w28260 & ~w28533;
assign w28535 = ~w28214 & ~w28534;
assign w28536 = ~w28214 & ~w28235;
assign w28537 = ~w28232 & ~w28536;
assign w28538 = w28532 & w28537;
assign w28539 = w28525 & w28538;
assign w28540 = ~w28530 & ~w28539;
assign w28541 = ~w28535 & w28540;
assign w28542 = pi1525 & w28541;
assign w28543 = ~pi1525 & ~w28541;
assign w28544 = ~w28542 & ~w28543;
assign w28545 = ~w28001 & w28016;
assign w28546 = ~w28030 & ~w28545;
assign w28547 = ~w28057 & w28546;
assign w28548 = w28061 & ~w28547;
assign w28549 = ~w28042 & ~w28045;
assign w28550 = ~w28027 & w28549;
assign w28551 = w27989 & ~w28550;
assign w28552 = w27989 & ~w28024;
assign w28553 = w27989 & w28015;
assign w28554 = w28028 & ~w28553;
assign w28555 = ~w28552 & w28554;
assign w28556 = ~w28551 & ~w28555;
assign w28557 = ~w28037 & ~w28556;
assign w28558 = ~w28014 & w28061;
assign w28559 = w28008 & w28014;
assign w28560 = ~w28061 & w28559;
assign w28561 = ~w28001 & ~w28558;
assign w28562 = ~w28560 & w28561;
assign w28563 = w28001 & ~w28019;
assign w28564 = ~w28026 & w28563;
assign w28565 = w28037 & ~w28562;
assign w28566 = ~w28564 & w28565;
assign w28567 = ~w28002 & ~w28045;
assign w28568 = ~w28017 & w28567;
assign w28569 = w28059 & ~w28568;
assign w28570 = ~w27989 & ~w28545;
assign w28571 = ~w28569 & w28570;
assign w28572 = ~w28548 & ~w28571;
assign w28573 = ~w28566 & w28572;
assign w28574 = ~w28557 & w28573;
assign w28575 = pi1553 & ~w28574;
assign w28576 = ~pi1553 & w28574;
assign w28577 = ~w28575 & ~w28576;
assign w28578 = ~w27876 & w27898;
assign w28579 = ~w27906 & w27922;
assign w28580 = ~w28578 & w28579;
assign w28581 = ~w28078 & ~w28580;
assign w28582 = w27936 & ~w28581;
assign w28583 = ~w27907 & ~w27911;
assign w28584 = ~w27922 & ~w28080;
assign w28585 = ~w28583 & w28584;
assign w28586 = (~w27936 & w27916) | (~w27936 & w65802) | (w27916 & w65802);
assign w28587 = ~w27927 & ~w28324;
assign w28588 = ~w27941 & ~w27950;
assign w28589 = w27899 & ~w28588;
assign w28590 = ~w28582 & ~w28589;
assign w28591 = ~w28587 & w28590;
assign w28592 = ~w28586 & w28591;
assign w28593 = pi1537 & w28592;
assign w28594 = ~pi1537 & ~w28592;
assign w28595 = ~w28593 & ~w28594;
assign w28596 = w28017 & ~w28041;
assign w28597 = ~w28044 & ~w28568;
assign w28598 = ~w28596 & w28597;
assign w28599 = w28037 & ~w28598;
assign w28600 = w28025 & w65803;
assign w28601 = ~w28014 & ~w28569;
assign w28602 = w28020 & w28049;
assign w28603 = ~w28002 & ~w28041;
assign w28604 = w28559 & ~w28603;
assign w28605 = ~w28602 & ~w28604;
assign w28606 = (w28049 & w28604) | (w28049 & w65804) | (w28604 & w65804);
assign w28607 = ~w28037 & ~w28057;
assign w28608 = ~w28600 & w28607;
assign w28609 = ~w28601 & ~w28606;
assign w28610 = w28608 & w28609;
assign w28611 = ~w28599 & ~w28610;
assign w28612 = w28016 & w28045;
assign w28613 = w27995 & w28020;
assign w28614 = ~w28037 & ~w28613;
assign w28615 = w28059 & w28614;
assign w28616 = w27989 & ~w28615;
assign w28617 = ~w28612 & ~w28616;
assign w28618 = ~w28056 & ~w28058;
assign w28619 = w28037 & ~w28545;
assign w28620 = w28047 & w28619;
assign w28621 = w28618 & w28620;
assign w28622 = ~w28617 & ~w28621;
assign w28623 = (pi1527 & w28611) | (pi1527 & w65805) | (w28611 & w65805);
assign w28624 = ~w28611 & w65806;
assign w28625 = ~w28623 & ~w28624;
assign w28626 = w27611 & ~w28130;
assign w28627 = (~w27584 & ~w28130) | (~w27584 & w63845) | (~w28130 & w63845);
assign w28628 = ~w27631 & ~w28627;
assign w28629 = ~w28626 & ~w28628;
assign w28630 = ~w27570 & ~w27593;
assign w28631 = (w27584 & ~w27605) | (w27584 & w65807) | (~w27605 & w65807);
assign w28632 = ~w28630 & w28631;
assign w28633 = w27592 & w28133;
assign w28634 = (~w28633 & w28629) | (~w28633 & w65808) | (w28629 & w65808);
assign w28635 = w27600 & ~w28634;
assign w28636 = w27625 & w28129;
assign w28637 = w27584 & ~w28636;
assign w28638 = w27570 & w27605;
assign w28639 = w28138 & ~w28638;
assign w28640 = ~w28637 & ~w28639;
assign w28641 = ~w27622 & w27629;
assign w28642 = ~w27570 & ~w28132;
assign w28643 = w28632 & ~w28642;
assign w28644 = w28278 & ~w28626;
assign w28645 = ~w27607 & ~w28641;
assign w28646 = ~w28644 & w28645;
assign w28647 = ~w28643 & w28646;
assign w28648 = (~w28640 & w28647) | (~w28640 & w65809) | (w28647 & w65809);
assign w28649 = ~w28635 & w28648;
assign w28650 = ~pi1530 & w28649;
assign w28651 = pi1530 & ~w28649;
assign w28652 = ~w28650 & ~w28651;
assign w28653 = ~w27740 & ~w27742;
assign w28654 = w27709 & ~w28653;
assign w28655 = ~w27709 & ~w27736;
assign w28656 = (~w27718 & ~w28655) | (~w27718 & w63846) | (~w28655 & w63846);
assign w28657 = ~w27741 & ~w28656;
assign w28658 = (~w27690 & w28657) | (~w27690 & w65810) | (w28657 & w65810);
assign w28659 = ~w28104 & ~w28107;
assign w28660 = ~w28307 & ~w28659;
assign w28661 = ~w27709 & ~w28660;
assign w28662 = ~w27739 & w28104;
assign w28663 = w27756 & w28662;
assign w28664 = ~w27736 & ~w27758;
assign w28665 = ~w28116 & w28664;
assign w28666 = ~w28663 & w28665;
assign w28667 = w27690 & ~w28666;
assign w28668 = ~w27696 & ~w28112;
assign w28669 = w27761 & w28668;
assign w28670 = ~w28667 & ~w28669;
assign w28671 = ~w28658 & w28670;
assign w28672 = (pi1540 & ~w28671) | (pi1540 & w65811) | (~w28671 & w65811);
assign w28673 = w28671 & w65812;
assign w28674 = ~w28672 & ~w28673;
assign w28675 = w28429 & w28505;
assign w28676 = w28416 & w28446;
assign w28677 = ~w28474 & w28676;
assign w28678 = ~w28444 & ~w28504;
assign w28679 = ~w28449 & w28678;
assign w28680 = ~w28431 & ~w28678;
assign w28681 = ~w28410 & ~w28677;
assign w28682 = ~w28680 & w28681;
assign w28683 = ~w28679 & w28682;
assign w28684 = ~w28429 & ~w28470;
assign w28685 = w28446 & ~w28678;
assign w28686 = ~w28684 & ~w28685;
assign w28687 = w28475 & ~w28686;
assign w28688 = ~w28429 & w28515;
assign w28689 = w28686 & w28688;
assign w28690 = w28416 & w28495;
assign w28691 = ~w28512 & ~w28675;
assign w28692 = ~w28690 & w28691;
assign w28693 = ~w28687 & w28692;
assign w28694 = ~w28689 & w28693;
assign w28695 = ~w28683 & w28694;
assign w28696 = pi1531 & ~w28695;
assign w28697 = ~pi1531 & w28695;
assign w28698 = ~w28696 & ~w28697;
assign w28699 = w28429 & w65813;
assign w28700 = (~w28437 & w28471) | (~w28437 & w65814) | (w28471 & w65814);
assign w28701 = ~w28685 & ~w28700;
assign w28702 = w28410 & ~w28701;
assign w28703 = (~w28464 & w28458) | (~w28464 & w65815) | (w28458 & w65815);
assign w28704 = ~w28416 & ~w28703;
assign w28705 = ~w28428 & w28511;
assign w28706 = w28466 & w28705;
assign w28707 = ~w28471 & w28483;
assign w28708 = ~w28495 & ~w28707;
assign w28709 = w28461 & w28708;
assign w28710 = ~w28410 & ~w28709;
assign w28711 = ~w28704 & ~w28706;
assign w28712 = ~w28702 & w28711;
assign w28713 = ~w28710 & w28712;
assign w28714 = pi1523 & ~w28713;
assign w28715 = ~pi1523 & w28713;
assign w28716 = ~w28714 & ~w28715;
assign w28717 = ~w28613 & w28618;
assign w28718 = ~w27989 & ~w28717;
assign w28719 = ~w28549 & w28552;
assign w28720 = w28547 & ~w28719;
assign w28721 = ~w28718 & w28720;
assign w28722 = w28037 & ~w28721;
assign w28723 = ~w28001 & w28553;
assign w28724 = ~w28025 & w28051;
assign w28725 = w28605 & ~w28724;
assign w28726 = ~w28037 & ~w28725;
assign w28727 = ~w28043 & ~w28723;
assign w28728 = ~w28600 & w28727;
assign w28729 = ~w28726 & w28728;
assign w28730 = ~w28722 & w28729;
assign w28731 = ~pi1543 & w28730;
assign w28732 = pi1543 & ~w28730;
assign w28733 = ~w28731 & ~w28732;
assign w28734 = ~w28232 & ~w28349;
assign w28735 = w28214 & w28224;
assign w28736 = w28194 & ~w28253;
assign w28737 = w28188 & ~w28214;
assign w28738 = ~w28221 & w28737;
assign w28739 = ~w28251 & ~w28738;
assign w28740 = ~w28736 & ~w28739;
assign w28741 = ~w28735 & ~w28740;
assign w28742 = w28232 & ~w28741;
assign w28743 = w28195 & w28201;
assign w28744 = w28214 & ~w28743;
assign w28745 = ~w28262 & w28744;
assign w28746 = ~w28536 & ~w28745;
assign w28747 = ~w28734 & ~w28746;
assign w28748 = ~w28742 & w28747;
assign w28749 = ~pi1557 & w28748;
assign w28750 = pi1557 & ~w28748;
assign w28751 = ~w28749 & ~w28750;
assign w28752 = ~pi5151 & pi9040;
assign w28753 = ~pi5065 & ~pi9040;
assign w28754 = ~w28752 & ~w28753;
assign w28755 = pi1539 & ~w28754;
assign w28756 = ~pi1539 & w28754;
assign w28757 = ~w28755 & ~w28756;
assign w28758 = ~pi5075 & pi9040;
assign w28759 = ~pi5245 & ~pi9040;
assign w28760 = ~w28758 & ~w28759;
assign w28761 = pi1528 & ~w28760;
assign w28762 = ~pi1528 & w28760;
assign w28763 = ~w28761 & ~w28762;
assign w28764 = ~w28757 & ~w28763;
assign w28765 = ~pi5255 & pi9040;
assign w28766 = ~pi5067 & ~pi9040;
assign w28767 = ~w28765 & ~w28766;
assign w28768 = pi1558 & ~w28767;
assign w28769 = ~pi1558 & w28767;
assign w28770 = ~w28768 & ~w28769;
assign w28771 = ~w28757 & w28770;
assign w28772 = ~w28764 & ~w28771;
assign w28773 = ~pi5065 & pi9040;
assign w28774 = ~pi5262 & ~pi9040;
assign w28775 = ~w28773 & ~w28774;
assign w28776 = pi1560 & ~w28775;
assign w28777 = ~pi1560 & w28775;
assign w28778 = ~w28776 & ~w28777;
assign w28779 = ~w28772 & w28778;
assign w28780 = w28763 & ~w28778;
assign w28781 = ~w28771 & w28780;
assign w28782 = ~w28779 & ~w28781;
assign w28783 = w28763 & w28778;
assign w28784 = ~w28763 & ~w28778;
assign w28785 = ~w28783 & ~w28784;
assign w28786 = ~pi5262 & pi9040;
assign w28787 = ~pi5194 & ~pi9040;
assign w28788 = ~w28786 & ~w28787;
assign w28789 = pi1542 & ~w28788;
assign w28790 = ~pi1542 & w28788;
assign w28791 = ~w28789 & ~w28790;
assign w28792 = ~w28785 & ~w28791;
assign w28793 = ~w28778 & w28791;
assign w28794 = (~w28770 & ~w28793) | (~w28770 & w28815) | (~w28793 & w28815);
assign w28795 = ~w28792 & w28794;
assign w28796 = w28782 & w28795;
assign w28797 = ~w28782 & ~w28791;
assign w28798 = ~pi5194 & pi9040;
assign w28799 = ~pi5112 & ~pi9040;
assign w28800 = ~w28798 & ~w28799;
assign w28801 = pi1551 & ~w28800;
assign w28802 = ~pi1551 & w28800;
assign w28803 = ~w28801 & ~w28802;
assign w28804 = w28757 & w28763;
assign w28805 = w28778 & w28791;
assign w28806 = w28804 & w28805;
assign w28807 = ~w28803 & ~w28806;
assign w28808 = ~w28796 & w28807;
assign w28809 = ~w28797 & w28808;
assign w28810 = ~w28757 & w28791;
assign w28811 = w28780 & w28810;
assign w28812 = ~w28757 & w28783;
assign w28813 = w28783 & w28810;
assign w28814 = ~w28770 & ~w28813;
assign w28815 = ~w28757 & ~w28770;
assign w28816 = ~w28764 & ~w28804;
assign w28817 = ~w28778 & ~w28815;
assign w28818 = ~w28816 & w28817;
assign w28819 = ~w28812 & ~w28818;
assign w28820 = w28814 & ~w28819;
assign w28821 = w28770 & w28778;
assign w28822 = ~w28791 & w28804;
assign w28823 = ~w28810 & ~w28822;
assign w28824 = w28821 & ~w28823;
assign w28825 = ~w28757 & ~w28791;
assign w28826 = w28784 & w28825;
assign w28827 = w28803 & ~w28811;
assign w28828 = ~w28826 & w28827;
assign w28829 = ~w28824 & w28828;
assign w28830 = ~w28820 & w28829;
assign w28831 = w28793 & w28816;
assign w28832 = w28764 & ~w28793;
assign w28833 = ~w28831 & ~w28832;
assign w28834 = w28770 & ~w28833;
assign w28835 = w28778 & ~w28791;
assign w28836 = ~w28793 & ~w28835;
assign w28837 = w28757 & ~w28770;
assign w28838 = w28836 & w28837;
assign w28839 = ~w28834 & ~w28838;
assign w28840 = (w28839 & w28809) | (w28839 & w65816) | (w28809 & w65816);
assign w28841 = ~pi1571 & w28840;
assign w28842 = pi1571 & ~w28840;
assign w28843 = ~w28841 & ~w28842;
assign w28844 = ~pi5312 & pi9040;
assign w28845 = ~pi5078 & ~pi9040;
assign w28846 = ~w28844 & ~w28845;
assign w28847 = pi1547 & ~w28846;
assign w28848 = ~pi1547 & w28846;
assign w28849 = ~w28847 & ~w28848;
assign w28850 = ~pi5314 & pi9040;
assign w28851 = ~pi5117 & ~pi9040;
assign w28852 = ~w28850 & ~w28851;
assign w28853 = pi1529 & ~w28852;
assign w28854 = ~pi1529 & w28852;
assign w28855 = ~w28853 & ~w28854;
assign w28856 = ~w28849 & ~w28855;
assign w28857 = w28849 & w28855;
assign w28858 = ~w28856 & ~w28857;
assign w28859 = ~pi5144 & pi9040;
assign w28860 = ~pi5302 & ~pi9040;
assign w28861 = ~w28859 & ~w28860;
assign w28862 = pi1564 & ~w28861;
assign w28863 = ~pi1564 & w28861;
assign w28864 = ~w28862 & ~w28863;
assign w28865 = ~pi5064 & pi9040;
assign w28866 = ~pi5069 & ~pi9040;
assign w28867 = ~w28865 & ~w28866;
assign w28868 = pi1562 & ~w28867;
assign w28869 = ~pi1562 & w28867;
assign w28870 = ~w28868 & ~w28869;
assign w28871 = w28864 & w28870;
assign w28872 = w28855 & ~w28870;
assign w28873 = ~w28855 & w28870;
assign w28874 = ~w28872 & ~w28873;
assign w28875 = ~w28864 & ~w28874;
assign w28876 = (~w28871 & w28874) | (~w28871 & w63847) | (w28874 & w63847);
assign w28877 = ~w28858 & ~w28876;
assign w28878 = ~pi5066 & pi9040;
assign w28879 = ~pi5193 & ~pi9040;
assign w28880 = ~w28878 & ~w28879;
assign w28881 = pi1548 & ~w28880;
assign w28882 = ~pi1548 & w28880;
assign w28883 = ~w28881 & ~w28882;
assign w28884 = w28849 & ~w28870;
assign w28885 = ~w28855 & w28864;
assign w28886 = w28884 & w28885;
assign w28887 = ~w28849 & ~w28864;
assign w28888 = ~w28872 & w28887;
assign w28889 = ~w28886 & ~w28888;
assign w28890 = ~w28883 & ~w28889;
assign w28891 = ~w28877 & ~w28890;
assign w28892 = ~pi5193 & pi9040;
assign w28893 = ~pi5267 & ~pi9040;
assign w28894 = ~w28892 & ~w28893;
assign w28895 = pi1563 & ~w28894;
assign w28896 = ~pi1563 & w28894;
assign w28897 = ~w28895 & ~w28896;
assign w28898 = ~w28891 & ~w28897;
assign w28899 = w28872 & w28897;
assign w28900 = w28871 & ~w28897;
assign w28901 = ~w28864 & w28897;
assign w28902 = w28858 & w28901;
assign w28903 = w28855 & w28864;
assign w28904 = ~w28870 & ~w28903;
assign w28905 = w28889 & w28904;
assign w28906 = ~w28899 & ~w28900;
assign w28907 = ~w28902 & w28906;
assign w28908 = ~w28905 & w28907;
assign w28909 = w28883 & ~w28908;
assign w28910 = w28864 & w28897;
assign w28911 = ~w28849 & ~w28870;
assign w28912 = w28910 & w28911;
assign w28913 = ~w28855 & ~w28864;
assign w28914 = ~w28903 & ~w28913;
assign w28915 = w28849 & w28870;
assign w28916 = w28897 & w28915;
assign w28917 = w28914 & w28916;
assign w28918 = w28903 & w28911;
assign w28919 = ~w28917 & ~w28918;
assign w28920 = ~w28873 & ~w28910;
assign w28921 = ~w28849 & ~w28885;
assign w28922 = ~w28920 & w28921;
assign w28923 = w28919 & ~w28922;
assign w28924 = ~w28883 & ~w28923;
assign w28925 = w28884 & ~w28914;
assign w28926 = w28901 & w28925;
assign w28927 = ~w28912 & ~w28926;
assign w28928 = ~w28909 & w28927;
assign w28929 = w28928 & w65817;
assign w28930 = pi1575 & ~w28929;
assign w28931 = ~pi1575 & w28929;
assign w28932 = ~w28930 & ~w28931;
assign w28933 = ~pi5155 & pi9040;
assign w28934 = ~pi5250 & ~pi9040;
assign w28935 = ~w28933 & ~w28934;
assign w28936 = pi1561 & ~w28935;
assign w28937 = ~pi1561 & w28935;
assign w28938 = ~w28936 & ~w28937;
assign w28939 = ~pi5253 & pi9040;
assign w28940 = ~pi5192 & ~pi9040;
assign w28941 = ~w28939 & ~w28940;
assign w28942 = pi1551 & ~w28941;
assign w28943 = ~pi1551 & w28941;
assign w28944 = ~w28942 & ~w28943;
assign w28945 = ~w28938 & w28944;
assign w28946 = ~pi5440 & pi9040;
assign w28947 = ~pi5164 & ~pi9040;
assign w28948 = ~w28946 & ~w28947;
assign w28949 = pi1562 & ~w28948;
assign w28950 = ~pi1562 & w28948;
assign w28951 = ~w28949 & ~w28950;
assign w28952 = ~pi5156 & pi9040;
assign w28953 = ~pi5076 & ~pi9040;
assign w28954 = ~w28952 & ~w28953;
assign w28955 = pi1528 & ~w28954;
assign w28956 = ~pi1528 & w28954;
assign w28957 = ~w28955 & ~w28956;
assign w28958 = ~w28951 & w28957;
assign w28959 = ~w28945 & ~w28958;
assign w28960 = w28938 & w28951;
assign w28961 = w28951 & ~w28957;
assign w28962 = w28938 & ~w28944;
assign w28963 = w28958 & w28962;
assign w28964 = ~w28960 & ~w28961;
assign w28965 = ~w28963 & w28964;
assign w28966 = ~w28959 & ~w28965;
assign w28967 = ~w28944 & ~w28957;
assign w28968 = w28938 & ~w28951;
assign w28969 = w28944 & w28957;
assign w28970 = ~w28967 & ~w28969;
assign w28971 = w28968 & ~w28970;
assign w28972 = w28951 & w28967;
assign w28973 = w28967 & w65818;
assign w28974 = ~w28971 & w65819;
assign w28975 = ~w28966 & ~w28974;
assign w28976 = ~pi5182 & pi9040;
assign w28977 = ~pi5439 & ~pi9040;
assign w28978 = ~w28976 & ~w28977;
assign w28979 = pi1534 & ~w28978;
assign w28980 = ~pi1534 & w28978;
assign w28981 = ~w28979 & ~w28980;
assign w28982 = ~w28975 & w28981;
assign w28983 = ~w28957 & ~w28981;
assign w28984 = ~w28945 & ~w28962;
assign w28985 = w28983 & w28984;
assign w28986 = ~pi5112 & pi9040;
assign w28987 = ~pi5058 & ~pi9040;
assign w28988 = ~w28986 & ~w28987;
assign w28989 = pi1564 & ~w28988;
assign w28990 = ~pi1564 & w28988;
assign w28991 = ~w28989 & ~w28990;
assign w28992 = w28938 & ~w28957;
assign w28993 = ~w28958 & ~w28992;
assign w28994 = w28962 & w28993;
assign w28995 = (w28991 & ~w28993) | (w28991 & w65820) | (~w28993 & w65820);
assign w28996 = w28944 & w28958;
assign w28997 = w28981 & ~w28996;
assign w28998 = w28945 & ~w28997;
assign w28999 = ~w28959 & w28981;
assign w29000 = ~w28998 & w28999;
assign w29001 = ~w28985 & w28995;
assign w29002 = ~w29000 & w29001;
assign w29003 = ~w28951 & ~w28981;
assign w29004 = w28962 & w29003;
assign w29005 = w28944 & ~w28957;
assign w29006 = w28968 & w29005;
assign w29007 = ~w28972 & ~w29006;
assign w29008 = w28981 & ~w29007;
assign w29009 = w28951 & ~w28981;
assign w29010 = w28944 & w28960;
assign w29011 = ~w29009 & ~w29010;
assign w29012 = w28957 & ~w29011;
assign w29013 = ~w28991 & ~w29004;
assign w29014 = ~w28998 & w29013;
assign w29015 = ~w29008 & ~w29012;
assign w29016 = w29014 & w29015;
assign w29017 = ~w29002 & ~w29016;
assign w29018 = w28945 & w28957;
assign w29019 = w29003 & w29018;
assign w29020 = ~w28982 & ~w29019;
assign w29021 = ~w29017 & w29020;
assign w29022 = pi1568 & w29021;
assign w29023 = ~pi1568 & ~w29021;
assign w29024 = ~w29022 & ~w29023;
assign w29025 = ~pi5192 & pi9040;
assign w29026 = ~pi5182 & ~pi9040;
assign w29027 = ~w29025 & ~w29026;
assign w29028 = pi1565 & ~w29027;
assign w29029 = ~pi1565 & w29027;
assign w29030 = ~w29028 & ~w29029;
assign w29031 = ~pi5439 & pi9040;
assign w29032 = ~pi5072 & ~pi9040;
assign w29033 = ~w29031 & ~w29032;
assign w29034 = pi1567 & ~w29033;
assign w29035 = ~pi1567 & w29033;
assign w29036 = ~w29034 & ~w29035;
assign w29037 = ~w29030 & ~w29036;
assign w29038 = ~w29030 & w29036;
assign w29039 = ~pi5164 & pi9040;
assign w29040 = ~pi5155 & ~pi9040;
assign w29041 = ~w29039 & ~w29040;
assign w29042 = pi1556 & ~w29041;
assign w29043 = ~pi1556 & w29041;
assign w29044 = ~w29042 & ~w29043;
assign w29045 = ~pi5058 & pi9040;
assign w29046 = ~pi5083 & ~pi9040;
assign w29047 = ~w29045 & ~w29046;
assign w29048 = pi1536 & ~w29047;
assign w29049 = ~pi1536 & w29047;
assign w29050 = ~w29048 & ~w29049;
assign w29051 = ~w29044 & ~w29050;
assign w29052 = w29038 & w29051;
assign w29053 = w29030 & ~w29036;
assign w29054 = ~w29044 & w29050;
assign w29055 = w29053 & w29054;
assign w29056 = ~w29052 & ~w29055;
assign w29057 = ~pi5076 & pi9040;
assign w29058 = ~pi5440 & ~pi9040;
assign w29059 = ~w29057 & ~w29058;
assign w29060 = pi1538 & ~w29059;
assign w29061 = ~pi1538 & w29059;
assign w29062 = ~w29060 & ~w29061;
assign w29063 = ~w29056 & w29062;
assign w29064 = (~w29037 & w29056) | (~w29037 & w65821) | (w29056 & w65821);
assign w29065 = w29030 & w29036;
assign w29066 = w29054 & w29065;
assign w29067 = ~w29030 & ~w29050;
assign w29068 = w29030 & w29050;
assign w29069 = ~w29044 & ~w29068;
assign w29070 = ~w29038 & ~w29053;
assign w29071 = w29069 & ~w29070;
assign w29072 = w29044 & w29068;
assign w29073 = ~w29067 & ~w29072;
assign w29074 = ~w29071 & w29073;
assign w29075 = w29062 & ~w29074;
assign w29076 = w29037 & w29050;
assign w29077 = w29030 & ~w29050;
assign w29078 = w29044 & w29077;
assign w29079 = ~w29076 & ~w29078;
assign w29080 = ~w29062 & ~w29079;
assign w29081 = w29044 & w29050;
assign w29082 = ~w29036 & w29081;
assign w29083 = ~w29066 & ~w29082;
assign w29084 = ~w29080 & w29083;
assign w29085 = ~w29075 & w29084;
assign w29086 = ~w29038 & ~w29051;
assign w29087 = w29062 & ~w29081;
assign w29088 = ~w29067 & ~w29086;
assign w29089 = ~w29087 & w29088;
assign w29090 = ~pi5083 & pi9040;
assign w29091 = ~pi5156 & ~pi9040;
assign w29092 = ~w29090 & ~w29091;
assign w29093 = pi1546 & ~w29092;
assign w29094 = ~pi1546 & w29092;
assign w29095 = ~w29093 & ~w29094;
assign w29096 = (w29085 & w65822) | (w29085 & w65823) | (w65822 & w65823);
assign w29097 = w29053 & w29081;
assign w29098 = ~w29085 & w29095;
assign w29099 = (w29062 & ~w29037) | (w29062 & w65824) | (~w29037 & w65824);
assign w29100 = w29037 & w29044;
assign w29101 = ~w29030 & ~w29062;
assign w29102 = w29081 & w29101;
assign w29103 = ~w29052 & ~w29066;
assign w29104 = ~w29076 & ~w29102;
assign w29105 = w29103 & w29104;
assign w29106 = (w29099 & ~w29105) | (w29099 & w65825) | (~w29105 & w65825);
assign w29107 = w29036 & ~w29050;
assign w29108 = w29030 & ~w29062;
assign w29109 = w29107 & w29108;
assign w29110 = ~w29097 & ~w29109;
assign w29111 = ~w29106 & w29110;
assign w29112 = ~w29098 & w29111;
assign w29113 = w29112 & w65826;
assign w29114 = (~pi1570 & ~w29112) | (~pi1570 & w65827) | (~w29112 & w65827);
assign w29115 = ~w29113 & ~w29114;
assign w29116 = ~pi5068 & pi9040;
assign w29117 = ~pi5312 & ~pi9040;
assign w29118 = ~w29116 & ~w29117;
assign w29119 = pi1549 & ~w29118;
assign w29120 = ~pi1549 & w29118;
assign w29121 = ~w29119 & ~w29120;
assign w29122 = ~pi5061 & pi9040;
assign w29123 = ~pi5062 & ~pi9040;
assign w29124 = ~w29122 & ~w29123;
assign w29125 = pi1536 & ~w29124;
assign w29126 = ~pi1536 & w29124;
assign w29127 = ~w29125 & ~w29126;
assign w29128 = ~w29121 & w29127;
assign w29129 = ~pi5089 & pi9040;
assign w29130 = ~pi5074 & ~pi9040;
assign w29131 = ~w29129 & ~w29130;
assign w29132 = pi1550 & ~w29131;
assign w29133 = ~pi1550 & w29131;
assign w29134 = ~w29132 & ~w29133;
assign w29135 = ~w29128 & ~w29134;
assign w29136 = w29121 & ~w29127;
assign w29137 = ~pi5315 & pi9040;
assign w29138 = ~pi5061 & ~pi9040;
assign w29139 = ~w29137 & ~w29138;
assign w29140 = pi1554 & ~w29139;
assign w29141 = ~pi1554 & w29139;
assign w29142 = ~w29140 & ~w29141;
assign w29143 = ~pi5070 & pi9040;
assign w29144 = ~pi5195 & ~pi9040;
assign w29145 = ~w29143 & ~w29144;
assign w29146 = pi1566 & ~w29145;
assign w29147 = ~pi1566 & w29145;
assign w29148 = ~w29146 & ~w29147;
assign w29149 = ~w29142 & ~w29148;
assign w29150 = w29134 & ~w29148;
assign w29151 = ~w29149 & ~w29150;
assign w29152 = w29136 & ~w29151;
assign w29153 = ~w29128 & w29134;
assign w29154 = ~w29136 & w29142;
assign w29155 = ~w29153 & w29154;
assign w29156 = ~w29148 & w29155;
assign w29157 = ~w29152 & ~w29156;
assign w29158 = w29135 & ~w29157;
assign w29159 = ~pi5355 & pi9040;
assign w29160 = ~pi5073 & ~pi9040;
assign w29161 = ~w29159 & ~w29160;
assign w29162 = pi1565 & ~w29161;
assign w29163 = ~pi1565 & w29161;
assign w29164 = ~w29162 & ~w29163;
assign w29165 = ~w29121 & ~w29127;
assign w29166 = w29121 & ~w29142;
assign w29167 = ~w29121 & w29142;
assign w29168 = ~w29166 & ~w29167;
assign w29169 = ~w29134 & ~w29168;
assign w29170 = ~w29165 & w29169;
assign w29171 = w29142 & w29148;
assign w29172 = ~w29155 & w29171;
assign w29173 = ~w29121 & w29134;
assign w29174 = w29127 & ~w29173;
assign w29175 = w29149 & ~w29174;
assign w29176 = ~w29164 & ~w29175;
assign w29177 = ~w29170 & w29176;
assign w29178 = ~w29172 & w29177;
assign w29179 = ~w29127 & w29134;
assign w29180 = ~w29173 & ~w29179;
assign w29181 = ~w29135 & w29180;
assign w29182 = ~w29151 & w29181;
assign w29183 = ~w29134 & w29165;
assign w29184 = w29142 & w29183;
assign w29185 = ~w29142 & w29148;
assign w29186 = w29165 & w29185;
assign w29187 = ~w29165 & ~w29166;
assign w29188 = ~w29149 & ~w29180;
assign w29189 = w29187 & w29188;
assign w29190 = w29164 & ~w29186;
assign w29191 = ~w29184 & w29190;
assign w29192 = ~w29182 & w29191;
assign w29193 = ~w29189 & w29192;
assign w29194 = ~w29178 & ~w29193;
assign w29195 = w29127 & ~w29134;
assign w29196 = w29148 & w29195;
assign w29197 = ~w29168 & w29196;
assign w29198 = ~w29158 & ~w29197;
assign w29199 = ~w29194 & w29198;
assign w29200 = pi1573 & ~w29199;
assign w29201 = ~pi1573 & w29199;
assign w29202 = ~w29200 & ~w29201;
assign w29203 = w28757 & w28791;
assign w29204 = w28785 & w29203;
assign w29205 = ~w28813 & ~w29204;
assign w29206 = w28763 & ~w29205;
assign w29207 = w28771 & w28780;
assign w29208 = ~w28805 & w28816;
assign w29209 = ~w28770 & ~w29208;
assign w29210 = ~w28757 & ~w28836;
assign w29211 = ~w28764 & w28792;
assign w29212 = ~w29210 & ~w29211;
assign w29213 = ~w28763 & ~w29212;
assign w29214 = ~w28803 & ~w29207;
assign w29215 = ~w29209 & w29214;
assign w29216 = ~w29206 & w29215;
assign w29217 = ~w29213 & w29216;
assign w29218 = w28757 & w28784;
assign w29219 = ~w28832 & ~w29218;
assign w29220 = w28791 & ~w29219;
assign w29221 = ~w28791 & ~w28819;
assign w29222 = ~w28811 & ~w28821;
assign w29223 = ~w28771 & ~w29222;
assign w29224 = w28803 & ~w29220;
assign w29225 = ~w29223 & w29224;
assign w29226 = ~w29221 & w29225;
assign w29227 = ~w29217 & ~w29226;
assign w29228 = pi1572 & w29227;
assign w29229 = ~pi1572 & ~w29227;
assign w29230 = ~w29228 & ~w29229;
assign w29231 = ~pi5250 & pi9040;
assign w29232 = ~pi5189 & ~pi9040;
assign w29233 = ~w29231 & ~w29232;
assign w29234 = pi1541 & ~w29233;
assign w29235 = ~pi1541 & w29233;
assign w29236 = ~w29234 & ~w29235;
assign w29237 = ~pi5067 & pi9040;
assign w29238 = ~pi5253 & ~pi9040;
assign w29239 = ~w29237 & ~w29238;
assign w29240 = pi1535 & ~w29239;
assign w29241 = ~pi1535 & w29239;
assign w29242 = ~w29240 & ~w29241;
assign w29243 = ~pi5188 & pi9040;
assign w29244 = ~pi5075 & ~pi9040;
assign w29245 = ~w29243 & ~w29244;
assign w29246 = pi1546 & ~w29245;
assign w29247 = ~pi1546 & w29245;
assign w29248 = ~w29246 & ~w29247;
assign w29249 = ~w29242 & ~w29248;
assign w29250 = ~pi5245 & pi9040;
assign w29251 = ~pi5143 & ~pi9040;
assign w29252 = ~w29250 & ~w29251;
assign w29253 = pi1539 & ~w29252;
assign w29254 = ~pi1539 & w29252;
assign w29255 = ~w29253 & ~w29254;
assign w29256 = ~pi5189 & pi9040;
assign w29257 = ~pi5079 & ~pi9040;
assign w29258 = ~w29256 & ~w29257;
assign w29259 = pi1556 & ~w29258;
assign w29260 = ~pi1556 & w29258;
assign w29261 = ~w29259 & ~w29260;
assign w29262 = ~w29255 & w29261;
assign w29263 = w29255 & ~w29261;
assign w29264 = ~w29262 & ~w29263;
assign w29265 = w29249 & ~w29264;
assign w29266 = w29242 & w29248;
assign w29267 = w29255 & w29266;
assign w29268 = ~w29265 & ~w29267;
assign w29269 = ~w29242 & ~w29255;
assign w29270 = ~w29249 & ~w29262;
assign w29271 = ~w29248 & ~w29255;
assign w29272 = ~w29270 & ~w29271;
assign w29273 = (w29261 & w29270) | (w29261 & w65828) | (w29270 & w65828);
assign w29274 = ~w29269 & ~w29273;
assign w29275 = w29248 & w29264;
assign w29276 = (~w29242 & ~w29264) | (~w29242 & w29249) | (~w29264 & w29249);
assign w29277 = ~pi5326 & pi9040;
assign w29278 = ~pi5255 & ~pi9040;
assign w29279 = ~w29277 & ~w29278;
assign w29280 = pi1560 & ~w29279;
assign w29281 = ~pi1560 & w29279;
assign w29282 = ~w29280 & ~w29281;
assign w29283 = ~w29276 & w29282;
assign w29284 = ~w29274 & w29283;
assign w29285 = w29268 & ~w29284;
assign w29286 = w29236 & ~w29285;
assign w29287 = ~w29236 & w29282;
assign w29288 = ~w29265 & w65829;
assign w29289 = w29274 & w29288;
assign w29290 = ~w29236 & ~w29242;
assign w29291 = ~w29270 & w29290;
assign w29292 = ~w29236 & w29248;
assign w29293 = w29269 & w29292;
assign w29294 = w29248 & w29255;
assign w29295 = w29242 & ~w29261;
assign w29296 = w29294 & w29295;
assign w29297 = ~w29293 & ~w29296;
assign w29298 = ~w29242 & w29261;
assign w29299 = w29271 & ~w29298;
assign w29300 = ~w29267 & ~w29299;
assign w29301 = ~w29236 & ~w29300;
assign w29302 = w29297 & ~w29301;
assign w29303 = (w29291 & w29301) | (w29291 & w65830) | (w29301 & w65830);
assign w29304 = w29236 & ~w29248;
assign w29305 = w29248 & w29262;
assign w29306 = ~w29304 & ~w29305;
assign w29307 = ~w29242 & ~w29306;
assign w29308 = ~w29249 & ~w29266;
assign w29309 = ~w29236 & w29261;
assign w29310 = w29308 & w29309;
assign w29311 = w29263 & w29304;
assign w29312 = w29248 & ~w29261;
assign w29313 = w29236 & w29242;
assign w29314 = w29312 & w29313;
assign w29315 = ~w29311 & ~w29314;
assign w29316 = w29297 & w29315;
assign w29317 = ~w29310 & w29316;
assign w29318 = (~w29282 & ~w29317) | (~w29282 & w65831) | (~w29317 & w65831);
assign w29319 = ~w29289 & ~w29303;
assign w29320 = ~w29318 & w29319;
assign w29321 = ~w29286 & w29320;
assign w29322 = ~pi1588 & ~w29321;
assign w29323 = pi1588 & w29321;
assign w29324 = ~w29322 & ~w29323;
assign w29325 = w29164 & w29187;
assign w29326 = ~w29134 & w29136;
assign w29327 = (w29142 & w29181) | (w29142 & w63399) | (w29181 & w63399);
assign w29328 = (~w29148 & ~w29136) | (~w29148 & w29150) | (~w29136 & w29150);
assign w29329 = w29127 & w29166;
assign w29330 = w29328 & ~w29329;
assign w29331 = w29166 & w29179;
assign w29332 = (w29148 & ~w29165) | (w29148 & w63400) | (~w29165 & w63400);
assign w29333 = ~w29331 & w29332;
assign w29334 = ~w29330 & ~w29333;
assign w29335 = ~w29327 & ~w29334;
assign w29336 = (w29148 & ~w63401) | (w29148 & w63849) | (~w63401 & w63849);
assign w29337 = ~w29164 & ~w29165;
assign w29338 = w29328 & w29337;
assign w29339 = (~w29154 & w29336) | (~w29154 & w65832) | (w29336 & w65832);
assign w29340 = ~w29127 & w29173;
assign w29341 = w29149 & w29340;
assign w29342 = w29142 & w29181;
assign w29343 = ~w29168 & w65833;
assign w29344 = w29164 & ~w29341;
assign w29345 = ~w29342 & w29344;
assign w29346 = ~w29343 & w29345;
assign w29347 = w29121 & w29195;
assign w29348 = ~w29340 & ~w29347;
assign w29349 = ~w29168 & ~w29348;
assign w29350 = w29128 & w29343;
assign w29351 = w29165 & w65834;
assign w29352 = w29148 & w29154;
assign w29353 = ~w29169 & w29352;
assign w29354 = ~w29164 & ~w29186;
assign w29355 = ~w29351 & w29354;
assign w29356 = ~w29349 & w29355;
assign w29357 = w29356 & w65835;
assign w29358 = ~w29346 & ~w29357;
assign w29359 = ~w29339 & ~w29358;
assign w29360 = ~pi1582 & w29359;
assign w29361 = pi1582 & ~w29359;
assign w29362 = ~w29360 & ~w29361;
assign w29363 = w29127 & w29134;
assign w29364 = w29168 & w29363;
assign w29365 = ~w29351 & ~w29364;
assign w29366 = ~w29148 & ~w29365;
assign w29367 = ~w29173 & ~w29326;
assign w29368 = w29171 & ~w29367;
assign w29369 = w29135 & w29168;
assign w29370 = ~w29148 & ~w29348;
assign w29371 = ~w29166 & ~w29195;
assign w29372 = w29148 & ~w29347;
assign w29373 = ~w29371 & w29372;
assign w29374 = w29167 & w29179;
assign w29375 = ~w29164 & ~w29374;
assign w29376 = ~w29369 & w29375;
assign w29377 = ~w29370 & w29376;
assign w29378 = ~w29373 & w29377;
assign w29379 = (w29148 & w29349) | (w29148 & w65836) | (w29349 & w65836);
assign w29380 = ~w29152 & w29164;
assign w29381 = ~w29364 & w29380;
assign w29382 = ~w29350 & w29381;
assign w29383 = ~w29379 & w29382;
assign w29384 = ~w29366 & ~w29368;
assign w29385 = (w29384 & w29383) | (w29384 & w65837) | (w29383 & w65837);
assign w29386 = pi1584 & ~w29385;
assign w29387 = ~pi1584 & w29385;
assign w29388 = ~w29386 & ~w29387;
assign w29389 = w28870 & w28902;
assign w29390 = ~w28856 & w28870;
assign w29391 = ~w28897 & ~w28914;
assign w29392 = ~w29390 & w29391;
assign w29393 = ~w28874 & w28914;
assign w29394 = w28849 & w29393;
assign w29395 = w28874 & w28910;
assign w29396 = ~w28883 & ~w29395;
assign w29397 = ~w29392 & w29396;
assign w29398 = ~w29394 & w29397;
assign w29399 = w28856 & w28871;
assign w29400 = w28883 & ~w29399;
assign w29401 = ~w28864 & ~w28911;
assign w29402 = ~w28849 & w28864;
assign w29403 = ~w28897 & ~w29402;
assign w29404 = ~w29401 & w29403;
assign w29405 = ~w28918 & ~w29401;
assign w29406 = w28897 & ~w29405;
assign w29407 = w28857 & w28870;
assign w29408 = w29400 & ~w29407;
assign w29409 = ~w29404 & w29408;
assign w29410 = ~w29406 & w29409;
assign w29411 = ~w29398 & ~w29410;
assign w29412 = ~w29389 & ~w29411;
assign w29413 = ~pi1576 & w29412;
assign w29414 = pi1576 & ~w29412;
assign w29415 = ~w29413 & ~w29414;
assign w29416 = ~pi5190 & pi9040;
assign w29417 = ~pi5314 & ~pi9040;
assign w29418 = ~w29416 & ~w29417;
assign w29419 = pi1545 & ~w29418;
assign w29420 = ~pi1545 & w29418;
assign w29421 = ~w29419 & ~w29420;
assign w29422 = ~pi5195 & pi9040;
assign w29423 = ~pi5190 & ~pi9040;
assign w29424 = ~w29422 & ~w29423;
assign w29425 = pi1559 & ~w29424;
assign w29426 = ~pi1559 & w29424;
assign w29427 = ~w29425 & ~w29426;
assign w29428 = ~w29421 & ~w29427;
assign w29429 = ~pi5196 & pi9040;
assign w29430 = ~pi5154 & ~pi9040;
assign w29431 = ~w29429 & ~w29430;
assign w29432 = pi1548 & ~w29431;
assign w29433 = ~pi1548 & w29431;
assign w29434 = ~w29432 & ~w29433;
assign w29435 = w29428 & ~w29434;
assign w29436 = w29421 & ~w29434;
assign w29437 = ~pi5117 & pi9040;
assign w29438 = ~pi5416 & ~pi9040;
assign w29439 = ~w29437 & ~w29438;
assign w29440 = pi1529 & ~w29439;
assign w29441 = ~pi1529 & w29439;
assign w29442 = ~w29440 & ~w29441;
assign w29443 = w29436 & w29442;
assign w29444 = ~w29435 & ~w29443;
assign w29445 = ~pi5078 & pi9040;
assign w29446 = ~pi5066 & ~pi9040;
assign w29447 = ~w29445 & ~w29446;
assign w29448 = pi1552 & ~w29447;
assign w29449 = ~pi1552 & w29447;
assign w29450 = ~w29448 & ~w29449;
assign w29451 = ~w29444 & w29450;
assign w29452 = ~w29421 & w29434;
assign w29453 = ~w29436 & ~w29452;
assign w29454 = w29427 & ~w29442;
assign w29455 = w29453 & w29454;
assign w29456 = ~w29421 & w29442;
assign w29457 = w29427 & w29434;
assign w29458 = w29456 & w29457;
assign w29459 = ~pi5252 & pi9040;
assign w29460 = ~pi5068 & ~pi9040;
assign w29461 = ~w29459 & ~w29460;
assign w29462 = pi1544 & ~w29461;
assign w29463 = ~pi1544 & w29461;
assign w29464 = ~w29462 & ~w29463;
assign w29465 = ~w29458 & ~w29464;
assign w29466 = ~w29455 & w29465;
assign w29467 = ~w29451 & w29466;
assign w29468 = w29427 & ~w29434;
assign w29469 = ~w29442 & w29468;
assign w29470 = w29421 & w29469;
assign w29471 = w29442 & w29450;
assign w29472 = ~w29468 & w29471;
assign w29473 = w29444 & ~w29450;
assign w29474 = w29450 & ~w29456;
assign w29475 = ~w29452 & w29474;
assign w29476 = ~w29472 & ~w29475;
assign w29477 = ~w29473 & w29476;
assign w29478 = ~w29427 & w29434;
assign w29479 = w29421 & ~w29442;
assign w29480 = w29434 & w29479;
assign w29481 = ~w29450 & ~w29480;
assign w29482 = w29478 & ~w29481;
assign w29483 = w29421 & w29442;
assign w29484 = w29434 & w29450;
assign w29485 = w29483 & w29484;
assign w29486 = w29464 & ~w29485;
assign w29487 = ~w29470 & w29486;
assign w29488 = ~w29482 & w29487;
assign w29489 = ~w29477 & w29488;
assign w29490 = ~w29467 & ~w29489;
assign w29491 = w29453 & ~w29483;
assign w29492 = ~w29421 & w29454;
assign w29493 = ~w29443 & ~w29464;
assign w29494 = ~w29492 & w29493;
assign w29495 = ~w29491 & w29494;
assign w29496 = ~w29458 & ~w29469;
assign w29497 = ~w29495 & w29496;
assign w29498 = ~w29450 & ~w29497;
assign w29499 = ~w29490 & ~w29498;
assign w29500 = ~pi1569 & w29499;
assign w29501 = pi1569 & ~w29499;
assign w29502 = ~w29500 & ~w29501;
assign w29503 = ~w29265 & ~w29271;
assign w29504 = w29274 & ~w29503;
assign w29505 = ~w29248 & w29261;
assign w29506 = ~w29299 & w29505;
assign w29507 = w29262 & w29266;
assign w29508 = (w29236 & w29506) | (w29236 & w65838) | (w29506 & w65838);
assign w29509 = w29302 & ~w29508;
assign w29510 = (w29282 & ~w29509) | (w29282 & w65839) | (~w29509 & w65839);
assign w29511 = ~w29294 & ~w29505;
assign w29512 = ~w29242 & ~w29511;
assign w29513 = ~w29507 & ~w29512;
assign w29514 = ~w29236 & ~w29282;
assign w29515 = ~w29513 & w29514;
assign w29516 = w29242 & w29255;
assign w29517 = ~w29282 & w29516;
assign w29518 = w29511 & w29517;
assign w29519 = w29269 & w29312;
assign w29520 = w29255 & ~w29290;
assign w29521 = w29298 & w29520;
assign w29522 = ~w29295 & ~w29300;
assign w29523 = ~w29275 & ~w29522;
assign w29524 = w29236 & ~w29282;
assign w29525 = ~w29523 & w29524;
assign w29526 = ~w29518 & ~w29519;
assign w29527 = ~w29521 & w29526;
assign w29528 = ~w29515 & w29527;
assign w29529 = ~w29525 & w29528;
assign w29530 = ~w29510 & w29529;
assign w29531 = pi1577 & w29530;
assign w29532 = ~pi1577 & ~w29530;
assign w29533 = ~w29531 & ~w29532;
assign w29534 = w29044 & ~w29067;
assign w29535 = ~w29534 & w65840;
assign w29536 = w29062 & w29535;
assign w29537 = w29037 & w29051;
assign w29538 = ~w29078 & ~w29537;
assign w29539 = w29062 & ~w29538;
assign w29540 = ~w29108 & ~w29535;
assign w29541 = ~w29065 & ~w29540;
assign w29542 = ~w29539 & ~w29541;
assign w29543 = w29095 & ~w29542;
assign w29544 = (~w29062 & ~w29037) | (~w29062 & w65841) | (~w29037 & w65841);
assign w29545 = ~w29078 & w29544;
assign w29546 = (w29062 & ~w29068) | (w29062 & w65842) | (~w29068 & w65842);
assign w29547 = w29051 & w29053;
assign w29548 = w29546 & ~w29547;
assign w29549 = ~w29545 & ~w29548;
assign w29550 = w29105 & ~w29549;
assign w29551 = ~w29095 & ~w29550;
assign w29552 = ~w29068 & ~w29100;
assign w29553 = w29546 & ~w29552;
assign w29554 = w29051 & w29065;
assign w29555 = (~w29554 & w29552) | (~w29554 & w65843) | (w29552 & w65843);
assign w29556 = ~w29099 & ~w29555;
assign w29557 = ~w29536 & ~w29556;
assign w29558 = ~w29551 & w29557;
assign w29559 = ~w29543 & w29558;
assign w29560 = pi1580 & ~w29559;
assign w29561 = ~pi1580 & w29559;
assign w29562 = ~w29560 & ~w29561;
assign w29563 = ~pi5073 & pi9040;
assign w29564 = ~pi5196 & ~pi9040;
assign w29565 = ~w29563 & ~w29564;
assign w29566 = pi1554 & ~w29565;
assign w29567 = ~pi1554 & w29565;
assign w29568 = ~w29566 & ~w29567;
assign w29569 = ~pi5416 & pi9040;
assign w29570 = ~pi5071 & ~pi9040;
assign w29571 = ~w29569 & ~w29570;
assign w29572 = pi1544 & ~w29571;
assign w29573 = ~pi1544 & w29571;
assign w29574 = ~w29572 & ~w29573;
assign w29575 = w29568 & ~w29574;
assign w29576 = ~pi5267 & pi9040;
assign w29577 = ~pi5144 & ~pi9040;
assign w29578 = ~w29576 & ~w29577;
assign w29579 = pi1545 & ~w29578;
assign w29580 = ~pi1545 & w29578;
assign w29581 = ~w29579 & ~w29580;
assign w29582 = ~pi5069 & pi9040;
assign w29583 = ~pi5315 & ~pi9040;
assign w29584 = ~w29582 & ~w29583;
assign w29585 = pi1555 & ~w29584;
assign w29586 = ~pi1555 & w29584;
assign w29587 = ~w29585 & ~w29586;
assign w29588 = w29581 & w29587;
assign w29589 = ~pi5154 & pi9040;
assign w29590 = ~pi5252 & ~pi9040;
assign w29591 = ~w29589 & ~w29590;
assign w29592 = pi1549 & ~w29591;
assign w29593 = ~pi1549 & w29591;
assign w29594 = ~w29592 & ~w29593;
assign w29595 = w29588 & w29594;
assign w29596 = w29575 & w29595;
assign w29597 = ~w29574 & ~w29581;
assign w29598 = w29574 & w29581;
assign w29599 = ~w29597 & ~w29598;
assign w29600 = w29568 & ~w29599;
assign w29601 = ~w29568 & ~w29574;
assign w29602 = ~w29587 & w29601;
assign w29603 = ~pi5152 & pi9040;
assign w29604 = ~pi5089 & ~pi9040;
assign w29605 = ~w29603 & ~w29604;
assign w29606 = pi1524 & ~w29605;
assign w29607 = ~pi1524 & w29605;
assign w29608 = ~w29606 & ~w29607;
assign w29609 = (~w29608 & w29600) | (~w29608 & w65844) | (w29600 & w65844);
assign w29610 = ~w29568 & w29608;
assign w29611 = ~w29568 & w29574;
assign w29612 = ~w29610 & ~w29611;
assign w29613 = w29599 & ~w29612;
assign w29614 = ~w29600 & ~w29613;
assign w29615 = w29587 & w29601;
assign w29616 = ~w29597 & ~w29608;
assign w29617 = ~w29615 & ~w29616;
assign w29618 = w29614 & w29617;
assign w29619 = ~w29609 & ~w29618;
assign w29620 = ~w29594 & ~w29619;
assign w29621 = ~w29587 & w29594;
assign w29622 = ~w29614 & w29621;
assign w29623 = ~w29599 & w29610;
assign w29624 = ~w29581 & w29616;
assign w29625 = ~w29623 & ~w29624;
assign w29626 = w29587 & ~w29625;
assign w29627 = w29574 & w29587;
assign w29628 = w29594 & ~w29608;
assign w29629 = ~w29568 & ~w29627;
assign w29630 = w29628 & w29629;
assign w29631 = ~w29602 & w29630;
assign w29632 = ~w29596 & ~w29631;
assign w29633 = ~w29622 & w29632;
assign w29634 = ~w29626 & w29633;
assign w29635 = ~w29620 & w29634;
assign w29636 = pi1597 & ~w29635;
assign w29637 = ~pi1597 & w29635;
assign w29638 = ~w29636 & ~w29637;
assign w29639 = ~w29575 & ~w29611;
assign w29640 = w29568 & w29587;
assign w29641 = ~w29598 & ~w29640;
assign w29642 = ~w29639 & ~w29641;
assign w29643 = ~w29581 & ~w29587;
assign w29644 = w29639 & w29643;
assign w29645 = ~w29642 & ~w29644;
assign w29646 = ~w29608 & ~w29645;
assign w29647 = ~w29574 & w29608;
assign w29648 = ~w29568 & w29581;
assign w29649 = ~w29627 & ~w29648;
assign w29650 = ~w29598 & ~w29649;
assign w29651 = ~w29647 & ~w29650;
assign w29652 = ~w29608 & ~w29643;
assign w29653 = w29639 & w29652;
assign w29654 = ~w29639 & ~w29647;
assign w29655 = ~w29639 & w63850;
assign w29656 = ~w29575 & ~w29643;
assign w29657 = ~w29602 & ~w29640;
assign w29658 = ~w29602 & w63851;
assign w29659 = (w29608 & ~w29656) | (w29608 & w63852) | (~w29656 & w63852);
assign w29660 = ~w29658 & w29659;
assign w29661 = ~w29653 & ~w29655;
assign w29662 = ~w29660 & w29661;
assign w29663 = ~w29651 & w29662;
assign w29664 = (~w29594 & w29663) | (~w29594 & w65845) | (w29663 & w65845);
assign w29665 = w29609 & w29627;
assign w29666 = w29594 & ~w29662;
assign w29667 = ~w29581 & ~w29645;
assign w29668 = ~w29608 & ~w29649;
assign w29669 = w29587 & w29648;
assign w29670 = ~w29649 & ~w29669;
assign w29671 = ~w29616 & ~w29670;
assign w29672 = ~w29668 & ~w29671;
assign w29673 = ~w29667 & ~w29672;
assign w29674 = w29568 & ~w29581;
assign w29675 = ~w29642 & ~w29674;
assign w29676 = ~w29656 & w29675;
assign w29677 = w29673 & w29676;
assign w29678 = ~w29665 & ~w29666;
assign w29679 = ~w29677 & w29678;
assign w29680 = (pi1581 & ~w29679) | (pi1581 & w65846) | (~w29679 & w65846);
assign w29681 = w29679 & w65847;
assign w29682 = ~w29680 & ~w29681;
assign w29683 = w29595 & ~w29600;
assign w29684 = ~w29594 & ~w29673;
assign w29685 = w29594 & w29608;
assign w29686 = ~w29655 & ~w29658;
assign w29687 = w29685 & ~w29686;
assign w29688 = ~w29581 & w29608;
assign w29689 = ~w29657 & w29688;
assign w29690 = ~w29669 & ~w29689;
assign w29691 = ~w29671 & ~w29690;
assign w29692 = (~w29627 & w29649) | (~w29627 & w65848) | (w29649 & w65848);
assign w29693 = w29628 & ~w29692;
assign w29694 = ~w29683 & ~w29693;
assign w29695 = ~w29687 & w29694;
assign w29696 = ~w29691 & w29695;
assign w29697 = ~w29684 & w29696;
assign w29698 = pi1587 & ~w29697;
assign w29699 = ~pi1587 & w29697;
assign w29700 = ~w29698 & ~w29699;
assign w29701 = w29101 & w29535;
assign w29702 = w29077 & w65849;
assign w29703 = ~w29547 & ~w29702;
assign w29704 = ~w29534 & w65850;
assign w29705 = ~w29062 & ~w29704;
assign w29706 = ~w29097 & w29703;
assign w29707 = w29705 & w29706;
assign w29708 = w29030 & ~w29044;
assign w29709 = ~w29051 & ~w29065;
assign w29710 = ~w29708 & ~w29709;
assign w29711 = w29099 & ~w29710;
assign w29712 = ~w29095 & ~w29711;
assign w29713 = ~w29707 & w29712;
assign w29714 = ~w29055 & ~w29077;
assign w29715 = w29703 & ~w29714;
assign w29716 = ~w29710 & w65851;
assign w29717 = w29070 & ~w29107;
assign w29718 = w29705 & w29717;
assign w29719 = ~w29715 & ~w29716;
assign w29720 = ~w29718 & w29719;
assign w29721 = w29095 & ~w29720;
assign w29722 = ~w29063 & ~w29701;
assign w29723 = ~w29713 & w29722;
assign w29724 = ~w29721 & w29723;
assign w29725 = ~pi1583 & ~w29724;
assign w29726 = pi1583 & w29724;
assign w29727 = ~w29725 & ~w29726;
assign w29728 = ~w29165 & ~w29179;
assign w29729 = w29185 & w29728;
assign w29730 = ~w29156 & ~w29729;
assign w29731 = w29164 & ~w29730;
assign w29732 = ~w29127 & ~w29148;
assign w29733 = ~w29164 & ~w29732;
assign w29734 = w29168 & ~w29180;
assign w29735 = ~w29733 & w29734;
assign w29736 = ~w29164 & ~w29335;
assign w29737 = ~w29364 & ~w29374;
assign w29738 = w29148 & ~w29737;
assign w29739 = ~w29735 & ~w29738;
assign w29740 = ~w29731 & w29739;
assign w29741 = ~w29736 & w29740;
assign w29742 = pi1589 & ~w29741;
assign w29743 = ~pi1589 & w29741;
assign w29744 = ~w29742 & ~w29743;
assign w29745 = ~w29442 & ~w29450;
assign w29746 = ~w29468 & ~w29745;
assign w29747 = w29421 & ~w29454;
assign w29748 = ~w29746 & w29747;
assign w29749 = w29427 & ~w29450;
assign w29750 = w29442 & ~w29749;
assign w29751 = ~w29434 & ~w29750;
assign w29752 = w29748 & w29751;
assign w29753 = ~w29457 & ~w29464;
assign w29754 = (~w29464 & w29456) | (~w29464 & w65852) | (w29456 & w65852);
assign w29755 = ~w29753 & ~w29754;
assign w29756 = ~w29466 & w29755;
assign w29757 = ~w29436 & ~w29442;
assign w29758 = ~w29483 & ~w29757;
assign w29759 = ~w29757 & w65853;
assign w29760 = ~w29748 & ~w29759;
assign w29761 = ~w29491 & w29749;
assign w29762 = ~w29756 & w65854;
assign w29763 = ~w29450 & w29491;
assign w29764 = w29760 & w29763;
assign w29765 = ~w29456 & w29478;
assign w29766 = ~w29479 & w29765;
assign w29767 = w29464 & ~w29472;
assign w29768 = ~w29766 & w29767;
assign w29769 = ~w29764 & w29768;
assign w29770 = ~w29762 & ~w29769;
assign w29771 = w29456 & w29478;
assign w29772 = ~w29442 & w29453;
assign w29773 = ~w29771 & ~w29772;
assign w29774 = w29450 & ~w29773;
assign w29775 = w29492 & w29774;
assign w29776 = w29471 & w29478;
assign w29777 = ~w29752 & ~w29776;
assign w29778 = ~w29775 & w29777;
assign w29779 = ~w29770 & w29778;
assign w29780 = pi1578 & ~w29779;
assign w29781 = ~pi1578 & w29779;
assign w29782 = ~w29780 & ~w29781;
assign w29783 = w28857 & w28900;
assign w29784 = ~w28897 & w29393;
assign w29785 = w28873 & w28901;
assign w29786 = ~w29784 & ~w29785;
assign w29787 = ~w28849 & ~w29786;
assign w29788 = ~w28901 & ~w29391;
assign w29789 = w28857 & ~w29788;
assign w29790 = ~w28883 & ~w29785;
assign w29791 = ~w28900 & ~w29407;
assign w29792 = w28856 & ~w28870;
assign w29793 = w29790 & ~w29792;
assign w29794 = w29791 & w29793;
assign w29795 = ~w29789 & w29794;
assign w29796 = ~w28875 & ~w28886;
assign w29797 = ~w28897 & ~w29796;
assign w29798 = w28874 & w28902;
assign w29799 = ~w28917 & w65855;
assign w29800 = ~w29798 & w29799;
assign w29801 = ~w29797 & w29800;
assign w29802 = ~w29795 & ~w29801;
assign w29803 = ~w28912 & ~w29783;
assign w29804 = ~w29787 & w29803;
assign w29805 = ~w29802 & w29804;
assign w29806 = pi1596 & w29805;
assign w29807 = ~pi1596 & ~w29805;
assign w29808 = ~w29806 & ~w29807;
assign w29809 = w29595 & w29601;
assign w29810 = ~w29588 & ~w29643;
assign w29811 = ~w29642 & ~w29654;
assign w29812 = w29810 & ~w29811;
assign w29813 = ~w29654 & ~w29810;
assign w29814 = ~w29594 & ~w29813;
assign w29815 = ~w29812 & w29814;
assign w29816 = ~w29601 & w29628;
assign w29817 = w29675 & w29816;
assign w29818 = ~w29675 & w29685;
assign w29819 = ~w29689 & ~w29809;
assign w29820 = ~w29817 & w29819;
assign w29821 = ~w29818 & w29820;
assign w29822 = ~w29815 & w29821;
assign w29823 = ~pi1586 & ~w29822;
assign w29824 = pi1586 & w29822;
assign w29825 = ~w29823 & ~w29824;
assign w29826 = w28764 & w28793;
assign w29827 = ~w28770 & w28803;
assign w29828 = w28770 & ~w28803;
assign w29829 = (w29828 & ~w29205) | (w29828 & w65856) | (~w29205 & w65856);
assign w29830 = w29205 & ~w29828;
assign w29831 = ~w29211 & w29830;
assign w29832 = ~w29826 & ~w29827;
assign w29833 = (w29832 & w29831) | (w29832 & w65857) | (w29831 & w65857);
assign w29834 = ~w28783 & w29212;
assign w29835 = w29205 & w29827;
assign w29836 = ~w29834 & w29835;
assign w29837 = ~w29833 & ~w29836;
assign w29838 = pi1595 & w29837;
assign w29839 = ~pi1595 & ~w29837;
assign w29840 = ~w29838 & ~w29839;
assign w29841 = w28944 & w28981;
assign w29842 = ~w28993 & w29841;
assign w29843 = w28944 & ~w28981;
assign w29844 = ~w28967 & ~w29843;
assign w29845 = (~w28991 & ~w29844) | (~w28991 & w65858) | (~w29844 & w65858);
assign w29846 = ~w28938 & ~w28951;
assign w29847 = w28957 & w29846;
assign w29848 = ~w28969 & ~w29847;
assign w29849 = ~w28972 & w29848;
assign w29850 = w29848 & w65859;
assign w29851 = ~w28951 & w29850;
assign w29852 = w28957 & ~w29846;
assign w29853 = ~w29009 & ~w29852;
assign w29854 = ~w28984 & ~w29853;
assign w29855 = ~w29842 & w29845;
assign w29856 = ~w29854 & w29855;
assign w29857 = ~w29851 & w29856;
assign w29858 = w28981 & ~w29846;
assign w29859 = ~w28951 & w28981;
assign w29860 = w28967 & w29859;
assign w29861 = ~w28963 & ~w29018;
assign w29862 = ~w29860 & w29861;
assign w29863 = ~w28992 & w29858;
assign w29864 = w29862 & w29863;
assign w29865 = (w28992 & w29010) | (w28992 & w65860) | (w29010 & w65860);
assign w29866 = ~w29846 & ~w29865;
assign w29867 = w29843 & ~w29866;
assign w29868 = ~w28971 & w65861;
assign w29869 = ~w29864 & w29868;
assign w29870 = ~w29867 & w29869;
assign w29871 = ~w28938 & ~w28958;
assign w29872 = ~w28983 & w29871;
assign w29873 = ~w29844 & w29872;
assign w29874 = (~w29873 & w29870) | (~w29873 & w65862) | (w29870 & w65862);
assign w29875 = pi1590 & w29874;
assign w29876 = ~pi1590 & ~w29874;
assign w29877 = ~w29875 & ~w29876;
assign w29878 = w29249 & w29262;
assign w29879 = ~w29249 & ~w29295;
assign w29880 = w29520 & w29879;
assign w29881 = ~w29291 & ~w29878;
assign w29882 = (w29282 & ~w29881) | (w29282 & w65863) | (~w29881 & w65863);
assign w29883 = ~w29272 & ~w29296;
assign w29884 = w29236 & ~w29883;
assign w29885 = ~w29519 & ~w29884;
assign w29886 = ~w29282 & ~w29885;
assign w29887 = ~w29248 & ~w29262;
assign w29888 = ~w29263 & w29887;
assign w29889 = ~w29305 & ~w29888;
assign w29890 = w29313 & ~w29889;
assign w29891 = w29264 & ~w29298;
assign w29892 = ~w29282 & ~w29891;
assign w29893 = w29308 & ~w29892;
assign w29894 = ~w29236 & w29883;
assign w29895 = ~w29893 & w29894;
assign w29896 = ~w29882 & ~w29890;
assign w29897 = ~w29895 & w29896;
assign w29898 = ~w29886 & w29897;
assign w29899 = pi1585 & ~w29898;
assign w29900 = ~pi1585 & w29898;
assign w29901 = ~w29899 & ~w29900;
assign w29902 = w29514 & w29888;
assign w29903 = ~w29292 & ~w29311;
assign w29904 = ~w29261 & ~w29903;
assign w29905 = w29308 & w29520;
assign w29906 = (w29261 & w29905) | (w29261 & w65864) | (w29905 & w65864);
assign w29907 = ~w29904 & ~w29906;
assign w29908 = ~w29504 & w29907;
assign w29909 = w29282 & ~w29908;
assign w29910 = w29517 & w29522;
assign w29911 = w29276 & ~w29903;
assign w29912 = w29248 & w29298;
assign w29913 = w29524 & ~w29887;
assign w29914 = ~w29912 & w29913;
assign w29915 = ~w29902 & ~w29914;
assign w29916 = ~w29910 & w29915;
assign w29917 = ~w29911 & w29916;
assign w29918 = ~w29909 & w29917;
assign w29919 = pi1592 & ~w29918;
assign w29920 = ~pi1592 & w29918;
assign w29921 = ~w29919 & ~w29920;
assign w29922 = w28992 & w29859;
assign w29923 = ~w28944 & w28993;
assign w29924 = ~w28996 & ~w29923;
assign w29925 = ~w28981 & ~w29924;
assign w29926 = w28997 & ~w29848;
assign w29927 = ~w28938 & w28961;
assign w29928 = ~w29006 & ~w29927;
assign w29929 = w28995 & w29928;
assign w29930 = ~w29926 & w29929;
assign w29931 = ~w29925 & w29930;
assign w29932 = w28960 & ~w29844;
assign w29933 = w28981 & ~w29847;
assign w29934 = w28965 & w29933;
assign w29935 = w29845 & ~w29932;
assign w29936 = ~w29934 & w29935;
assign w29937 = ~w29931 & ~w29936;
assign w29938 = w28966 & ~w28981;
assign w29939 = ~w29019 & ~w29922;
assign w29940 = ~w29938 & w29939;
assign w29941 = ~w29937 & w29940;
assign w29942 = ~pi1606 & ~w29941;
assign w29943 = pi1606 & w29941;
assign w29944 = ~w29942 & ~w29943;
assign w29945 = w28770 & ~w28811;
assign w29946 = w28804 & w28835;
assign w29947 = w28794 & ~w29946;
assign w29948 = ~w29945 & ~w29947;
assign w29949 = ~w28763 & w29204;
assign w29950 = w28785 & w28825;
assign w29951 = w28814 & ~w29950;
assign w29952 = ~w29218 & w29951;
assign w29953 = w28764 & ~w28835;
assign w29954 = w28770 & ~w28822;
assign w29955 = ~w29953 & w29954;
assign w29956 = ~w29952 & ~w29955;
assign w29957 = w28803 & ~w29949;
assign w29958 = ~w29956 & w29957;
assign w29959 = ~w28816 & w29951;
assign w29960 = ~w28763 & w28835;
assign w29961 = ~w28812 & ~w29960;
assign w29962 = ~w28815 & ~w29961;
assign w29963 = w28807 & ~w28831;
assign w29964 = ~w29962 & w29963;
assign w29965 = ~w29959 & w29964;
assign w29966 = (~w29948 & w29958) | (~w29948 & w65865) | (w29958 & w65865);
assign w29967 = ~pi1594 & w29966;
assign w29968 = pi1594 & ~w29966;
assign w29969 = ~w29967 & ~w29968;
assign w29970 = w28897 & ~w28903;
assign w29971 = w28874 & ~w29970;
assign w29972 = ~w28877 & w29971;
assign w29973 = ~w29791 & w29972;
assign w29974 = ~w28849 & w28874;
assign w29975 = w29970 & w29974;
assign w29976 = ~w28877 & w29796;
assign w29977 = w28849 & ~w29976;
assign w29978 = w29400 & ~w29975;
assign w29979 = ~w29977 & w29978;
assign w29980 = w28885 & w28916;
assign w29981 = ~w28899 & ~w28925;
assign w29982 = w29790 & ~w29980;
assign w29983 = w29981 & w29982;
assign w29984 = ~w29972 & w29983;
assign w29985 = (~w29973 & w29979) | (~w29973 & w65866) | (w29979 & w65866);
assign w29986 = ~pi1574 & w29985;
assign w29987 = pi1574 & ~w29985;
assign w29988 = ~w29986 & ~w29987;
assign w29989 = w29478 & w29483;
assign w29990 = ~w29458 & ~w29989;
assign w29991 = ~w29747 & w29753;
assign w29992 = w29773 & w29991;
assign w29993 = w29990 & ~w29992;
assign w29994 = ~w29450 & ~w29993;
assign w29995 = w29481 & ~w29492;
assign w29996 = w29428 & ~w29442;
assign w29997 = w29421 & w29468;
assign w29998 = w29450 & ~w29996;
assign w29999 = ~w29997 & w29998;
assign w30000 = ~w29995 & ~w29999;
assign w30001 = w29435 & w29442;
assign w30002 = w29464 & ~w29748;
assign w30003 = w29990 & ~w30001;
assign w30004 = w30002 & w30003;
assign w30005 = ~w30000 & w30004;
assign w30006 = w29436 & w29746;
assign w30007 = ~w29755 & ~w30006;
assign w30008 = ~w29774 & w30007;
assign w30009 = ~w30005 & ~w30008;
assign w30010 = ~w29994 & ~w30009;
assign w30011 = ~pi1579 & w30010;
assign w30012 = pi1579 & ~w30010;
assign w30013 = ~w30011 & ~w30012;
assign w30014 = ~w29107 & ~w29544;
assign w30015 = ~w29097 & ~w29708;
assign w30016 = ~w30014 & w30015;
assign w30017 = ~w29547 & ~w30016;
assign w30018 = w29711 & ~w30017;
assign w30019 = ~w29553 & ~w30016;
assign w30020 = ~w29095 & ~w30019;
assign w30021 = ~w29055 & ~w29537;
assign w30022 = ~w29702 & w30021;
assign w30023 = ~w29062 & ~w30022;
assign w30024 = ~w29053 & ~w29054;
assign w30025 = w29062 & ~w29708;
assign w30026 = ~w30024 & w30025;
assign w30027 = ~w29097 & ~w29102;
assign w30028 = ~w29554 & w30027;
assign w30029 = (w29095 & ~w30028) | (w29095 & w65867) | (~w30028 & w65867);
assign w30030 = ~w30023 & ~w30029;
assign w30031 = ~w30018 & w30030;
assign w30032 = ~w30020 & w30031;
assign w30033 = pi1601 & ~w30032;
assign w30034 = ~pi1601 & w30032;
assign w30035 = ~w30033 & ~w30034;
assign w30036 = ~w28963 & ~w29850;
assign w30037 = ~w28981 & ~w30036;
assign w30038 = w28981 & ~w29849;
assign w30039 = w29005 & ~w29858;
assign w30040 = ~w30038 & ~w30039;
assign w30041 = ~w28991 & ~w30040;
assign w30042 = (w28991 & ~w29862) | (w28991 & w65868) | (~w29862 & w65868);
assign w30043 = ~w28973 & ~w28994;
assign w30044 = w28981 & ~w30043;
assign w30045 = ~w30042 & ~w30044;
assign w30046 = ~w30037 & w30045;
assign w30047 = ~w30041 & w30046;
assign w30048 = pi1619 & ~w30047;
assign w30049 = ~pi1619 & w30047;
assign w30050 = ~w30048 & ~w30049;
assign w30051 = ~w29454 & w29751;
assign w30052 = ~w29466 & ~w29753;
assign w30053 = ~w29485 & ~w29996;
assign w30054 = ~w30051 & w30053;
assign w30055 = ~w30052 & w30054;
assign w30056 = ~w29492 & ~w29765;
assign w30057 = ~w29484 & ~w30056;
assign w30058 = w29450 & w29758;
assign w30059 = w29464 & ~w30057;
assign w30060 = ~w30058 & w30059;
assign w30061 = ~w30055 & ~w30060;
assign w30062 = w29421 & w29457;
assign w30063 = ~w30001 & ~w30062;
assign w30064 = w29450 & ~w30063;
assign w30065 = w29443 & ~w29450;
assign w30066 = ~w30064 & ~w30065;
assign w30067 = ~w30061 & w30066;
assign w30068 = ~pi1602 & w30067;
assign w30069 = pi1602 & ~w30067;
assign w30070 = ~w30068 & ~w30069;
assign w30071 = ~pi5514 & pi9040;
assign w30072 = ~pi5317 & ~pi9040;
assign w30073 = ~w30071 & ~w30072;
assign w30074 = pi1621 & ~w30073;
assign w30075 = ~pi1621 & w30073;
assign w30076 = ~w30074 & ~w30075;
assign w30077 = ~pi5400 & pi9040;
assign w30078 = ~pi5401 & ~pi9040;
assign w30079 = ~w30077 & ~w30078;
assign w30080 = pi1624 & ~w30079;
assign w30081 = ~pi1624 & w30079;
assign w30082 = ~w30080 & ~w30081;
assign w30083 = ~pi5513 & pi9040;
assign w30084 = ~pi5407 & ~pi9040;
assign w30085 = ~w30083 & ~w30084;
assign w30086 = pi1612 & ~w30085;
assign w30087 = ~pi1612 & w30085;
assign w30088 = ~w30086 & ~w30087;
assign w30089 = ~pi5509 & pi9040;
assign w30090 = ~pi5443 & ~pi9040;
assign w30091 = ~w30089 & ~w30090;
assign w30092 = pi1593 & ~w30091;
assign w30093 = ~pi1593 & w30091;
assign w30094 = ~w30092 & ~w30093;
assign w30095 = ~w30088 & ~w30094;
assign w30096 = w30088 & w30094;
assign w30097 = w30076 & w30096;
assign w30098 = ~w30095 & ~w30097;
assign w30099 = ~pi5396 & pi9040;
assign w30100 = ~pi5510 & ~pi9040;
assign w30101 = ~w30099 & ~w30100;
assign w30102 = pi1598 & ~w30101;
assign w30103 = ~pi1598 & w30101;
assign w30104 = ~w30102 & ~w30103;
assign w30105 = w30076 & ~w30104;
assign w30106 = ~w30076 & w30104;
assign w30107 = ~w30105 & ~w30106;
assign w30108 = ~w30082 & w30107;
assign w30109 = ~w30098 & w30108;
assign w30110 = ~w30076 & w30109;
assign w30111 = w30088 & w30104;
assign w30112 = w30094 & w30111;
assign w30113 = w30095 & w30105;
assign w30114 = ~w30112 & ~w30113;
assign w30115 = w30082 & ~w30114;
assign w30116 = ~w30094 & ~w30104;
assign w30117 = ~w30082 & w30088;
assign w30118 = w30116 & w30117;
assign w30119 = w30096 & w30106;
assign w30120 = ~w30118 & ~w30119;
assign w30121 = ~pi5570 & pi9040;
assign w30122 = ~pi5402 & ~pi9040;
assign w30123 = ~w30121 & ~w30122;
assign w30124 = pi1611 & ~w30123;
assign w30125 = ~pi1611 & w30123;
assign w30126 = ~w30124 & ~w30125;
assign w30127 = w30088 & w30105;
assign w30128 = ~w30088 & ~w30104;
assign w30129 = ~w30106 & ~w30128;
assign w30130 = (~w30082 & ~w30129) | (~w30082 & w30117) | (~w30129 & w30117);
assign w30131 = ~w30127 & w30130;
assign w30132 = ~w30076 & w30094;
assign w30133 = ~w30088 & w30132;
assign w30134 = w30082 & ~w30128;
assign w30135 = ~w30133 & w30134;
assign w30136 = ~w30131 & ~w30135;
assign w30137 = w30082 & w30106;
assign w30138 = ~w30094 & w30105;
assign w30139 = ~w30137 & ~w30138;
assign w30140 = w30088 & ~w30139;
assign w30141 = w30120 & ~w30126;
assign w30142 = ~w30140 & w30141;
assign w30143 = ~w30136 & w30142;
assign w30144 = w30094 & w30104;
assign w30145 = ~w30076 & w30088;
assign w30146 = ~w30144 & ~w30145;
assign w30147 = ~w30076 & ~w30116;
assign w30148 = w30146 & w30147;
assign w30149 = w30120 & ~w30148;
assign w30150 = w30136 & ~w30149;
assign w30151 = ~w30082 & ~w30104;
assign w30152 = ~w30127 & ~w30133;
assign w30153 = (w30151 & ~w30152) | (w30151 & w65869) | (~w30152 & w65869);
assign w30154 = ~w30112 & w30130;
assign w30155 = w30076 & ~w30094;
assign w30156 = ~w30132 & ~w30155;
assign w30157 = w30088 & ~w30156;
assign w30158 = w30082 & w30129;
assign w30159 = ~w30157 & w30158;
assign w30160 = ~w30154 & ~w30159;
assign w30161 = ~w30153 & ~w30160;
assign w30162 = (w30126 & ~w30136) | (w30126 & w63853) | (~w30136 & w63853);
assign w30163 = ~w30161 & w30162;
assign w30164 = ~w30110 & ~w30115;
assign w30165 = (w30164 & w30163) | (w30164 & w65870) | (w30163 & w65870);
assign w30166 = pi1656 & w30165;
assign w30167 = ~pi1656 & ~w30165;
assign w30168 = ~w30166 & ~w30167;
assign w30169 = w30129 & w65871;
assign w30170 = ~w30111 & ~w30128;
assign w30171 = w30076 & ~w30096;
assign w30172 = ~w30170 & w30171;
assign w30173 = ~w30169 & ~w30172;
assign w30174 = w30082 & ~w30173;
assign w30175 = ~w30109 & w30149;
assign w30176 = ~w30174 & w30175;
assign w30177 = w30126 & ~w30176;
assign w30178 = w30096 & w30151;
assign w30179 = ~w30172 & ~w30178;
assign w30180 = ~w30082 & ~w30126;
assign w30181 = ~w30179 & w30180;
assign w30182 = w30094 & ~w30151;
assign w30183 = w30105 & w30182;
assign w30184 = w30116 & w30145;
assign w30185 = (~w30088 & ~w30107) | (~w30088 & w65871) | (~w30107 & w65871);
assign w30186 = w30082 & ~w30126;
assign w30187 = ~w30185 & w30186;
assign w30188 = w30104 & ~w30126;
assign w30189 = w30132 & w30188;
assign w30190 = ~w30187 & ~w30189;
assign w30191 = ~w30157 & ~w30190;
assign w30192 = ~w30183 & ~w30184;
assign w30193 = ~w30181 & w30192;
assign w30194 = ~w30191 & w30193;
assign w30195 = ~w30177 & w30194;
assign w30196 = ~pi1646 & w30195;
assign w30197 = pi1646 & ~w30195;
assign w30198 = ~w30196 & ~w30197;
assign w30199 = ~pi5316 & pi9040;
assign w30200 = ~pi5400 & ~pi9040;
assign w30201 = ~w30199 & ~w30200;
assign w30202 = pi1600 & ~w30201;
assign w30203 = ~pi1600 & w30201;
assign w30204 = ~w30202 & ~w30203;
assign w30205 = ~pi5510 & pi9040;
assign w30206 = ~pi5320 & ~pi9040;
assign w30207 = ~w30205 & ~w30206;
assign w30208 = pi1617 & ~w30207;
assign w30209 = ~pi1617 & w30207;
assign w30210 = ~w30208 & ~w30209;
assign w30211 = w30204 & ~w30210;
assign w30212 = ~w30204 & w30210;
assign w30213 = ~w30211 & ~w30212;
assign w30214 = ~pi5438 & pi9040;
assign w30215 = ~pi5511 & ~pi9040;
assign w30216 = ~w30214 & ~w30215;
assign w30217 = pi1608 & ~w30216;
assign w30218 = ~pi1608 & w30216;
assign w30219 = ~w30217 & ~w30218;
assign w30220 = ~pi5402 & pi9040;
assign w30221 = ~pi5392 & ~pi9040;
assign w30222 = ~w30220 & ~w30221;
assign w30223 = pi1620 & ~w30222;
assign w30224 = ~pi1620 & w30222;
assign w30225 = ~w30223 & ~w30224;
assign w30226 = ~w30219 & ~w30225;
assign w30227 = w30213 & w30226;
assign w30228 = w30212 & w30219;
assign w30229 = ~w30227 & ~w30228;
assign w30230 = w30210 & ~w30219;
assign w30231 = ~w30204 & w30219;
assign w30232 = w30225 & w30231;
assign w30233 = ~w30230 & ~w30232;
assign w30234 = ~w30229 & w30233;
assign w30235 = ~w30219 & w30225;
assign w30236 = ~w30213 & w30235;
assign w30237 = (~w30236 & w30229) | (~w30236 & w65872) | (w30229 & w65872);
assign w30238 = ~pi5441 & pi9040;
assign w30239 = ~pi5435 & ~pi9040;
assign w30240 = ~w30238 & ~w30239;
assign w30241 = pi1603 & ~w30240;
assign w30242 = ~pi1603 & w30240;
assign w30243 = ~w30241 & ~w30242;
assign w30244 = ~w30237 & w30243;
assign w30245 = w30219 & ~w30225;
assign w30246 = w30204 & w30245;
assign w30247 = ~w30219 & w30243;
assign w30248 = ~w30210 & ~w30225;
assign w30249 = w30243 & ~w30248;
assign w30250 = ~w30247 & ~w30249;
assign w30251 = ~w30249 & w65873;
assign w30252 = ~w30204 & w30243;
assign w30253 = w30210 & w30225;
assign w30254 = ~w30219 & ~w30252;
assign w30255 = w30253 & w30254;
assign w30256 = ~w30251 & ~w30255;
assign w30257 = ~w30230 & ~w30245;
assign w30258 = w30204 & w30243;
assign w30259 = ~w30257 & w30258;
assign w30260 = ~w30248 & w30252;
assign w30261 = ~w30247 & ~w30260;
assign w30262 = ~w30213 & w30225;
assign w30263 = w30261 & w30262;
assign w30264 = w30229 & ~w30259;
assign w30265 = ~w30263 & w30264;
assign w30266 = w30264 & w65874;
assign w30267 = w30265 & w63854;
assign w30268 = ~w30219 & ~w30243;
assign w30269 = w30213 & w30268;
assign w30270 = ~w30211 & ~w30245;
assign w30271 = ~w30249 & w63855;
assign w30272 = ~w30270 & ~w30271;
assign w30273 = ~pi5407 & pi9040;
assign w30274 = ~pi5308 & ~pi9040;
assign w30275 = ~w30273 & ~w30274;
assign w30276 = pi1628 & ~w30275;
assign w30277 = ~pi1628 & w30275;
assign w30278 = ~w30276 & ~w30277;
assign w30279 = w30231 & w30253;
assign w30280 = w30278 & ~w30279;
assign w30281 = ~w30269 & w30280;
assign w30282 = ~w30272 & w30281;
assign w30283 = ~w30259 & w30261;
assign w30284 = ~w30212 & ~w30225;
assign w30285 = ~w30235 & ~w30284;
assign w30286 = w30283 & w30285;
assign w30287 = ~w30272 & w30286;
assign w30288 = (~w30251 & ~w30286) | (~w30251 & w63856) | (~w30286 & w63856);
assign w30289 = w30226 & w30252;
assign w30290 = ~w30255 & ~w30289;
assign w30291 = ~w30211 & w30247;
assign w30292 = ~w30255 & w65875;
assign w30293 = ~w30278 & ~w30292;
assign w30294 = (~w30282 & ~w30288) | (~w30282 & w65876) | (~w30288 & w65876);
assign w30295 = ~w30244 & ~w30267;
assign w30296 = w30295 & w65877;
assign w30297 = (pi1635 & ~w30295) | (pi1635 & w65878) | (~w30295 & w65878);
assign w30298 = ~w30296 & ~w30297;
assign w30299 = ~pi5436 & pi9040;
assign w30300 = ~pi5303 & ~pi9040;
assign w30301 = ~w30299 & ~w30300;
assign w30302 = pi1591 & ~w30301;
assign w30303 = ~pi1591 & w30301;
assign w30304 = ~w30302 & ~w30303;
assign w30305 = ~pi5322 & pi9040;
assign w30306 = ~pi5502 & ~pi9040;
assign w30307 = ~w30305 & ~w30306;
assign w30308 = pi1629 & ~w30307;
assign w30309 = ~pi1629 & w30307;
assign w30310 = ~w30308 & ~w30309;
assign w30311 = ~w30304 & w30310;
assign w30312 = ~pi5325 & pi9040;
assign w30313 = ~pi5505 & ~pi9040;
assign w30314 = ~w30312 & ~w30313;
assign w30315 = pi1628 & ~w30314;
assign w30316 = ~pi1628 & w30314;
assign w30317 = ~w30315 & ~w30316;
assign w30318 = ~pi5566 & pi9040;
assign w30319 = ~pi5299 & ~pi9040;
assign w30320 = ~w30318 & ~w30319;
assign w30321 = pi1607 & ~w30320;
assign w30322 = ~pi1607 & w30320;
assign w30323 = ~w30321 & ~w30322;
assign w30324 = ~w30304 & ~w30323;
assign w30325 = ~pi5437 & pi9040;
assign w30326 = ~pi5408 & ~pi9040;
assign w30327 = ~w30325 & ~w30326;
assign w30328 = pi1620 & ~w30327;
assign w30329 = ~pi1620 & w30327;
assign w30330 = ~w30328 & ~w30329;
assign w30331 = ~w30317 & ~w30330;
assign w30332 = ~w30324 & w30331;
assign w30333 = w30311 & w30332;
assign w30334 = w30304 & w30317;
assign w30335 = ~w30304 & ~w30317;
assign w30336 = ~w30334 & ~w30335;
assign w30337 = ~w30330 & ~w30336;
assign w30338 = ~w30336 & w65879;
assign w30339 = ~w30304 & w30330;
assign w30340 = ~w30323 & ~w30339;
assign w30341 = w30304 & ~w30330;
assign w30342 = w30323 & ~w30334;
assign w30343 = ~w30341 & w30342;
assign w30344 = ~w30310 & ~w30340;
assign w30345 = ~w30343 & w30344;
assign w30346 = ~w30338 & w30345;
assign w30347 = ~pi5310 & pi9040;
assign w30348 = ~pi5304 & ~pi9040;
assign w30349 = ~w30347 & ~w30348;
assign w30350 = pi1622 & ~w30349;
assign w30351 = ~pi1622 & w30349;
assign w30352 = ~w30350 & ~w30351;
assign w30353 = w30317 & w30330;
assign w30354 = ~w30310 & w30353;
assign w30355 = ~w30332 & ~w30354;
assign w30356 = w30310 & ~w30353;
assign w30357 = w30340 & w30356;
assign w30358 = ~w30323 & ~w30330;
assign w30359 = ~w30304 & w30358;
assign w30360 = (w30336 & w30357) | (w30336 & w65880) | (w30357 & w65880);
assign w30361 = ~w30339 & ~w30341;
assign w30362 = w30324 & w30353;
assign w30363 = w30310 & ~w30361;
assign w30364 = ~w30362 & w30363;
assign w30365 = ~w30338 & ~w30364;
assign w30366 = ~w30324 & w30356;
assign w30367 = (w30366 & w30364) | (w30366 & w65881) | (w30364 & w65881);
assign w30368 = w30355 & ~w30360;
assign w30369 = ~w30367 & w30368;
assign w30370 = w30352 & ~w30369;
assign w30371 = w30310 & w30317;
assign w30372 = w30358 & w30371;
assign w30373 = w30361 & ~w30371;
assign w30374 = ~w30323 & ~w30336;
assign w30375 = ~w30373 & w30374;
assign w30376 = w30330 & w30336;
assign w30377 = w30336 & w30485;
assign w30378 = w30323 & w30377;
assign w30379 = w30317 & ~w30323;
assign w30380 = ~w30310 & ~w30334;
assign w30381 = w30323 & w30330;
assign w30382 = ~w30379 & ~w30381;
assign w30383 = w30380 & w30382;
assign w30384 = w30355 & w30383;
assign w30385 = ~w30375 & ~w30384;
assign w30386 = (~w30352 & ~w30385) | (~w30352 & w65882) | (~w30385 & w65882);
assign w30387 = ~w30333 & ~w30372;
assign w30388 = ~w30346 & w30387;
assign w30389 = ~w30386 & w30388;
assign w30390 = ~w30370 & w30389;
assign w30391 = pi1634 & ~w30390;
assign w30392 = ~pi1634 & w30390;
assign w30393 = ~w30391 & ~w30392;
assign w30394 = ~pi5317 & pi9040;
assign w30395 = ~pi5434 & ~pi9040;
assign w30396 = ~w30394 & ~w30395;
assign w30397 = pi1599 & ~w30396;
assign w30398 = ~pi1599 & w30396;
assign w30399 = ~w30397 & ~w30398;
assign w30400 = ~pi5401 & pi9040;
assign w30401 = ~pi5442 & ~pi9040;
assign w30402 = ~w30400 & ~w30401;
assign w30403 = pi1611 & ~w30402;
assign w30404 = ~pi1611 & w30402;
assign w30405 = ~w30403 & ~w30404;
assign w30406 = w30399 & ~w30405;
assign w30407 = ~pi5320 & pi9040;
assign w30408 = ~pi5509 & ~pi9040;
assign w30409 = ~w30407 & ~w30408;
assign w30410 = pi1593 & ~w30409;
assign w30411 = ~pi1593 & w30409;
assign w30412 = ~w30410 & ~w30411;
assign w30413 = ~pi5309 & pi9040;
assign w30414 = ~pi5415 & ~pi9040;
assign w30415 = ~w30413 & ~w30414;
assign w30416 = pi1608 & ~w30415;
assign w30417 = ~pi1608 & w30415;
assign w30418 = ~w30416 & ~w30417;
assign w30419 = w30412 & w30418;
assign w30420 = w30406 & ~w30419;
assign w30421 = ~w30412 & ~w30418;
assign w30422 = ~w30420 & ~w30421;
assign w30423 = w30406 & w30421;
assign w30424 = ~pi5308 & pi9040;
assign w30425 = ~pi5323 & ~pi9040;
assign w30426 = ~w30424 & ~w30425;
assign w30427 = pi1625 & ~w30426;
assign w30428 = ~pi1625 & w30426;
assign w30429 = ~w30427 & ~w30428;
assign w30430 = ~w30423 & w30429;
assign w30431 = ~w30422 & w30430;
assign w30432 = ~w30399 & ~w30412;
assign w30433 = ~w30405 & ~w30418;
assign w30434 = w30405 & w30418;
assign w30435 = ~w30433 & ~w30434;
assign w30436 = w30432 & w30435;
assign w30437 = w30405 & ~w30412;
assign w30438 = w30399 & w30418;
assign w30439 = w30437 & w30438;
assign w30440 = w30412 & w30433;
assign w30441 = ~w30429 & ~w30439;
assign w30442 = ~w30440 & w30441;
assign w30443 = ~w30436 & w30442;
assign w30444 = ~w30399 & w30405;
assign w30445 = ~w30412 & ~w30444;
assign w30446 = ~w30406 & ~w30438;
assign w30447 = w30445 & w30446;
assign w30448 = ~w30418 & ~w30447;
assign w30449 = w30443 & w30448;
assign w30450 = w30418 & ~w30429;
assign w30451 = ~w30412 & ~w30450;
assign w30452 = w30444 & w30451;
assign w30453 = ~w30406 & ~w30444;
assign w30454 = ~w30419 & ~w30450;
assign w30455 = w30453 & ~w30454;
assign w30456 = ~pi5565 & pi9040;
assign w30457 = ~pi5570 & ~pi9040;
assign w30458 = ~w30456 & ~w30457;
assign w30459 = pi1600 & ~w30458;
assign w30460 = ~pi1600 & w30458;
assign w30461 = ~w30459 & ~w30460;
assign w30462 = ~w30452 & ~w30461;
assign w30463 = ~w30455 & w30462;
assign w30464 = ~w30449 & w30463;
assign w30465 = ~w30399 & ~w30419;
assign w30466 = ~w30437 & ~w30444;
assign w30467 = w30429 & ~w30466;
assign w30468 = ~w30465 & w30467;
assign w30469 = w30418 & w30420;
assign w30470 = w30432 & w30433;
assign w30471 = w30405 & w30412;
assign w30472 = w30450 & ~w30471;
assign w30473 = ~w30445 & w30472;
assign w30474 = ~w30470 & ~w30473;
assign w30475 = w30461 & ~w30469;
assign w30476 = ~w30468 & w30475;
assign w30477 = w30474 & w30476;
assign w30478 = w30412 & ~w30429;
assign w30479 = w30453 & w30478;
assign w30480 = ~w30431 & ~w30479;
assign w30481 = (w30480 & w30464) | (w30480 & w65883) | (w30464 & w65883);
assign w30482 = pi1639 & ~w30481;
assign w30483 = ~pi1639 & w30481;
assign w30484 = ~w30482 & ~w30483;
assign w30485 = w30310 & w30330;
assign w30486 = ~w30369 & w30485;
assign w30487 = w30361 & w30371;
assign w30488 = ~w30341 & ~w30353;
assign w30489 = w30342 & ~w30488;
assign w30490 = (~w30310 & w30375) | (~w30310 & w65884) | (w30375 & w65884);
assign w30491 = ~w30352 & ~w30487;
assign w30492 = ~w30489 & w30491;
assign w30493 = ~w30490 & w30492;
assign w30494 = w30304 & w30381;
assign w30495 = w30352 & ~w30494;
assign w30496 = ~w30317 & ~w30358;
assign w30497 = ~w30310 & ~w30379;
assign w30498 = ~w30496 & w30497;
assign w30499 = w30334 & w30358;
assign w30500 = ~w30496 & ~w30499;
assign w30501 = w30310 & ~w30500;
assign w30502 = ~w30362 & w30495;
assign w30503 = ~w30498 & w30502;
assign w30504 = ~w30501 & w30503;
assign w30505 = ~w30493 & ~w30504;
assign w30506 = ~w30486 & ~w30505;
assign w30507 = ~pi1640 & w30506;
assign w30508 = pi1640 & ~w30506;
assign w30509 = ~w30507 & ~w30508;
assign w30510 = w30082 & ~w30152;
assign w30511 = ~w30138 & ~w30148;
assign w30512 = ~w30169 & w30511;
assign w30513 = ~w30510 & w30512;
assign w30514 = w30126 & ~w30513;
assign w30515 = w30117 & w30126;
assign w30516 = ~w30178 & ~w30515;
assign w30517 = ~w30076 & ~w30516;
assign w30518 = ~w30088 & w30156;
assign w30519 = w30180 & w30518;
assign w30520 = w30097 & w30188;
assign w30521 = w30152 & w30186;
assign w30522 = ~w30518 & w30521;
assign w30523 = ~w30517 & ~w30520;
assign w30524 = ~w30519 & w30523;
assign w30525 = ~w30522 & w30524;
assign w30526 = ~w30150 & w30525;
assign w30527 = (pi1660 & ~w30526) | (pi1660 & w65885) | (~w30526 & w65885);
assign w30528 = w30526 & w65886;
assign w30529 = ~w30527 & ~w30528;
assign w30530 = ~pi5392 & pi9040;
assign w30531 = ~pi5513 & ~pi9040;
assign w30532 = ~w30530 & ~w30531;
assign w30533 = pi1630 & ~w30532;
assign w30534 = ~pi1630 & w30532;
assign w30535 = ~w30533 & ~w30534;
assign w30536 = ~pi5415 & pi9040;
assign w30537 = ~pi5396 & ~pi9040;
assign w30538 = ~w30536 & ~w30537;
assign w30539 = pi1605 & ~w30538;
assign w30540 = ~pi1605 & w30538;
assign w30541 = ~w30539 & ~w30540;
assign w30542 = w30535 & ~w30541;
assign w30543 = ~pi5511 & pi9040;
assign w30544 = ~pi5514 & ~pi9040;
assign w30545 = ~w30543 & ~w30544;
assign w30546 = pi1627 & ~w30545;
assign w30547 = ~pi1627 & w30545;
assign w30548 = ~w30546 & ~w30547;
assign w30549 = ~w30541 & ~w30548;
assign w30550 = ~pi5443 & pi9040;
assign w30551 = ~pi5316 & ~pi9040;
assign w30552 = ~w30550 & ~w30551;
assign w30553 = pi1612 & ~w30552;
assign w30554 = ~pi1612 & w30552;
assign w30555 = ~w30553 & ~w30554;
assign w30556 = w30549 & ~w30555;
assign w30557 = ~w30542 & ~w30556;
assign w30558 = w30535 & ~w30548;
assign w30559 = ~pi5311 & pi9040;
assign w30560 = ~pi5441 & ~pi9040;
assign w30561 = ~w30559 & ~w30560;
assign w30562 = pi1623 & ~w30561;
assign w30563 = ~pi1623 & w30561;
assign w30564 = ~w30562 & ~w30563;
assign w30565 = ~w30558 & ~w30564;
assign w30566 = ~w30557 & w30565;
assign w30567 = ~pi5323 & pi9040;
assign w30568 = ~pi5318 & ~pi9040;
assign w30569 = ~w30567 & ~w30568;
assign w30570 = pi1621 & ~w30569;
assign w30571 = ~pi1621 & w30569;
assign w30572 = ~w30570 & ~w30571;
assign w30573 = ~w30541 & w30572;
assign w30574 = w30548 & ~w30572;
assign w30575 = w30535 & w30541;
assign w30576 = w30574 & w30575;
assign w30577 = ~w30541 & ~w30572;
assign w30578 = w30558 & w30577;
assign w30579 = ~w30576 & ~w30578;
assign w30580 = ~w30573 & w30579;
assign w30581 = w30548 & w30572;
assign w30582 = ~w30558 & ~w30581;
assign w30583 = w30541 & ~w30572;
assign w30584 = ~w30573 & ~w30583;
assign w30585 = ~w30582 & ~w30584;
assign w30586 = w30564 & ~w30585;
assign w30587 = ~w30580 & w30586;
assign w30588 = ~w30541 & ~w30564;
assign w30589 = w30581 & w30588;
assign w30590 = ~w30535 & w30541;
assign w30591 = ~w30548 & ~w30564;
assign w30592 = ~w30572 & ~w30591;
assign w30593 = w30590 & ~w30592;
assign w30594 = ~w30558 & ~w30577;
assign w30595 = ~w30535 & w30548;
assign w30596 = ~w30583 & ~w30595;
assign w30597 = ~w30594 & ~w30596;
assign w30598 = w30541 & w30572;
assign w30599 = w30548 & w30598;
assign w30600 = ~w30549 & ~w30599;
assign w30601 = ~w30597 & w30600;
assign w30602 = w30564 & ~w30601;
assign w30603 = w30555 & ~w30576;
assign w30604 = ~w30589 & w30603;
assign w30605 = ~w30593 & w30604;
assign w30606 = ~w30602 & w30605;
assign w30607 = w30564 & ~w30598;
assign w30608 = w30590 & w30607;
assign w30609 = ~w30549 & ~w30594;
assign w30610 = ~w30607 & w30609;
assign w30611 = ~w30555 & ~w30608;
assign w30612 = ~w30610 & w30611;
assign w30613 = ~w30606 & ~w30612;
assign w30614 = w30581 & w30590;
assign w30615 = ~w30566 & ~w30614;
assign w30616 = ~w30587 & w30615;
assign w30617 = ~w30613 & w30616;
assign w30618 = ~pi1637 & w30617;
assign w30619 = pi1637 & ~w30617;
assign w30620 = ~w30618 & ~w30619;
assign w30621 = w30354 & ~w30495;
assign w30622 = ~w30337 & ~w30376;
assign w30623 = w30380 & w30622;
assign w30624 = ~w30333 & ~w30499;
assign w30625 = (~w30623 & w65887) | (~w30623 & w65888) | (w65887 & w65888);
assign w30626 = w30352 & ~w30625;
assign w30627 = w30335 & w30485;
assign w30628 = w30323 & ~w30380;
assign w30629 = ~w30311 & ~w30371;
assign w30630 = w30628 & w30629;
assign w30631 = ~w30359 & ~w30494;
assign w30632 = ~w30627 & w30631;
assign w30633 = ~w30630 & w30632;
assign w30634 = ~w30352 & ~w30633;
assign w30635 = w30380 & ~w30488;
assign w30636 = ~w30627 & ~w30635;
assign w30637 = ~w30323 & ~w30636;
assign w30638 = ~w30372 & ~w30621;
assign w30639 = ~w30637 & w30638;
assign w30640 = ~w30634 & w30639;
assign w30641 = ~w30626 & w30640;
assign w30642 = pi1644 & ~w30641;
assign w30643 = ~pi1644 & w30641;
assign w30644 = ~w30642 & ~w30643;
assign w30645 = ~pi5505 & pi9040;
assign w30646 = ~pi5399 & ~pi9040;
assign w30647 = ~w30645 & ~w30646;
assign w30648 = pi1627 & ~w30647;
assign w30649 = ~pi1627 & w30647;
assign w30650 = ~w30648 & ~w30649;
assign w30651 = ~pi5576 & pi9040;
assign w30652 = ~pi5398 & ~pi9040;
assign w30653 = ~w30651 & ~w30652;
assign w30654 = pi1609 & ~w30653;
assign w30655 = ~pi1609 & w30653;
assign w30656 = ~w30654 & ~w30655;
assign w30657 = ~pi5305 & pi9040;
assign w30658 = ~pi5313 & ~pi9040;
assign w30659 = ~w30657 & ~w30658;
assign w30660 = pi1631 & ~w30659;
assign w30661 = ~pi1631 & w30659;
assign w30662 = ~w30660 & ~w30661;
assign w30663 = w30656 & w30662;
assign w30664 = ~pi5408 & pi9040;
assign w30665 = ~pi5665 & ~pi9040;
assign w30666 = ~w30664 & ~w30665;
assign w30667 = pi1614 & ~w30666;
assign w30668 = ~pi1614 & w30666;
assign w30669 = ~w30667 & ~w30668;
assign w30670 = ~pi5403 & pi9040;
assign w30671 = ~pi5310 & ~pi9040;
assign w30672 = ~w30670 & ~w30671;
assign w30673 = pi1605 & ~w30672;
assign w30674 = ~pi1605 & w30672;
assign w30675 = ~w30673 & ~w30674;
assign w30676 = ~w30669 & w30675;
assign w30677 = ~pi5306 & pi9040;
assign w30678 = ~pi5328 & ~pi9040;
assign w30679 = ~w30677 & ~w30678;
assign w30680 = pi1615 & ~w30679;
assign w30681 = ~pi1615 & w30679;
assign w30682 = ~w30680 & ~w30681;
assign w30683 = ~w30676 & w30682;
assign w30684 = w30663 & w30683;
assign w30685 = w30669 & ~w30675;
assign w30686 = w30663 & w30685;
assign w30687 = w30656 & ~w30682;
assign w30688 = w30676 & w30687;
assign w30689 = ~w30686 & ~w30688;
assign w30690 = w30669 & ~w30682;
assign w30691 = ~w30656 & w30690;
assign w30692 = ~w30656 & ~w30662;
assign w30693 = ~w30669 & w30682;
assign w30694 = w30675 & ~w30693;
assign w30695 = w30692 & ~w30694;
assign w30696 = ~w30684 & ~w30691;
assign w30697 = w30689 & ~w30695;
assign w30698 = w30696 & w30697;
assign w30699 = ~w30650 & ~w30698;
assign w30700 = w30656 & w30669;
assign w30701 = ~w30656 & ~w30669;
assign w30702 = ~w30700 & ~w30701;
assign w30703 = w30682 & ~w30702;
assign w30704 = ~w30702 & w63329;
assign w30705 = ~w30702 & w63402;
assign w30706 = ~w30692 & ~w30705;
assign w30707 = w30698 & ~w30706;
assign w30708 = w30675 & w30693;
assign w30709 = ~w30675 & ~w30690;
assign w30710 = ~w30693 & w30709;
assign w30711 = w30709 & w63403;
assign w30712 = ~w30669 & ~w30675;
assign w30713 = ~w30656 & w30712;
assign w30714 = ~w30708 & ~w30713;
assign w30715 = ~w30711 & w30714;
assign w30716 = ~w30692 & ~w30715;
assign w30717 = ~w30707 & ~w30716;
assign w30718 = (w30650 & w30707) | (w30650 & w65889) | (w30707 & w65889);
assign w30719 = ~w30662 & ~w30675;
assign w30720 = w30662 & w30675;
assign w30721 = ~w30719 & ~w30720;
assign w30722 = w30702 & ~w30721;
assign w30723 = w30669 & w30675;
assign w30724 = w30656 & ~w30662;
assign w30725 = w30723 & w30724;
assign w30726 = ~w30722 & ~w30725;
assign w30727 = ~w30682 & ~w30726;
assign w30728 = ~w30699 & ~w30727;
assign w30729 = ~w30718 & w30728;
assign w30730 = pi1642 & w30729;
assign w30731 = ~pi1642 & ~w30729;
assign w30732 = ~w30730 & ~w30731;
assign w30733 = w30564 & ~w30578;
assign w30734 = ~w30548 & w30590;
assign w30735 = ~w30535 & w30572;
assign w30736 = ~w30574 & ~w30735;
assign w30737 = ~w30558 & w30736;
assign w30738 = ~w30734 & ~w30737;
assign w30739 = w30733 & w30738;
assign w30740 = ~w30542 & w30564;
assign w30741 = w30736 & ~w30740;
assign w30742 = w30738 & w65890;
assign w30743 = w30564 & ~w30583;
assign w30744 = ~w30734 & w30743;
assign w30745 = w30542 & w30574;
assign w30746 = ~w30564 & ~w30745;
assign w30747 = ~w30608 & ~w30744;
assign w30748 = ~w30746 & w30747;
assign w30749 = w30736 & w65891;
assign w30750 = w30586 & ~w30749;
assign w30751 = ~w30564 & w30584;
assign w30752 = ~w30565 & ~w30751;
assign w30753 = (~w30595 & w30751) | (~w30595 & w65892) | (w30751 & w65892);
assign w30754 = (w30555 & w30750) | (w30555 & w65893) | (w30750 & w65893);
assign w30755 = w30548 & w30564;
assign w30756 = ~w30591 & ~w30755;
assign w30757 = w30598 & ~w30756;
assign w30758 = w30597 & w30755;
assign w30759 = w30565 & w30573;
assign w30760 = ~w30555 & ~w30734;
assign w30761 = w30579 & w30760;
assign w30762 = ~w30757 & ~w30759;
assign w30763 = w30761 & w30762;
assign w30764 = ~w30758 & w30763;
assign w30765 = ~w30754 & ~w30764;
assign w30766 = ~w30742 & ~w30748;
assign w30767 = ~w30765 & w30766;
assign w30768 = pi1632 & ~w30767;
assign w30769 = ~pi1632 & w30767;
assign w30770 = ~w30768 & ~w30769;
assign w30771 = ~w30352 & ~w30365;
assign w30772 = ~w30341 & w30357;
assign w30773 = w30323 & w30622;
assign w30774 = ~w30362 & ~w30772;
assign w30775 = ~w30773 & w30774;
assign w30776 = w30352 & ~w30775;
assign w30777 = ~w30354 & w30495;
assign w30778 = ~w30357 & w30361;
assign w30779 = ~w30628 & w30778;
assign w30780 = ~w30777 & w30779;
assign w30781 = ~w30771 & ~w30780;
assign w30782 = ~w30776 & w30781;
assign w30783 = ~pi1633 & w30782;
assign w30784 = pi1633 & ~w30782;
assign w30785 = ~w30783 & ~w30784;
assign w30786 = ~w30702 & w63858;
assign w30787 = ~w30687 & w30712;
assign w30788 = ~w30786 & w30787;
assign w30789 = w30662 & ~w30690;
assign w30790 = ~w30700 & w30789;
assign w30791 = w30675 & ~w30724;
assign w30792 = ~w30790 & w30791;
assign w30793 = ~w30788 & ~w30792;
assign w30794 = w30663 & w30693;
assign w30795 = w30669 & w30719;
assign w30796 = w30682 & w30795;
assign w30797 = ~w30794 & ~w30796;
assign w30798 = (~w30650 & ~w30793) | (~w30650 & w65894) | (~w30793 & w65894);
assign w30799 = w30701 & w30793;
assign w30800 = ~w30662 & ~w30682;
assign w30801 = w30702 & w30800;
assign w30802 = w30689 & ~w30801;
assign w30803 = ~w30705 & w30802;
assign w30804 = (w30650 & w30799) | (w30650 & w65895) | (w30799 & w65895);
assign w30805 = ~w30682 & w30686;
assign w30806 = ~w30656 & w30662;
assign w30807 = w30709 & w63859;
assign w30808 = ~w30662 & w30688;
assign w30809 = ~w30805 & ~w30808;
assign w30810 = ~w30807 & w30809;
assign w30811 = ~w30798 & w30810;
assign w30812 = ~w30804 & w30811;
assign w30813 = pi1645 & w30812;
assign w30814 = ~pi1645 & ~w30812;
assign w30815 = ~w30813 & ~w30814;
assign w30816 = ~pi5405 & pi9040;
assign w30817 = ~pi5305 & ~pi9040;
assign w30818 = ~w30816 & ~w30817;
assign w30819 = pi1610 & ~w30818;
assign w30820 = ~pi1610 & w30818;
assign w30821 = ~w30819 & ~w30820;
assign w30822 = ~pi5398 & pi9040;
assign w30823 = ~pi5436 & ~pi9040;
assign w30824 = ~w30822 & ~w30823;
assign w30825 = pi1626 & ~w30824;
assign w30826 = ~pi1626 & w30824;
assign w30827 = ~w30825 & ~w30826;
assign w30828 = ~pi5304 & pi9040;
assign w30829 = ~pi5306 & ~pi9040;
assign w30830 = ~w30828 & ~w30829;
assign w30831 = pi1591 & ~w30830;
assign w30832 = ~pi1591 & w30830;
assign w30833 = ~w30831 & ~w30832;
assign w30834 = ~pi5299 & pi9040;
assign w30835 = ~pi5573 & ~pi9040;
assign w30836 = ~w30834 & ~w30835;
assign w30837 = pi1618 & ~w30836;
assign w30838 = ~pi1618 & w30836;
assign w30839 = ~w30837 & ~w30838;
assign w30840 = ~w30833 & w30839;
assign w30841 = ~pi5665 & pi9040;
assign w30842 = ~pi5325 & ~pi9040;
assign w30843 = ~w30841 & ~w30842;
assign w30844 = pi1616 & ~w30843;
assign w30845 = ~pi1616 & w30843;
assign w30846 = ~w30844 & ~w30845;
assign w30847 = ~pi5321 & pi9040;
assign w30848 = ~pi5403 & ~pi9040;
assign w30849 = ~w30847 & ~w30848;
assign w30850 = pi1622 & ~w30849;
assign w30851 = ~pi1622 & w30849;
assign w30852 = ~w30850 & ~w30851;
assign w30853 = w30846 & w30852;
assign w30854 = w30840 & w30853;
assign w30855 = w30827 & w30854;
assign w30856 = ~w30840 & w30853;
assign w30857 = w30840 & ~w30852;
assign w30858 = ~w30856 & ~w30857;
assign w30859 = ~w30827 & ~w30858;
assign w30860 = w30833 & ~w30839;
assign w30861 = ~w30840 & ~w30860;
assign w30862 = w30839 & w30852;
assign w30863 = ~w30861 & ~w30862;
assign w30864 = ~w30846 & w30863;
assign w30865 = ~w30855 & ~w30859;
assign w30866 = ~w30864 & w30865;
assign w30867 = ~w30821 & ~w30866;
assign w30868 = w30827 & w30833;
assign w30869 = w30846 & ~w30852;
assign w30870 = w30868 & ~w30869;
assign w30871 = ~w30839 & ~w30852;
assign w30872 = w30833 & ~w30846;
assign w30873 = w30871 & ~w30872;
assign w30874 = ~w30854 & ~w30873;
assign w30875 = ~w30827 & ~w30874;
assign w30876 = ~w30846 & w30852;
assign w30877 = w30861 & w30876;
assign w30878 = ~w30870 & ~w30877;
assign w30879 = ~w30875 & w30878;
assign w30880 = w30821 & ~w30879;
assign w30881 = ~w30852 & ~w30868;
assign w30882 = w30821 & ~w30881;
assign w30883 = ~w30827 & ~w30833;
assign w30884 = ~w30846 & ~w30883;
assign w30885 = w30839 & ~w30846;
assign w30886 = w30839 & ~w30852;
assign w30887 = w30833 & w30886;
assign w30888 = ~w30885 & ~w30887;
assign w30889 = ~w30884 & ~w30888;
assign w30890 = ~w30882 & w30889;
assign w30891 = ~w30833 & ~w30839;
assign w30892 = w30869 & w30891;
assign w30893 = w30852 & w30872;
assign w30894 = ~w30892 & ~w30893;
assign w30895 = w30827 & ~w30894;
assign w30896 = ~w30890 & ~w30895;
assign w30897 = ~w30880 & w30896;
assign w30898 = ~w30867 & w30897;
assign w30899 = pi1641 & ~w30898;
assign w30900 = ~pi1641 & w30898;
assign w30901 = ~w30899 & ~w30900;
assign w30902 = ~w30178 & ~w30184;
assign w30903 = ~w30119 & ~w30146;
assign w30904 = ~w30097 & w65896;
assign w30905 = ~w30903 & w30904;
assign w30906 = w30902 & ~w30905;
assign w30907 = ~w30126 & ~w30906;
assign w30908 = ~w30172 & ~w30518;
assign w30909 = w30135 & ~w30908;
assign w30910 = w30129 & w30182;
assign w30911 = w30151 & w30902;
assign w30912 = ~w30113 & ~w30910;
assign w30913 = ~w30911 & w30912;
assign w30914 = w30126 & ~w30913;
assign w30915 = ~w30156 & w30188;
assign w30916 = ~w30116 & ~w30915;
assign w30917 = ~w30088 & ~w30916;
assign w30918 = ~w30111 & ~w30917;
assign w30919 = ~w30082 & ~w30157;
assign w30920 = ~w30918 & w30919;
assign w30921 = ~w30909 & ~w30914;
assign w30922 = ~w30907 & w30921;
assign w30923 = w30922 & w65897;
assign w30924 = (~pi1658 & ~w30922) | (~pi1658 & w65898) | (~w30922 & w65898);
assign w30925 = ~w30923 & ~w30924;
assign w30926 = w30399 & ~w30429;
assign w30927 = ~w30440 & ~w30926;
assign w30928 = ~w30406 & ~w30927;
assign w30929 = ~w30419 & ~w30421;
assign w30930 = ~w30429 & ~w30929;
assign w30931 = w30399 & ~w30437;
assign w30932 = ~w30435 & ~w30931;
assign w30933 = w30446 & ~w30465;
assign w30934 = w30451 & ~w30932;
assign w30935 = ~w30933 & w30934;
assign w30936 = w30412 & w30435;
assign w30937 = w30435 & w65899;
assign w30938 = ~w30439 & ~w30937;
assign w30939 = w30438 & ~w30938;
assign w30940 = ~w30461 & ~w30930;
assign w30941 = ~w30928 & w30940;
assign w30942 = ~w30935 & w30941;
assign w30943 = ~w30939 & w30942;
assign w30944 = w30420 & w30450;
assign w30945 = ~w30470 & ~w30471;
assign w30946 = w30429 & ~w30945;
assign w30947 = w30406 & w30412;
assign w30948 = ~w30434 & ~w30947;
assign w30949 = ~w30933 & w30948;
assign w30950 = ~w30438 & ~w30471;
assign w30951 = ~w30949 & w30950;
assign w30952 = w30461 & ~w30944;
assign w30953 = ~w30946 & w30952;
assign w30954 = ~w30951 & w30953;
assign w30955 = ~w30943 & ~w30954;
assign w30956 = ~pi1643 & w30955;
assign w30957 = pi1643 & ~w30955;
assign w30958 = ~w30956 & ~w30957;
assign w30959 = ~w30743 & ~w30755;
assign w30960 = ~w30577 & ~w30959;
assign w30961 = w30738 & w30960;
assign w30962 = ~w30738 & w30751;
assign w30963 = ~w30584 & w30595;
assign w30964 = ~w30745 & ~w30963;
assign w30965 = ~w30962 & w30964;
assign w30966 = (w30555 & ~w30965) | (w30555 & w65900) | (~w30965 & w65900);
assign w30967 = ~w30555 & ~w30739;
assign w30968 = w30574 & w30590;
assign w30969 = w30733 & ~w30968;
assign w30970 = w30752 & ~w30969;
assign w30971 = ~w30967 & ~w30970;
assign w30972 = (~w30752 & w30962) | (~w30752 & w65901) | (w30962 & w65901);
assign w30973 = ~w30971 & ~w30972;
assign w30974 = ~w30973 & w65902;
assign w30975 = (~pi1636 & w30973) | (~pi1636 & w65903) | (w30973 & w65903);
assign w30976 = ~w30974 & ~w30975;
assign w30977 = w30853 & ~w30861;
assign w30978 = ~w30846 & w30871;
assign w30979 = ~w30887 & ~w30978;
assign w30980 = w30827 & ~w30979;
assign w30981 = ~w30892 & ~w30977;
assign w30982 = ~w30980 & w30981;
assign w30983 = ~w30821 & w30982;
assign w30984 = ~w30827 & ~w30979;
assign w30985 = w30827 & ~w30886;
assign w30986 = w30982 & w30985;
assign w30987 = ~w30869 & ~w30876;
assign w30988 = w30840 & ~w30987;
assign w30989 = w30821 & ~w30988;
assign w30990 = ~w30984 & w30989;
assign w30991 = ~w30986 & w30990;
assign w30992 = ~w30983 & ~w30991;
assign w30993 = w30833 & w30852;
assign w30994 = ~w30833 & ~w30846;
assign w30995 = ~w30886 & ~w30994;
assign w30996 = ~w30885 & ~w30995;
assign w30997 = w30979 & w30996;
assign w30998 = ~w30857 & ~w30993;
assign w30999 = (~w30821 & w30997) | (~w30821 & w65904) | (w30997 & w65904);
assign w31000 = w30853 & w30860;
assign w31001 = ~w30833 & w30846;
assign w31002 = ~w30852 & w31001;
assign w31003 = ~w31000 & ~w31002;
assign w31004 = ~w30999 & w31003;
assign w31005 = ~w30827 & ~w31004;
assign w31006 = ~w30992 & w65905;
assign w31007 = (pi1638 & w30992) | (pi1638 & w65906) | (w30992 & w65906);
assign w31008 = ~w31006 & ~w31007;
assign w31009 = (w30429 & ~w30932) | (w30429 & w65907) | (~w30932 & w65907);
assign w31010 = ~w30429 & ~w30947;
assign w31011 = ~w30447 & ~w30936;
assign w31012 = w31010 & w31011;
assign w31013 = (w30938 & w31012) | (w30938 & w65908) | (w31012 & w65908);
assign w31014 = w30461 & ~w31013;
assign w31015 = ~w30461 & ~w30932;
assign w31016 = ~w30937 & w31015;
assign w31017 = w30430 & ~w31016;
assign w31018 = (~w30423 & ~w30932) | (~w30423 & w65909) | (~w30932 & w65909);
assign w31019 = ~w30461 & ~w31018;
assign w31020 = ~w30429 & w30938;
assign w31021 = ~w31019 & w31020;
assign w31022 = ~w31017 & ~w31021;
assign w31023 = ~w31014 & ~w31022;
assign w31024 = ~pi1655 & w31023;
assign w31025 = pi1655 & ~w31023;
assign w31026 = ~w31024 & ~w31025;
assign w31027 = ~w30852 & w30860;
assign w31028 = ~w30997 & ~w31027;
assign w31029 = (~w30821 & w30997) | (~w30821 & w65910) | (w30997 & w65910);
assign w31030 = w30872 & w30862;
assign w31031 = ~w31000 & ~w31030;
assign w31032 = ~w31029 & w31031;
assign w31033 = ~w30827 & ~w31032;
assign w31034 = ~w30827 & ~w30995;
assign w31035 = ~w30883 & ~w30996;
assign w31036 = ~w31034 & ~w31035;
assign w31037 = w30871 & w30872;
assign w31038 = w30821 & ~w31037;
assign w31039 = ~w30889 & w65911;
assign w31040 = ~w31036 & w31039;
assign w31041 = w30884 & w30886;
assign w31042 = w30985 & w31031;
assign w31043 = ~w30821 & ~w31041;
assign w31044 = (w31043 & ~w31028) | (w31043 & w65912) | (~w31028 & w65912);
assign w31045 = ~w31040 & ~w31044;
assign w31046 = ~w31033 & ~w31045;
assign w31047 = pi1647 & w31046;
assign w31048 = ~pi1647 & ~w31046;
assign w31049 = ~w31047 & ~w31048;
assign w31050 = ~w30687 & w30795;
assign w31051 = w30663 & w30712;
assign w31052 = ~w30704 & ~w31051;
assign w31053 = w30691 & w30720;
assign w31054 = ~w30808 & ~w31050;
assign w31055 = ~w31053 & w31054;
assign w31056 = w31052 & w31055;
assign w31057 = w31055 & w63404;
assign w31058 = w30662 & w30682;
assign w31059 = w30713 & ~w31058;
assign w31060 = ~w30669 & ~w30800;
assign w31061 = (~w31059 & ~w30715) | (~w31059 & w63861) | (~w30715 & w63861);
assign w31062 = (w31061 & ~w30717) | (w31061 & w63405) | (~w30717 & w63405);
assign w31063 = ~w30650 & ~w31062;
assign w31064 = ~w30662 & w30704;
assign w31065 = w30650 & ~w31056;
assign w31066 = w30713 & w30800;
assign w31067 = ~w30794 & ~w30805;
assign w31068 = ~w31066 & w31067;
assign w31069 = ~w31064 & w31068;
assign w31070 = (pi1648 & w31063) | (pi1648 & w63862) | (w31063 & w63862);
assign w31071 = ~w31063 & w63863;
assign w31072 = ~w31070 & ~w31071;
assign w31073 = w30251 & w30287;
assign w31074 = (~w30243 & ~w30231) | (~w30243 & w63864) | (~w30231 & w63864);
assign w31075 = ~w30246 & w31074;
assign w31076 = (~w30278 & ~w31075) | (~w30278 & w65913) | (~w31075 & w65913);
assign w31077 = w30265 & w31076;
assign w31078 = ~w30248 & ~w30253;
assign w31079 = w30204 & ~w30245;
assign w31080 = ~w30231 & w31078;
assign w31081 = ~w31079 & w31080;
assign w31082 = w30219 & ~w30253;
assign w31083 = ~w30213 & w31082;
assign w31084 = ~w30230 & w30249;
assign w31085 = ~w31083 & w31084;
assign w31086 = w30278 & ~w31081;
assign w31087 = ~w31085 & w31086;
assign w31088 = ~w30266 & w31087;
assign w31089 = ~w31077 & ~w31088;
assign w31090 = ~w30204 & ~w30210;
assign w31091 = w30247 & w31090;
assign w31092 = ~w31089 & w63865;
assign w31093 = (~pi1651 & w31089) | (~pi1651 & w63866) | (w31089 & w63866);
assign w31094 = ~w31092 & ~w31093;
assign w31095 = w30226 & w30249;
assign w31096 = ~w30237 & ~w30288;
assign w31097 = ~w30231 & w30253;
assign w31098 = ~w30258 & w31097;
assign w31099 = ~w30235 & ~w30253;
assign w31100 = ~w30228 & w31099;
assign w31101 = ~w30250 & w31100;
assign w31102 = ~w31098 & ~w31101;
assign w31103 = w31076 & w31102;
assign w31104 = ~w30212 & ~w30219;
assign w31105 = w31078 & w31104;
assign w31106 = w30283 & ~w31075;
assign w31107 = w30268 & w31090;
assign w31108 = ~w31105 & ~w31107;
assign w31109 = w30280 & w31108;
assign w31110 = ~w31106 & w31109;
assign w31111 = ~w31103 & ~w31110;
assign w31112 = (~w31095 & ~w30265) | (~w31095 & w65914) | (~w30265 & w65914);
assign w31113 = ~w31096 & ~w31111;
assign w31114 = (pi1671 & ~w31113) | (pi1671 & w65915) | (~w31113 & w65915);
assign w31115 = w31113 & w65916;
assign w31116 = ~w31114 & ~w31115;
assign w31117 = ~pi5303 & pi9040;
assign w31118 = ~pi5321 & ~pi9040;
assign w31119 = ~w31117 & ~w31118;
assign w31120 = pi1604 & ~w31119;
assign w31121 = ~pi1604 & w31119;
assign w31122 = ~w31120 & ~w31121;
assign w31123 = ~pi5502 & pi9040;
assign w31124 = ~pi5324 & ~pi9040;
assign w31125 = ~w31123 & ~w31124;
assign w31126 = pi1610 & ~w31125;
assign w31127 = ~pi1610 & w31125;
assign w31128 = ~w31126 & ~w31127;
assign w31129 = w31122 & ~w31128;
assign w31130 = ~pi5313 & pi9040;
assign w31131 = ~pi5319 & ~pi9040;
assign w31132 = ~w31130 & ~w31131;
assign w31133 = pi1618 & ~w31132;
assign w31134 = ~pi1618 & w31132;
assign w31135 = ~w31133 & ~w31134;
assign w31136 = ~pi5399 & pi9040;
assign w31137 = ~pi5566 & ~pi9040;
assign w31138 = ~w31136 & ~w31137;
assign w31139 = pi1613 & ~w31138;
assign w31140 = ~pi1613 & w31138;
assign w31141 = ~w31139 & ~w31140;
assign w31142 = w31135 & ~w31141;
assign w31143 = ~pi5293 & pi9040;
assign w31144 = ~pi5576 & ~pi9040;
assign w31145 = ~w31143 & ~w31144;
assign w31146 = pi1609 & ~w31145;
assign w31147 = ~pi1609 & w31145;
assign w31148 = ~w31146 & ~w31147;
assign w31149 = ~w31128 & ~w31148;
assign w31150 = w31141 & w31149;
assign w31151 = ~w31128 & ~w31141;
assign w31152 = w31148 & w31151;
assign w31153 = ~w31150 & ~w31152;
assign w31154 = w31128 & w31141;
assign w31155 = ~w31135 & w31154;
assign w31156 = w31135 & w31149;
assign w31157 = ~w31155 & ~w31156;
assign w31158 = w31153 & w31157;
assign w31159 = w31128 & ~w31148;
assign w31160 = w31135 & w31141;
assign w31161 = ~w31159 & ~w31160;
assign w31162 = w31158 & w63867;
assign w31163 = w31129 & w31162;
assign w31164 = w31122 & ~w31149;
assign w31165 = w31128 & w31148;
assign w31166 = ~w31149 & ~w31165;
assign w31167 = ~w31135 & w31141;
assign w31168 = ~w31166 & w31167;
assign w31169 = w31164 & w31168;
assign w31170 = w31141 & w31156;
assign w31171 = w31135 & ~w31148;
assign w31172 = ~w31142 & ~w31159;
assign w31173 = ~w31171 & ~w31172;
assign w31174 = w31135 & w31165;
assign w31175 = ~w31173 & ~w31174;
assign w31176 = ~w31122 & ~w31175;
assign w31177 = ~pi5328 & pi9040;
assign w31178 = ~pi5508 & ~pi9040;
assign w31179 = ~w31177 & ~w31178;
assign w31180 = pi1614 & ~w31179;
assign w31181 = ~pi1614 & w31179;
assign w31182 = ~w31180 & ~w31181;
assign w31183 = w31164 & ~w31174;
assign w31184 = ~w31173 & w31183;
assign w31185 = ~w31170 & w31182;
assign w31186 = ~w31184 & w31185;
assign w31187 = ~w31176 & w31186;
assign w31188 = ~w31129 & w31166;
assign w31189 = w31160 & w31188;
assign w31190 = ~w31168 & ~w31189;
assign w31191 = (w31142 & ~w31166) | (w31142 & w65917) | (~w31166 & w65917);
assign w31192 = ~w31135 & ~w31141;
assign w31193 = w31166 & w65918;
assign w31194 = ~w31182 & ~w31191;
assign w31195 = ~w31193 & w31194;
assign w31196 = w31190 & w31195;
assign w31197 = ~w31187 & ~w31196;
assign w31198 = ~w31163 & ~w31169;
assign w31199 = ~w31197 & w31198;
assign w31200 = ~pi1681 & w31199;
assign w31201 = pi1681 & ~w31199;
assign w31202 = ~w31200 & ~w31201;
assign w31203 = ~w31173 & w63868;
assign w31204 = w31158 & ~w31203;
assign w31205 = ~w31122 & ~w31159;
assign w31206 = ~w31158 & w31205;
assign w31207 = ~w31204 & ~w31206;
assign w31208 = ~w31182 & ~w31207;
assign w31209 = ~w31122 & ~w31192;
assign w31210 = ~w31166 & w31209;
assign w31211 = w31158 & w65919;
assign w31212 = w31182 & ~w31210;
assign w31213 = ~w31193 & w31212;
assign w31214 = ~w31211 & w31213;
assign w31215 = ~w31208 & ~w31214;
assign w31216 = w31160 & ~w31165;
assign w31217 = w31153 & ~w31193;
assign w31218 = w31122 & ~w31217;
assign w31219 = ~w31154 & ~w31171;
assign w31220 = ~w31122 & ~w31219;
assign w31221 = ~w31151 & ~w31154;
assign w31222 = w31220 & ~w31221;
assign w31223 = ~w31216 & ~w31222;
assign w31224 = ~w31218 & w31223;
assign w31225 = w31157 & ~w31175;
assign w31226 = ~w31224 & w31225;
assign w31227 = ~w31215 & w65920;
assign w31228 = (~pi1673 & w31215) | (~pi1673 & w65921) | (w31215 & w65921);
assign w31229 = ~w31227 & ~w31228;
assign w31230 = ~w31128 & ~w31135;
assign w31231 = ~w31122 & ~w31230;
assign w31232 = w31219 & ~w31231;
assign w31233 = ~w31148 & w31160;
assign w31234 = ~w31220 & ~w31233;
assign w31235 = ~w31232 & w31234;
assign w31236 = ~w31162 & ~w31235;
assign w31237 = ~w31122 & ~w31148;
assign w31238 = w31160 & w31237;
assign w31239 = ~w31182 & ~w31238;
assign w31240 = ~w31224 & ~w31239;
assign w31241 = (~w31169 & w31236) | (~w31169 & w65922) | (w31236 & w65922);
assign w31242 = ~w31240 & w31241;
assign w31243 = ~pi1674 & ~w31242;
assign w31244 = pi1674 & w31242;
assign w31245 = ~w31243 & ~w31244;
assign w31246 = ~w31052 & w31058;
assign w31247 = ~w30709 & w30806;
assign w31248 = w30703 & ~w30723;
assign w31249 = ~w30685 & w30724;
assign w31250 = ~w30683 & w31249;
assign w31251 = ~w31247 & ~w31250;
assign w31252 = ~w31248 & w31251;
assign w31253 = w30650 & ~w31252;
assign w31254 = (w30723 & w30705) | (w30723 & w65923) | (w30705 & w65923);
assign w31255 = w30809 & w63869;
assign w31256 = w30685 & ~w31255;
assign w31257 = w30710 & w31060;
assign w31258 = ~w30688 & ~w30786;
assign w31259 = ~w31257 & w31258;
assign w31260 = ~w31254 & w31259;
assign w31261 = ~w31256 & w31260;
assign w31262 = ~w30650 & ~w31261;
assign w31263 = ~w31246 & ~w31253;
assign w31264 = ~w31262 & w65924;
assign w31265 = (~pi1650 & w31262) | (~pi1650 & w65925) | (w31262 & w65925);
assign w31266 = ~w31264 & ~w31265;
assign w31267 = ~w30749 & ~w30968;
assign w31268 = ~w30564 & ~w31267;
assign w31269 = w30582 & w30960;
assign w31270 = ~w30555 & ~w30589;
assign w31271 = ~w30741 & w31270;
assign w31272 = ~w31269 & w31271;
assign w31273 = ~w30591 & ~w30595;
assign w31274 = w30598 & ~w31273;
assign w31275 = w30564 & ~w30574;
assign w31276 = ~w30596 & w31275;
assign w31277 = w30555 & ~w30745;
assign w31278 = ~w31274 & w31277;
assign w31279 = ~w31276 & w31278;
assign w31280 = ~w30742 & w31279;
assign w31281 = ~w31272 & ~w31280;
assign w31282 = ~w30758 & ~w31268;
assign w31283 = ~w31281 & w31282;
assign w31284 = ~pi1654 & w31283;
assign w31285 = pi1654 & ~w31283;
assign w31286 = ~w31284 & ~w31285;
assign w31287 = w30405 & w30937;
assign w31288 = w30430 & ~w30933;
assign w31289 = w30474 & w31288;
assign w31290 = ~w30443 & ~w31289;
assign w31291 = (w30461 & w31290) | (w30461 & w65926) | (w31290 & w65926);
assign w31292 = w30419 & w30444;
assign w31293 = w31010 & ~w31292;
assign w31294 = w30429 & ~w30469;
assign w31295 = ~w31293 & ~w31294;
assign w31296 = w30420 & ~w30421;
assign w31297 = ~w30452 & w30930;
assign w31298 = (~w30471 & w30466) | (~w30471 & w65927) | (w30466 & w65927);
assign w31299 = ~w30933 & ~w31298;
assign w31300 = ~w31296 & ~w31297;
assign w31301 = (~w30461 & ~w31300) | (~w30461 & w65928) | (~w31300 & w65928);
assign w31302 = ~w31295 & ~w31301;
assign w31303 = ~w31291 & w31302;
assign w31304 = ~pi1653 & w31303;
assign w31305 = pi1653 & ~w31303;
assign w31306 = ~w31304 & ~w31305;
assign w31307 = ~w31122 & w31155;
assign w31308 = w31221 & w31237;
assign w31309 = w31148 & w31230;
assign w31310 = ~w31174 & ~w31309;
assign w31311 = w31129 & w31171;
assign w31312 = w31310 & ~w31311;
assign w31313 = ~w31141 & ~w31312;
assign w31314 = ~w31161 & w31219;
assign w31315 = w31182 & ~w31308;
assign w31316 = ~w31314 & w31315;
assign w31317 = ~w31313 & w31316;
assign w31318 = ~w31148 & w31151;
assign w31319 = w31312 & w31318;
assign w31320 = ~w31135 & ~w31165;
assign w31321 = ~w31122 & ~w31310;
assign w31322 = (~w31182 & ~w31183) | (~w31182 & w65929) | (~w31183 & w65929);
assign w31323 = ~w31321 & w31322;
assign w31324 = ~w31319 & w31323;
assign w31325 = ~w31317 & ~w31324;
assign w31326 = w31122 & ~w31148;
assign w31327 = ~w31190 & w31326;
assign w31328 = ~w31307 & ~w31327;
assign w31329 = ~w31325 & w31328;
assign w31330 = pi1649 & ~w31329;
assign w31331 = ~pi1649 & w31329;
assign w31332 = ~w31330 & ~w31331;
assign w31333 = ~w30212 & ~w30233;
assign w31334 = (~w30243 & w30234) | (~w30243 & w65930) | (w30234 & w65930);
assign w31335 = (w30278 & ~w30290) | (w30278 & w65931) | (~w30290 & w65931);
assign w31336 = ~w30204 & w30235;
assign w31337 = ~w30261 & ~w31336;
assign w31338 = w30243 & ~w31337;
assign w31339 = w30204 & ~w30219;
assign w31340 = ~w30249 & w31339;
assign w31341 = ~w31338 & ~w31340;
assign w31342 = ~w30278 & ~w31341;
assign w31343 = ~w30279 & ~w31105;
assign w31344 = w30252 & ~w31343;
assign w31345 = ~w31335 & ~w31344;
assign w31346 = ~w31334 & w31345;
assign w31347 = ~w31342 & w31346;
assign w31348 = pi1682 & w31347;
assign w31349 = ~pi1682 & ~w31347;
assign w31350 = ~w31348 & ~w31349;
assign w31351 = ~w30885 & ~w30891;
assign w31352 = w30821 & w30852;
assign w31353 = ~w31351 & w31352;
assign w31354 = ~w30887 & ~w31353;
assign w31355 = ~w30827 & ~w31354;
assign w31356 = w30827 & w30863;
assign w31357 = ~w30892 & ~w31356;
assign w31358 = w30821 & ~w31357;
assign w31359 = w30862 & w30868;
assign w31360 = ~w30977 & ~w31359;
assign w31361 = ~w31037 & w31360;
assign w31362 = w31042 & ~w31361;
assign w31363 = ~w30881 & ~w30891;
assign w31364 = ~w30872 & ~w31001;
assign w31365 = ~w31363 & w31364;
assign w31366 = w31360 & ~w31365;
assign w31367 = ~w30821 & ~w31366;
assign w31368 = ~w31355 & ~w31358;
assign w31369 = ~w31362 & ~w31367;
assign w31370 = w31368 & w31369;
assign w31371 = pi1666 & ~w31370;
assign w31372 = ~pi1666 & w31370;
assign w31373 = ~w31371 & ~w31372;
assign w31374 = ~pi5666 & pi9040;
assign w31375 = ~pi5572 & ~pi9040;
assign w31376 = ~w31374 & ~w31375;
assign w31377 = pi1684 & ~w31376;
assign w31378 = ~pi1684 & w31376;
assign w31379 = ~w31377 & ~w31378;
assign w31380 = ~pi5669 & pi9040;
assign w31381 = ~pi5579 & ~pi9040;
assign w31382 = ~w31380 & ~w31381;
assign w31383 = pi1665 & ~w31382;
assign w31384 = ~pi1665 & w31382;
assign w31385 = ~w31383 & ~w31384;
assign w31386 = w31379 & ~w31385;
assign w31387 = ~pi5783 & pi9040;
assign w31388 = ~pi5695 & ~pi9040;
assign w31389 = ~w31387 & ~w31388;
assign w31390 = pi1668 & ~w31389;
assign w31391 = ~pi1668 & w31389;
assign w31392 = ~w31390 & ~w31391;
assign w31393 = ~pi5577 & pi9040;
assign w31394 = ~pi5782 & ~pi9040;
assign w31395 = ~w31393 & ~w31394;
assign w31396 = pi1694 & ~w31395;
assign w31397 = ~pi1694 & w31395;
assign w31398 = ~w31396 & ~w31397;
assign w31399 = ~w31392 & w31398;
assign w31400 = w31386 & w31399;
assign w31401 = ~w31379 & w31385;
assign w31402 = ~w31386 & ~w31401;
assign w31403 = ~w31379 & ~w31398;
assign w31404 = ~w31385 & w31392;
assign w31405 = ~w31403 & w31404;
assign w31406 = ~w31386 & ~w31392;
assign w31407 = ~w31405 & ~w31406;
assign w31408 = w31402 & ~w31407;
assign w31409 = ~w31407 & w65932;
assign w31410 = ~w31400 & ~w31409;
assign w31411 = ~pi5704 & pi9040;
assign w31412 = ~pi5697 & ~pi9040;
assign w31413 = ~w31411 & ~w31412;
assign w31414 = pi1657 & ~w31413;
assign w31415 = ~pi1657 & w31413;
assign w31416 = ~w31414 & ~w31415;
assign w31417 = ~w31410 & w31416;
assign w31418 = ~pi5555 & pi9040;
assign w31419 = ~pi5672 & ~pi9040;
assign w31420 = ~w31418 & ~w31419;
assign w31421 = pi1689 & ~w31420;
assign w31422 = ~pi1689 & w31420;
assign w31423 = ~w31421 & ~w31422;
assign w31424 = ~w31385 & ~w31398;
assign w31425 = ~w31392 & w31424;
assign w31426 = w31385 & ~w31392;
assign w31427 = w31398 & w31426;
assign w31428 = ~w31425 & ~w31427;
assign w31429 = w31379 & w31392;
assign w31430 = ~w31385 & w31398;
assign w31431 = w31429 & w31430;
assign w31432 = ~w31416 & ~w31431;
assign w31433 = w31428 & w31432;
assign w31434 = w31385 & ~w31398;
assign w31435 = ~w31379 & w31392;
assign w31436 = w31434 & ~w31435;
assign w31437 = w31416 & ~w31436;
assign w31438 = ~w31434 & w31435;
assign w31439 = ~w31431 & ~w31438;
assign w31440 = w31437 & w31439;
assign w31441 = w31423 & ~w31433;
assign w31442 = ~w31379 & w31398;
assign w31443 = ~w31401 & ~w31427;
assign w31444 = ~w31416 & ~w31442;
assign w31445 = ~w31443 & w31444;
assign w31446 = ~w31443 & w65933;
assign w31447 = ~w31379 & ~w31416;
assign w31448 = w31430 & w31447;
assign w31449 = ~w31429 & ~w31448;
assign w31450 = w31385 & w31398;
assign w31451 = w31416 & ~w31450;
assign w31452 = ~w31449 & ~w31451;
assign w31453 = w31435 & ~w31450;
assign w31454 = w31416 & ~w31453;
assign w31455 = w31434 & ~w31454;
assign w31456 = ~w31392 & w31416;
assign w31457 = ~w31403 & w31456;
assign w31458 = ~w31402 & w31457;
assign w31459 = ~w31452 & ~w31458;
assign w31460 = ~w31455 & w31459;
assign w31461 = ~w31423 & ~w31460;
assign w31462 = (~w31446 & ~w31441) | (~w31446 & w65934) | (~w31441 & w65934);
assign w31463 = ~w31417 & w31462;
assign w31464 = ~w31461 & w31463;
assign w31465 = pi1696 & ~w31464;
assign w31466 = ~pi1696 & w31464;
assign w31467 = ~w31465 & ~w31466;
assign w31468 = ~pi5664 & pi9040;
assign w31469 = ~pi5588 & ~pi9040;
assign w31470 = ~w31468 & ~w31469;
assign w31471 = pi1659 & ~w31470;
assign w31472 = ~pi1659 & w31470;
assign w31473 = ~w31471 & ~w31472;
assign w31474 = ~pi5785 & pi9040;
assign w31475 = ~pi5783 & ~pi9040;
assign w31476 = ~w31474 & ~w31475;
assign w31477 = pi1690 & ~w31476;
assign w31478 = ~pi1690 & w31476;
assign w31479 = ~w31477 & ~w31478;
assign w31480 = w31473 & w31479;
assign w31481 = ~pi5571 & pi9040;
assign w31482 = ~pi5557 & ~pi9040;
assign w31483 = ~w31481 & ~w31482;
assign w31484 = pi1685 & ~w31483;
assign w31485 = ~pi1685 & w31483;
assign w31486 = ~w31484 & ~w31485;
assign w31487 = ~w31479 & w31486;
assign w31488 = ~pi5697 & pi9040;
assign w31489 = ~pi5582 & ~pi9040;
assign w31490 = ~w31488 & ~w31489;
assign w31491 = pi1680 & ~w31490;
assign w31492 = ~pi1680 & w31490;
assign w31493 = ~w31491 & ~w31492;
assign w31494 = ~w31487 & w31493;
assign w31495 = ~w31480 & ~w31494;
assign w31496 = ~pi5780 & pi9040;
assign w31497 = ~pi5666 & ~pi9040;
assign w31498 = ~w31496 & ~w31497;
assign w31499 = pi1691 & ~w31498;
assign w31500 = ~pi1691 & w31498;
assign w31501 = ~w31499 & ~w31500;
assign w31502 = w31479 & w31501;
assign w31503 = w31495 & w31502;
assign w31504 = ~w31479 & ~w31501;
assign w31505 = w31473 & w31504;
assign w31506 = (w31493 & ~w31504) | (w31493 & w65935) | (~w31504 & w65935);
assign w31507 = ~w31473 & ~w31486;
assign w31508 = ~w31479 & w31501;
assign w31509 = w31507 & w31508;
assign w31510 = w31479 & ~w31486;
assign w31511 = w31473 & w31501;
assign w31512 = w31510 & w31511;
assign w31513 = ~w31505 & ~w31512;
assign w31514 = w31473 & ~w31493;
assign w31515 = w31487 & w31514;
assign w31516 = ~w31509 & ~w31515;
assign w31517 = w31513 & w31516;
assign w31518 = w31486 & w31504;
assign w31519 = ~pi5579 & pi9040;
assign w31520 = ~pi5696 & ~pi9040;
assign w31521 = ~w31519 & ~w31520;
assign w31522 = pi1676 & ~w31521;
assign w31523 = ~pi1676 & w31521;
assign w31524 = ~w31522 & ~w31523;
assign w31525 = w31480 & w31486;
assign w31526 = w31479 & ~w31501;
assign w31527 = w31507 & w31526;
assign w31528 = w31493 & ~w31527;
assign w31529 = ~w31525 & w31528;
assign w31530 = w31528 & w65936;
assign w31531 = ~w31510 & ~w31511;
assign w31532 = w31495 & ~w31531;
assign w31533 = (w31524 & ~w31495) | (w31524 & w65937) | (~w31495 & w65937);
assign w31534 = ~w31530 & w31533;
assign w31535 = w31517 & ~w31518;
assign w31536 = ~w31534 & w31535;
assign w31537 = w31506 & ~w31536;
assign w31538 = w31494 & ~w31510;
assign w31539 = ~w31473 & w31486;
assign w31540 = w31479 & w31539;
assign w31541 = w31513 & ~w31540;
assign w31542 = w31524 & ~w31538;
assign w31543 = ~w31541 & w31542;
assign w31544 = w31473 & ~w31486;
assign w31545 = ~w31501 & w31544;
assign w31546 = ~w31493 & w31504;
assign w31547 = ~w31545 & ~w31546;
assign w31548 = ~w31514 & ~w31547;
assign w31549 = ~w31532 & ~w31548;
assign w31550 = ~w31524 & ~w31549;
assign w31551 = w31480 & w63870;
assign w31552 = ~w31503 & ~w31551;
assign w31553 = ~w31543 & w31552;
assign w31554 = ~w31550 & w31553;
assign w31555 = ~w31537 & w31554;
assign w31556 = pi1703 & ~w31555;
assign w31557 = ~pi1703 & w31555;
assign w31558 = ~w31556 & ~w31557;
assign w31559 = ~pi5784 & pi9040;
assign w31560 = ~pi5577 & ~pi9040;
assign w31561 = ~w31559 & ~w31560;
assign w31562 = pi1664 & ~w31561;
assign w31563 = ~pi1664 & w31561;
assign w31564 = ~w31562 & ~w31563;
assign w31565 = ~pi5588 & pi9040;
assign w31566 = ~pi5574 & ~pi9040;
assign w31567 = ~w31565 & ~w31566;
assign w31568 = pi1668 & ~w31567;
assign w31569 = ~pi1668 & w31567;
assign w31570 = ~w31568 & ~w31569;
assign w31571 = ~w31564 & ~w31570;
assign w31572 = ~pi5701 & pi9040;
assign w31573 = ~pi5661 & ~pi9040;
assign w31574 = ~w31572 & ~w31573;
assign w31575 = pi1693 & ~w31574;
assign w31576 = ~pi1693 & w31574;
assign w31577 = ~w31575 & ~w31576;
assign w31578 = ~pi5699 & pi9040;
assign w31579 = ~pi5554 & ~pi9040;
assign w31580 = ~w31578 & ~w31579;
assign w31581 = pi1670 & ~w31580;
assign w31582 = ~pi1670 & w31580;
assign w31583 = ~w31581 & ~w31582;
assign w31584 = ~w31577 & w31583;
assign w31585 = w31564 & w31570;
assign w31586 = ~w31571 & ~w31585;
assign w31587 = w31584 & w31586;
assign w31588 = (~w31571 & ~w31586) | (~w31571 & w65938) | (~w31586 & w65938);
assign w31589 = w31571 & w31584;
assign w31590 = ~pi5557 & pi9040;
assign w31591 = ~pi5555 & ~pi9040;
assign w31592 = ~w31590 & ~w31591;
assign w31593 = pi1686 & ~w31592;
assign w31594 = ~pi1686 & w31592;
assign w31595 = ~w31593 & ~w31594;
assign w31596 = ~w31589 & w31595;
assign w31597 = ~w31588 & w31596;
assign w31598 = ~pi5702 & pi9040;
assign w31599 = ~pi5705 & ~pi9040;
assign w31600 = ~w31598 & ~w31599;
assign w31601 = pi1665 & ~w31600;
assign w31602 = ~pi1665 & w31600;
assign w31603 = ~w31601 & ~w31602;
assign w31604 = ~w31570 & w31577;
assign w31605 = w31564 & w31604;
assign w31606 = ~w31589 & ~w31605;
assign w31607 = ~w31595 & ~w31606;
assign w31608 = ~w31564 & ~w31583;
assign w31609 = w31570 & ~w31595;
assign w31610 = w31577 & w31608;
assign w31611 = ~w31609 & w31610;
assign w31612 = ~w31607 & ~w31611;
assign w31613 = ~w31603 & ~w31612;
assign w31614 = ~w31577 & ~w31583;
assign w31615 = w31577 & w31583;
assign w31616 = ~w31614 & ~w31615;
assign w31617 = ~w31585 & ~w31609;
assign w31618 = ~w31603 & ~w31617;
assign w31619 = w31564 & ~w31595;
assign w31620 = ~w31618 & ~w31619;
assign w31621 = ~w31616 & ~w31620;
assign w31622 = w31577 & w31595;
assign w31623 = ~w31564 & w31583;
assign w31624 = ~w31583 & w31585;
assign w31625 = ~w31623 & ~w31624;
assign w31626 = w31622 & ~w31625;
assign w31627 = w31570 & ~w31577;
assign w31628 = ~w31577 & w31608;
assign w31629 = ~w31627 & ~w31628;
assign w31630 = ~w31588 & ~w31629;
assign w31631 = ~w31604 & ~w31627;
assign w31632 = w31564 & ~w31631;
assign w31633 = w31570 & w31577;
assign w31634 = ~w31564 & w31633;
assign w31635 = ~w31632 & ~w31634;
assign w31636 = w31609 & ~w31623;
assign w31637 = ~w31635 & w31636;
assign w31638 = ~w31626 & ~w31630;
assign w31639 = ~w31637 & w31638;
assign w31640 = w31603 & ~w31639;
assign w31641 = ~w31597 & ~w31621;
assign w31642 = ~w31613 & w31641;
assign w31643 = ~w31640 & w31642;
assign w31644 = pi1697 & ~w31643;
assign w31645 = ~pi1697 & w31643;
assign w31646 = ~w31644 & ~w31645;
assign w31647 = ~pi5663 & pi9040;
assign w31648 = ~pi5578 & ~pi9040;
assign w31649 = ~w31647 & ~w31648;
assign w31650 = pi1663 & ~w31649;
assign w31651 = ~pi1663 & w31649;
assign w31652 = ~w31650 & ~w31651;
assign w31653 = ~pi5671 & pi9040;
assign w31654 = ~pi5834 & ~pi9040;
assign w31655 = ~w31653 & ~w31654;
assign w31656 = pi1678 & ~w31655;
assign w31657 = ~pi1678 & w31655;
assign w31658 = ~w31656 & ~w31657;
assign w31659 = ~w31652 & w31658;
assign w31660 = ~pi5575 & pi9040;
assign w31661 = ~pi5677 & ~pi9040;
assign w31662 = ~w31660 & ~w31661;
assign w31663 = pi1659 & ~w31662;
assign w31664 = ~pi1659 & w31662;
assign w31665 = ~w31663 & ~w31664;
assign w31666 = ~pi5919 & pi9040;
assign w31667 = ~pi5667 & ~pi9040;
assign w31668 = ~w31666 & ~w31667;
assign w31669 = pi1677 & ~w31668;
assign w31670 = ~pi1677 & w31668;
assign w31671 = ~w31669 & ~w31670;
assign w31672 = ~w31665 & w31671;
assign w31673 = ~w31659 & w31672;
assign w31674 = w31659 & ~w31672;
assign w31675 = ~w31673 & ~w31674;
assign w31676 = w31665 & ~w31671;
assign w31677 = ~pi5553 & pi9040;
assign w31678 = ~pi5564 & ~pi9040;
assign w31679 = ~w31677 & ~w31678;
assign w31680 = pi1692 & ~w31679;
assign w31681 = ~pi1692 & w31679;
assign w31682 = ~w31680 & ~w31681;
assign w31683 = ~w31676 & ~w31682;
assign w31684 = ~w31652 & w31683;
assign w31685 = ~w31675 & w31684;
assign w31686 = w31665 & w31682;
assign w31687 = ~w31658 & w31671;
assign w31688 = ~w31652 & w31687;
assign w31689 = w31658 & ~w31671;
assign w31690 = ~w31652 & w31689;
assign w31691 = ~w31688 & ~w31690;
assign w31692 = w31686 & ~w31691;
assign w31693 = w31658 & ~w31676;
assign w31694 = ~w31658 & w31665;
assign w31695 = ~w31682 & w31694;
assign w31696 = ~w31693 & ~w31695;
assign w31697 = ~w31652 & ~w31671;
assign w31698 = ~w31696 & w31697;
assign w31699 = ~pi5561 & pi9040;
assign w31700 = ~pi5700 & ~pi9040;
assign w31701 = ~w31699 & ~w31700;
assign w31702 = pi1690 & ~w31701;
assign w31703 = ~pi1690 & w31701;
assign w31704 = ~w31702 & ~w31703;
assign w31705 = ~w31676 & w31682;
assign w31706 = ~w31658 & ~w31671;
assign w31707 = w31705 & w31706;
assign w31708 = w31658 & w31671;
assign w31709 = ~w31665 & w31708;
assign w31710 = w31665 & w31689;
assign w31711 = ~w31709 & ~w31710;
assign w31712 = w31676 & w31682;
assign w31713 = ~w31683 & ~w31712;
assign w31714 = w31665 & ~w31713;
assign w31715 = (w31652 & w31714) | (w31652 & w65939) | (w31714 & w65939);
assign w31716 = w31704 & ~w31707;
assign w31717 = ~w31698 & w31716;
assign w31718 = ~w31715 & w31717;
assign w31719 = w31689 & w63884;
assign w31720 = ~w31682 & ~w31719;
assign w31721 = ~w31709 & ~w31719;
assign w31722 = ~w31720 & ~w31721;
assign w31723 = ~w31682 & ~w31710;
assign w31724 = w31652 & ~w31658;
assign w31725 = w31676 & w31724;
assign w31726 = ~w31696 & ~w31725;
assign w31727 = w31723 & ~w31726;
assign w31728 = w31652 & w31682;
assign w31729 = w31693 & w31728;
assign w31730 = ~w31688 & ~w31704;
assign w31731 = ~w31729 & w31730;
assign w31732 = ~w31722 & w31731;
assign w31733 = ~w31727 & w31732;
assign w31734 = ~w31718 & ~w31733;
assign w31735 = ~w31685 & ~w31692;
assign w31736 = ~w31734 & w31735;
assign w31737 = pi1712 & ~w31736;
assign w31738 = ~pi1712 & w31736;
assign w31739 = ~w31737 & ~w31738;
assign w31740 = ~pi5564 & pi9040;
assign w31741 = pi5567 & ~pi9040;
assign w31742 = ~w31740 & ~w31741;
assign w31743 = pi1662 & ~w31742;
assign w31744 = ~pi1662 & w31742;
assign w31745 = ~w31743 & ~w31744;
assign w31746 = ~pi5826 & pi9040;
assign w31747 = ~pi5569 & ~pi9040;
assign w31748 = ~w31746 & ~w31747;
assign w31749 = pi1672 & ~w31748;
assign w31750 = ~pi1672 & w31748;
assign w31751 = ~w31749 & ~w31750;
assign w31752 = ~pi5568 & pi9040;
assign w31753 = ~pi5919 & ~pi9040;
assign w31754 = ~w31752 & ~w31753;
assign w31755 = pi1695 & ~w31754;
assign w31756 = ~pi1695 & w31754;
assign w31757 = ~w31755 & ~w31756;
assign w31758 = ~w31751 & ~w31757;
assign w31759 = ~pi5578 & pi9040;
assign w31760 = ~pi5563 & ~pi9040;
assign w31761 = ~w31759 & ~w31760;
assign w31762 = pi1652 & ~w31761;
assign w31763 = ~pi1652 & w31761;
assign w31764 = ~w31762 & ~w31763;
assign w31765 = w31751 & w31764;
assign w31766 = ~w31758 & ~w31765;
assign w31767 = ~pi5698 & pi9040;
assign w31768 = ~pi5671 & ~pi9040;
assign w31769 = ~w31767 & ~w31768;
assign w31770 = pi1688 & ~w31769;
assign w31771 = ~pi1688 & w31769;
assign w31772 = ~w31770 & ~w31771;
assign w31773 = ~pi5677 & pi9040;
assign w31774 = ~pi5559 & ~pi9040;
assign w31775 = ~w31773 & ~w31774;
assign w31776 = pi1683 & ~w31775;
assign w31777 = ~pi1683 & w31775;
assign w31778 = ~w31776 & ~w31777;
assign w31779 = ~w31772 & ~w31778;
assign w31780 = ~w31766 & w31779;
assign w31781 = w31751 & w31778;
assign w31782 = ~w31764 & w31781;
assign w31783 = ~w31751 & w31764;
assign w31784 = w31778 & ~w31783;
assign w31785 = ~w31782 & w31784;
assign w31786 = ~w31778 & w31783;
assign w31787 = w31783 & w65940;
assign w31788 = (w31772 & w31785) | (w31772 & w65941) | (w31785 & w65941);
assign w31789 = ~w31772 & ~w31782;
assign w31790 = ~w31757 & w31778;
assign w31791 = (w31790 & w31782) | (w31790 & w65942) | (w31782 & w65942);
assign w31792 = w31751 & ~w31778;
assign w31793 = ~w31764 & w31792;
assign w31794 = w31792 & w31801;
assign w31795 = ~w31780 & ~w31794;
assign w31796 = ~w31791 & w31795;
assign w31797 = (w31745 & ~w31796) | (w31745 & w65943) | (~w31796 & w65943);
assign w31798 = w31772 & ~w31778;
assign w31799 = ~w31766 & w31798;
assign w31800 = ~w31778 & ~w31793;
assign w31801 = w31757 & ~w31764;
assign w31802 = ~w31751 & w31801;
assign w31803 = w31789 & ~w31802;
assign w31804 = ~w31800 & w31803;
assign w31805 = w31757 & w31778;
assign w31806 = w31783 & w31805;
assign w31807 = ~w31778 & w31802;
assign w31808 = w31757 & w31782;
assign w31809 = ~w31799 & ~w31806;
assign w31810 = ~w31807 & ~w31808;
assign w31811 = w31809 & w31810;
assign w31812 = ~w31804 & w31811;
assign w31813 = ~w31745 & ~w31812;
assign w31814 = ~w31801 & ~w31805;
assign w31815 = ~w31772 & ~w31784;
assign w31816 = ~w31814 & w31815;
assign w31817 = ~w31797 & ~w31816;
assign w31818 = ~w31813 & w31817;
assign w31819 = pi1700 & w31818;
assign w31820 = ~pi1700 & ~w31818;
assign w31821 = ~w31819 & ~w31820;
assign w31822 = ~pi5563 & pi9040;
assign w31823 = ~pi5575 & ~pi9040;
assign w31824 = ~w31822 & ~w31823;
assign w31825 = pi1683 & ~w31824;
assign w31826 = ~pi1683 & w31824;
assign w31827 = ~w31825 & ~w31826;
assign w31828 = ~pi5667 & pi9040;
assign w31829 = ~pi5706 & ~pi9040;
assign w31830 = ~w31828 & ~w31829;
assign w31831 = pi1684 & ~w31830;
assign w31832 = ~pi1684 & w31830;
assign w31833 = ~w31831 & ~w31832;
assign w31834 = ~pi5569 & pi9040;
assign w31835 = ~pi5830 & ~pi9040;
assign w31836 = ~w31834 & ~w31835;
assign w31837 = pi1661 & ~w31836;
assign w31838 = ~pi1661 & w31836;
assign w31839 = ~w31837 & ~w31838;
assign w31840 = ~pi5581 & pi9040;
assign w31841 = ~pi5698 & ~pi9040;
assign w31842 = ~w31840 & ~w31841;
assign w31843 = pi1652 & ~w31842;
assign w31844 = ~pi1652 & w31842;
assign w31845 = ~w31843 & ~w31844;
assign w31846 = ~w31839 & ~w31845;
assign w31847 = ~pi5700 & pi9040;
assign w31848 = ~pi5568 & ~pi9040;
assign w31849 = ~w31847 & ~w31848;
assign w31850 = pi1689 & ~w31849;
assign w31851 = ~pi1689 & w31849;
assign w31852 = ~w31850 & ~w31851;
assign w31853 = ~w31833 & ~w31852;
assign w31854 = ~w31846 & w31853;
assign w31855 = ~w31833 & w31845;
assign w31856 = ~pi5779 & pi9040;
assign w31857 = ~pi5558 & ~pi9040;
assign w31858 = ~w31856 & ~w31857;
assign w31859 = pi1687 & ~w31858;
assign w31860 = ~pi1687 & w31858;
assign w31861 = ~w31859 & ~w31860;
assign w31862 = ~w31855 & w31861;
assign w31863 = w31833 & w31852;
assign w31864 = ~w31861 & ~w31863;
assign w31865 = ~w31862 & ~w31864;
assign w31866 = ~w31845 & ~w31852;
assign w31867 = w31839 & w31861;
assign w31868 = w31866 & w31867;
assign w31869 = ~w31854 & ~w31868;
assign w31870 = ~w31865 & w31869;
assign w31871 = ~w31839 & w31852;
assign w31872 = ~w31861 & ~w31871;
assign w31873 = w31833 & ~w31845;
assign w31874 = ~w31855 & ~w31873;
assign w31875 = w31852 & w31874;
assign w31876 = w31839 & ~w31875;
assign w31877 = w31870 & w31872;
assign w31878 = ~w31876 & w31877;
assign w31879 = ~w31852 & w31861;
assign w31880 = w31845 & w31879;
assign w31881 = w31845 & w31852;
assign w31882 = ~w31866 & ~w31881;
assign w31883 = ~w31874 & w31882;
assign w31884 = w31839 & w31883;
assign w31885 = (w31883 & w63871) | (w31883 & w63872) | (w63871 & w63872);
assign w31886 = w31839 & w31885;
assign w31887 = w31839 & w31845;
assign w31888 = (w31833 & w31865) | (w31833 & w63873) | (w31865 & w63873);
assign w31889 = ~w31839 & w31845;
assign w31890 = ~w31833 & ~w31839;
assign w31891 = ~w31880 & ~w31890;
assign w31892 = ~w31889 & ~w31891;
assign w31893 = ~w31888 & ~w31892;
assign w31894 = ~w31839 & ~w31882;
assign w31895 = ~w31878 & ~w31886;
assign w31896 = (~w31827 & ~w31895) | (~w31827 & w63874) | (~w31895 & w63874);
assign w31897 = ~w31833 & w31868;
assign w31898 = ~w31852 & ~w31874;
assign w31899 = ~w31863 & ~w31898;
assign w31900 = ~w31846 & ~w31887;
assign w31901 = ~w31861 & ~w31900;
assign w31902 = ~w31899 & w31901;
assign w31903 = w31874 & w63875;
assign w31904 = (~w31839 & w31903) | (~w31839 & w65944) | (w31903 & w65944);
assign w31905 = w31870 & ~w31904;
assign w31906 = w31827 & ~w31905;
assign w31907 = w31852 & w31861;
assign w31908 = w31890 & w31907;
assign w31909 = ~w31897 & ~w31908;
assign w31910 = ~w31902 & w31909;
assign w31911 = ~w31906 & w31910;
assign w31912 = ~w31896 & w65945;
assign w31913 = (pi1708 & w31896) | (pi1708 & w65946) | (w31896 & w65946);
assign w31914 = ~w31912 & ~w31913;
assign w31915 = ~pi5554 & pi9040;
assign w31916 = ~pi5785 & ~pi9040;
assign w31917 = ~w31915 & ~w31916;
assign w31918 = pi1685 & ~w31917;
assign w31919 = ~pi1685 & w31917;
assign w31920 = ~w31918 & ~w31919;
assign w31921 = ~pi5672 & pi9040;
assign w31922 = ~pi5780 & ~pi9040;
assign w31923 = ~w31921 & ~w31922;
assign w31924 = pi1676 & ~w31923;
assign w31925 = ~pi1676 & w31923;
assign w31926 = ~w31924 & ~w31925;
assign w31927 = w31920 & ~w31926;
assign w31928 = ~pi5782 & pi9040;
assign w31929 = ~pi5664 & ~pi9040;
assign w31930 = ~w31928 & ~w31929;
assign w31931 = pi1667 & ~w31930;
assign w31932 = ~pi1667 & w31930;
assign w31933 = ~w31931 & ~w31932;
assign w31934 = ~pi5661 & pi9040;
assign w31935 = ~pi5669 & ~pi9040;
assign w31936 = ~w31934 & ~w31935;
assign w31937 = pi1669 & ~w31936;
assign w31938 = ~pi1669 & w31936;
assign w31939 = ~w31937 & ~w31938;
assign w31940 = (w31939 & ~w31927) | (w31939 & w65947) | (~w31927 & w65947);
assign w31941 = ~w31920 & w31926;
assign w31942 = ~pi5696 & pi9040;
assign w31943 = ~pi5784 & ~pi9040;
assign w31944 = ~w31942 & ~w31943;
assign w31945 = pi1664 & ~w31944;
assign w31946 = ~pi1664 & w31944;
assign w31947 = ~w31945 & ~w31946;
assign w31948 = ~w31933 & ~w31947;
assign w31949 = w31941 & w31948;
assign w31950 = w31920 & w31926;
assign w31951 = w31947 & w31950;
assign w31952 = ~w31949 & ~w31951;
assign w31953 = ~pi5572 & pi9040;
assign w31954 = ~pi5702 & ~pi9040;
assign w31955 = ~w31953 & ~w31954;
assign w31956 = pi1693 & ~w31955;
assign w31957 = ~pi1693 & w31955;
assign w31958 = ~w31956 & ~w31957;
assign w31959 = w31926 & w31947;
assign w31960 = ~w31927 & w31933;
assign w31961 = ~w31920 & ~w31926;
assign w31962 = w31947 & ~w31961;
assign w31963 = ~w31933 & ~w31950;
assign w31964 = w31962 & w31963;
assign w31965 = (~w31939 & ~w31960) | (~w31939 & w65948) | (~w31960 & w65948);
assign w31966 = ~w31964 & w31965;
assign w31967 = (w31958 & ~w31952) | (w31958 & w65949) | (~w31952 & w65949);
assign w31968 = ~w31966 & w31967;
assign w31969 = w31920 & ~w31933;
assign w31970 = ~w31947 & ~w31969;
assign w31971 = ~w31933 & ~w31961;
assign w31972 = (~w31939 & w31961) | (~w31939 & w63876) | (w31961 & w63876);
assign w31973 = ~w31962 & ~w31970;
assign w31974 = ~w31972 & w31973;
assign w31975 = w31973 & w65950;
assign w31976 = w31933 & w31947;
assign w31977 = w31941 & w31976;
assign w31978 = ~w31933 & ~w31939;
assign w31979 = ~w31959 & w31978;
assign w31980 = w31926 & w31979;
assign w31981 = ~w31977 & ~w31980;
assign w31982 = w31926 & ~w31933;
assign w31983 = w31939 & ~w31982;
assign w31984 = w31933 & ~w31941;
assign w31985 = w31983 & ~w31984;
assign w31986 = w31981 & ~w31985;
assign w31987 = ~w31975 & w31986;
assign w31988 = ~w31958 & ~w31987;
assign w31989 = ~w31926 & ~w31947;
assign w31990 = ~w31959 & ~w31989;
assign w31991 = ~w31970 & w31983;
assign w31992 = ~w31990 & w31991;
assign w31993 = ~w31939 & ~w31958;
assign w31994 = ~w31960 & ~w31963;
assign w31995 = w31993 & w31994;
assign w31996 = w31975 & ~w31986;
assign w31997 = w31978 & w31989;
assign w31998 = ~w31920 & w31997;
assign w31999 = ~w31992 & ~w31998;
assign w32000 = ~w31995 & w31999;
assign w32001 = ~w31968 & w32000;
assign w32002 = ~w31996 & w32001;
assign w32003 = (pi1710 & ~w32002) | (pi1710 & w65951) | (~w32002 & w65951);
assign w32004 = w32002 & w65952;
assign w32005 = ~w32003 & ~w32004;
assign w32006 = w31833 & w31879;
assign w32007 = w31900 & w32006;
assign w32008 = ~w31839 & ~w31852;
assign w32009 = w31833 & ~w32008;
assign w32010 = ~w31861 & ~w31882;
assign w32011 = ~w32009 & w32010;
assign w32012 = w31861 & w31875;
assign w32013 = ~w31827 & ~w31884;
assign w32014 = ~w32011 & ~w32012;
assign w32015 = w32013 & w32014;
assign w32016 = ~w31852 & ~w31890;
assign w32017 = w31872 & ~w32016;
assign w32018 = ~w31900 & w32009;
assign w32019 = w31881 & w31890;
assign w32020 = ~w32016 & ~w32019;
assign w32021 = w31861 & ~w32020;
assign w32022 = w31827 & ~w32017;
assign w32023 = ~w32018 & w32022;
assign w32024 = ~w32021 & w32023;
assign w32025 = ~w32015 & ~w32024;
assign w32026 = ~w32007 & ~w32025;
assign w32027 = ~pi1715 & w32026;
assign w32028 = pi1715 & ~w32026;
assign w32029 = ~w32027 & ~w32028;
assign w32030 = ~w31757 & w31764;
assign w32031 = ~w31807 & ~w32030;
assign w32032 = w31772 & ~w31792;
assign w32033 = w31758 & ~w31764;
assign w32034 = w31758 & w65953;
assign w32035 = ~w31786 & ~w32034;
assign w32036 = w32032 & w32035;
assign w32037 = ~w32031 & w32036;
assign w32038 = ~w31783 & ~w31793;
assign w32039 = (~w31757 & w31793) | (~w31757 & w63877) | (w31793 & w63877);
assign w32040 = ~w31757 & w31772;
assign w32041 = ~w32030 & ~w32040;
assign w32042 = w31751 & w31814;
assign w32043 = w32041 & w32042;
assign w32044 = w31783 & w65954;
assign w32045 = w31757 & w31781;
assign w32046 = ~w32044 & ~w32045;
assign w32047 = w31772 & ~w32046;
assign w32048 = ~w31764 & w32047;
assign w32049 = ~w31782 & w65955;
assign w32050 = ~w31800 & w32049;
assign w32051 = ~w31745 & ~w32039;
assign w32052 = ~w32043 & w32051;
assign w32053 = ~w32050 & w32052;
assign w32054 = ~w32048 & w32053;
assign w32055 = w31781 & w32030;
assign w32056 = w32042 & w65956;
assign w32057 = ~w31778 & ~w32030;
assign w32058 = ~w31751 & w32057;
assign w32059 = ~w31808 & ~w32058;
assign w32060 = ~w31772 & ~w32059;
assign w32061 = w31764 & w31772;
assign w32062 = ~w32057 & w32061;
assign w32063 = w31745 & ~w32055;
assign w32064 = ~w32034 & w32063;
assign w32065 = ~w32062 & w32064;
assign w32066 = ~w32056 & w32065;
assign w32067 = ~w32060 & w32066;
assign w32068 = ~w32054 & ~w32067;
assign w32069 = ~w32068 & w65957;
assign w32070 = (pi1716 & w32068) | (pi1716 & w65958) | (w32068 & w65958);
assign w32071 = ~w32069 & ~w32070;
assign w32072 = ~w31948 & w31961;
assign w32073 = ~w31976 & w32072;
assign w32074 = ~w31960 & w31970;
assign w32075 = w31941 & ~w31947;
assign w32076 = ~w31951 & ~w32075;
assign w32077 = w31939 & ~w32074;
assign w32078 = w32076 & w32077;
assign w32079 = w32077 & w63878;
assign w32080 = w31920 & w32079;
assign w32081 = w31972 & ~w31990;
assign w32082 = w31981 & w65959;
assign w32083 = (w31958 & w32080) | (w31958 & w65960) | (w32080 & w65960);
assign w32084 = w31939 & w31947;
assign w32085 = w31969 & w32084;
assign w32086 = w31961 & w31976;
assign w32087 = ~w31947 & w31950;
assign w32088 = w31972 & ~w32087;
assign w32089 = ~w31980 & ~w32088;
assign w32090 = (~w32086 & w32078) | (~w32086 & w63879) | (w32078 & w63879);
assign w32091 = ~w31949 & ~w32085;
assign w32092 = (w32091 & w32090) | (w32091 & w65961) | (w32090 & w65961);
assign w32093 = ~w32083 & w32092;
assign w32094 = pi1701 & ~w32093;
assign w32095 = ~pi1701 & w32093;
assign w32096 = ~w32094 & ~w32095;
assign w32097 = ~w31806 & ~w32055;
assign w32098 = ~w31794 & w32097;
assign w32099 = (~w31772 & ~w32098) | (~w31772 & w65962) | (~w32098 & w65962);
assign w32100 = w32036 & w32097;
assign w32101 = w31792 & ~w32041;
assign w32102 = ~w31745 & ~w32101;
assign w32103 = ~w32099 & w32102;
assign w32104 = ~w32100 & w32103;
assign w32105 = ~w32032 & ~w32040;
assign w32106 = ~w32033 & ~w32105;
assign w32107 = ~w31803 & ~w32106;
assign w32108 = w31745 & ~w32044;
assign w32109 = w32097 & w32108;
assign w32110 = ~w32043 & w32109;
assign w32111 = ~w32107 & w32110;
assign w32112 = ~w32104 & ~w32111;
assign w32113 = ~pi1722 & w32112;
assign w32114 = pi1722 & ~w32112;
assign w32115 = ~w32113 & ~w32114;
assign w32116 = ~w31493 & ~w31518;
assign w32117 = ~w31540 & w32116;
assign w32118 = ~w31529 & ~w32117;
assign w32119 = w31517 & ~w32118;
assign w32120 = ~w31524 & ~w32119;
assign w32121 = ~w31510 & ~w31518;
assign w32122 = (w31493 & w31480) | (w31493 & w65963) | (w31480 & w65963);
assign w32123 = ~w32121 & w32122;
assign w32124 = w31502 & w31507;
assign w32125 = (~w32124 & w32121) | (~w32124 & w65964) | (w32121 & w65964);
assign w32126 = ~w31506 & ~w32125;
assign w32127 = w31493 & ~w31509;
assign w32128 = ~w31539 & ~w31544;
assign w32129 = w31508 & ~w32128;
assign w32130 = ~w31512 & ~w32129;
assign w32131 = w32127 & ~w32130;
assign w32132 = ~w31473 & ~w31508;
assign w32133 = w31538 & w32132;
assign w32134 = ~w31493 & w31526;
assign w32135 = ~w32129 & ~w32134;
assign w32136 = ~w32133 & w32135;
assign w32137 = w31524 & ~w32136;
assign w32138 = ~w32126 & ~w32131;
assign w32139 = ~w32137 & w32138;
assign w32140 = ~w32120 & w32139;
assign w32141 = ~pi1707 & w32140;
assign w32142 = pi1707 & ~w32140;
assign w32143 = ~w32141 & ~w32142;
assign w32144 = ~pi5830 & pi9040;
assign w32145 = ~pi5561 & ~pi9040;
assign w32146 = ~w32144 & ~w32145;
assign w32147 = pi1679 & ~w32146;
assign w32148 = ~pi1679 & w32146;
assign w32149 = ~w32147 & ~w32148;
assign w32150 = ~pi5580 & pi9040;
assign w32151 = ~pi5553 & ~pi9040;
assign w32152 = ~w32150 & ~w32151;
assign w32153 = pi1672 & ~w32152;
assign w32154 = ~pi1672 & w32152;
assign w32155 = ~w32153 & ~w32154;
assign w32156 = ~w32149 & ~w32155;
assign w32157 = ~pi5556 & pi9040;
assign w32158 = ~pi5779 & ~pi9040;
assign w32159 = ~w32157 & ~w32158;
assign w32160 = pi1662 & ~w32159;
assign w32161 = ~pi1662 & w32159;
assign w32162 = ~w32160 & ~w32161;
assign w32163 = ~pi5834 & pi9040;
assign w32164 = ~pi5560 & ~pi9040;
assign w32165 = ~w32163 & ~w32164;
assign w32166 = pi1678 & ~w32165;
assign w32167 = ~pi1678 & w32165;
assign w32168 = ~w32166 & ~w32167;
assign w32169 = w32162 & w32168;
assign w32170 = ~w32162 & ~w32168;
assign w32171 = ~w32169 & ~w32170;
assign w32172 = ~w32156 & ~w32171;
assign w32173 = ~pi5675 & pi9040;
assign w32174 = ~pi5663 & ~pi9040;
assign w32175 = ~w32173 & ~w32174;
assign w32176 = pi1677 & ~w32175;
assign w32177 = ~pi1677 & w32175;
assign w32178 = ~w32176 & ~w32177;
assign w32179 = ~pi5559 & pi9040;
assign w32180 = ~pi5581 & ~pi9040;
assign w32181 = ~w32179 & ~w32180;
assign w32182 = pi1675 & ~w32181;
assign w32183 = ~pi1675 & w32181;
assign w32184 = ~w32182 & ~w32183;
assign w32185 = w32178 & ~w32184;
assign w32186 = w32172 & w32185;
assign w32187 = ~w32155 & w32168;
assign w32188 = ~w32184 & w32187;
assign w32189 = ~w32149 & ~w32162;
assign w32190 = w32188 & w32189;
assign w32191 = w32162 & ~w32168;
assign w32192 = w32156 & w32191;
assign w32193 = ~w32155 & w32162;
assign w32194 = w32149 & w32193;
assign w32195 = ~w32149 & w32168;
assign w32196 = w32149 & ~w32168;
assign w32197 = ~w32195 & ~w32196;
assign w32198 = ~w32162 & ~w32197;
assign w32199 = w32155 & w32170;
assign w32200 = ~w32194 & ~w32199;
assign w32201 = ~w32198 & w32200;
assign w32202 = ~w32149 & w32155;
assign w32203 = w32184 & ~w32202;
assign w32204 = w32201 & w32203;
assign w32205 = (w32178 & w32204) | (w32178 & w63880) | (w32204 & w63880);
assign w32206 = ~w32155 & w32171;
assign w32207 = ~w32171 & ~w32187;
assign w32208 = ~w32206 & ~w32207;
assign w32209 = w32184 & w32208;
assign w32210 = w32170 & w63881;
assign w32211 = ~w32206 & ~w32210;
assign w32212 = (~w32149 & w32206) | (~w32149 & w63882) | (w32206 & w63882);
assign w32213 = ~w32193 & ~w32195;
assign w32214 = w32171 & w32213;
assign w32215 = ~w32187 & ~w32214;
assign w32216 = (w32215 & w32209) | (w32215 & w63883) | (w32209 & w63883);
assign w32217 = w32155 & ~w32168;
assign w32218 = w32149 & w32162;
assign w32219 = ~w32217 & ~w32218;
assign w32220 = ~w32155 & ~w32162;
assign w32221 = ~w32184 & ~w32220;
assign w32222 = w32219 & w32221;
assign w32223 = w32149 & w32155;
assign w32224 = ~w32168 & w32223;
assign w32225 = w32184 & ~w32219;
assign w32226 = ~w32224 & w32225;
assign w32227 = ~w32222 & ~w32226;
assign w32228 = w32216 & w32227;
assign w32229 = w32169 & w32223;
assign w32230 = ~w32169 & ~w32213;
assign w32231 = (~w32178 & w32171) | (~w32178 & w65965) | (w32171 & w65965);
assign w32232 = ~w32230 & w32231;
assign w32233 = ~w32229 & ~w32232;
assign w32234 = ~w32184 & ~w32233;
assign w32235 = (~w32184 & ~w32193) | (~w32184 & w65966) | (~w32193 & w65966);
assign w32236 = (~w32178 & ~w32187) | (~w32178 & w65967) | (~w32187 & w65967);
assign w32237 = ~w32235 & w32236;
assign w32238 = ~w32201 & w32237;
assign w32239 = ~w32186 & ~w32238;
assign w32240 = ~w32205 & w32239;
assign w32241 = ~w32234 & w32240;
assign w32242 = w32241 & w65968;
assign w32243 = (~pi1727 & ~w32241) | (~pi1727 & w65969) | (~w32241 & w65969);
assign w32244 = ~w32242 & ~w32243;
assign w32245 = w31687 & w63884;
assign w32246 = w31652 & ~w31682;
assign w32247 = w31672 & w32246;
assign w32248 = ~w31672 & ~w31690;
assign w32249 = ~w31665 & ~w31724;
assign w32250 = w32248 & w32249;
assign w32251 = w31682 & ~w31694;
assign w32252 = w32248 & w32251;
assign w32253 = ~w31695 & ~w32247;
assign w32254 = ~w32245 & w32253;
assign w32255 = ~w32250 & w32254;
assign w32256 = (~w31704 & ~w32255) | (~w31704 & w65970) | (~w32255 & w65970);
assign w32257 = w31652 & w31665;
assign w32258 = w31708 & w32257;
assign w32259 = w32255 & w63885;
assign w32260 = (~w32258 & w31691) | (~w32258 & w65971) | (w31691 & w65971);
assign w32261 = ~w31722 & w32260;
assign w32262 = (w31704 & w32259) | (w31704 & w65972) | (w32259 & w65972);
assign w32263 = ~w31652 & ~w31711;
assign w32264 = ~w31672 & ~w31682;
assign w32265 = ~w31687 & w32264;
assign w32266 = ~w32247 & ~w32265;
assign w32267 = w31682 & ~w31697;
assign w32268 = w31671 & w31724;
assign w32269 = w32267 & ~w32268;
assign w32270 = ~w31686 & ~w32269;
assign w32271 = w32266 & w32270;
assign w32272 = (~w32258 & w31711) | (~w32258 & w65973) | (w31711 & w65973);
assign w32273 = ~w32271 & w32272;
assign w32274 = w31689 & w31705;
assign w32275 = ~w31725 & ~w32258;
assign w32276 = ~w32274 & w32275;
assign w32277 = w31713 & w32276;
assign w32278 = ~w32273 & w32277;
assign w32279 = ~w32256 & ~w32278;
assign w32280 = w32279 & w65974;
assign w32281 = (~pi1711 & ~w32279) | (~pi1711 & w65975) | (~w32279 & w65975);
assign w32282 = ~w32280 & ~w32281;
assign w32283 = w31706 & w32249;
assign w32284 = w32276 & ~w32283;
assign w32285 = ~w32266 & ~w32284;
assign w32286 = ~w31689 & ~w32263;
assign w32287 = w32267 & ~w32286;
assign w32288 = (~w31708 & w31713) | (~w31708 & w65976) | (w31713 & w65976);
assign w32289 = ~w31652 & ~w32288;
assign w32290 = w31682 & ~w32245;
assign w32291 = w31687 & w32290;
assign w32292 = ~w31665 & ~w31682;
assign w32293 = w31706 & w32292;
assign w32294 = ~w31704 & ~w32293;
assign w32295 = ~w32250 & w32294;
assign w32296 = ~w32291 & w32295;
assign w32297 = ~w32289 & w32296;
assign w32298 = ~w31673 & w31720;
assign w32299 = ~w32290 & ~w32298;
assign w32300 = w31704 & w32276;
assign w32301 = ~w32299 & w32300;
assign w32302 = ~w32297 & ~w32301;
assign w32303 = ~w32285 & ~w32287;
assign w32304 = (~pi1721 & w32302) | (~pi1721 & w65977) | (w32302 & w65977);
assign w32305 = ~w32302 & w65978;
assign w32306 = ~w32304 & ~w32305;
assign w32307 = w31608 & w31633;
assign w32308 = w31564 & w31584;
assign w32309 = w31583 & w31604;
assign w32310 = ~w32308 & ~w32309;
assign w32311 = ~w31588 & ~w32310;
assign w32312 = (~w31595 & ~w31608) | (~w31595 & w65979) | (~w31608 & w65979);
assign w32313 = w32310 & w32312;
assign w32314 = ~w31624 & ~w32313;
assign w32315 = w31627 & ~w32314;
assign w32316 = w31564 & ~w31614;
assign w32317 = ~w31570 & w31628;
assign w32318 = ~w32316 & ~w32317;
assign w32319 = w31595 & ~w32308;
assign w32320 = ~w32318 & w32319;
assign w32321 = w31603 & ~w32307;
assign w32322 = ~w32311 & w32321;
assign w32323 = ~w32320 & w32322;
assign w32324 = ~w32315 & w32323;
assign w32325 = w31570 & w31617;
assign w32326 = ~w31615 & ~w32325;
assign w32327 = ~w31622 & ~w32326;
assign w32328 = ~w31586 & ~w32319;
assign w32329 = ~w31608 & w31631;
assign w32330 = ~w31583 & w31604;
assign w32331 = ~w32329 & ~w32330;
assign w32332 = w32318 & ~w32331;
assign w32333 = ~w31603 & ~w32328;
assign w32334 = ~w32327 & w32333;
assign w32335 = ~w32332 & w32334;
assign w32336 = ~w32324 & ~w32335;
assign w32337 = pi1698 & w32336;
assign w32338 = ~pi1698 & ~w32336;
assign w32339 = ~w32337 & ~w32338;
assign w32340 = ~w31502 & ~w31507;
assign w32341 = ~w31510 & ~w32340;
assign w32342 = w31506 & ~w32341;
assign w32343 = ~w31493 & ~w31551;
assign w32344 = ~w31526 & ~w32128;
assign w32345 = ~w31527 & ~w32344;
assign w32346 = w32343 & w32345;
assign w32347 = ~w32346 & w65980;
assign w32348 = ~w31493 & ~w32129;
assign w32349 = w31479 & w31545;
assign w32350 = w32127 & ~w32349;
assign w32351 = ~w32348 & ~w32350;
assign w32352 = ~w31546 & w32128;
assign w32353 = ~w32344 & ~w32352;
assign w32354 = ~w31525 & ~w32122;
assign w32355 = (~w32354 & w32346) | (~w32354 & w63886) | (w32346 & w63886);
assign w32356 = ~w32124 & ~w32353;
assign w32357 = (w31524 & w32355) | (w31524 & w65981) | (w32355 & w65981);
assign w32358 = ~w32347 & ~w32351;
assign w32359 = ~w32357 & w32358;
assign w32360 = ~pi1714 & w32359;
assign w32361 = pi1714 & ~w32359;
assign w32362 = ~w32360 & ~w32361;
assign w32363 = w32178 & w32223;
assign w32364 = w32170 & w32363;
assign w32365 = ~w32172 & ~w32190;
assign w32366 = ~w32223 & ~w32365;
assign w32367 = (w32223 & w32222) | (w32223 & w65982) | (w32222 & w65982);
assign w32368 = ~w32366 & ~w32367;
assign w32369 = ~w32216 & w32368;
assign w32370 = ~w32178 & ~w32369;
assign w32371 = (w32178 & w32214) | (w32178 & w65983) | (w32214 & w65983);
assign w32372 = ~w32155 & ~w32191;
assign w32373 = w32197 & w32372;
assign w32374 = ~w32371 & ~w32373;
assign w32375 = w32184 & ~w32374;
assign w32376 = ~w32170 & w32185;
assign w32377 = w32215 & w32376;
assign w32378 = ~w32364 & ~w32377;
assign w32379 = ~w32375 & w32378;
assign w32380 = ~w32370 & w65984;
assign w32381 = (~pi1726 & w32370) | (~pi1726 & w65985) | (w32370 & w65985);
assign w32382 = ~w32380 & ~w32381;
assign w32383 = ~w32184 & w32224;
assign w32384 = ~w32192 & ~w32198;
assign w32385 = w32178 & ~w32384;
assign w32386 = w32168 & w32194;
assign w32387 = ~w32385 & ~w32386;
assign w32388 = w32184 & ~w32387;
assign w32389 = ~w32155 & w32232;
assign w32390 = ~w32178 & ~w32227;
assign w32391 = ~w32199 & ~w32218;
assign w32392 = w32185 & ~w32391;
assign w32393 = ~w32169 & w32363;
assign w32394 = ~w32383 & ~w32393;
assign w32395 = ~w32392 & w32394;
assign w32396 = ~w32389 & w32395;
assign w32397 = ~w32390 & w32396;
assign w32398 = ~w32388 & w32397;
assign w32399 = pi1729 & ~w32398;
assign w32400 = ~pi1729 & w32398;
assign w32401 = ~w32399 & ~w32400;
assign w32402 = w31864 & w31874;
assign w32403 = w31833 & ~w31871;
assign w32404 = ~w31882 & ~w31890;
assign w32405 = ~w32403 & w32404;
assign w32406 = ~w32402 & ~w32405;
assign w32407 = ~w31874 & ~w32018;
assign w32408 = ~w31827 & w31861;
assign w32409 = w32407 & w32408;
assign w32410 = w32406 & ~w32409;
assign w32411 = w31827 & ~w31888;
assign w32412 = ~w32410 & ~w32411;
assign w32413 = w31876 & ~w31898;
assign w32414 = (~w31839 & ~w32406) | (~w31839 & w65986) | (~w32406 & w65986);
assign w32415 = w31827 & ~w32413;
assign w32416 = ~w32414 & w32415;
assign w32417 = ~w32412 & ~w32416;
assign w32418 = ~pi1719 & w32417;
assign w32419 = pi1719 & ~w32417;
assign w32420 = ~w32418 & ~w32419;
assign w32421 = w31728 & ~w32276;
assign w32422 = ~w31704 & ~w32273;
assign w32423 = ~w31704 & ~w32292;
assign w32424 = ~w31706 & ~w31709;
assign w32425 = w31652 & ~w32423;
assign w32426 = ~w32424 & w32425;
assign w32427 = ~w31688 & w32251;
assign w32428 = ~w31674 & w31723;
assign w32429 = w31704 & ~w32427;
assign w32430 = ~w32428 & w32429;
assign w32431 = ~w32421 & ~w32426;
assign w32432 = ~w32430 & w32431;
assign w32433 = ~w32422 & w32432;
assign w32434 = pi1730 & ~w32433;
assign w32435 = ~pi1730 & w32433;
assign w32436 = ~w32434 & ~w32435;
assign w32437 = w31434 & w31452;
assign w32438 = w31424 & w31456;
assign w32439 = ~w31423 & ~w32438;
assign w32440 = w31425 & ~w31447;
assign w32441 = w31398 & ~w31404;
assign w32442 = ~w31379 & ~w32441;
assign w32443 = ~w31379 & w31428;
assign w32444 = w31392 & w31434;
assign w32445 = ~w31399 & w31416;
assign w32446 = ~w32444 & w32445;
assign w32447 = (~w32442 & w32443) | (~w32442 & w65987) | (w32443 & w65987);
assign w32448 = ~w31445 & ~w32440;
assign w32449 = ~w32447 & w32448;
assign w32450 = ~w32439 & ~w32449;
assign w32451 = w31399 & w31401;
assign w32452 = w31437 & ~w31443;
assign w32453 = w31424 & w65988;
assign w32454 = ~w31430 & ~w31436;
assign w32455 = w31379 & ~w31416;
assign w32456 = ~w31392 & ~w32455;
assign w32457 = ~w32454 & ~w32456;
assign w32458 = w31404 & w31447;
assign w32459 = ~w32451 & ~w32458;
assign w32460 = ~w32453 & w32459;
assign w32461 = ~w32452 & w32460;
assign w32462 = (~w31423 & ~w32461) | (~w31423 & w65989) | (~w32461 & w65989);
assign w32463 = ~w32437 & ~w32462;
assign w32464 = ~w32450 & w32463;
assign w32465 = pi1699 & ~w32464;
assign w32466 = ~pi1699 & w32464;
assign w32467 = ~w32465 & ~w32466;
assign w32468 = w31987 & w32079;
assign w32469 = w31959 & w31978;
assign w32470 = w31947 & w31985;
assign w32471 = w31939 & ~w32087;
assign w32472 = w31920 & w31989;
assign w32473 = ~w31939 & ~w32086;
assign w32474 = ~w32472 & w32473;
assign w32475 = ~w32471 & ~w32474;
assign w32476 = ~w31949 & ~w32469;
assign w32477 = ~w32470 & w32476;
assign w32478 = ~w32475 & w32477;
assign w32479 = ~w31958 & ~w32478;
assign w32480 = w31972 & ~w32076;
assign w32481 = w31920 & w31976;
assign w32482 = w31979 & ~w32075;
assign w32483 = w31971 & ~w31990;
assign w32484 = ~w32469 & w32483;
assign w32485 = ~w32481 & ~w32482;
assign w32486 = ~w32484 & w32485;
assign w32487 = w31958 & ~w32486;
assign w32488 = ~w31997 & ~w32480;
assign w32489 = ~w32487 & w32488;
assign w32490 = ~w32468 & w32489;
assign w32491 = (pi1717 & ~w32490) | (pi1717 & w65990) | (~w32490 & w65990);
assign w32492 = w32490 & w65991;
assign w32493 = ~w32491 & ~w32492;
assign w32494 = ~w31920 & w32469;
assign w32495 = ~w31927 & ~w31989;
assign w32496 = w31993 & ~w32495;
assign w32497 = ~w32494 & ~w32496;
assign w32498 = ~w32472 & ~w32497;
assign w32499 = w31926 & ~w31969;
assign w32500 = ~w32472 & ~w32499;
assign w32501 = w31939 & ~w32500;
assign w32502 = w31926 & w32481;
assign w32503 = ~w32501 & ~w32502;
assign w32504 = (~w31958 & w31996) | (~w31958 & w65992) | (w31996 & w65992);
assign w32505 = ~w31940 & ~w32481;
assign w32506 = w31994 & ~w32505;
assign w32507 = ~w31939 & w31941;
assign w32508 = ~w32073 & ~w32507;
assign w32509 = ~w31974 & w32508;
assign w32510 = (w31958 & ~w32509) | (w31958 & w65993) | (~w32509 & w65993);
assign w32511 = ~w32498 & ~w32510;
assign w32512 = ~w32504 & w32511;
assign w32513 = pi1704 & w32512;
assign w32514 = ~pi1704 & ~w32512;
assign w32515 = ~w32513 & ~w32514;
assign w32516 = ~w31898 & ~w31903;
assign w32517 = w31872 & ~w32516;
assign w32518 = ~w31897 & ~w32019;
assign w32519 = ~w31885 & w32518;
assign w32520 = ~w32517 & w32519;
assign w32521 = w31827 & ~w32520;
assign w32522 = ~w31839 & ~w31861;
assign w32523 = w31883 & w32522;
assign w32524 = ~w31827 & ~w31893;
assign w32525 = w31833 & ~w31867;
assign w32526 = w31827 & ~w32525;
assign w32527 = ~w32006 & ~w32017;
assign w32528 = w32404 & ~w32526;
assign w32529 = ~w32527 & w32528;
assign w32530 = ~w31908 & ~w32523;
assign w32531 = ~w32529 & w32530;
assign w32532 = ~w32524 & w32531;
assign w32533 = ~w32521 & w32532;
assign w32534 = pi1718 & w32533;
assign w32535 = ~pi1718 & ~w32533;
assign w32536 = ~w32534 & ~w32535;
assign w32537 = w31442 & w31456;
assign w32538 = w31392 & ~w31402;
assign w32539 = (~w31416 & w32538) | (~w31416 & w65994) | (w32538 & w65994);
assign w32540 = w31407 & w31416;
assign w32541 = w31402 & w32540;
assign w32542 = w31392 & ~w31398;
assign w32543 = w31379 & ~w32542;
assign w32544 = ~w32441 & w32543;
assign w32545 = ~w32451 & ~w32544;
assign w32546 = ~w32539 & w32545;
assign w32547 = ~w32541 & w32546;
assign w32548 = w31423 & ~w32547;
assign w32549 = w31409 & w31433;
assign w32550 = w31454 & ~w32543;
assign w32551 = w31450 & w32455;
assign w32552 = ~w31400 & ~w32458;
assign w32553 = ~w32551 & w32552;
assign w32554 = ~w32550 & w32553;
assign w32555 = ~w31423 & ~w32554;
assign w32556 = ~w31446 & ~w32537;
assign w32557 = ~w32549 & w32556;
assign w32558 = ~w32555 & w32557;
assign w32559 = ~w32548 & w32558;
assign w32560 = ~pi1713 & w32559;
assign w32561 = pi1713 & ~w32559;
assign w32562 = ~w32560 & ~w32561;
assign w32563 = ~w31632 & w32313;
assign w32564 = ~w31583 & w31631;
assign w32565 = w31631 & w65995;
assign w32566 = w31595 & ~w32565;
assign w32567 = (w31583 & w31632) | (w31583 & w65996) | (w31632 & w65996);
assign w32568 = (~w32567 & w32563) | (~w32567 & w65997) | (w32563 & w65997);
assign w32569 = w31603 & ~w32568;
assign w32570 = ~w31603 & ~w32564;
assign w32571 = ~w32567 & w32570;
assign w32572 = w31596 & ~w32571;
assign w32573 = ~w31589 & ~w32565;
assign w32574 = ~w31603 & ~w32573;
assign w32575 = ~w31595 & ~w32567;
assign w32576 = ~w32574 & w32575;
assign w32577 = ~w32572 & ~w32576;
assign w32578 = ~w32569 & ~w32577;
assign w32579 = ~pi1706 & w32578;
assign w32580 = pi1706 & ~w32578;
assign w32581 = ~w32579 & ~w32580;
assign w32582 = w32196 & w32211;
assign w32583 = w32184 & ~w32582;
assign w32584 = ~w32235 & ~w32583;
assign w32585 = ~w32189 & ~w32218;
assign w32586 = ~w32168 & w32585;
assign w32587 = w32235 & ~w32586;
assign w32588 = ~w32208 & w32587;
assign w32589 = w32156 & w32170;
assign w32590 = ~w32178 & ~w32589;
assign w32591 = (w32590 & ~w32208) | (w32590 & w65998) | (~w32208 & w65998);
assign w32592 = ~w32588 & w32591;
assign w32593 = ~w32168 & w32184;
assign w32594 = ~w32187 & ~w32593;
assign w32595 = w32585 & w32594;
assign w32596 = w32178 & ~w32595;
assign w32597 = ~w32212 & w32596;
assign w32598 = ~w32592 & ~w32597;
assign w32599 = ~w32584 & ~w32598;
assign w32600 = ~pi1733 & w32599;
assign w32601 = pi1733 & ~w32599;
assign w32602 = ~w32600 & ~w32601;
assign w32603 = (~w31595 & w31631) | (~w31595 & w65999) | (w31631 & w65999);
assign w32604 = w31586 & w32329;
assign w32605 = w31585 & w31615;
assign w32606 = w32316 & ~w32330;
assign w32607 = ~w32605 & w32606;
assign w32608 = w32603 & ~w32604;
assign w32609 = ~w32607 & w32608;
assign w32610 = ~w31624 & ~w32309;
assign w32611 = w31596 & w32610;
assign w32612 = ~w31630 & w32611;
assign w32613 = (w31603 & w32609) | (w31603 & w66000) | (w32609 & w66000);
assign w32614 = ~w31634 & ~w32330;
assign w32615 = ~w32563 & ~w32614;
assign w32616 = ~w31586 & w32603;
assign w32617 = ~w31603 & ~w32605;
assign w32618 = ~w31587 & w32617;
assign w32619 = ~w32616 & w32618;
assign w32620 = ~w32615 & w32619;
assign w32621 = ~w32613 & ~w32620;
assign w32622 = pi1705 & ~w32621;
assign w32623 = ~pi1705 & w32621;
assign w32624 = ~w32622 & ~w32623;
assign w32625 = ~w31473 & w31501;
assign w32626 = ~w32343 & ~w32625;
assign w32627 = w32121 & ~w32626;
assign w32628 = ~w32123 & ~w32627;
assign w32629 = ~w31524 & ~w32628;
assign w32630 = w31538 & w32340;
assign w32631 = ~w31515 & ~w32124;
assign w32632 = ~w31551 & w32631;
assign w32633 = ~w32630 & w32632;
assign w32634 = w31524 & ~w32633;
assign w32635 = w31487 & w32625;
assign w32636 = w31528 & ~w32635;
assign w32637 = w32132 & w32341;
assign w32638 = ~w31493 & ~w32349;
assign w32639 = ~w32637 & w32638;
assign w32640 = ~w32636 & ~w32639;
assign w32641 = ~w32634 & ~w32640;
assign w32642 = ~w32629 & w32641;
assign w32643 = ~pi1735 & w32642;
assign w32644 = pi1735 & ~w32642;
assign w32645 = ~w32643 & ~w32644;
assign w32646 = w31772 & ~w32038;
assign w32647 = ~w31772 & w31784;
assign w32648 = ~w32045 & w32647;
assign w32649 = ~w31807 & ~w32646;
assign w32650 = ~w32648 & w32649;
assign w32651 = w31745 & ~w32650;
assign w32652 = ~w31801 & ~w32061;
assign w32653 = w32057 & w32652;
assign w32654 = w31781 & ~w32652;
assign w32655 = ~w31806 & ~w32033;
assign w32656 = ~w32653 & w32655;
assign w32657 = ~w32654 & w32656;
assign w32658 = ~w31745 & ~w32657;
assign w32659 = w31765 & w31779;
assign w32660 = ~w32047 & ~w32659;
assign w32661 = ~w32658 & w32660;
assign w32662 = ~w32651 & w32661;
assign w32663 = pi1737 & w32662;
assign w32664 = ~pi1737 & ~w32662;
assign w32665 = ~w32663 & ~w32664;
assign w32666 = (~w31427 & ~w31454) | (~w31427 & w66001) | (~w31454 & w66001);
assign w32667 = w31408 & ~w32666;
assign w32668 = w31398 & ~w31401;
assign w32669 = ~w31429 & w32668;
assign w32670 = ~w32456 & w32669;
assign w32671 = w31423 & ~w32444;
assign w32672 = ~w32670 & w32671;
assign w32673 = ~w32667 & w32672;
assign w32674 = w31426 & ~w31457;
assign w32675 = ~w31423 & ~w32674;
assign w32676 = ~w32540 & w32675;
assign w32677 = ~w32673 & ~w32676;
assign w32678 = w31437 & w32544;
assign w32679 = ~w31405 & ~w31427;
assign w32680 = ~w32453 & w32679;
assign w32681 = w31432 & ~w32680;
assign w32682 = ~w32678 & ~w32681;
assign w32683 = ~w32677 & w32682;
assign w32684 = ~pi1720 & w32683;
assign w32685 = pi1720 & ~w32683;
assign w32686 = ~w32684 & ~w32685;
assign w32687 = ~pi5943 & pi9040;
assign w32688 = ~pi6012 & ~pi9040;
assign w32689 = ~w32687 & ~w32688;
assign w32690 = pi1732 & ~w32689;
assign w32691 = ~pi1732 & w32689;
assign w32692 = ~w32690 & ~w32691;
assign w32693 = ~pi5940 & pi9040;
assign w32694 = ~pi5909 & ~pi9040;
assign w32695 = ~w32693 & ~w32694;
assign w32696 = pi1754 & ~w32695;
assign w32697 = ~pi1754 & w32695;
assign w32698 = ~w32696 & ~w32697;
assign w32699 = ~w32692 & w32698;
assign w32700 = ~pi5824 & pi9040;
assign w32701 = ~pi5929 & ~pi9040;
assign w32702 = ~w32700 & ~w32701;
assign w32703 = pi1725 & ~w32702;
assign w32704 = ~pi1725 & w32702;
assign w32705 = ~w32703 & ~w32704;
assign w32706 = w32699 & w32705;
assign w32707 = ~pi5913 & pi9040;
assign w32708 = ~pi5945 & ~pi9040;
assign w32709 = ~w32707 & ~w32708;
assign w32710 = pi1756 & ~w32709;
assign w32711 = ~pi1756 & w32709;
assign w32712 = ~w32710 & ~w32711;
assign w32713 = ~w32705 & w32712;
assign w32714 = ~w32698 & w32713;
assign w32715 = ~w32706 & ~w32714;
assign w32716 = w32705 & ~w32712;
assign w32717 = w32698 & ~w32705;
assign w32718 = ~w32716 & ~w32717;
assign w32719 = ~w32692 & w32718;
assign w32720 = ~w32715 & ~w32719;
assign w32721 = ~w32692 & ~w32705;
assign w32722 = ~w32698 & ~w32712;
assign w32723 = w32712 & w32717;
assign w32724 = ~w32722 & ~w32723;
assign w32725 = w32721 & ~w32724;
assign w32726 = ~w32720 & ~w32725;
assign w32727 = ~pi5941 & pi9040;
assign w32728 = ~pi5938 & ~pi9040;
assign w32729 = ~w32727 & ~w32728;
assign w32730 = pi1738 & ~w32729;
assign w32731 = ~pi1738 & w32729;
assign w32732 = ~w32730 & ~w32731;
assign w32733 = ~w32726 & w32732;
assign w32734 = w32692 & ~w32732;
assign w32735 = w32705 & w32722;
assign w32736 = w32734 & w32735;
assign w32737 = w32692 & ~w32698;
assign w32738 = ~w32699 & ~w32737;
assign w32739 = ~w32732 & w32738;
assign w32740 = ~w32705 & w32739;
assign w32741 = w32732 & ~w32735;
assign w32742 = w32737 & ~w32741;
assign w32743 = w32716 & w32732;
assign w32744 = ~w32737 & ~w32743;
assign w32745 = ~w32742 & ~w32744;
assign w32746 = w32699 & w66002;
assign w32747 = ~pi5843 & pi9040;
assign w32748 = pi5835 & ~pi9040;
assign w32749 = ~w32747 & ~w32748;
assign w32750 = pi1742 & ~w32749;
assign w32751 = ~pi1742 & w32749;
assign w32752 = ~w32750 & ~w32751;
assign w32753 = ~w32746 & w32752;
assign w32754 = ~w32740 & w32753;
assign w32755 = ~w32745 & w32754;
assign w32756 = ~w32699 & ~w32712;
assign w32757 = (~w32732 & w32756) | (~w32732 & w63407) | (w32756 & w63407);
assign w32758 = w32698 & ~w32712;
assign w32759 = w32692 & ~w32705;
assign w32760 = w32758 & w32759;
assign w32761 = ~w32692 & w32713;
assign w32762 = w32732 & ~w32760;
assign w32763 = ~w32761 & w32762;
assign w32764 = ~w32757 & ~w32763;
assign w32765 = w32698 & w32712;
assign w32766 = w32692 & w32705;
assign w32767 = w32765 & w32766;
assign w32768 = ~w32752 & ~w32767;
assign w32769 = ~w32742 & w32768;
assign w32770 = ~w32764 & w32769;
assign w32771 = ~w32755 & ~w32770;
assign w32772 = ~w32733 & ~w32736;
assign w32773 = ~w32771 & w32772;
assign w32774 = ~pi1761 & w32773;
assign w32775 = pi1761 & ~w32773;
assign w32776 = ~w32774 & ~w32775;
assign w32777 = ~pi5921 & pi9040;
assign w32778 = ~pi5832 & ~pi9040;
assign w32779 = ~w32777 & ~w32778;
assign w32780 = pi1748 & ~w32779;
assign w32781 = ~pi1748 & w32779;
assign w32782 = ~w32780 & ~w32781;
assign w32783 = ~pi5823 & pi9040;
assign w32784 = ~pi5937 & ~pi9040;
assign w32785 = ~w32783 & ~w32784;
assign w32786 = pi1747 & ~w32785;
assign w32787 = ~pi1747 & w32785;
assign w32788 = ~w32786 & ~w32787;
assign w32789 = ~pi6080 & pi9040;
assign w32790 = ~pi5918 & ~pi9040;
assign w32791 = ~w32789 & ~w32790;
assign w32792 = pi1742 & ~w32791;
assign w32793 = ~pi1742 & w32791;
assign w32794 = ~w32792 & ~w32793;
assign w32795 = ~pi5923 & pi9040;
assign w32796 = ~pi6069 & ~pi9040;
assign w32797 = ~w32795 & ~w32796;
assign w32798 = pi1702 & ~w32797;
assign w32799 = ~pi1702 & w32797;
assign w32800 = ~w32798 & ~w32799;
assign w32801 = ~w32794 & ~w32800;
assign w32802 = ~pi5833 & pi9040;
assign w32803 = ~pi5921 & ~pi9040;
assign w32804 = ~w32802 & ~w32803;
assign w32805 = pi1758 & ~w32804;
assign w32806 = ~pi1758 & w32804;
assign w32807 = ~w32805 & ~w32806;
assign w32808 = w32788 & w32807;
assign w32809 = w32801 & w32808;
assign w32810 = ~pi5827 & pi9040;
assign w32811 = ~pi5840 & ~pi9040;
assign w32812 = ~w32810 & ~w32811;
assign w32813 = pi1756 & ~w32812;
assign w32814 = ~pi1756 & w32812;
assign w32815 = ~w32813 & ~w32814;
assign w32816 = w32794 & w32815;
assign w32817 = w32800 & w32807;
assign w32818 = w32788 & w32815;
assign w32819 = w32817 & ~w32818;
assign w32820 = ~w32788 & w32794;
assign w32821 = w32800 & ~w32815;
assign w32822 = w32820 & ~w32821;
assign w32823 = ~w32819 & ~w32822;
assign w32824 = ~w32816 & ~w32823;
assign w32825 = ~w32788 & ~w32800;
assign w32826 = ~w32794 & ~w32815;
assign w32827 = ~w32825 & w32826;
assign w32828 = ~w32807 & w32816;
assign w32829 = ~w32827 & ~w32828;
assign w32830 = ~w32809 & w32829;
assign w32831 = ~w32824 & w32830;
assign w32832 = w32809 & ~w32815;
assign w32833 = w32794 & w32807;
assign w32834 = ~w32788 & ~w32815;
assign w32835 = w32833 & w32834;
assign w32836 = w32815 & w32825;
assign w32837 = ~w32816 & ~w32826;
assign w32838 = w32800 & ~w32837;
assign w32839 = ~w32837 & w66003;
assign w32840 = ~w32836 & ~w32839;
assign w32841 = ~w32807 & ~w32840;
assign w32842 = w32788 & w32817;
assign w32843 = ~w32825 & ~w32842;
assign w32844 = ~w32794 & w32815;
assign w32845 = (w32844 & w32842) | (w32844 & w66004) | (w32842 & w66004);
assign w32846 = ~w32817 & ~w32821;
assign w32847 = w32820 & ~w32846;
assign w32848 = w32794 & w32800;
assign w32849 = ~w32801 & ~w32848;
assign w32850 = w32788 & ~w32837;
assign w32851 = w32849 & w32850;
assign w32852 = w32850 & w66005;
assign w32853 = ~w32807 & ~w32820;
assign w32854 = ~w32848 & w32853;
assign w32855 = ~w32818 & ~w32827;
assign w32856 = w32854 & w32855;
assign w32857 = ~w32845 & ~w32847;
assign w32858 = ~w32856 & w32857;
assign w32859 = ~w32852 & w32858;
assign w32860 = ~w32782 & ~w32859;
assign w32861 = ~w32832 & ~w32835;
assign w32862 = (w32861 & w32831) | (w32861 & w66006) | (w32831 & w66006);
assign w32863 = ~w32841 & w32862;
assign w32864 = ~w32860 & w32863;
assign w32865 = pi1764 & w32864;
assign w32866 = ~pi1764 & ~w32864;
assign w32867 = ~w32865 & ~w32866;
assign w32868 = ~w32831 & w32844;
assign w32869 = ~w32794 & ~w32834;
assign w32870 = w32834 & w32848;
assign w32871 = ~w32869 & ~w32870;
assign w32872 = w32807 & ~w32871;
assign w32873 = w32800 & w32818;
assign w32874 = w32782 & ~w32873;
assign w32875 = w32853 & ~w32869;
assign w32876 = w32816 & w32825;
assign w32877 = ~w32875 & ~w32876;
assign w32878 = ~w32872 & w32874;
assign w32879 = w32877 & w32878;
assign w32880 = ~w32800 & w32837;
assign w32881 = ~w32838 & ~w32880;
assign w32882 = w32833 & ~w32881;
assign w32883 = w32815 & ~w32825;
assign w32884 = ~w32807 & ~w32849;
assign w32885 = ~w32883 & w32884;
assign w32886 = (~w32782 & ~w32850) | (~w32782 & w66007) | (~w32850 & w66007);
assign w32887 = ~w32885 & w32886;
assign w32888 = ~w32882 & w32887;
assign w32889 = ~w32879 & ~w32888;
assign w32890 = ~w32868 & ~w32889;
assign w32891 = ~pi1770 & w32890;
assign w32892 = pi1770 & ~w32890;
assign w32893 = ~w32891 & ~w32892;
assign w32894 = ~pi5911 & pi9040;
assign w32895 = ~pi5923 & ~pi9040;
assign w32896 = ~w32894 & ~w32895;
assign w32897 = pi1702 & ~w32896;
assign w32898 = ~pi1702 & w32896;
assign w32899 = ~w32897 & ~w32898;
assign w32900 = ~pi5818 & pi9040;
assign w32901 = ~pi5948 & ~pi9040;
assign w32902 = ~w32900 & ~w32901;
assign w32903 = pi1752 & ~w32902;
assign w32904 = ~pi1752 & w32902;
assign w32905 = ~w32903 & ~w32904;
assign w32906 = w32899 & ~w32905;
assign w32907 = ~w32899 & w32905;
assign w32908 = ~pi6069 & pi9040;
assign w32909 = ~pi5818 & ~pi9040;
assign w32910 = ~w32908 & ~w32909;
assign w32911 = pi1755 & ~w32910;
assign w32912 = ~pi1755 & w32910;
assign w32913 = ~w32911 & ~w32912;
assign w32914 = w32907 & ~w32913;
assign w32915 = ~pi5836 & pi9040;
assign w32916 = ~pi5946 & ~pi9040;
assign w32917 = ~w32915 & ~w32916;
assign w32918 = pi1748 & ~w32917;
assign w32919 = ~pi1748 & w32917;
assign w32920 = ~w32918 & ~w32919;
assign w32921 = w32907 & w63887;
assign w32922 = ~w32906 & ~w32921;
assign w32923 = ~w32905 & ~w32920;
assign w32924 = w32913 & ~w32920;
assign w32925 = ~w32923 & ~w32924;
assign w32926 = ~pi5832 & pi9040;
assign w32927 = ~pi5823 & ~pi9040;
assign w32928 = ~w32926 & ~w32927;
assign w32929 = pi1736 & ~w32928;
assign w32930 = ~pi1736 & w32928;
assign w32931 = ~w32929 & ~w32930;
assign w32932 = w32925 & w32931;
assign w32933 = ~w32922 & w32932;
assign w32934 = ~w32899 & w32913;
assign w32935 = w32905 & w32920;
assign w32936 = w32934 & w32935;
assign w32937 = w32931 & w32936;
assign w32938 = w32899 & ~w32913;
assign w32939 = ~w32920 & w32934;
assign w32940 = ~w32938 & ~w32939;
assign w32941 = (~w32905 & w32939) | (~w32905 & w66008) | (w32939 & w66008);
assign w32942 = ~w32934 & ~w32935;
assign w32943 = w32905 & w32913;
assign w32944 = w32942 & w32943;
assign w32945 = ~w32905 & ~w32931;
assign w32946 = w32934 & w32945;
assign w32947 = ~w32944 & ~w32946;
assign w32948 = ~pi5819 & pi9040;
assign w32949 = ~pi5917 & ~pi9040;
assign w32950 = ~w32948 & ~w32949;
assign w32951 = pi1743 & ~w32950;
assign w32952 = ~pi1743 & w32950;
assign w32953 = ~w32951 & ~w32952;
assign w32954 = ~w32944 & w66009;
assign w32955 = w32920 & w32934;
assign w32956 = ~w32931 & ~w32955;
assign w32957 = ~w32942 & w32956;
assign w32958 = ~w32937 & ~w32941;
assign w32959 = ~w32957 & w32958;
assign w32960 = w32954 & w32959;
assign w32961 = w32899 & w32920;
assign w32962 = ~w32905 & w32913;
assign w32963 = w32961 & w32962;
assign w32964 = ~w32906 & ~w32961;
assign w32965 = w32931 & ~w32964;
assign w32966 = ~w32931 & ~w32934;
assign w32967 = ~w32899 & ~w32920;
assign w32968 = w32966 & w32967;
assign w32969 = w32905 & ~w32931;
assign w32970 = w32899 & ~w32969;
assign w32971 = ~w32907 & ~w32920;
assign w32972 = ~w32970 & w32971;
assign w32973 = ~w32947 & w32972;
assign w32974 = w32920 & ~w32934;
assign w32975 = ~w32924 & w32969;
assign w32976 = ~w32974 & w32975;
assign w32977 = ~w32899 & ~w32905;
assign w32978 = w32974 & w32977;
assign w32979 = w32953 & ~w32963;
assign w32980 = ~w32965 & w32979;
assign w32981 = ~w32968 & ~w32976;
assign w32982 = ~w32978 & w32981;
assign w32983 = w32980 & w32982;
assign w32984 = ~w32973 & w32983;
assign w32985 = (~w32933 & w32984) | (~w32933 & w66010) | (w32984 & w66010);
assign w32986 = ~pi1771 & w32985;
assign w32987 = pi1771 & ~w32985;
assign w32988 = ~w32986 & ~w32987;
assign w32989 = ~pi5929 & pi9040;
assign w32990 = ~pi5842 & ~pi9040;
assign w32991 = ~w32989 & ~w32990;
assign w32992 = pi1744 & ~w32991;
assign w32993 = ~pi1744 & w32991;
assign w32994 = ~w32992 & ~w32993;
assign w32995 = ~pi5842 & pi9040;
assign w32996 = ~pi5843 & ~pi9040;
assign w32997 = ~w32995 & ~w32996;
assign w32998 = pi1746 & ~w32997;
assign w32999 = ~pi1746 & w32997;
assign w33000 = ~w32998 & ~w32999;
assign w33001 = ~pi5938 & pi9040;
assign w33002 = ~pi5943 & ~pi9040;
assign w33003 = ~w33001 & ~w33002;
assign w33004 = pi1757 & ~w33003;
assign w33005 = ~pi1757 & w33003;
assign w33006 = ~w33004 & ~w33005;
assign w33007 = w33000 & w33006;
assign w33008 = ~pi5909 & pi9040;
assign w33009 = ~pi5913 & ~pi9040;
assign w33010 = ~w33008 & ~w33009;
assign w33011 = pi1724 & ~w33010;
assign w33012 = ~pi1724 & w33010;
assign w33013 = ~w33011 & ~w33012;
assign w33014 = ~w33006 & w33013;
assign w33015 = w33006 & ~w33013;
assign w33016 = ~w33014 & ~w33015;
assign w33017 = ~pi5945 & pi9040;
assign w33018 = ~pi5824 & ~pi9040;
assign w33019 = ~w33017 & ~w33018;
assign w33020 = pi1734 & ~w33019;
assign w33021 = ~pi1734 & w33019;
assign w33022 = ~w33020 & ~w33021;
assign w33023 = w33016 & w33022;
assign w33024 = w33007 & w33023;
assign w33025 = ~pi5837 & pi9040;
assign w33026 = ~pi5941 & ~pi9040;
assign w33027 = ~w33025 & ~w33026;
assign w33028 = pi1759 & ~w33027;
assign w33029 = ~pi1759 & w33027;
assign w33030 = ~w33028 & ~w33029;
assign w33031 = w33006 & ~w33030;
assign w33032 = ~w33000 & ~w33013;
assign w33033 = w33031 & w33032;
assign w33034 = w33022 & ~w33033;
assign w33035 = ~w33000 & w33006;
assign w33036 = (~w33022 & ~w33035) | (~w33022 & w66011) | (~w33035 & w66011);
assign w33037 = w33014 & ~w33030;
assign w33038 = w33036 & ~w33037;
assign w33039 = ~w33034 & ~w33038;
assign w33040 = w33000 & w33013;
assign w33041 = ~w33022 & w33040;
assign w33042 = w33040 & w66012;
assign w33043 = ~w33006 & ~w33030;
assign w33044 = w33000 & w33043;
assign w33045 = ~w33000 & ~w33006;
assign w33046 = ~w33007 & ~w33045;
assign w33047 = ~w33013 & w33030;
assign w33048 = ~w33046 & w33047;
assign w33049 = ~w33042 & ~w33044;
assign w33050 = ~w33048 & w33049;
assign w33051 = ~w33024 & w33050;
assign w33052 = ~w33039 & w33051;
assign w33053 = ~w32994 & ~w33052;
assign w33054 = ~w33006 & w33030;
assign w33055 = ~w33032 & ~w33040;
assign w33056 = w33054 & w33055;
assign w33057 = ~w33037 & ~w33048;
assign w33058 = w33000 & ~w33057;
assign w33059 = ~w33000 & ~w33054;
assign w33060 = w33016 & w33059;
assign w33061 = w32994 & w33060;
assign w33062 = w33022 & ~w33056;
assign w33063 = ~w33061 & w33062;
assign w33064 = ~w33058 & w33063;
assign w33065 = ~w33031 & ~w33056;
assign w33066 = w32994 & ~w33065;
assign w33067 = ~w33000 & w33030;
assign w33068 = w33015 & w33067;
assign w33069 = ~w33022 & ~w33068;
assign w33070 = ~w33066 & w33069;
assign w33071 = ~w33064 & ~w33070;
assign w33072 = ~w33053 & ~w33071;
assign w33073 = ~pi1768 & w33072;
assign w33074 = pi1768 & ~w33072;
assign w33075 = ~w33073 & ~w33074;
assign w33076 = ~w33031 & w33055;
assign w33077 = (~w33022 & ~w33055) | (~w33022 & w66013) | (~w33055 & w66013);
assign w33078 = w33043 & w33077;
assign w33079 = w33031 & w33055;
assign w33080 = (w33022 & ~w33043) | (w33022 & w66014) | (~w33043 & w66014);
assign w33081 = w33013 & ~w33030;
assign w33082 = w33000 & ~w33013;
assign w33083 = ~w33081 & ~w33082;
assign w33084 = w33016 & w33083;
assign w33085 = w33080 & ~w33084;
assign w33086 = ~w33007 & ~w33013;
assign w33087 = w33085 & ~w33086;
assign w33088 = w33041 & w33084;
assign w33089 = ~w33068 & ~w33079;
assign w33090 = ~w33088 & w33089;
assign w33091 = ~w33078 & w33090;
assign w33092 = (w32994 & ~w33091) | (w32994 & w66015) | (~w33091 & w66015);
assign w33093 = ~w33022 & w33056;
assign w33094 = w33031 & ~w33055;
assign w33095 = w33077 & ~w33094;
assign w33096 = (~w32994 & w33084) | (~w32994 & w66016) | (w33084 & w66016);
assign w33097 = ~w33095 & w33096;
assign w33098 = ~w33015 & w33067;
assign w33099 = w33022 & ~w33082;
assign w33100 = ~w33043 & w33099;
assign w33101 = ~w33015 & ~w33081;
assign w33102 = w33036 & ~w33101;
assign w33103 = ~w33023 & ~w33100;
assign w33104 = (~w33098 & ~w33103) | (~w33098 & w66017) | (~w33103 & w66017);
assign w33105 = ~w33076 & w33080;
assign w33106 = ~w33104 & w33105;
assign w33107 = ~w33093 & ~w33097;
assign w33108 = ~w33106 & w33107;
assign w33109 = ~w33092 & w33108;
assign w33110 = pi1779 & ~w33109;
assign w33111 = ~pi1779 & w33109;
assign w33112 = ~w33110 & ~w33111;
assign w33113 = w33031 & w33040;
assign w33114 = ~w33032 & ~w33054;
assign w33115 = w33046 & w33114;
assign w33116 = ~w33022 & ~w33115;
assign w33117 = w33016 & ~w33115;
assign w33118 = ~w33033 & w66018;
assign w33119 = ~w33117 & w33118;
assign w33120 = ~w33116 & ~w33119;
assign w33121 = (w32994 & w33120) | (w32994 & w66019) | (w33120 & w66019);
assign w33122 = ~w33057 & w33080;
assign w33123 = ~w33022 & ~w33045;
assign w33124 = ~w33040 & ~w33123;
assign w33125 = ~w33114 & ~w33124;
assign w33126 = ~w33030 & ~w33099;
assign w33127 = ~w33123 & w33126;
assign w33128 = ~w33125 & ~w33127;
assign w33129 = ~w32994 & ~w33128;
assign w33130 = w33067 & w33123;
assign w33131 = ~w33113 & ~w33130;
assign w33132 = ~w33122 & w33131;
assign w33133 = ~w33129 & w33132;
assign w33134 = ~w33121 & w33133;
assign w33135 = pi1763 & ~w33134;
assign w33136 = ~pi1763 & w33134;
assign w33137 = ~w33135 & ~w33136;
assign w33138 = w32935 & w32938;
assign w33139 = ~w32921 & ~w33138;
assign w33140 = w32943 & w32967;
assign w33141 = w32953 & ~w33140;
assign w33142 = ~w32939 & ~w32961;
assign w33143 = ~w32978 & w33142;
assign w33144 = ~w33141 & ~w33143;
assign w33145 = w33139 & ~w33144;
assign w33146 = ~w32931 & ~w33145;
assign w33147 = ~w32925 & w32966;
assign w33148 = w32932 & w33139;
assign w33149 = (~w32936 & w33148) | (~w32936 & w66020) | (w33148 & w66020);
assign w33150 = w33141 & ~w33147;
assign w33151 = ~w33149 & w33150;
assign w33152 = ~w32936 & ~w32953;
assign w33153 = w32931 & ~w32934;
assign w33154 = ~w32925 & w33153;
assign w33155 = w33152 & ~w33154;
assign w33156 = w33139 & w33155;
assign w33157 = ~w33151 & ~w33156;
assign w33158 = ~w33146 & ~w33157;
assign w33159 = ~pi1776 & w33158;
assign w33160 = pi1776 & ~w33158;
assign w33161 = ~w33159 & ~w33160;
assign w33162 = ~pi5796 & pi9040;
assign w33163 = ~pi5916 & ~pi9040;
assign w33164 = ~w33162 & ~w33163;
assign w33165 = pi1731 & ~w33164;
assign w33166 = ~pi1731 & w33164;
assign w33167 = ~w33165 & ~w33166;
assign w33168 = ~pi6013 & pi9040;
assign w33169 = ~pi5792 & ~pi9040;
assign w33170 = ~w33168 & ~w33169;
assign w33171 = pi1725 & ~w33170;
assign w33172 = ~pi1725 & w33170;
assign w33173 = ~w33171 & ~w33172;
assign w33174 = ~w33167 & ~w33173;
assign w33175 = ~pi5942 & pi9040;
assign w33176 = ~pi6015 & ~pi9040;
assign w33177 = ~w33175 & ~w33176;
assign w33178 = pi1741 & ~w33177;
assign w33179 = ~pi1741 & w33177;
assign w33180 = ~w33178 & ~w33179;
assign w33181 = ~pi6015 & pi9040;
assign w33182 = ~pi5796 & ~pi9040;
assign w33183 = ~w33181 & ~w33182;
assign w33184 = pi1753 & ~w33183;
assign w33185 = ~pi1753 & w33183;
assign w33186 = ~w33184 & ~w33185;
assign w33187 = w33180 & ~w33186;
assign w33188 = w33167 & ~w33173;
assign w33189 = ~w33167 & w33173;
assign w33190 = ~w33188 & ~w33189;
assign w33191 = w33187 & ~w33190;
assign w33192 = ~w33174 & ~w33191;
assign w33193 = ~pi5825 & pi9040;
assign w33194 = ~pi5939 & ~pi9040;
assign w33195 = ~w33193 & ~w33194;
assign w33196 = pi1728 & ~w33195;
assign w33197 = ~pi1728 & w33195;
assign w33198 = ~w33196 & ~w33197;
assign w33199 = w33174 & ~w33186;
assign w33200 = w33180 & w33199;
assign w33201 = w33198 & ~w33200;
assign w33202 = ~w33192 & w33201;
assign w33203 = ~w33167 & w33198;
assign w33204 = w33180 & w33186;
assign w33205 = ~w33180 & ~w33186;
assign w33206 = ~w33204 & ~w33205;
assign w33207 = w33167 & ~w33198;
assign w33208 = ~pi5835 & pi9040;
assign w33209 = pi5942 & ~pi9040;
assign w33210 = ~w33208 & ~w33209;
assign w33211 = pi1732 & ~w33210;
assign w33212 = ~pi1732 & w33210;
assign w33213 = ~w33211 & ~w33212;
assign w33214 = w33173 & w33213;
assign w33215 = ~w33207 & ~w33214;
assign w33216 = ~w33203 & ~w33206;
assign w33217 = ~w33215 & w33216;
assign w33218 = ~w33167 & ~w33180;
assign w33219 = ~w33173 & w33186;
assign w33220 = w33186 & w33198;
assign w33221 = ~w33219 & ~w33220;
assign w33222 = w33218 & ~w33221;
assign w33223 = ~w33188 & ~w33200;
assign w33224 = w33186 & w33189;
assign w33225 = w33189 & w33204;
assign w33226 = ~w33198 & ~w33225;
assign w33227 = w33173 & ~w33186;
assign w33228 = ~w33219 & ~w33227;
assign w33229 = w33218 & ~w33228;
assign w33230 = w33226 & ~w33229;
assign w33231 = ~w33186 & w33188;
assign w33232 = w33230 & ~w33231;
assign w33233 = w33213 & ~w33222;
assign w33234 = (w33233 & ~w33232) | (w33233 & w66021) | (~w33232 & w66021);
assign w33235 = w33187 & w33189;
assign w33236 = w33167 & w33227;
assign w33237 = ~w33224 & ~w33236;
assign w33238 = w33226 & ~w33237;
assign w33239 = w33173 & ~w33180;
assign w33240 = w33167 & ~w33239;
assign w33241 = ~w33218 & w33220;
assign w33242 = ~w33240 & w33241;
assign w33243 = ~w33186 & w33218;
assign w33244 = ~w33173 & w33243;
assign w33245 = ~w33213 & ~w33235;
assign w33246 = ~w33242 & w33245;
assign w33247 = ~w33244 & w33246;
assign w33248 = ~w33238 & w33247;
assign w33249 = ~w33234 & ~w33248;
assign w33250 = ~w33202 & ~w33217;
assign w33251 = ~w33249 & w33250;
assign w33252 = pi1765 & ~w33251;
assign w33253 = ~pi1765 & w33251;
assign w33254 = ~w33252 & ~w33253;
assign w33255 = ~pi5821 & pi9040;
assign w33256 = ~pi5947 & ~pi9040;
assign w33257 = ~w33255 & ~w33256;
assign w33258 = pi1724 & ~w33257;
assign w33259 = ~pi1724 & w33257;
assign w33260 = ~w33258 & ~w33259;
assign w33261 = ~pi6012 & pi9040;
assign w33262 = ~pi5825 & ~pi9040;
assign w33263 = ~w33261 & ~w33262;
assign w33264 = pi1709 & ~w33263;
assign w33265 = ~pi1709 & w33263;
assign w33266 = ~w33264 & ~w33265;
assign w33267 = ~pi5792 & pi9040;
assign w33268 = ~pi5831 & ~pi9040;
assign w33269 = ~w33267 & ~w33268;
assign w33270 = pi1744 & ~w33269;
assign w33271 = ~pi1744 & w33269;
assign w33272 = ~w33270 & ~w33271;
assign w33273 = ~w33266 & w33272;
assign w33274 = ~pi5920 & pi9040;
assign w33275 = ~pi6013 & ~pi9040;
assign w33276 = ~w33274 & ~w33275;
assign w33277 = pi1731 & ~w33276;
assign w33278 = ~pi1731 & w33276;
assign w33279 = ~w33277 & ~w33278;
assign w33280 = w33273 & ~w33279;
assign w33281 = ~w33260 & w33280;
assign w33282 = w33260 & ~w33266;
assign w33283 = ~pi5947 & pi9040;
assign w33284 = ~pi5940 & ~pi9040;
assign w33285 = ~w33283 & ~w33284;
assign w33286 = pi1749 & ~w33285;
assign w33287 = ~pi1749 & w33285;
assign w33288 = ~w33286 & ~w33287;
assign w33289 = w33279 & w33288;
assign w33290 = w33282 & w33289;
assign w33291 = ~pi5939 & pi9040;
assign w33292 = ~pi5816 & ~pi9040;
assign w33293 = ~w33291 & ~w33292;
assign w33294 = pi1753 & ~w33293;
assign w33295 = ~pi1753 & w33293;
assign w33296 = ~w33294 & ~w33295;
assign w33297 = ~w33266 & ~w33272;
assign w33298 = w33279 & w33297;
assign w33299 = ~w33260 & w33298;
assign w33300 = w33296 & ~w33299;
assign w33301 = ~w33282 & ~w33288;
assign w33302 = ~w33260 & ~w33272;
assign w33303 = w33266 & ~w33279;
assign w33304 = w33302 & w33303;
assign w33305 = ~w33301 & ~w33304;
assign w33306 = w33272 & ~w33279;
assign w33307 = w33266 & w33272;
assign w33308 = w33279 & ~w33307;
assign w33309 = ~w33306 & ~w33308;
assign w33310 = ~w33305 & w33309;
assign w33311 = w33260 & ~w33272;
assign w33312 = ~w33303 & w33311;
assign w33313 = w33260 & ~w33279;
assign w33314 = w33272 & w33313;
assign w33315 = w33313 & w33307;
assign w33316 = ~w33312 & ~w33315;
assign w33317 = w33288 & ~w33316;
assign w33318 = ~w33310 & ~w33317;
assign w33319 = ~w33260 & w33279;
assign w33320 = w33307 & w33319;
assign w33321 = w33273 & w63888;
assign w33322 = ~w33320 & ~w33321;
assign w33323 = w33300 & w33322;
assign w33324 = w33318 & w33323;
assign w33325 = w33266 & ~w33272;
assign w33326 = w33319 & w33325;
assign w33327 = ~w33302 & ~w33306;
assign w33328 = ~w33266 & w33327;
assign w33329 = (~w33288 & w33328) | (~w33288 & w66022) | (w33328 & w66022);
assign w33330 = ~w33279 & w33282;
assign w33331 = ~w33313 & ~w33319;
assign w33332 = w33325 & w33331;
assign w33333 = w33289 & w33302;
assign w33334 = ~w33330 & ~w33333;
assign w33335 = ~w33332 & w33334;
assign w33336 = ~w33298 & ~w33314;
assign w33337 = ~w33320 & w33336;
assign w33338 = w33336 & w63408;
assign w33339 = ~w33319 & w33335;
assign w33340 = w33338 & w33339;
assign w33341 = ~w33296 & ~w33326;
assign w33342 = ~w33329 & w33341;
assign w33343 = ~w33340 & w33342;
assign w33344 = ~w33281 & ~w33290;
assign w33345 = (w33344 & w33343) | (w33344 & w66023) | (w33343 & w66023);
assign w33346 = pi1760 & ~w33345;
assign w33347 = ~pi1760 & w33345;
assign w33348 = ~w33346 & ~w33347;
assign w33349 = w32801 & w32815;
assign w33350 = ~w32875 & ~w33349;
assign w33351 = ~w32854 & ~w33350;
assign w33352 = ~w32836 & ~w32848;
assign w33353 = ~w32843 & w33352;
assign w33354 = ~w32828 & ~w32873;
assign w33355 = ~w33353 & w33354;
assign w33356 = ~w33351 & w33355;
assign w33357 = ~w32782 & ~w33356;
assign w33358 = ~w32788 & ~w32829;
assign w33359 = ~w32877 & w33358;
assign w33360 = ~w32840 & w33351;
assign w33361 = ~w32847 & ~w32872;
assign w33362 = w32881 & ~w33361;
assign w33363 = w32854 & ~w32881;
assign w33364 = ~w32852 & ~w33363;
assign w33365 = ~w33362 & w33364;
assign w33366 = w32782 & ~w33365;
assign w33367 = ~w32835 & ~w33359;
assign w33368 = ~w33360 & w33367;
assign w33369 = ~w33357 & w33368;
assign w33370 = ~w33366 & w33369;
assign w33371 = pi1780 & w33370;
assign w33372 = ~pi1780 & ~w33370;
assign w33373 = ~w33371 & ~w33372;
assign w33374 = ~pi5815 & pi9040;
assign w33375 = ~pi6076 & ~pi9040;
assign w33376 = ~w33374 & ~w33375;
assign w33377 = pi1751 & ~w33376;
assign w33378 = ~pi1751 & w33376;
assign w33379 = ~w33377 & ~w33378;
assign w33380 = ~pi5937 & pi9040;
assign w33381 = ~pi5819 & ~pi9040;
assign w33382 = ~w33380 & ~w33381;
assign w33383 = pi1723 & ~w33382;
assign w33384 = ~pi1723 & w33382;
assign w33385 = ~w33383 & ~w33384;
assign w33386 = ~w33379 & w33385;
assign w33387 = ~pi5829 & pi9040;
assign w33388 = ~pi5838 & ~pi9040;
assign w33389 = ~w33387 & ~w33388;
assign w33390 = pi1745 & ~w33389;
assign w33391 = ~pi1745 & w33389;
assign w33392 = ~w33390 & ~w33391;
assign w33393 = w33386 & ~w33392;
assign w33394 = ~pi5948 & pi9040;
assign w33395 = ~pi5820 & ~pi9040;
assign w33396 = ~w33394 & ~w33395;
assign w33397 = pi1740 & ~w33396;
assign w33398 = ~pi1740 & w33396;
assign w33399 = ~w33397 & ~w33398;
assign w33400 = w33379 & w33399;
assign w33401 = ~pi5817 & pi9040;
assign w33402 = ~pi5815 & ~pi9040;
assign w33403 = ~w33401 & ~w33402;
assign w33404 = pi1746 & ~w33403;
assign w33405 = ~pi1746 & w33403;
assign w33406 = ~w33404 & ~w33405;
assign w33407 = w33385 & ~w33406;
assign w33408 = w33400 & w33407;
assign w33409 = ~w33385 & w33406;
assign w33410 = w33379 & ~w33392;
assign w33411 = w33409 & w33410;
assign w33412 = ~w33408 & ~w33411;
assign w33413 = ~w33393 & w33412;
assign w33414 = w33399 & w33406;
assign w33415 = ~w33413 & w33414;
assign w33416 = ~w33379 & ~w33399;
assign w33417 = ~w33385 & ~w33406;
assign w33418 = ~w33392 & w33417;
assign w33419 = w33379 & ~w33385;
assign w33420 = ~w33386 & ~w33419;
assign w33421 = ~w33406 & ~w33420;
assign w33422 = w33385 & w33406;
assign w33423 = w33392 & ~w33422;
assign w33424 = (~w33418 & w33421) | (~w33418 & w66024) | (w33421 & w66024);
assign w33425 = ~w33416 & ~w33424;
assign w33426 = w33379 & w33422;
assign w33427 = w33392 & w33426;
assign w33428 = ~w33416 & ~w33427;
assign w33429 = ~w33392 & w33406;
assign w33430 = w33416 & ~w33422;
assign w33431 = ~w33429 & w33430;
assign w33432 = w33392 & ~w33409;
assign w33433 = w33400 & w33432;
assign w33434 = ~w33431 & ~w33433;
assign w33435 = w33413 & w33434;
assign w33436 = ~w33428 & w33435;
assign w33437 = ~pi5822 & pi9040;
assign w33438 = ~pi5949 & ~pi9040;
assign w33439 = ~w33437 & ~w33438;
assign w33440 = pi1757 & ~w33439;
assign w33441 = ~pi1757 & w33439;
assign w33442 = ~w33440 & ~w33441;
assign w33443 = (w33442 & w33436) | (w33442 & w66025) | (w33436 & w66025);
assign w33444 = ~w33435 & ~w33442;
assign w33445 = ~w33421 & ~w33426;
assign w33446 = ~w33392 & ~w33399;
assign w33447 = ~w33445 & w33446;
assign w33448 = ~w33415 & ~w33447;
assign w33449 = ~w33444 & w33448;
assign w33450 = ~w33443 & w33449;
assign w33451 = pi1772 & ~w33450;
assign w33452 = ~pi1772 & w33450;
assign w33453 = ~w33451 & ~w33452;
assign w33454 = ~w32821 & ~w33349;
assign w33455 = w32820 & w32883;
assign w33456 = w32788 & w32881;
assign w33457 = w32881 & w63409;
assign w33458 = ~w32807 & ~w32816;
assign w33459 = w33454 & w33458;
assign w33460 = ~w33455 & ~w33459;
assign w33461 = ~w33457 & w33460;
assign w33462 = (~w32788 & ~w33461) | (~w32788 & w63889) | (~w33461 & w63889);
assign w33463 = w32782 & ~w33456;
assign w33464 = ~w33462 & w33463;
assign w33465 = ~w32828 & w32874;
assign w33466 = ~w33461 & ~w33465;
assign w33467 = ~w32851 & w33454;
assign w33468 = ~w32782 & w32807;
assign w33469 = ~w33467 & w33468;
assign w33470 = ~w33466 & ~w33469;
assign w33471 = ~w33464 & w33470;
assign w33472 = pi1769 & ~w33471;
assign w33473 = ~pi1769 & w33471;
assign w33474 = ~w33472 & ~w33473;
assign w33475 = ~w33273 & ~w33288;
assign w33476 = ~w33297 & ~w33330;
assign w33477 = ~w33475 & ~w33476;
assign w33478 = ~w33325 & w33475;
assign w33479 = w33260 & ~w33288;
assign w33480 = (w33479 & ~w33475) | (w33479 & w63890) | (~w33475 & w63890);
assign w33481 = ~w33260 & w33288;
assign w33482 = w33307 & w33481;
assign w33483 = ~w33333 & ~w33482;
assign w33484 = w33322 & w33483;
assign w33485 = ~w33477 & ~w33480;
assign w33486 = w33484 & w33485;
assign w33487 = w33266 & w33311;
assign w33488 = (~w33487 & ~w33339) | (~w33487 & w63410) | (~w33339 & w63410);
assign w33489 = w33486 & ~w33488;
assign w33490 = w33266 & ~w33327;
assign w33491 = w33273 & ~w33289;
assign w33492 = w33319 & w33491;
assign w33493 = w33260 & w33279;
assign w33494 = w33297 & w33493;
assign w33495 = ~w33490 & ~w33494;
assign w33496 = ~w33492 & w33495;
assign w33497 = (w33296 & w33489) | (w33296 & w63891) | (w33489 & w63891);
assign w33498 = w33272 & ~w33282;
assign w33499 = ~w33279 & w33311;
assign w33500 = ~w33498 & ~w33499;
assign w33501 = w33288 & ~w33500;
assign w33502 = ~w33272 & ~w33288;
assign w33503 = w33331 & w33502;
assign w33504 = ~w33501 & ~w33503;
assign w33505 = ~w33303 & w33309;
assign w33506 = ~w33504 & w33505;
assign w33507 = (~w33296 & ~w33485) | (~w33296 & w66026) | (~w33485 & w66026);
assign w33508 = ~w33476 & ~w33484;
assign w33509 = ~w33506 & ~w33508;
assign w33510 = ~w33507 & w33509;
assign w33511 = ~w33497 & w33510;
assign w33512 = pi1783 & w33511;
assign w33513 = ~pi1783 & ~w33511;
assign w33514 = ~w33512 & ~w33513;
assign w33515 = ~w33386 & ~w33418;
assign w33516 = ~w33379 & w33406;
assign w33517 = w33399 & ~w33516;
assign w33518 = ~w33393 & w33517;
assign w33519 = ~w33515 & w33518;
assign w33520 = ~w33411 & ~w33519;
assign w33521 = ~w33400 & ~w33520;
assign w33522 = ~w33392 & w33408;
assign w33523 = ~w33420 & w33446;
assign w33524 = w33392 & ~w33399;
assign w33525 = ~w33516 & ~w33524;
assign w33526 = ~w33379 & w33417;
assign w33527 = w33399 & w33409;
assign w33528 = ~w33526 & ~w33527;
assign w33529 = ~w33525 & ~w33528;
assign w33530 = w33412 & w33442;
assign w33531 = ~w33427 & ~w33523;
assign w33532 = w33530 & w33531;
assign w33533 = ~w33529 & w33532;
assign w33534 = w33407 & w33524;
assign w33535 = ~w33393 & ~w33400;
assign w33536 = w33422 & ~w33535;
assign w33537 = w33392 & w33399;
assign w33538 = w33419 & w33537;
assign w33539 = ~w33524 & w33526;
assign w33540 = w33392 & ~w33406;
assign w33541 = w33419 & w33540;
assign w33542 = ~w33399 & w33516;
assign w33543 = ~w33442 & ~w33534;
assign w33544 = ~w33538 & ~w33541;
assign w33545 = ~w33542 & w33544;
assign w33546 = ~w33539 & w33543;
assign w33547 = w33545 & w33546;
assign w33548 = ~w33536 & w33547;
assign w33549 = ~w33533 & ~w33548;
assign w33550 = ~w33521 & ~w33522;
assign w33551 = ~w33549 & w33550;
assign w33552 = pi1766 & ~w33551;
assign w33553 = ~pi1766 & w33551;
assign w33554 = ~w33552 & ~w33553;
assign w33555 = w33213 & ~w33225;
assign w33556 = ~w33180 & w33228;
assign w33557 = w33228 & w66027;
assign w33558 = ~w33200 & ~w33557;
assign w33559 = ~w33173 & ~w33558;
assign w33560 = ~w33229 & ~w33236;
assign w33561 = ~w33205 & ~w33560;
assign w33562 = ~w33190 & ~w33204;
assign w33563 = ~w33198 & ~w33562;
assign w33564 = w33203 & w33227;
assign w33565 = w33555 & ~w33564;
assign w33566 = ~w33563 & w33565;
assign w33567 = ~w33561 & w33566;
assign w33568 = ~w33559 & w33567;
assign w33569 = ~w33198 & w33235;
assign w33570 = ~w33180 & ~w33237;
assign w33571 = ~w33167 & ~w33204;
assign w33572 = ~w33192 & ~w33571;
assign w33573 = w33167 & w33186;
assign w33574 = ~w33244 & ~w33573;
assign w33575 = w33198 & ~w33574;
assign w33576 = ~w33213 & ~w33569;
assign w33577 = ~w33570 & w33576;
assign w33578 = ~w33572 & w33577;
assign w33579 = ~w33575 & w33578;
assign w33580 = ~w33568 & ~w33579;
assign w33581 = ~pi1774 & w33580;
assign w33582 = pi1774 & ~w33580;
assign w33583 = ~w33581 & ~w33582;
assign w33584 = ~w32963 & ~w33138;
assign w33585 = ~w32920 & w32938;
assign w33586 = ~w33140 & ~w33585;
assign w33587 = ~w32978 & w33586;
assign w33588 = (w33584 & w33587) | (w33584 & w66028) | (w33587 & w66028);
assign w33589 = ~w32931 & ~w33588;
assign w33590 = ~w32905 & w32924;
assign w33591 = w32954 & w33590;
assign w33592 = w32931 & ~w32953;
assign w33593 = ~w32924 & w33592;
assign w33594 = w33584 & w33593;
assign w33595 = w33587 & w33594;
assign w33596 = ~w32924 & ~w32977;
assign w33597 = ~w32962 & ~w33596;
assign w33598 = w32931 & ~w33597;
assign w33599 = ~w32914 & w32956;
assign w33600 = ~w33598 & ~w33599;
assign w33601 = w32923 & w32938;
assign w33602 = w33584 & ~w33601;
assign w33603 = w32947 & w33602;
assign w33604 = ~w33600 & w33603;
assign w33605 = w32953 & ~w33604;
assign w33606 = ~w33591 & ~w33595;
assign w33607 = ~w33589 & w33606;
assign w33608 = ~w33605 & w33607;
assign w33609 = pi1778 & ~w33608;
assign w33610 = ~pi1778 & w33608;
assign w33611 = ~w33609 & ~w33610;
assign w33612 = w33422 & w33446;
assign w33613 = ~w33528 & ~w33537;
assign w33614 = ~w33379 & w33399;
assign w33615 = ~w33429 & w33614;
assign w33616 = ~w33410 & ~w33615;
assign w33617 = w33385 & ~w33616;
assign w33618 = ~w33541 & ~w33612;
assign w33619 = ~w33613 & w33618;
assign w33620 = ~w33617 & w33619;
assign w33621 = ~w33442 & ~w33620;
assign w33622 = w33407 & ~w33410;
assign w33623 = ~w33411 & ~w33622;
assign w33624 = w33442 & ~w33623;
assign w33625 = w33392 & w33406;
assign w33626 = w33420 & w33625;
assign w33627 = ~w33539 & ~w33626;
assign w33628 = ~w33624 & w33627;
assign w33629 = w33393 & w33414;
assign w33630 = w33400 & w33417;
assign w33631 = ~w33626 & ~w33630;
assign w33632 = ~w33629 & w33631;
assign w33633 = w33442 & ~w33632;
assign w33634 = ~w33522 & ~w33538;
assign w33635 = (w33634 & w33628) | (w33634 & w66029) | (w33628 & w66029);
assign w33636 = ~w33633 & w33635;
assign w33637 = ~w33621 & w33636;
assign w33638 = pi1773 & ~w33637;
assign w33639 = ~pi1773 & w33637;
assign w33640 = ~w33638 & ~w33639;
assign w33641 = w33307 & w33493;
assign w33642 = ~w33296 & ~w33641;
assign w33643 = w33504 & w33642;
assign w33644 = ~w33282 & w33288;
assign w33645 = w33272 & ~w33479;
assign w33646 = ~w33644 & w33645;
assign w33647 = w33300 & ~w33646;
assign w33648 = w33335 & w33647;
assign w33649 = ~w33643 & ~w33648;
assign w33650 = ~w33492 & ~w33508;
assign w33651 = ~w33649 & w33650;
assign w33652 = pi1762 & ~w33651;
assign w33653 = ~pi1762 & w33651;
assign w33654 = ~w33652 & ~w33653;
assign w33655 = ~w33318 & w33644;
assign w33656 = (~w33288 & w33330) | (~w33288 & w66030) | (w33330 & w66030);
assign w33657 = w33266 & w33493;
assign w33658 = ~w33298 & ~w33491;
assign w33659 = w33328 & w33658;
assign w33660 = ~w33656 & ~w33657;
assign w33661 = ~w33659 & w33660;
assign w33662 = w33296 & ~w33661;
assign w33663 = ~w33313 & w33491;
assign w33664 = ~w33288 & ~w33326;
assign w33665 = ~w33499 & w33664;
assign w33666 = ~w33338 & ~w33665;
assign w33667 = ~w33663 & ~w33666;
assign w33668 = ~w33296 & ~w33667;
assign w33669 = w33337 & w33478;
assign w33670 = ~w33655 & ~w33669;
assign w33671 = ~w33662 & w33670;
assign w33672 = (pi1767 & ~w33671) | (pi1767 & w66031) | (~w33671 & w66031);
assign w33673 = w33671 & w66032;
assign w33674 = ~w33672 & ~w33673;
assign w33675 = w33537 & ~w33631;
assign w33676 = w33379 & ~w33407;
assign w33677 = ~w33432 & w33676;
assign w33678 = ~w33399 & ~w33677;
assign w33679 = w33420 & w33423;
assign w33680 = (~w33679 & w33678) | (~w33679 & w66033) | (w33678 & w66033);
assign w33681 = w33442 & ~w33680;
assign w33682 = w33379 & w33429;
assign w33683 = w33385 & ~w33540;
assign w33684 = ~w33614 & w33683;
assign w33685 = ~w33682 & w33684;
assign w33686 = w33520 & ~w33685;
assign w33687 = ~w33442 & ~w33686;
assign w33688 = ~w33399 & w33540;
assign w33689 = w33420 & w33688;
assign w33690 = ~w33675 & ~w33689;
assign w33691 = ~w33681 & w33690;
assign w33692 = ~w33687 & w33691;
assign w33693 = pi1784 & ~w33692;
assign w33694 = ~pi1784 & w33692;
assign w33695 = ~w33693 & ~w33694;
assign w33696 = ~w32721 & ~w32734;
assign w33697 = ~w32757 & ~w33696;
assign w33698 = w32752 & w32761;
assign w33699 = ~w33697 & ~w33698;
assign w33700 = ~w32698 & ~w33699;
assign w33701 = (w32734 & w32723) | (w32734 & w66034) | (w32723 & w66034);
assign w33702 = (w32699 & w32757) | (w32699 & w63892) | (w32757 & w63892);
assign w33703 = ~w32705 & ~w32737;
assign w33704 = w32756 & w33703;
assign w33705 = ~w33702 & ~w33704;
assign w33706 = ~w33702 & w66035;
assign w33707 = ~w32722 & w32732;
assign w33708 = ~w32717 & w33707;
assign w33709 = w32705 & ~w32765;
assign w33710 = ~w32738 & w33709;
assign w33711 = w33708 & ~w33710;
assign w33712 = w32752 & ~w33701;
assign w33713 = ~w33711 & w33712;
assign w33714 = ~w33706 & w33713;
assign w33715 = ~w32692 & ~w32732;
assign w33716 = w32716 & w33715;
assign w33717 = ~w32752 & ~w33716;
assign w33718 = ~w32718 & w32732;
assign w33719 = ~w32705 & w32732;
assign w33720 = ~w32698 & w32712;
assign w33721 = ~w33719 & w33720;
assign w33722 = (w32692 & w33718) | (w32692 & w66036) | (w33718 & w66036);
assign w33723 = w33717 & ~w33722;
assign w33724 = w33705 & w33723;
assign w33725 = ~w33714 & ~w33724;
assign w33726 = ~w33700 & ~w33725;
assign w33727 = ~pi1793 & w33726;
assign w33728 = pi1793 & ~w33726;
assign w33729 = ~w33727 & ~w33728;
assign w33730 = w32758 & w33719;
assign w33731 = w32692 & w32716;
assign w33732 = ~w32735 & ~w32766;
assign w33733 = w32732 & ~w33731;
assign w33734 = ~w33732 & w33733;
assign w33735 = ~w32719 & ~w33731;
assign w33736 = ~w32732 & ~w33735;
assign w33737 = ~w32714 & ~w32760;
assign w33738 = w32753 & w33737;
assign w33739 = ~w33734 & w33738;
assign w33740 = ~w33736 & w33739;
assign w33741 = w32765 & ~w33696;
assign w33742 = w32715 & ~w32765;
assign w33743 = w32741 & w33742;
assign w33744 = w33717 & ~w33741;
assign w33745 = ~w33743 & w33744;
assign w33746 = ~w33740 & ~w33745;
assign w33747 = w32720 & ~w32732;
assign w33748 = ~w32736 & ~w33730;
assign w33749 = ~w33747 & w33748;
assign w33750 = ~w33746 & w33749;
assign w33751 = pi1810 & w33750;
assign w33752 = ~pi1810 & ~w33750;
assign w33753 = ~w33751 & ~w33752;
assign w33754 = w33014 & w33067;
assign w33755 = w33034 & ~w33754;
assign w33756 = ~w33060 & ~w33079;
assign w33757 = (~w33022 & w33756) | (~w33022 & w66037) | (w33756 & w66037);
assign w33758 = ~w33755 & ~w33757;
assign w33759 = ~w32994 & ~w33104;
assign w33760 = w33023 & ~w33083;
assign w33761 = ~w33068 & ~w33113;
assign w33762 = ~w33042 & w33761;
assign w33763 = ~w33760 & w33762;
assign w33764 = w32994 & ~w33763;
assign w33765 = ~w33758 & ~w33764;
assign w33766 = ~w33759 & w33765;
assign w33767 = ~pi1795 & w33766;
assign w33768 = pi1795 & ~w33766;
assign w33769 = ~w33767 & ~w33768;
assign w33770 = w33198 & ~w33557;
assign w33771 = (~w33198 & ~w33187) | (~w33198 & w66038) | (~w33187 & w66038);
assign w33772 = w33167 & ~w33228;
assign w33773 = w33180 & w33219;
assign w33774 = ~w33243 & ~w33773;
assign w33775 = w33771 & w33774;
assign w33776 = ~w33772 & w33775;
assign w33777 = ~w33228 & w66039;
assign w33778 = ~w33225 & ~w33777;
assign w33779 = (w33778 & w33776) | (w33778 & w66040) | (w33776 & w66040);
assign w33780 = ~w33213 & ~w33779;
assign w33781 = w33555 & ~w33556;
assign w33782 = ~w33777 & w33781;
assign w33783 = w33201 & ~w33782;
assign w33784 = w33213 & ~w33558;
assign w33785 = ~w33198 & w33778;
assign w33786 = ~w33784 & w33785;
assign w33787 = ~w33783 & ~w33786;
assign w33788 = ~w33780 & ~w33787;
assign w33789 = ~pi1789 & w33788;
assign w33790 = pi1789 & ~w33788;
assign w33791 = ~w33789 & ~w33790;
assign w33792 = w33167 & w33239;
assign w33793 = ~w33773 & ~w33792;
assign w33794 = ~w33220 & ~w33573;
assign w33795 = w33793 & ~w33794;
assign w33796 = w33190 & w33230;
assign w33797 = ~w33191 & w33213;
assign w33798 = ~w33795 & w33797;
assign w33799 = ~w33796 & w33798;
assign w33800 = w33198 & ~w33199;
assign w33801 = w33793 & w33800;
assign w33802 = ~w33232 & ~w33801;
assign w33803 = w33198 & ~w33235;
assign w33804 = w33239 & w33573;
assign w33805 = w33771 & ~w33804;
assign w33806 = ~w33803 & ~w33805;
assign w33807 = w33167 & w33773;
assign w33808 = ~w33213 & ~w33807;
assign w33809 = ~w33806 & w33808;
assign w33810 = ~w33802 & w33809;
assign w33811 = ~w33799 & ~w33810;
assign w33812 = pi1788 & w33811;
assign w33813 = ~pi1788 & ~w33811;
assign w33814 = ~w33812 & ~w33813;
assign w33815 = ~pi5917 & pi9040;
assign w33816 = ~pi5836 & ~pi9040;
assign w33817 = ~w33815 & ~w33816;
assign w33818 = pi1723 & ~w33817;
assign w33819 = ~pi1723 & w33817;
assign w33820 = ~w33818 & ~w33819;
assign w33821 = ~pi6076 & pi9040;
assign w33822 = ~pi5827 & ~pi9040;
assign w33823 = ~w33821 & ~w33822;
assign w33824 = pi1750 & ~w33823;
assign w33825 = ~pi1750 & w33823;
assign w33826 = ~w33824 & ~w33825;
assign w33827 = ~pi5918 & pi9040;
assign w33828 = ~pi5833 & ~pi9040;
assign w33829 = ~w33827 & ~w33828;
assign w33830 = pi1755 & ~w33829;
assign w33831 = ~pi1755 & w33829;
assign w33832 = ~w33830 & ~w33831;
assign w33833 = ~w33826 & ~w33832;
assign w33834 = ~pi5828 & pi9040;
assign w33835 = ~pi5911 & ~pi9040;
assign w33836 = ~w33834 & ~w33835;
assign w33837 = pi1743 & ~w33836;
assign w33838 = ~pi1743 & w33836;
assign w33839 = ~w33837 & ~w33838;
assign w33840 = ~pi5946 & pi9040;
assign w33841 = ~pi5822 & ~pi9040;
assign w33842 = ~w33840 & ~w33841;
assign w33843 = pi1751 & ~w33842;
assign w33844 = ~pi1751 & w33842;
assign w33845 = ~w33843 & ~w33844;
assign w33846 = w33839 & ~w33845;
assign w33847 = w33833 & w33846;
assign w33848 = w33826 & w33839;
assign w33849 = w33832 & ~w33845;
assign w33850 = ~w33848 & ~w33849;
assign w33851 = ~w33832 & ~w33839;
assign w33852 = ~pi5838 & pi9040;
assign w33853 = ~pi5922 & ~pi9040;
assign w33854 = ~w33852 & ~w33853;
assign w33855 = pi1739 & ~w33854;
assign w33856 = ~pi1739 & w33854;
assign w33857 = ~w33855 & ~w33856;
assign w33858 = w33826 & ~w33845;
assign w33859 = w33832 & w33858;
assign w33860 = ~w33851 & w33857;
assign w33861 = ~w33859 & w33860;
assign w33862 = ~w33850 & w33861;
assign w33863 = ~w33845 & ~w33857;
assign w33864 = w33832 & w33839;
assign w33865 = ~w33851 & ~w33864;
assign w33866 = w33845 & ~w33865;
assign w33867 = ~w33839 & ~w33845;
assign w33868 = (~w33867 & w33865) | (~w33867 & w63411) | (w33865 & w63411);
assign w33869 = (w33826 & w33868) | (w33826 & w63893) | (w33868 & w63893);
assign w33870 = ~w33862 & ~w33869;
assign w33871 = ~w33839 & ~w33870;
assign w33872 = w33839 & w33863;
assign w33873 = (~w33826 & w33866) | (~w33826 & w66041) | (w33866 & w66041);
assign w33874 = ~w33847 & ~w33873;
assign w33875 = (w33820 & w33871) | (w33820 & w66042) | (w33871 & w66042);
assign w33876 = ~w33826 & w33845;
assign w33877 = ~w33858 & ~w33876;
assign w33878 = w33826 & w33857;
assign w33879 = ~w33847 & ~w33878;
assign w33880 = ~w33850 & ~w33864;
assign w33881 = ~w33879 & ~w33880;
assign w33882 = ~w33877 & w33881;
assign w33883 = ~w33832 & ~w33857;
assign w33884 = w33848 & w33883;
assign w33885 = ~w33857 & ~w33858;
assign w33886 = ~w33868 & w33885;
assign w33887 = w33833 & w33867;
assign w33888 = ~w33845 & ~w33864;
assign w33889 = (w33857 & w33864) | (w33857 & w66043) | (w33864 & w66043);
assign w33890 = (~w33887 & w33866) | (~w33887 & w66044) | (w33866 & w66044);
assign w33891 = ~w33886 & w33890;
assign w33892 = ~w33820 & ~w33891;
assign w33893 = ~w33882 & ~w33884;
assign w33894 = ~w33892 & w33893;
assign w33895 = ~w33875 & w33894;
assign w33896 = ~pi1777 & w33895;
assign w33897 = pi1777 & ~w33895;
assign w33898 = ~w33896 & ~w33897;
assign w33899 = w32920 & w32931;
assign w33900 = ~w32938 & ~w33899;
assign w33901 = ~w32923 & ~w32943;
assign w33902 = w33900 & w33901;
assign w33903 = w32931 & ~w32940;
assign w33904 = w32953 & ~w33902;
assign w33905 = ~w33903 & w33904;
assign w33906 = w32961 & ~w33900;
assign w33907 = ~w32941 & w33906;
assign w33908 = ~w32972 & ~w32978;
assign w33909 = w33152 & w33908;
assign w33910 = ~w33907 & w33909;
assign w33911 = ~w33905 & ~w33910;
assign w33912 = w32924 & w32966;
assign w33913 = ~w32943 & ~w33601;
assign w33914 = w33598 & ~w33913;
assign w33915 = ~w33912 & ~w33914;
assign w33916 = ~w33911 & w33915;
assign w33917 = pi1796 & ~w33916;
assign w33918 = ~pi1796 & w33916;
assign w33919 = ~w33917 & ~w33918;
assign w33920 = ~w32721 & ~w32746;
assign w33921 = w33708 & ~w33920;
assign w33922 = ~w32761 & w33732;
assign w33923 = ~w32739 & ~w33716;
assign w33924 = w33922 & ~w33923;
assign w33925 = w32732 & ~w33922;
assign w33926 = w32759 & ~w33707;
assign w33927 = ~w32752 & ~w33926;
assign w33928 = ~w33925 & w33927;
assign w33929 = (~w32723 & w32757) | (~w32723 & w66045) | (w32757 & w66045);
assign w33930 = w32752 & ~w33710;
assign w33931 = (w33930 & w32764) | (w33930 & w66046) | (w32764 & w66046);
assign w33932 = ~w33928 & ~w33931;
assign w33933 = ~w33921 & ~w33924;
assign w33934 = ~w33932 & w33933;
assign w33935 = ~pi1814 & ~w33934;
assign w33936 = pi1814 & w33934;
assign w33937 = ~w33935 & ~w33936;
assign w33938 = w33826 & w33832;
assign w33939 = w33886 & w33938;
assign w33940 = w33826 & ~w33839;
assign w33941 = w33845 & ~w33940;
assign w33942 = ~w33888 & ~w33941;
assign w33943 = ~w33839 & w33845;
assign w33944 = w33833 & ~w33943;
assign w33945 = ~w33846 & w33944;
assign w33946 = ~w33942 & ~w33945;
assign w33947 = ~w33820 & ~w33946;
assign w33948 = ~w33857 & w33947;
assign w33949 = ~w33839 & ~w33877;
assign w33950 = ~w33847 & ~w33949;
assign w33951 = w33861 & ~w33950;
assign w33952 = w33881 & ~w33949;
assign w33953 = ~w33846 & ~w33943;
assign w33954 = ~w33833 & ~w33953;
assign w33955 = ~w33857 & ~w33944;
assign w33956 = ~w33954 & w33955;
assign w33957 = w33857 & w33944;
assign w33958 = ~w33956 & ~w33957;
assign w33959 = ~w33952 & w33958;
assign w33960 = w33820 & ~w33959;
assign w33961 = ~w33839 & w33857;
assign w33962 = ~w33880 & ~w33961;
assign w33963 = ~w33820 & ~w33962;
assign w33964 = w33959 & w33963;
assign w33965 = ~w33939 & ~w33951;
assign w33966 = ~w33948 & w33965;
assign w33967 = ~w33960 & ~w33964;
assign w33968 = (pi1782 & ~w33967) | (pi1782 & w66047) | (~w33967 & w66047);
assign w33969 = w33967 & w66048;
assign w33970 = ~w33968 & ~w33969;
assign w33971 = (w33820 & w33949) | (w33820 & w66049) | (w33949 & w66049);
assign w33972 = ~w33832 & w33845;
assign w33973 = w33848 & w33972;
assign w33974 = ~w33971 & ~w33973;
assign w33975 = w33857 & ~w33974;
assign w33976 = ~w33851 & ~w33857;
assign w33977 = w33850 & w33976;
assign w33978 = (~w33820 & w33862) | (~w33820 & w66050) | (w33862 & w66050);
assign w33979 = ~w33832 & w33947;
assign w33980 = ~w33820 & ~w33863;
assign w33981 = w33938 & ~w33941;
assign w33982 = ~w33980 & w33981;
assign w33983 = w33820 & ~w33857;
assign w33984 = (~w33848 & w33850) | (~w33848 & w66051) | (w33850 & w66051);
assign w33985 = w33983 & ~w33984;
assign w33986 = ~w33982 & ~w33985;
assign w33987 = ~w33978 & w33986;
assign w33988 = ~w33979 & w33987;
assign w33989 = ~w33975 & w33988;
assign w33990 = pi1790 & ~w33989;
assign w33991 = ~pi1790 & w33989;
assign w33992 = ~w33990 & ~w33991;
assign w33993 = w33971 & w33981;
assign w33994 = ~w33942 & ~w33972;
assign w33995 = w33820 & ~w33994;
assign w33996 = ~w33832 & ~w33846;
assign w33997 = w33877 & w33996;
assign w33998 = ~w33995 & ~w33997;
assign w33999 = w33857 & ~w33998;
assign w34000 = ~w33953 & ~w33961;
assign w34001 = ~w33833 & ~w33938;
assign w34002 = ~w33942 & w34001;
assign w34003 = ~w34000 & ~w34002;
assign w34004 = w34000 & w34001;
assign w34005 = ~w33820 & ~w34004;
assign w34006 = ~w34003 & w34005;
assign w34007 = ~w33867 & w33983;
assign w34008 = w33994 & w34007;
assign w34009 = ~w33993 & ~w34008;
assign w34010 = ~w34006 & w34009;
assign w34011 = ~w33999 & w34010;
assign w34012 = pi1781 & ~w34011;
assign w34013 = ~pi1781 & w34011;
assign w34014 = ~w34012 & ~w34013;
assign w34015 = ~pi6031 & pi9040;
assign w34016 = ~pi6050 & ~pi9040;
assign w34017 = ~w34015 & ~w34016;
assign w34018 = pi1775 & ~w34017;
assign w34019 = ~pi1775 & w34017;
assign w34020 = ~w34018 & ~w34019;
assign w34021 = ~pi6063 & pi9040;
assign w34022 = ~pi6150 & ~pi9040;
assign w34023 = ~w34021 & ~w34022;
assign w34024 = pi1791 & ~w34023;
assign w34025 = ~pi1791 & w34023;
assign w34026 = ~w34024 & ~w34025;
assign w34027 = ~pi6257 & pi9040;
assign w34028 = ~pi6233 & ~pi9040;
assign w34029 = ~w34027 & ~w34028;
assign w34030 = pi1803 & ~w34029;
assign w34031 = ~pi1803 & w34029;
assign w34032 = ~w34030 & ~w34031;
assign w34033 = ~w34026 & w34032;
assign w34034 = ~pi6152 & pi9040;
assign w34035 = ~pi6027 & ~pi9040;
assign w34036 = ~w34034 & ~w34035;
assign w34037 = pi1817 & ~w34036;
assign w34038 = ~pi1817 & w34036;
assign w34039 = ~w34037 & ~w34038;
assign w34040 = ~pi6058 & pi9040;
assign w34041 = ~pi6168 & ~pi9040;
assign w34042 = ~w34040 & ~w34041;
assign w34043 = pi1815 & ~w34042;
assign w34044 = ~pi1815 & w34042;
assign w34045 = ~w34043 & ~w34044;
assign w34046 = w34039 & w34045;
assign w34047 = ~w34020 & w34032;
assign w34048 = w34046 & w34047;
assign w34049 = ~w34039 & ~w34045;
assign w34050 = (w34033 & w34048) | (w34033 & w66052) | (w34048 & w66052);
assign w34051 = w34020 & w34050;
assign w34052 = ~pi6148 & pi9040;
assign w34053 = ~pi6083 & ~pi9040;
assign w34054 = ~w34052 & ~w34053;
assign w34055 = pi1820 & ~w34054;
assign w34056 = ~pi1820 & w34054;
assign w34057 = ~w34055 & ~w34056;
assign w34058 = w34020 & w34045;
assign w34059 = ~w34026 & w34058;
assign w34060 = ~w34032 & ~w34045;
assign w34061 = ~w34026 & w34060;
assign w34062 = w34060 & w66053;
assign w34063 = w34020 & w34032;
assign w34064 = ~w34046 & ~w34049;
assign w34065 = w34063 & ~w34064;
assign w34066 = w34033 & ~w34039;
assign w34067 = ~w34059 & ~w34066;
assign w34068 = ~w34062 & w34067;
assign w34069 = ~w34065 & w34068;
assign w34070 = ~w34020 & w34026;
assign w34071 = w34032 & w34045;
assign w34072 = ~w34060 & ~w34071;
assign w34073 = ~w34049 & w34070;
assign w34074 = w34072 & w34073;
assign w34075 = w34068 & w66054;
assign w34076 = ~w34057 & ~w34075;
assign w34077 = ~w34020 & ~w34032;
assign w34078 = w34046 & w34077;
assign w34079 = ~w34020 & ~w34039;
assign w34080 = w34020 & w34039;
assign w34081 = ~w34071 & w34080;
assign w34082 = ~w34079 & ~w34081;
assign w34083 = (~w34078 & w34082) | (~w34078 & w66055) | (w34082 & w66055);
assign w34084 = w34026 & ~w34083;
assign w34085 = w34032 & w34039;
assign w34086 = ~w34032 & w34045;
assign w34087 = ~w34085 & ~w34086;
assign w34088 = ~w34063 & ~w34077;
assign w34089 = ~w34058 & ~w34088;
assign w34090 = w34087 & ~w34089;
assign w34091 = w34026 & ~w34081;
assign w34092 = (w34057 & w34090) | (w34057 & w66056) | (w34090 & w66056);
assign w34093 = ~w34084 & ~w34092;
assign w34094 = ~w34058 & ~w34085;
assign w34095 = w34039 & ~w34071;
assign w34096 = w34088 & w34095;
assign w34097 = ~w34094 & w34096;
assign w34098 = ~w34032 & w34079;
assign w34099 = ~w34026 & ~w34048;
assign w34100 = ~w34098 & w34099;
assign w34101 = ~w34097 & w34100;
assign w34102 = ~w34093 & ~w34101;
assign w34103 = ~w34051 & ~w34076;
assign w34104 = ~w34102 & w34103;
assign w34105 = ~pi1824 & w34104;
assign w34106 = pi1824 & ~w34104;
assign w34107 = ~w34105 & ~w34106;
assign w34108 = ~pi6153 & pi9040;
assign w34109 = ~pi6056 & ~pi9040;
assign w34110 = ~w34108 & ~w34109;
assign w34111 = pi1787 & ~w34110;
assign w34112 = ~pi1787 & w34110;
assign w34113 = ~w34111 & ~w34112;
assign w34114 = ~pi6225 & pi9040;
assign w34115 = ~pi6061 & ~pi9040;
assign w34116 = ~w34114 & ~w34115;
assign w34117 = pi1775 & ~w34116;
assign w34118 = ~pi1775 & w34116;
assign w34119 = ~w34117 & ~w34118;
assign w34120 = ~w34113 & ~w34119;
assign w34121 = ~pi6026 & pi9040;
assign w34122 = ~pi6225 & ~pi9040;
assign w34123 = ~w34121 & ~w34122;
assign w34124 = pi1813 & ~w34123;
assign w34125 = ~pi1813 & w34123;
assign w34126 = ~w34124 & ~w34125;
assign w34127 = ~pi6175 & pi9040;
assign w34128 = ~pi6174 & ~pi9040;
assign w34129 = ~w34127 & ~w34128;
assign w34130 = pi1802 & ~w34129;
assign w34131 = ~pi1802 & w34129;
assign w34132 = ~w34130 & ~w34131;
assign w34133 = ~w34126 & w34132;
assign w34134 = w34120 & w34133;
assign w34135 = ~pi6133 & pi9040;
assign w34136 = ~pi6066 & ~pi9040;
assign w34137 = ~w34135 & ~w34136;
assign w34138 = pi1819 & ~w34137;
assign w34139 = ~pi1819 & w34137;
assign w34140 = ~w34138 & ~w34139;
assign w34141 = ~w34134 & w34140;
assign w34142 = w34113 & w34119;
assign w34143 = w34133 & ~w34142;
assign w34144 = ~w34120 & ~w34143;
assign w34145 = w34141 & ~w34144;
assign w34146 = ~w34113 & ~w34132;
assign w34147 = ~w34119 & w34126;
assign w34148 = w34126 & w34140;
assign w34149 = ~w34147 & ~w34148;
assign w34150 = w34146 & ~w34149;
assign w34151 = ~w34113 & w34140;
assign w34152 = w34126 & ~w34132;
assign w34153 = ~w34133 & ~w34152;
assign w34154 = w34119 & ~w34151;
assign w34155 = w34153 & w34154;
assign w34156 = w34113 & w34147;
assign w34157 = ~w34134 & ~w34156;
assign w34158 = ~w34140 & ~w34157;
assign w34159 = ~pi6061 & pi9040;
assign w34160 = ~pi6049 & ~pi9040;
assign w34161 = ~w34159 & ~w34160;
assign w34162 = pi1803 & ~w34161;
assign w34163 = ~pi1803 & w34161;
assign w34164 = ~w34162 & ~w34163;
assign w34165 = ~w34150 & ~w34164;
assign w34166 = ~w34155 & w34165;
assign w34167 = ~w34158 & w34166;
assign w34168 = ~w34113 & w34132;
assign w34169 = w34119 & ~w34126;
assign w34170 = w34168 & w34169;
assign w34171 = ~w34132 & w34142;
assign w34172 = ~w34168 & ~w34171;
assign w34173 = (w34148 & w34171) | (w34148 & w66057) | (w34171 & w66057);
assign w34174 = w34113 & ~w34126;
assign w34175 = w34119 & w34126;
assign w34176 = ~w34113 & w34175;
assign w34177 = ~w34132 & w34176;
assign w34178 = ~w34174 & ~w34177;
assign w34179 = ~w34147 & ~w34169;
assign w34180 = ~w34120 & ~w34142;
assign w34181 = ~w34146 & w34180;
assign w34182 = (~w34140 & ~w34181) | (~w34140 & w63894) | (~w34181 & w63894);
assign w34183 = ~w34178 & w34182;
assign w34184 = ~w34119 & ~w34152;
assign w34185 = ~w34174 & w34184;
assign w34186 = ~w34132 & w34185;
assign w34187 = w34164 & ~w34170;
assign w34188 = ~w34173 & w34187;
assign w34189 = ~w34186 & w34188;
assign w34190 = ~w34183 & w34189;
assign w34191 = ~w34167 & ~w34190;
assign w34192 = w34113 & ~w34140;
assign w34193 = w34153 & w34192;
assign w34194 = ~w34145 & ~w34193;
assign w34195 = ~w34191 & w34194;
assign w34196 = pi1826 & ~w34195;
assign w34197 = ~pi1826 & w34195;
assign w34198 = ~w34196 & ~w34197;
assign w34199 = w34126 & w34132;
assign w34200 = w34120 & w34199;
assign w34201 = w34140 & w34186;
assign w34202 = w34140 & ~w34171;
assign w34203 = ~w34185 & w34202;
assign w34204 = w34169 & ~w34172;
assign w34205 = ~w34203 & w34204;
assign w34206 = ~w34143 & ~w34148;
assign w34207 = w34113 & ~w34206;
assign w34208 = w34164 & ~w34200;
assign w34209 = ~w34177 & w34208;
assign w34210 = ~w34207 & w34209;
assign w34211 = ~w34201 & w34210;
assign w34212 = ~w34205 & w34211;
assign w34213 = (w34140 & ~w34175) | (w34140 & w66058) | (~w34175 & w66058);
assign w34214 = w34199 & ~w34213;
assign w34215 = (~w34140 & ~w34174) | (~w34140 & w66059) | (~w34174 & w66059);
assign w34216 = ~w34155 & w34169;
assign w34217 = ~w34215 & w34216;
assign w34218 = w34146 & ~w34179;
assign w34219 = ~w34132 & w34179;
assign w34220 = w34179 & w66060;
assign w34221 = ~w34218 & ~w34220;
assign w34222 = ~w34119 & ~w34221;
assign w34223 = ~w34141 & ~w34180;
assign w34224 = ~w34164 & ~w34214;
assign w34225 = ~w34223 & w34224;
assign w34226 = ~w34217 & w34225;
assign w34227 = ~w34222 & w34226;
assign w34228 = ~w34212 & ~w34227;
assign w34229 = pi1828 & w34228;
assign w34230 = ~pi1828 & ~w34228;
assign w34231 = ~w34229 & ~w34230;
assign w34232 = w34026 & ~w34079;
assign w34233 = w34020 & ~w34039;
assign w34234 = w34071 & w34233;
assign w34235 = (~w34234 & w34090) | (~w34234 & w66061) | (w34090 & w66061);
assign w34236 = ~w34232 & ~w34235;
assign w34237 = w34045 & w34079;
assign w34238 = w34020 & ~w34087;
assign w34239 = (w34026 & w34238) | (w34026 & w66062) | (w34238 & w66062);
assign w34240 = w34064 & w34089;
assign w34241 = ~w34050 & ~w34240;
assign w34242 = (w34057 & ~w34241) | (w34057 & w66063) | (~w34241 & w66063);
assign w34243 = w34020 & w34061;
assign w34244 = ~w34078 & ~w34243;
assign w34245 = ~w34026 & ~w34244;
assign w34246 = ~w34066 & ~w34098;
assign w34247 = ~w34072 & ~w34246;
assign w34248 = w34032 & ~w34058;
assign w34249 = w34232 & w34248;
assign w34250 = ~w34096 & ~w34234;
assign w34251 = ~w34249 & w34250;
assign w34252 = ~w34247 & w34251;
assign w34253 = (~w34057 & ~w34252) | (~w34057 & w66064) | (~w34252 & w66064);
assign w34254 = ~w34236 & ~w34242;
assign w34255 = ~w34253 & w34254;
assign w34256 = ~pi1850 & w34255;
assign w34257 = pi1850 & ~w34255;
assign w34258 = ~w34256 & ~w34257;
assign w34259 = ~pi6057 & pi9040;
assign w34260 = ~pi6153 & ~pi9040;
assign w34261 = ~w34259 & ~w34260;
assign w34262 = pi1818 & ~w34261;
assign w34263 = ~pi1818 & w34261;
assign w34264 = ~w34262 & ~w34263;
assign w34265 = ~pi6050 & pi9040;
assign w34266 = ~pi6058 & ~pi9040;
assign w34267 = ~w34265 & ~w34266;
assign w34268 = pi1792 & ~w34267;
assign w34269 = ~pi1792 & w34267;
assign w34270 = ~w34268 & ~w34269;
assign w34271 = w34264 & ~w34270;
assign w34272 = ~pi6174 & pi9040;
assign w34273 = ~pi6148 & ~pi9040;
assign w34274 = ~w34272 & ~w34273;
assign w34275 = pi1787 & ~w34274;
assign w34276 = ~pi1787 & w34274;
assign w34277 = ~w34275 & ~w34276;
assign w34278 = ~pi6150 & pi9040;
assign w34279 = ~pi6067 & ~pi9040;
assign w34280 = ~w34278 & ~w34279;
assign w34281 = pi1809 & ~w34280;
assign w34282 = ~pi1809 & w34280;
assign w34283 = ~w34281 & ~w34282;
assign w34284 = w34277 & w34283;
assign w34285 = w34271 & w34284;
assign w34286 = ~pi6056 & pi9040;
assign w34287 = ~pi6175 & ~pi9040;
assign w34288 = ~w34286 & ~w34287;
assign w34289 = pi1799 & ~w34288;
assign w34290 = ~pi1799 & w34288;
assign w34291 = ~w34289 & ~w34290;
assign w34292 = ~w34264 & ~w34291;
assign w34293 = w34270 & w34277;
assign w34294 = ~w34270 & ~w34277;
assign w34295 = ~w34291 & w34294;
assign w34296 = ~w34293 & ~w34295;
assign w34297 = ~w34295 & w63895;
assign w34298 = ~w34283 & w34291;
assign w34299 = w34294 & w34298;
assign w34300 = ~w34264 & w34291;
assign w34301 = w34293 & w34300;
assign w34302 = ~w34299 & ~w34301;
assign w34303 = ~w34297 & w34302;
assign w34304 = w34264 & w34291;
assign w34305 = ~w34277 & w34304;
assign w34306 = w34304 & w63896;
assign w34307 = w34283 & ~w34306;
assign w34308 = w34264 & ~w34291;
assign w34309 = ~w34277 & ~w34291;
assign w34310 = ~w34271 & w34309;
assign w34311 = w34308 & ~w34310;
assign w34312 = w34307 & ~w34311;
assign w34313 = ~w34283 & ~w34310;
assign w34314 = w34291 & w34293;
assign w34315 = w34313 & ~w34314;
assign w34316 = ~w34312 & ~w34315;
assign w34317 = ~pi6081 & pi9040;
assign w34318 = ~pi6031 & ~pi9040;
assign w34319 = ~w34317 & ~w34318;
assign w34320 = pi1813 & ~w34319;
assign w34321 = ~pi1813 & w34319;
assign w34322 = ~w34320 & ~w34321;
assign w34323 = (w34322 & w34316) | (w34322 & w66065) | (w34316 & w66065);
assign w34324 = w34294 & w34300;
assign w34325 = w34277 & w34291;
assign w34326 = ~w34308 & ~w34325;
assign w34327 = ~w34270 & ~w34326;
assign w34328 = (~w34283 & w34327) | (~w34283 & w66066) | (w34327 & w66066);
assign w34329 = w34277 & ~w34304;
assign w34330 = ~w34300 & ~w34325;
assign w34331 = ~w34329 & ~w34330;
assign w34332 = ~w34310 & ~w34331;
assign w34333 = w34264 & w34309;
assign w34334 = ~w34308 & ~w34309;
assign w34335 = (w34270 & ~w34309) | (w34270 & w66067) | (~w34309 & w66067);
assign w34336 = ~w34334 & w34335;
assign w34337 = w34307 & ~w34336;
assign w34338 = ~w34332 & w34337;
assign w34339 = w34292 & w34293;
assign w34340 = ~w34328 & ~w34339;
assign w34341 = ~w34338 & w34340;
assign w34342 = ~w34322 & ~w34341;
assign w34343 = ~w34285 & ~w34324;
assign w34344 = ~w34323 & w34343;
assign w34345 = ~w34342 & w34344;
assign w34346 = pi1836 & ~w34345;
assign w34347 = ~pi1836 & w34345;
assign w34348 = ~w34346 & ~w34347;
assign w34349 = ~w34069 & ~w34083;
assign w34350 = ~w34020 & ~w34045;
assign w34351 = w34232 & w34350;
assign w34352 = w34020 & w34072;
assign w34353 = (~w34026 & w34352) | (~w34026 & w66068) | (w34352 & w66068);
assign w34354 = ~w34049 & w34088;
assign w34355 = w34026 & ~w34350;
assign w34356 = ~w34047 & ~w34355;
assign w34357 = ~w34354 & ~w34356;
assign w34358 = ~w34072 & w34357;
assign w34359 = w34057 & ~w34237;
assign w34360 = ~w34097 & w34359;
assign w34361 = ~w34353 & w34360;
assign w34362 = ~w34358 & w34361;
assign w34363 = w34094 & ~w34350;
assign w34364 = w34026 & ~w34046;
assign w34365 = ~w34363 & w34364;
assign w34366 = w34033 & w34046;
assign w34367 = ~w34057 & ~w34366;
assign w34368 = w34244 & w34367;
assign w34369 = ~w34365 & w34368;
assign w34370 = ~w34362 & ~w34369;
assign w34371 = ~w34051 & ~w34351;
assign w34372 = ~w34349 & w34371;
assign w34373 = ~w34370 & w66069;
assign w34374 = (pi1863 & w34370) | (pi1863 & w66070) | (w34370 & w66070);
assign w34375 = ~w34373 & ~w34374;
assign w34376 = ~pi6066 & pi9040;
assign w34377 = ~pi6257 & ~pi9040;
assign w34378 = ~w34376 & ~w34377;
assign w34379 = pi1786 & ~w34378;
assign w34380 = ~pi1786 & w34378;
assign w34381 = ~w34379 & ~w34380;
assign w34382 = ~pi6027 & pi9040;
assign w34383 = ~pi6057 & ~pi9040;
assign w34384 = ~w34382 & ~w34383;
assign w34385 = pi1822 & ~w34384;
assign w34386 = ~pi1822 & w34384;
assign w34387 = ~w34385 & ~w34386;
assign w34388 = ~pi6233 & pi9040;
assign w34389 = ~pi6063 & ~pi9040;
assign w34390 = ~w34388 & ~w34389;
assign w34391 = pi1818 & ~w34390;
assign w34392 = ~pi1818 & w34390;
assign w34393 = ~w34391 & ~w34392;
assign w34394 = w34387 & ~w34393;
assign w34395 = ~pi6169 & pi9040;
assign w34396 = ~pi6081 & ~pi9040;
assign w34397 = ~w34395 & ~w34396;
assign w34398 = pi1798 & ~w34397;
assign w34399 = ~pi1798 & w34397;
assign w34400 = ~w34398 & ~w34399;
assign w34401 = ~pi6168 & pi9040;
assign w34402 = ~pi6152 & ~pi9040;
assign w34403 = ~w34401 & ~w34402;
assign w34404 = pi1805 & ~w34403;
assign w34405 = ~pi1805 & w34403;
assign w34406 = ~w34404 & ~w34405;
assign w34407 = ~w34400 & w34406;
assign w34408 = w34400 & ~w34406;
assign w34409 = ~w34407 & ~w34408;
assign w34410 = w34394 & w34409;
assign w34411 = ~pi6065 & pi9040;
assign w34412 = ~pi6133 & ~pi9040;
assign w34413 = ~w34411 & ~w34412;
assign w34414 = pi1799 & ~w34413;
assign w34415 = ~pi1799 & w34413;
assign w34416 = ~w34414 & ~w34415;
assign w34417 = ~w34410 & ~w34416;
assign w34418 = w34393 & w34406;
assign w34419 = w34400 & w34418;
assign w34420 = ~w34393 & ~w34400;
assign w34421 = ~w34387 & w34420;
assign w34422 = ~w34419 & ~w34421;
assign w34423 = ~w34400 & ~w34406;
assign w34424 = ~w34394 & ~w34423;
assign w34425 = ~w34420 & ~w34424;
assign w34426 = w34422 & ~w34423;
assign w34427 = ~w34425 & w34426;
assign w34428 = w34381 & ~w34417;
assign w34429 = ~w34427 & w34428;
assign w34430 = ~w34387 & w34400;
assign w34431 = w34418 & w34430;
assign w34432 = ~w34387 & ~w34406;
assign w34433 = ~w34387 & w34408;
assign w34434 = (w34381 & ~w34408) | (w34381 & w34868) | (~w34408 & w34868);
assign w34435 = w34387 & w34393;
assign w34436 = ~w34393 & ~w34406;
assign w34437 = ~w34435 & ~w34436;
assign w34438 = ~w34406 & ~w34420;
assign w34439 = ~w34437 & ~w34438;
assign w34440 = w34434 & ~w34439;
assign w34441 = w34432 & w34440;
assign w34442 = ~w34381 & w34387;
assign w34443 = w34407 & w34442;
assign w34444 = ~w34393 & w34406;
assign w34445 = ~w34432 & ~w34444;
assign w34446 = ~w34381 & ~w34400;
assign w34447 = ~w34445 & w34446;
assign w34448 = ~w34435 & ~w34442;
assign w34449 = w34408 & ~w34448;
assign w34450 = ~w34387 & ~w34393;
assign w34451 = w34381 & ~w34420;
assign w34452 = w34450 & w34451;
assign w34453 = ~w34416 & ~w34447;
assign w34454 = ~w34449 & ~w34452;
assign w34455 = w34453 & w34454;
assign w34456 = w34400 & ~w34450;
assign w34457 = w34437 & w34456;
assign w34458 = w34393 & w34407;
assign w34459 = ~w34433 & ~w34458;
assign w34460 = ~w34381 & ~w34459;
assign w34461 = w34416 & ~w34457;
assign w34462 = ~w34460 & w34461;
assign w34463 = ~w34455 & ~w34462;
assign w34464 = ~w34431 & ~w34443;
assign w34465 = ~w34441 & w34464;
assign w34466 = ~w34429 & w34465;
assign w34467 = ~w34463 & w34466;
assign w34468 = pi1830 & ~w34467;
assign w34469 = ~pi1830 & w34467;
assign w34470 = ~w34468 & ~w34469;
assign w34471 = ~pi6147 & pi9040;
assign w34472 = ~pi6159 & ~pi9040;
assign w34473 = ~w34471 & ~w34472;
assign w34474 = pi1804 & ~w34473;
assign w34475 = ~pi1804 & w34473;
assign w34476 = ~w34474 & ~w34475;
assign w34477 = ~pi6176 & pi9040;
assign w34478 = ~pi6078 & ~pi9040;
assign w34479 = ~w34477 & ~w34478;
assign w34480 = pi1812 & ~w34479;
assign w34481 = ~pi1812 & w34479;
assign w34482 = ~w34480 & ~w34481;
assign w34483 = ~pi6143 & pi9040;
assign w34484 = ~pi6294 & ~pi9040;
assign w34485 = ~w34483 & ~w34484;
assign w34486 = pi1794 & ~w34485;
assign w34487 = ~pi1794 & w34485;
assign w34488 = ~w34486 & ~w34487;
assign w34489 = ~w34482 & w34488;
assign w34490 = ~pi6082 & pi9040;
assign w34491 = ~pi6064 & ~pi9040;
assign w34492 = ~w34490 & ~w34491;
assign w34493 = pi1811 & ~w34492;
assign w34494 = ~pi1811 & w34492;
assign w34495 = ~w34493 & ~w34494;
assign w34496 = ~pi6154 & pi9040;
assign w34497 = ~pi6038 & ~pi9040;
assign w34498 = ~w34496 & ~w34497;
assign w34499 = pi1785 & ~w34498;
assign w34500 = ~pi1785 & w34498;
assign w34501 = ~w34499 & ~w34500;
assign w34502 = w34495 & w34501;
assign w34503 = w34489 & w34502;
assign w34504 = ~w34482 & ~w34501;
assign w34505 = w34495 & w34504;
assign w34506 = w34504 & w34998;
assign w34507 = ~w34503 & ~w34506;
assign w34508 = w34482 & ~w34488;
assign w34509 = ~w34488 & ~w34495;
assign w34510 = ~w34508 & ~w34509;
assign w34511 = w34482 & ~w34501;
assign w34512 = ~pi6052 & pi9040;
assign w34513 = ~pi6082 & ~pi9040;
assign w34514 = ~w34512 & ~w34513;
assign w34515 = pi1816 & ~w34514;
assign w34516 = ~pi1816 & w34514;
assign w34517 = ~w34515 & ~w34516;
assign w34518 = ~w34511 & w34517;
assign w34519 = ~w34510 & w34518;
assign w34520 = w34482 & w34488;
assign w34521 = w34495 & w34520;
assign w34522 = w34520 & w66071;
assign w34523 = ~w34519 & ~w34522;
assign w34524 = w34507 & w34523;
assign w34525 = ~w34476 & ~w34524;
assign w34526 = ~w34511 & ~w34517;
assign w34527 = w34510 & w34526;
assign w34528 = ~w34488 & w34511;
assign w34529 = w34495 & w34528;
assign w34530 = w34488 & ~w34495;
assign w34531 = ~w34526 & ~w34530;
assign w34532 = ~w34529 & w34531;
assign w34533 = ~w34527 & ~w34532;
assign w34534 = ~w34482 & w34501;
assign w34535 = ~w34528 & ~w34534;
assign w34536 = (~w34495 & w34528) | (~w34495 & w66072) | (w34528 & w66072);
assign w34537 = w34518 & ~w34536;
assign w34538 = w34524 & w34537;
assign w34539 = (w34476 & w34538) | (w34476 & w66073) | (w34538 & w66073);
assign w34540 = w34488 & ~w34511;
assign w34541 = ~w34528 & ~w34540;
assign w34542 = ~w34476 & ~w34505;
assign w34543 = ~w34541 & w34542;
assign w34544 = w34507 & ~w34529;
assign w34545 = ~w34543 & w34544;
assign w34546 = ~w34517 & ~w34545;
assign w34547 = ~w34525 & ~w34546;
assign w34548 = ~w34539 & w34547;
assign w34549 = ~pi1829 & w34548;
assign w34550 = pi1829 & ~w34548;
assign w34551 = ~w34549 & ~w34550;
assign w34552 = ~w34283 & ~w34333;
assign w34553 = ~w34334 & w34552;
assign w34554 = w34271 & w34291;
assign w34555 = w34277 & w34304;
assign w34556 = w34277 & ~w34291;
assign w34557 = w34283 & ~w34292;
assign w34558 = ~w34556 & w34557;
assign w34559 = (~w34554 & w34558) | (~w34554 & w66074) | (w34558 & w66074);
assign w34560 = ~w34553 & ~w34559;
assign w34561 = ~w34322 & ~w34560;
assign w34562 = ~w34270 & ~w34283;
assign w34563 = w34325 & w34562;
assign w34564 = ~w34264 & w34563;
assign w34565 = ~w34270 & w34283;
assign w34566 = ~w34554 & ~w34565;
assign w34567 = w34330 & ~w34566;
assign w34568 = ~w34303 & w34567;
assign w34569 = w34325 & w34565;
assign w34570 = w34277 & ~w34569;
assign w34571 = w34271 & ~w34570;
assign w34572 = w34284 & w34292;
assign w34573 = ~w34270 & w34556;
assign w34574 = ~w34298 & ~w34573;
assign w34575 = ~w34264 & ~w34574;
assign w34576 = ~w34336 & ~w34572;
assign w34577 = ~w34571 & ~w34575;
assign w34578 = w34576 & w34577;
assign w34579 = w34322 & ~w34578;
assign w34580 = ~w34564 & ~w34568;
assign w34581 = ~w34561 & w34580;
assign w34582 = ~w34579 & w34581;
assign w34583 = pi1845 & w34582;
assign w34584 = ~pi1845 & ~w34582;
assign w34585 = ~w34583 & ~w34584;
assign w34586 = w34113 & ~w34179;
assign w34587 = (w34132 & w34586) | (w34132 & w66075) | (w34586 & w66075);
assign w34588 = w34140 & ~w34220;
assign w34589 = ~w34174 & ~w34175;
assign w34590 = w34153 & w34589;
assign w34591 = w34215 & ~w34586;
assign w34592 = ~w34590 & w34591;
assign w34593 = (~w34587 & w34592) | (~w34587 & w66076) | (w34592 & w66076);
assign w34594 = w34164 & ~w34593;
assign w34595 = ~w34164 & ~w34176;
assign w34596 = ~w34219 & w34595;
assign w34597 = ~w34587 & w34596;
assign w34598 = w34141 & ~w34597;
assign w34599 = ~w34134 & ~w34220;
assign w34600 = ~w34164 & ~w34599;
assign w34601 = ~w34140 & ~w34587;
assign w34602 = ~w34600 & w34601;
assign w34603 = ~w34598 & ~w34602;
assign w34604 = ~w34594 & ~w34603;
assign w34605 = ~pi1846 & w34604;
assign w34606 = pi1846 & ~w34604;
assign w34607 = ~w34605 & ~w34606;
assign w34608 = ~pi6064 & pi9040;
assign w34609 = ~pi6070 & ~pi9040;
assign w34610 = ~w34608 & ~w34609;
assign w34611 = pi1821 & ~w34610;
assign w34612 = ~pi1821 & w34610;
assign w34613 = ~w34611 & ~w34612;
assign w34614 = ~pi6298 & pi9040;
assign w34615 = ~pi6041 & ~pi9040;
assign w34616 = ~w34614 & ~w34615;
assign w34617 = pi1820 & ~w34616;
assign w34618 = ~pi1820 & w34616;
assign w34619 = ~w34617 & ~w34618;
assign w34620 = w34613 & w34619;
assign w34621 = ~pi6084 & pi9040;
assign w34622 = ~pi6051 & ~pi9040;
assign w34623 = ~w34621 & ~w34622;
assign w34624 = pi1815 & ~w34623;
assign w34625 = ~pi1815 & w34623;
assign w34626 = ~w34624 & ~w34625;
assign w34627 = ~pi6149 & pi9040;
assign w34628 = ~pi6259 & ~pi9040;
assign w34629 = ~w34627 & ~w34628;
assign w34630 = pi1800 & ~w34629;
assign w34631 = ~pi1800 & w34629;
assign w34632 = ~w34630 & ~w34631;
assign w34633 = ~w34626 & ~w34632;
assign w34634 = w34620 & w34633;
assign w34635 = w34619 & ~w34632;
assign w34636 = ~w34613 & ~w34635;
assign w34637 = ~pi6062 & pi9040;
assign w34638 = ~pi6176 & ~pi9040;
assign w34639 = ~w34637 & ~w34638;
assign w34640 = pi1794 & ~w34639;
assign w34641 = ~pi1794 & w34639;
assign w34642 = ~w34640 & ~w34641;
assign w34643 = ~pi6070 & pi9040;
assign w34644 = ~pi6298 & ~pi9040;
assign w34645 = ~w34643 & ~w34644;
assign w34646 = pi1785 & ~w34645;
assign w34647 = ~pi1785 & w34645;
assign w34648 = ~w34646 & ~w34647;
assign w34649 = w34626 & w34648;
assign w34650 = w34619 & ~w34648;
assign w34651 = ~w34632 & ~w34648;
assign w34652 = ~w34650 & ~w34651;
assign w34653 = ~w34649 & w34652;
assign w34654 = w34626 & w34632;
assign w34655 = ~w34642 & ~w34654;
assign w34656 = w34636 & w34655;
assign w34657 = ~w34653 & w34656;
assign w34658 = w34652 & w63897;
assign w34659 = (~w34648 & w34635) | (~w34648 & w66077) | (w34635 & w66077);
assign w34660 = w34658 & w34659;
assign w34661 = w34632 & w34648;
assign w34662 = ~w34651 & ~w34661;
assign w34663 = ~w34619 & w34648;
assign w34664 = w34626 & ~w34663;
assign w34665 = ~w34626 & w34663;
assign w34666 = ~w34664 & ~w34665;
assign w34667 = ~w34613 & ~w34662;
assign w34668 = ~w34666 & w34667;
assign w34669 = ~w34654 & ~w34663;
assign w34670 = w34613 & ~w34669;
assign w34671 = ~w34650 & w34666;
assign w34672 = w34626 & w34650;
assign w34673 = (~w34672 & ~w34666) | (~w34672 & w63898) | (~w34666 & w63898);
assign w34674 = w34632 & ~w34673;
assign w34675 = ~w34673 & w66078;
assign w34676 = ~w34619 & w34651;
assign w34677 = w34626 & w34676;
assign w34678 = ~w34613 & w34619;
assign w34679 = w34626 & w34678;
assign w34680 = w34632 & w34649;
assign w34681 = ~w34679 & ~w34680;
assign w34682 = w34635 & w34648;
assign w34683 = w34681 & w34682;
assign w34684 = ~w34642 & ~w34677;
assign w34685 = ~w34683 & w34684;
assign w34686 = ~w34675 & w34685;
assign w34687 = w34613 & ~w34619;
assign w34688 = w34626 & w34687;
assign w34689 = w34662 & w34688;
assign w34690 = w34642 & ~w34679;
assign w34691 = w34619 & ~w34651;
assign w34692 = ~w34626 & ~w34676;
assign w34693 = ~w34691 & w34692;
assign w34694 = ~w34689 & w34690;
assign w34695 = ~w34658 & w34694;
assign w34696 = ~w34693 & w34695;
assign w34697 = ~w34686 & ~w34696;
assign w34698 = ~w34634 & ~w34657;
assign w34699 = ~w34668 & w34698;
assign w34700 = ~w34660 & w34699;
assign w34701 = ~w34697 & w34700;
assign w34702 = pi1825 & w34701;
assign w34703 = ~pi1825 & ~w34701;
assign w34704 = ~w34702 & ~w34703;
assign w34705 = w34327 & w34329;
assign w34706 = (~w34283 & ~w34326) | (~w34283 & w34562) | (~w34326 & w34562);
assign w34707 = ~w34705 & w34706;
assign w34708 = w34270 & w34308;
assign w34709 = w34283 & ~w34324;
assign w34710 = ~w34555 & ~w34708;
assign w34711 = w34709 & w34710;
assign w34712 = ~w34707 & ~w34711;
assign w34713 = w34322 & ~w34568;
assign w34714 = ~w34712 & w34713;
assign w34715 = w34270 & w34283;
assign w34716 = w34300 & w34715;
assign w34717 = ~w34554 & ~w34708;
assign w34718 = ~w34283 & ~w34717;
assign w34719 = ~w34322 & ~w34572;
assign w34720 = ~w34716 & w34719;
assign w34721 = w34302 & w34720;
assign w34722 = ~w34567 & ~w34718;
assign w34723 = w34721 & w34722;
assign w34724 = ~w34296 & ~w34313;
assign w34725 = ~w34560 & w34724;
assign w34726 = (~w34725 & w34714) | (~w34725 & w66079) | (w34714 & w66079);
assign w34727 = pi1839 & w34726;
assign w34728 = ~pi1839 & ~w34726;
assign w34729 = ~w34727 & ~w34728;
assign w34730 = ~w34057 & w34357;
assign w34731 = ~w34079 & ~w34080;
assign w34732 = w34032 & ~w34350;
assign w34733 = w34731 & w34732;
assign w34734 = ~w34070 & ~w34080;
assign w34735 = w34060 & ~w34734;
assign w34736 = w34046 & w34734;
assign w34737 = ~w34733 & ~w34735;
assign w34738 = ~w34736 & w34737;
assign w34739 = w34057 & ~w34738;
assign w34740 = w34026 & w34086;
assign w34741 = ~w34061 & ~w34740;
assign w34742 = ~w34731 & ~w34741;
assign w34743 = ~w34039 & w34057;
assign w34744 = w34047 & ~w34743;
assign w34745 = w34086 & w34233;
assign w34746 = ~w34744 & ~w34745;
assign w34747 = ~w34026 & ~w34746;
assign w34748 = ~w34742 & ~w34747;
assign w34749 = ~w34730 & w34748;
assign w34750 = ~w34739 & w34749;
assign w34751 = ~pi1870 & w34750;
assign w34752 = pi1870 & ~w34750;
assign w34753 = ~w34751 & ~w34752;
assign w34754 = ~pi6297 & pi9040;
assign w34755 = ~pi6053 & ~pi9040;
assign w34756 = ~w34754 & ~w34755;
assign w34757 = pi1806 & ~w34756;
assign w34758 = ~pi1806 & w34756;
assign w34759 = ~w34757 & ~w34758;
assign w34760 = ~pi6159 & pi9040;
assign w34761 = ~pi6149 & ~pi9040;
assign w34762 = ~w34760 & ~w34761;
assign w34763 = pi1798 & ~w34762;
assign w34764 = ~pi1798 & w34762;
assign w34765 = ~w34763 & ~w34764;
assign w34766 = ~w34759 & w34765;
assign w34767 = ~pi6060 & pi9040;
assign w34768 = ~pi6059 & ~pi9040;
assign w34769 = ~w34767 & ~w34768;
assign w34770 = pi1808 & ~w34769;
assign w34771 = ~pi1808 & w34769;
assign w34772 = ~w34770 & ~w34771;
assign w34773 = ~w34766 & ~w34772;
assign w34774 = ~pi6151 & pi9040;
assign w34775 = ~pi6297 & ~pi9040;
assign w34776 = ~w34774 & ~w34775;
assign w34777 = pi1807 & ~w34776;
assign w34778 = ~pi1807 & w34776;
assign w34779 = ~w34777 & ~w34778;
assign w34780 = ~w34772 & w34779;
assign w34781 = ~pi6259 & pi9040;
assign w34782 = ~pi6062 & ~pi9040;
assign w34783 = ~w34781 & ~w34782;
assign w34784 = pi1823 & ~w34783;
assign w34785 = ~pi1823 & w34783;
assign w34786 = ~w34784 & ~w34785;
assign w34787 = ~w34780 & ~w34786;
assign w34788 = w34759 & ~w34765;
assign w34789 = w34787 & w34788;
assign w34790 = ~w34759 & w34779;
assign w34791 = w34765 & ~w34772;
assign w34792 = ~w34786 & w34791;
assign w34793 = w34790 & w34792;
assign w34794 = ~w34789 & ~w34793;
assign w34795 = ~w34766 & w34772;
assign w34796 = w34779 & ~w34788;
assign w34797 = ~w34795 & w34796;
assign w34798 = ~w34786 & w34797;
assign w34799 = w34794 & ~w34798;
assign w34800 = w34773 & ~w34799;
assign w34801 = ~w34759 & ~w34779;
assign w34802 = ~w34765 & w34801;
assign w34803 = w34786 & w34802;
assign w34804 = w34759 & w34765;
assign w34805 = w34772 & ~w34804;
assign w34806 = ~w34773 & ~w34805;
assign w34807 = w34787 & w34806;
assign w34808 = ~pi6071 & pi9040;
assign w34809 = ~pi6054 & ~pi9040;
assign w34810 = ~w34808 & ~w34809;
assign w34811 = pi1805 & ~w34810;
assign w34812 = ~pi1805 & w34810;
assign w34813 = ~w34811 & ~w34812;
assign w34814 = w34765 & w34786;
assign w34815 = w34801 & w34814;
assign w34816 = ~w34779 & ~w34815;
assign w34817 = ~w34765 & w34790;
assign w34818 = ~w34805 & ~w34817;
assign w34819 = w34790 & w66080;
assign w34820 = ~w34816 & ~w34818;
assign w34821 = ~w34819 & w34820;
assign w34822 = ~w34803 & w34813;
assign w34823 = ~w34807 & w34822;
assign w34824 = ~w34821 & w34823;
assign w34825 = ~w34765 & ~w34786;
assign w34826 = w34759 & ~w34779;
assign w34827 = ~w34790 & ~w34826;
assign w34828 = w34765 & w34772;
assign w34829 = w34827 & w34828;
assign w34830 = ~w34825 & ~w34829;
assign w34831 = w34816 & ~w34830;
assign w34832 = w34779 & w34786;
assign w34833 = ~w34797 & w34832;
assign w34834 = ~w34813 & ~w34833;
assign w34835 = ~w34831 & w34834;
assign w34836 = ~w34824 & ~w34835;
assign w34837 = ~w34772 & ~w34827;
assign w34838 = ~w34791 & ~w34826;
assign w34839 = w34813 & ~w34814;
assign w34840 = ~w34838 & ~w34839;
assign w34841 = w34837 & w34840;
assign w34842 = ~w34800 & ~w34841;
assign w34843 = ~w34836 & w34842;
assign w34844 = pi1835 & ~w34843;
assign w34845 = ~pi1835 & w34843;
assign w34846 = ~w34844 & ~w34845;
assign w34847 = w34142 & w34199;
assign w34848 = ~w34119 & w34152;
assign w34849 = ~w34180 & ~w34848;
assign w34850 = ~w34140 & ~w34849;
assign w34851 = w34213 & ~w34848;
assign w34852 = ~w34850 & ~w34851;
assign w34853 = (~w34847 & ~w34181) | (~w34847 & w66081) | (~w34181 & w66081);
assign w34854 = (~w34164 & w34852) | (~w34164 & w66082) | (w34852 & w66082);
assign w34855 = w34182 & ~w34218;
assign w34856 = w34132 & w34156;
assign w34857 = (~w34856 & w34855) | (~w34856 & w66083) | (w34855 & w66083);
assign w34858 = w34164 & ~w34857;
assign w34859 = w34140 & ~w34170;
assign w34860 = w34142 & w34152;
assign w34861 = w34215 & ~w34860;
assign w34862 = ~w34859 & ~w34861;
assign w34863 = ~w34854 & ~w34862;
assign w34864 = ~w34858 & w34863;
assign w34865 = ~pi1851 & w34864;
assign w34866 = pi1851 & ~w34864;
assign w34867 = ~w34865 & ~w34866;
assign w34868 = w34381 & w34387;
assign w34869 = w34425 & w34868;
assign w34870 = ~w34436 & w34451;
assign w34871 = ~w34445 & w34870;
assign w34872 = w34387 & ~w34400;
assign w34873 = w34444 & w34872;
assign w34874 = ~w34871 & ~w34873;
assign w34875 = ~w34434 & ~w34874;
assign w34876 = ~w34381 & w34393;
assign w34877 = ~w34430 & ~w34876;
assign w34878 = w34409 & ~w34432;
assign w34879 = ~w34877 & ~w34878;
assign w34880 = ~w34406 & w34421;
assign w34881 = w34381 & ~w34458;
assign w34882 = ~w34880 & w34881;
assign w34883 = ~w34422 & w34882;
assign w34884 = w34417 & ~w34879;
assign w34885 = ~w34883 & w34884;
assign w34886 = w34425 & ~w34437;
assign w34887 = ~w34381 & ~w34406;
assign w34888 = ~w34442 & ~w34887;
assign w34889 = ~w34882 & w34888;
assign w34890 = w34416 & ~w34886;
assign w34891 = ~w34889 & w34890;
assign w34892 = ~w34885 & ~w34891;
assign w34893 = ~w34869 & ~w34875;
assign w34894 = ~w34892 & w34893;
assign w34895 = pi1834 & ~w34894;
assign w34896 = ~pi1834 & w34894;
assign w34897 = ~w34895 & ~w34896;
assign w34898 = w34788 & w34832;
assign w34899 = ~w34772 & w34898;
assign w34900 = ~w34759 & ~w34772;
assign w34901 = w34786 & ~w34900;
assign w34902 = w34772 & w34826;
assign w34903 = w34901 & ~w34902;
assign w34904 = ~w34814 & ~w34903;
assign w34905 = ~w34772 & w34788;
assign w34906 = ~w34786 & ~w34905;
assign w34907 = ~w34779 & w34804;
assign w34908 = w34906 & ~w34907;
assign w34909 = w34904 & ~w34908;
assign w34910 = ~w34772 & w34802;
assign w34911 = w34772 & w34825;
assign w34912 = w34801 & w34911;
assign w34913 = w34796 & w34901;
assign w34914 = w34804 & w63899;
assign w34915 = ~w34913 & ~w34914;
assign w34916 = w34786 & ~w34838;
assign w34917 = (~w34912 & ~w34915) | (~w34912 & w63900) | (~w34915 & w63900);
assign w34918 = ~w34910 & w34917;
assign w34919 = w34813 & ~w34815;
assign w34920 = w34779 & w34806;
assign w34921 = ~w34786 & w34837;
assign w34922 = ~w34898 & ~w34912;
assign w34923 = w34919 & w34922;
assign w34924 = ~w34920 & ~w34921;
assign w34925 = w34923 & w34924;
assign w34926 = ~w34813 & ~w34819;
assign w34927 = ~w34910 & w34926;
assign w34928 = w34765 & ~w34779;
assign w34929 = ~w34789 & ~w34928;
assign w34930 = w34906 & ~w34929;
assign w34931 = ~w34803 & w34915;
assign w34932 = w34927 & w34931;
assign w34933 = ~w34930 & w34932;
assign w34934 = ~w34925 & ~w34933;
assign w34935 = ~w34793 & ~w34899;
assign w34936 = (w34935 & w34918) | (w34935 & w66084) | (w34918 & w66084);
assign w34937 = (pi1827 & w34934) | (pi1827 & w66085) | (w34934 & w66085);
assign w34938 = ~w34934 & w66086;
assign w34939 = ~w34937 & ~w34938;
assign w34940 = ~w34430 & ~w34872;
assign w34941 = w34444 & ~w34940;
assign w34942 = w34407 & w34435;
assign w34943 = ~w34450 & ~w34942;
assign w34944 = ~w34409 & ~w34943;
assign w34945 = ~w34381 & ~w34431;
assign w34946 = ~w34425 & w34945;
assign w34947 = ~w34944 & w34946;
assign w34948 = w34432 & w34947;
assign w34949 = w34440 & w34870;
assign w34950 = w34418 & ~w34868;
assign w34951 = w34940 & w34950;
assign w34952 = ~w34941 & ~w34951;
assign w34953 = ~w34949 & w34952;
assign w34954 = ~w34948 & w34953;
assign w34955 = w34416 & ~w34954;
assign w34956 = ~w34381 & w34886;
assign w34957 = w34394 & w34423;
assign w34958 = ~w34452 & ~w34957;
assign w34959 = w34434 & ~w34958;
assign w34960 = ~w34416 & ~w34440;
assign w34961 = ~w34947 & w34960;
assign w34962 = ~w34956 & ~w34959;
assign w34963 = ~w34961 & w34962;
assign w34964 = (pi1840 & w34955) | (pi1840 & w66087) | (w34955 & w66087);
assign w34965 = ~w34955 & w66088;
assign w34966 = ~w34964 & ~w34965;
assign w34967 = ~w34619 & ~w34633;
assign w34968 = ~w34626 & w34648;
assign w34969 = w34635 & w34968;
assign w34970 = ~w34967 & ~w34969;
assign w34971 = w34613 & ~w34970;
assign w34972 = w34636 & ~w34967;
assign w34973 = ~w34632 & w34672;
assign w34974 = w34642 & ~w34680;
assign w34975 = ~w34972 & w34974;
assign w34976 = ~w34973 & w34975;
assign w34977 = ~w34971 & w34976;
assign w34978 = w34620 & w34673;
assign w34979 = ~w34665 & ~w34672;
assign w34980 = w34619 & ~w34968;
assign w34981 = ~w34613 & w34669;
assign w34982 = ~w34980 & w34981;
assign w34983 = (~w34642 & w34979) | (~w34642 & w66089) | (w34979 & w66089);
assign w34984 = ~w34982 & w34983;
assign w34985 = ~w34978 & w34984;
assign w34986 = ~w34977 & ~w34985;
assign w34987 = ~w34689 & ~w34986;
assign w34988 = ~pi1831 & w34987;
assign w34989 = pi1831 & ~w34987;
assign w34990 = ~w34988 & ~w34989;
assign w34991 = ~w34506 & ~w34530;
assign w34992 = ~w34495 & ~w34501;
assign w34993 = ~w34526 & ~w34992;
assign w34994 = ~w34991 & w34993;
assign w34995 = w34495 & ~w34517;
assign w34996 = ~w34508 & w34995;
assign w34997 = ~w34540 & w34996;
assign w34998 = ~w34488 & w34495;
assign w34999 = ~w34495 & w34520;
assign w35000 = ~w34517 & ~w34999;
assign w35001 = w34501 & ~w34998;
assign w35002 = ~w35000 & w35001;
assign w35003 = ~w34488 & ~w34517;
assign w35004 = ~w34530 & ~w35003;
assign w35005 = w34504 & ~w35004;
assign w35006 = w34482 & ~w34495;
assign w35007 = ~w34501 & ~w34517;
assign w35008 = w35006 & w35007;
assign w35009 = w34502 & w34508;
assign w35010 = ~w35008 & ~w35009;
assign w35011 = ~w34509 & ~w35003;
assign w35012 = ~w35010 & ~w35011;
assign w35013 = w34476 & ~w34997;
assign w35014 = ~w35005 & w35013;
assign w35015 = ~w35002 & ~w35012;
assign w35016 = w35014 & w35015;
assign w35017 = w34517 & w34522;
assign w35018 = ~w34541 & w34995;
assign w35019 = ~w34476 & w35010;
assign w35020 = ~w34536 & w35019;
assign w35021 = ~w35017 & ~w35018;
assign w35022 = w35020 & w35021;
assign w35023 = ~w35016 & ~w35022;
assign w35024 = ~w34994 & ~w35023;
assign w35025 = ~pi1832 & ~w35024;
assign w35026 = pi1832 & w35024;
assign w35027 = ~w35025 & ~w35026;
assign w35028 = w34270 & w34331;
assign w35029 = ~w34283 & ~w34295;
assign w35030 = ~w35028 & w35029;
assign w35031 = ~w34337 & ~w35030;
assign w35032 = w34330 & w34562;
assign w35033 = w34264 & ~w34296;
assign w35034 = w34322 & ~w34569;
assign w35035 = ~w35032 & w35034;
assign w35036 = ~w35033 & w35035;
assign w35037 = ~w34339 & w34552;
assign w35038 = w34283 & ~w34301;
assign w35039 = ~w34305 & ~w34573;
assign w35040 = w35038 & w35039;
assign w35041 = ~w35037 & ~w35040;
assign w35042 = ~w34322 & ~w34324;
assign w35043 = ~w34563 & w35042;
assign w35044 = ~w35041 & w35043;
assign w35045 = ~w35036 & ~w35044;
assign w35046 = ~w35031 & ~w35045;
assign w35047 = ~pi1833 & w35046;
assign w35048 = pi1833 & ~w35046;
assign w35049 = ~w35047 & ~w35048;
assign w35050 = w34670 & ~w34673;
assign w35051 = w34636 & ~w34679;
assign w35052 = ~w34671 & w35051;
assign w35053 = (~w34969 & ~w34658) | (~w34969 & w66090) | (~w34658 & w66090);
assign w35054 = ~w35052 & w35053;
assign w35055 = (w34642 & ~w35054) | (w34642 & w66091) | (~w35054 & w66091);
assign w35056 = ~w34613 & ~w34632;
assign w35057 = ~w34979 & w35056;
assign w35058 = ~w34677 & w34690;
assign w35059 = ~w34678 & ~w34687;
assign w35060 = w34661 & ~w35059;
assign w35061 = ~w34642 & ~w34681;
assign w35062 = ~w34633 & ~w34688;
assign w35063 = ~w34648 & ~w35062;
assign w35064 = ~w35060 & ~w35061;
assign w35065 = (~w35058 & ~w35064) | (~w35058 & w66092) | (~w35064 & w66092);
assign w35066 = ~w34634 & ~w35057;
assign w35067 = ~w35065 & w35066;
assign w35068 = ~w35055 & w35067;
assign w35069 = ~pi1837 & w35068;
assign w35070 = pi1837 & ~w35068;
assign w35071 = ~w35069 & ~w35070;
assign w35072 = ~w34780 & ~w34792;
assign w35073 = w34759 & ~w35072;
assign w35074 = w34927 & ~w35073;
assign w35075 = w34917 & w35074;
assign w35076 = ~w34817 & ~w34914;
assign w35077 = w34786 & ~w35076;
assign w35078 = w34813 & ~w34829;
assign w35079 = w34794 & w35078;
assign w35080 = ~w35077 & w35079;
assign w35081 = ~w35075 & ~w35080;
assign w35082 = ~w34829 & ~w34910;
assign w35083 = ~w34786 & ~w35082;
assign w35084 = w34790 & w34901;
assign w35085 = ~w34899 & ~w35084;
assign w35086 = ~w35083 & w35085;
assign w35087 = ~w35081 & w35086;
assign w35088 = pi1841 & ~w35087;
assign w35089 = ~pi1841 & w35087;
assign w35090 = ~w35088 & ~w35089;
assign w35091 = ~w34495 & w34508;
assign w35092 = ~w35007 & w35091;
assign w35093 = ~w34508 & ~w34992;
assign w35094 = ~w35006 & ~w35093;
assign w35095 = ~w34541 & w35094;
assign w35096 = w34501 & w34999;
assign w35097 = ~w34503 & ~w35096;
assign w35098 = ~w34488 & w34534;
assign w35099 = ~w35095 & ~w35098;
assign w35100 = ~w34508 & w34517;
assign w35101 = w35099 & w66093;
assign w35102 = ~w34476 & ~w35092;
assign w35103 = (w35099 & w66094) | (w35099 & w66095) | (w66094 & w66095);
assign w35104 = ~w35101 & w35103;
assign w35105 = ~w34996 & ~w35098;
assign w35106 = ~w34502 & ~w35105;
assign w35107 = w34517 & w35094;
assign w35108 = w34476 & w35010;
assign w35109 = w35097 & w35108;
assign w35110 = ~w35106 & ~w35107;
assign w35111 = w35109 & w35110;
assign w35112 = ~w35104 & ~w35111;
assign w35113 = ~pi1844 & w35112;
assign w35114 = pi1844 & ~w35112;
assign w35115 = ~w35113 & ~w35114;
assign w35116 = ~pi6051 & pi9040;
assign w35117 = ~pi6151 & ~pi9040;
assign w35118 = ~w35116 & ~w35117;
assign w35119 = pi1806 & ~w35118;
assign w35120 = ~pi1806 & w35118;
assign w35121 = ~w35119 & ~w35120;
assign w35122 = ~pi6294 & pi9040;
assign w35123 = ~pi6147 & ~pi9040;
assign w35124 = ~w35122 & ~w35123;
assign w35125 = pi1801 & ~w35124;
assign w35126 = ~pi1801 & w35124;
assign w35127 = ~w35125 & ~w35126;
assign w35128 = ~pi6078 & pi9040;
assign w35129 = ~pi6154 & ~pi9040;
assign w35130 = ~w35128 & ~w35129;
assign w35131 = pi1812 & ~w35130;
assign w35132 = ~pi1812 & w35130;
assign w35133 = ~w35131 & ~w35132;
assign w35134 = ~w35127 & ~w35133;
assign w35135 = w35127 & w35133;
assign w35136 = ~w35134 & ~w35135;
assign w35137 = ~pi6059 & pi9040;
assign w35138 = ~pi6084 & ~pi9040;
assign w35139 = ~w35137 & ~w35138;
assign w35140 = pi1807 & ~w35139;
assign w35141 = ~pi1807 & w35139;
assign w35142 = ~w35140 & ~w35141;
assign w35143 = ~pi6041 & pi9040;
assign w35144 = ~pi6035 & ~pi9040;
assign w35145 = ~w35143 & ~w35144;
assign w35146 = pi1804 & ~w35145;
assign w35147 = ~pi1804 & w35145;
assign w35148 = ~w35146 & ~w35147;
assign w35149 = ~w35142 & w35148;
assign w35150 = w35142 & ~w35148;
assign w35151 = ~pi6035 & pi9040;
assign w35152 = ~pi6071 & ~pi9040;
assign w35153 = ~w35151 & ~w35152;
assign w35154 = pi1797 & ~w35153;
assign w35155 = ~pi1797 & w35153;
assign w35156 = ~w35154 & ~w35155;
assign w35157 = w35150 & ~w35156;
assign w35158 = ~w35149 & ~w35157;
assign w35159 = ~w35142 & ~w35148;
assign w35160 = ~w35127 & ~w35148;
assign w35161 = ~w35159 & ~w35160;
assign w35162 = w35133 & ~w35142;
assign w35163 = w35148 & ~w35162;
assign w35164 = w35161 & ~w35163;
assign w35165 = ~w35134 & ~w35164;
assign w35166 = w35134 & w35149;
assign w35167 = ~w35127 & w35159;
assign w35168 = ~w35161 & ~w35167;
assign w35169 = ~w35166 & ~w35168;
assign w35170 = ~w35165 & w35169;
assign w35171 = (w35136 & w35170) | (w35136 & w66096) | (w35170 & w66096);
assign w35172 = ~w35136 & w35158;
assign w35173 = ~w35121 & ~w35172;
assign w35174 = ~w35171 & w35173;
assign w35175 = ~w35133 & w35142;
assign w35176 = ~w35164 & ~w35175;
assign w35177 = w35121 & ~w35156;
assign w35178 = ~w35159 & w35177;
assign w35179 = w35176 & w35178;
assign w35180 = w35127 & w35175;
assign w35181 = w35134 & w35159;
assign w35182 = ~w35180 & ~w35181;
assign w35183 = w35156 & ~w35182;
assign w35184 = w35121 & w35156;
assign w35185 = ~w35176 & w35184;
assign w35186 = w35121 & w35135;
assign w35187 = w35159 & w35186;
assign w35188 = ~w35183 & ~w35187;
assign w35189 = ~w35179 & w35188;
assign w35190 = ~w35185 & w35189;
assign w35191 = ~w35174 & w35190;
assign w35192 = ~pi1865 & w35191;
assign w35193 = pi1865 & ~w35191;
assign w35194 = ~w35192 & ~w35193;
assign w35195 = w35133 & w35148;
assign w35196 = ~w35133 & ~w35148;
assign w35197 = ~w35195 & ~w35196;
assign w35198 = w35142 & ~w35197;
assign w35199 = (~w35156 & w35198) | (~w35156 & w63902) | (w35198 & w63902);
assign w35200 = (w35198 & w66097) | (w35198 & w66098) | (w66097 & w66098);
assign w35201 = ~w35156 & w35170;
assign w35202 = ~w35149 & ~w35156;
assign w35203 = ~w35166 & ~w35195;
assign w35204 = ~w35202 & w35203;
assign w35205 = ~w35170 & w35204;
assign w35206 = ~w35201 & ~w35205;
assign w35207 = ~w35121 & ~w35206;
assign w35208 = (w35134 & w35157) | (w35134 & w35166) | (w35157 & w35166);
assign w35209 = ~w35134 & ~w35202;
assign w35210 = ~w35133 & ~w35156;
assign w35211 = ~w35127 & w35210;
assign w35212 = ~w35150 & ~w35211;
assign w35213 = ~w35209 & w35212;
assign w35214 = (w35121 & w35213) | (w35121 & w66099) | (w35213 & w66099);
assign w35215 = w35156 & ~w35159;
assign w35216 = ~w35175 & w35215;
assign w35217 = ~w35169 & w35216;
assign w35218 = w35127 & w35184;
assign w35219 = (w35218 & w35170) | (w35218 & w66100) | (w35170 & w66100);
assign w35220 = ~w35200 & ~w35217;
assign w35221 = ~w35214 & w35220;
assign w35222 = ~w35219 & w35221;
assign w35223 = ~w35207 & w35222;
assign w35224 = pi1859 & w35223;
assign w35225 = ~pi1859 & ~w35223;
assign w35226 = ~w35224 & ~w35225;
assign w35227 = ~w35133 & w35170;
assign w35228 = w35127 & w35148;
assign w35229 = ~w35162 & ~w35228;
assign w35230 = w35127 & w35162;
assign w35231 = ~w35229 & ~w35230;
assign w35232 = w35156 & ~w35231;
assign w35233 = ~w35196 & w35229;
assign w35234 = ~w35156 & ~w35233;
assign w35235 = ~w35232 & ~w35234;
assign w35236 = (~w35121 & w35227) | (~w35121 & w66101) | (w35227 & w66101);
assign w35237 = w35133 & w35159;
assign w35238 = ~w35228 & ~w35237;
assign w35239 = w35177 & ~w35238;
assign w35240 = ~w35169 & w35184;
assign w35241 = w35183 & w35197;
assign w35242 = w35135 & w35150;
assign w35243 = ~w35230 & ~w35242;
assign w35244 = ~w35142 & ~w35156;
assign w35245 = ~w35121 & ~w35244;
assign w35246 = ~w35243 & ~w35245;
assign w35247 = ~w35239 & ~w35246;
assign w35248 = ~w35240 & w35247;
assign w35249 = ~w35241 & w35248;
assign w35250 = ~w35236 & w35249;
assign w35251 = pi1867 & w35250;
assign w35252 = ~pi1867 & ~w35250;
assign w35253 = ~w35251 & ~w35252;
assign w35254 = ~w34613 & ~w34968;
assign w35255 = ~w34664 & w35254;
assign w35256 = ~w34633 & w34652;
assign w35257 = w34669 & w35256;
assign w35258 = ~w35255 & ~w35257;
assign w35259 = ~w34680 & w34690;
assign w35260 = ~w35258 & ~w35259;
assign w35261 = ~w34649 & ~w34659;
assign w35262 = w34613 & ~w34642;
assign w35263 = w35261 & w35262;
assign w35264 = ~w35257 & w66102;
assign w35265 = ~w34632 & ~w35264;
assign w35266 = w34642 & ~w34674;
assign w35267 = ~w35265 & w35266;
assign w35268 = ~w35260 & ~w35263;
assign w35269 = ~w35267 & w35268;
assign w35270 = pi1838 & ~w35269;
assign w35271 = ~pi1838 & w35269;
assign w35272 = ~w35270 & ~w35271;
assign w35273 = ~w34819 & ~w34829;
assign w35274 = w34786 & ~w35273;
assign w35275 = w34805 & w34813;
assign w35276 = ~w34911 & ~w35275;
assign w35277 = w34827 & ~w35276;
assign w35278 = ~w34813 & ~w34899;
assign w35279 = ~w34920 & w35278;
assign w35280 = ~w34909 & w35279;
assign w35281 = w34826 & ~w34904;
assign w35282 = ~w34798 & w34919;
assign w35283 = ~w35281 & w35282;
assign w35284 = ~w35280 & ~w35283;
assign w35285 = ~w35274 & ~w35277;
assign w35286 = ~w35284 & w35285;
assign w35287 = pi1842 & ~w35286;
assign w35288 = ~pi1842 & w35286;
assign w35289 = ~w35287 & ~w35288;
assign w35290 = ~w35142 & w35156;
assign w35291 = ~w35197 & ~w35290;
assign w35292 = w35197 & ~w35210;
assign w35293 = w35127 & ~w35291;
assign w35294 = ~w35292 & w35293;
assign w35295 = ~w35149 & ~w35290;
assign w35296 = w35197 & ~w35295;
assign w35297 = ~w35198 & ~w35296;
assign w35298 = w35215 & w35297;
assign w35299 = ~w35181 & ~w35199;
assign w35300 = ~w35298 & w35299;
assign w35301 = ~w35121 & ~w35300;
assign w35302 = ~w35127 & ~w35297;
assign w35303 = ~w35160 & ~w35228;
assign w35304 = w35244 & w35303;
assign w35305 = ~w35242 & ~w35304;
assign w35306 = (w35121 & w35302) | (w35121 & w66103) | (w35302 & w66103);
assign w35307 = ~w35294 & ~w35306;
assign w35308 = ~w35301 & w35307;
assign w35309 = pi1852 & w35308;
assign w35310 = ~pi1852 & ~w35308;
assign w35311 = ~w35309 & ~w35310;
assign w35312 = (~w34943 & w34947) | (~w34943 & w66104) | (w34947 & w66104);
assign w35313 = ~w34444 & w34872;
assign w35314 = ~w34421 & ~w35313;
assign w35315 = w34440 & ~w35314;
assign w35316 = w34437 & ~w34458;
assign w35317 = ~w34381 & ~w35316;
assign w35318 = (~w35313 & ~w34870) | (~w35313 & w66105) | (~w34870 & w66105);
assign w35319 = ~w35317 & w35318;
assign w35320 = ~w34416 & ~w35319;
assign w35321 = w34408 & w34876;
assign w35322 = ~w34435 & w34451;
assign w35323 = ~w34871 & w35322;
assign w35324 = ~w34431 & ~w34873;
assign w35325 = ~w35321 & w35324;
assign w35326 = (w34416 & w35323) | (w34416 & w66106) | (w35323 & w66106);
assign w35327 = ~w35312 & ~w35315;
assign w35328 = ~w35320 & ~w35326;
assign w35329 = w35327 & w35328;
assign w35330 = ~pi1847 & ~w35329;
assign w35331 = pi1847 & w35329;
assign w35332 = ~w35330 & ~w35331;
assign w35333 = w34508 & w34526;
assign w35334 = w34489 & w35007;
assign w35335 = w34517 & w34535;
assign w35336 = ~w35000 & ~w35335;
assign w35337 = ~w34506 & ~w35334;
assign w35338 = ~w35336 & w35337;
assign w35339 = w34476 & ~w35338;
assign w35340 = (~w34521 & w35105) | (~w34521 & w66107) | (w35105 & w66107);
assign w35341 = w34517 & ~w35340;
assign w35342 = w34520 & w34993;
assign w35343 = ~w34502 & ~w34992;
assign w35344 = ~w34489 & w35011;
assign w35345 = ~w35343 & ~w35344;
assign w35346 = ~w35342 & ~w35345;
assign w35347 = ~w34476 & ~w35346;
assign w35348 = ~w35333 & ~w35341;
assign w35349 = ~w35347 & w35348;
assign w35350 = ~w35339 & w35349;
assign w35351 = ~pi1853 & ~w35350;
assign w35352 = pi1853 & w35350;
assign w35353 = ~w35351 & ~w35352;
assign w35354 = ~pi6293 & pi9040;
assign w35355 = ~pi6261 & ~pi9040;
assign w35356 = ~w35354 & ~w35355;
assign w35357 = pi1879 & ~w35356;
assign w35358 = ~pi1879 & w35356;
assign w35359 = ~w35357 & ~w35358;
assign w35360 = ~pi6369 & pi9040;
assign w35361 = ~pi6304 & ~pi9040;
assign w35362 = ~w35360 & ~w35361;
assign w35363 = pi1848 & ~w35362;
assign w35364 = ~pi1848 & w35362;
assign w35365 = ~w35363 & ~w35364;
assign w35366 = w35359 & ~w35365;
assign w35367 = ~pi6403 & pi9040;
assign w35368 = ~pi6311 & ~pi9040;
assign w35369 = ~w35367 & ~w35368;
assign w35370 = pi1861 & ~w35369;
assign w35371 = ~pi1861 & w35369;
assign w35372 = ~w35370 & ~w35371;
assign w35373 = ~pi6286 & pi9040;
assign w35374 = ~pi6372 & ~pi9040;
assign w35375 = ~w35373 & ~w35374;
assign w35376 = pi1866 & ~w35375;
assign w35377 = ~pi1866 & w35375;
assign w35378 = ~w35376 & ~w35377;
assign w35379 = w35372 & w35378;
assign w35380 = w35366 & w35379;
assign w35381 = w35365 & w35372;
assign w35382 = ~pi6372 & pi9040;
assign w35383 = ~pi6397 & ~pi9040;
assign w35384 = ~w35382 & ~w35383;
assign w35385 = pi1855 & ~w35384;
assign w35386 = ~pi1855 & w35384;
assign w35387 = ~w35385 & ~w35386;
assign w35388 = ~w35359 & ~w35387;
assign w35389 = w35381 & w35388;
assign w35390 = w35378 & w35387;
assign w35391 = ~w35359 & ~w35372;
assign w35392 = w35390 & w35391;
assign w35393 = ~w35359 & w35365;
assign w35394 = ~w35372 & ~w35387;
assign w35395 = ~w35366 & w35394;
assign w35396 = w35381 & w35387;
assign w35397 = ~w35395 & ~w35396;
assign w35398 = ~w35393 & ~w35397;
assign w35399 = w35359 & w35387;
assign w35400 = (w35378 & ~w35399) | (w35378 & w66108) | (~w35399 & w66108);
assign w35401 = ~w35398 & w35400;
assign w35402 = w35372 & w35387;
assign w35403 = w35359 & ~w35387;
assign w35404 = ~w35402 & ~w35403;
assign w35405 = ~w35365 & ~w35404;
assign w35406 = w35404 & w66109;
assign w35407 = (~w35378 & w35404) | (~w35378 & w66110) | (w35404 & w66110);
assign w35408 = ~w35406 & w35407;
assign w35409 = ~pi6311 & pi9040;
assign w35410 = ~pi6296 & ~pi9040;
assign w35411 = ~w35409 & ~w35410;
assign w35412 = pi1885 & ~w35411;
assign w35413 = ~pi1885 & w35411;
assign w35414 = ~w35412 & ~w35413;
assign w35415 = ~w35389 & ~w35414;
assign w35416 = ~w35392 & w35415;
assign w35417 = (w35416 & w35401) | (w35416 & w66111) | (w35401 & w66111);
assign w35418 = ~w35365 & w35399;
assign w35419 = w35378 & ~w35418;
assign w35420 = w35359 & w35397;
assign w35421 = w35419 & w35420;
assign w35422 = ~w35378 & ~w35397;
assign w35423 = ~w35365 & ~w35372;
assign w35424 = w35387 & w35423;
assign w35425 = w35423 & w63903;
assign w35426 = w35387 & w35393;
assign w35427 = w35393 & w35402;
assign w35428 = ~w35425 & ~w35427;
assign w35429 = ~w35381 & w35388;
assign w35430 = ~w35423 & w35429;
assign w35431 = w35428 & ~w35430;
assign w35432 = (w35414 & w35397) | (w35414 & w66112) | (w35397 & w66112);
assign w35433 = ~w35421 & w66113;
assign w35434 = ~w35417 & ~w35433;
assign w35435 = ~w35359 & w35424;
assign w35436 = ~w35380 & ~w35435;
assign w35437 = ~w35434 & w35436;
assign w35438 = ~pi1891 & w35437;
assign w35439 = pi1891 & ~w35437;
assign w35440 = ~w35438 & ~w35439;
assign w35441 = ~pi6304 & pi9040;
assign w35442 = ~pi6278 & ~pi9040;
assign w35443 = ~w35441 & ~w35442;
assign w35444 = pi1849 & ~w35443;
assign w35445 = ~pi1849 & w35443;
assign w35446 = ~w35444 & ~w35445;
assign w35447 = ~pi6300 & pi9040;
assign w35448 = ~pi6467 & ~pi9040;
assign w35449 = ~w35447 & ~w35448;
assign w35450 = pi1864 & ~w35449;
assign w35451 = ~pi1864 & w35449;
assign w35452 = ~w35450 & ~w35451;
assign w35453 = ~pi6314 & pi9040;
assign w35454 = ~pi6286 & ~pi9040;
assign w35455 = ~w35453 & ~w35454;
assign w35456 = pi1873 & ~w35455;
assign w35457 = ~pi1873 & w35455;
assign w35458 = ~w35456 & ~w35457;
assign w35459 = ~w35452 & w35458;
assign w35460 = ~pi6296 & pi9040;
assign w35461 = ~pi6322 & ~pi9040;
assign w35462 = ~w35460 & ~w35461;
assign w35463 = pi1857 & ~w35462;
assign w35464 = ~pi1857 & w35462;
assign w35465 = ~w35463 & ~w35464;
assign w35466 = w35459 & ~w35465;
assign w35467 = ~pi6396 & pi9040;
assign w35468 = ~pi6291 & ~pi9040;
assign w35469 = ~w35467 & ~w35468;
assign w35470 = pi1887 & ~w35469;
assign w35471 = ~pi1887 & w35469;
assign w35472 = ~w35470 & ~w35471;
assign w35473 = w35459 & w63904;
assign w35474 = w35452 & w35458;
assign w35475 = ~w35452 & w35472;
assign w35476 = ~w35458 & ~w35472;
assign w35477 = ~w35465 & ~w35472;
assign w35478 = w35465 & w35472;
assign w35479 = ~w35477 & ~w35478;
assign w35480 = ~w35475 & ~w35476;
assign w35481 = w35479 & w35480;
assign w35482 = ~w35474 & w35481;
assign w35483 = ~w35452 & ~w35458;
assign w35484 = w35477 & w35483;
assign w35485 = ~w35473 & ~w35484;
assign w35486 = ~w35482 & w35485;
assign w35487 = w35446 & ~w35486;
assign w35488 = ~w35446 & w35452;
assign w35489 = w35465 & ~w35472;
assign w35490 = ~w35458 & w35489;
assign w35491 = w35488 & w35490;
assign w35492 = ~w35446 & ~w35479;
assign w35493 = ~w35452 & w35492;
assign w35494 = w35452 & ~w35458;
assign w35495 = ~w35489 & ~w35494;
assign w35496 = w35465 & w35494;
assign w35497 = (w35446 & ~w35494) | (w35446 & w66114) | (~w35494 & w66114);
assign w35498 = w35446 & ~w35476;
assign w35499 = ~w35497 & ~w35498;
assign w35500 = ~w35495 & ~w35499;
assign w35501 = ~w35465 & w35474;
assign w35502 = w35472 & w35501;
assign w35503 = ~pi6466 & pi9040;
assign w35504 = ~pi6300 & ~pi9040;
assign w35505 = ~w35503 & ~w35504;
assign w35506 = pi1881 & ~w35505;
assign w35507 = ~pi1881 & w35505;
assign w35508 = ~w35506 & ~w35507;
assign w35509 = ~w35502 & w35508;
assign w35510 = ~w35493 & w35509;
assign w35511 = ~w35500 & w35510;
assign w35512 = w35478 & w35483;
assign w35513 = w35446 & ~w35512;
assign w35514 = ~w35466 & w35513;
assign w35515 = ~w35458 & ~w35465;
assign w35516 = w35472 & w35515;
assign w35517 = ~w35446 & ~w35474;
assign w35518 = ~w35516 & w35517;
assign w35519 = w35472 & ~w35474;
assign w35520 = w35465 & ~w35519;
assign w35521 = ~w35500 & w35520;
assign w35522 = (~w35508 & w35514) | (~w35508 & w66115) | (w35514 & w66115);
assign w35523 = ~w35521 & w35522;
assign w35524 = ~w35511 & ~w35523;
assign w35525 = ~w35487 & ~w35491;
assign w35526 = ~w35524 & w35525;
assign w35527 = pi1888 & w35526;
assign w35528 = ~pi1888 & ~w35526;
assign w35529 = ~w35527 & ~w35528;
assign w35530 = w35379 & w35388;
assign w35531 = ~w35394 & ~w35403;
assign w35532 = w35359 & w35394;
assign w35533 = ~w35531 & ~w35532;
assign w35534 = w35365 & w35533;
assign w35535 = w35372 & ~w35390;
assign w35536 = w35366 & ~w35535;
assign w35537 = ~w35530 & ~w35536;
assign w35538 = ~w35534 & w35537;
assign w35539 = ~w35365 & w35372;
assign w35540 = ~w35387 & ~w35539;
assign w35541 = ~w35365 & w35402;
assign w35542 = ~w35414 & ~w35541;
assign w35543 = ~w35359 & ~w35390;
assign w35544 = ~w35540 & w35543;
assign w35545 = ~w35542 & w35544;
assign w35546 = w35399 & w35423;
assign w35547 = ~w35530 & ~w35546;
assign w35548 = ~w35431 & ~w35547;
assign w35549 = w35419 & ~w35530;
assign w35550 = ~w35533 & w35549;
assign w35551 = ~w35378 & w35533;
assign w35552 = w35359 & w35396;
assign w35553 = ~w35551 & ~w35552;
assign w35554 = ~w35550 & w35553;
assign w35555 = ~w35414 & ~w35554;
assign w35556 = (~w35545 & w35538) | (~w35545 & w66116) | (w35538 & w66116);
assign w35557 = ~w35548 & w35556;
assign w35558 = ~w35555 & w35557;
assign w35559 = ~pi1907 & ~w35558;
assign w35560 = pi1907 & w35558;
assign w35561 = ~w35559 & ~w35560;
assign w35562 = ~pi6322 & pi9040;
assign w35563 = ~pi6260 & ~pi9040;
assign w35564 = ~w35562 & ~w35563;
assign w35565 = pi1883 & ~w35564;
assign w35566 = ~pi1883 & w35564;
assign w35567 = ~w35565 & ~w35566;
assign w35568 = ~pi6467 & pi9040;
assign w35569 = ~pi6293 & ~pi9040;
assign w35570 = ~w35568 & ~w35569;
assign w35571 = pi1879 & ~w35570;
assign w35572 = ~pi1879 & w35570;
assign w35573 = ~w35571 & ~w35572;
assign w35574 = ~pi6375 & pi9040;
assign w35575 = ~pi6277 & ~pi9040;
assign w35576 = ~w35574 & ~w35575;
assign w35577 = pi1856 & ~w35576;
assign w35578 = ~pi1856 & w35576;
assign w35579 = ~w35577 & ~w35578;
assign w35580 = w35573 & w35579;
assign w35581 = ~pi6395 & pi9040;
assign w35582 = ~pi6402 & ~pi9040;
assign w35583 = ~w35581 & ~w35582;
assign w35584 = pi1882 & ~w35583;
assign w35585 = ~pi1882 & w35583;
assign w35586 = ~w35584 & ~w35585;
assign w35587 = w35580 & w35586;
assign w35588 = ~w35567 & w35587;
assign w35589 = ~w35567 & ~w35586;
assign w35590 = w35579 & w35589;
assign w35591 = ~pi6277 & pi9040;
assign w35592 = ~pi6396 & ~pi9040;
assign w35593 = ~w35591 & ~w35592;
assign w35594 = pi1876 & ~w35593;
assign w35595 = ~pi1876 & w35593;
assign w35596 = ~w35594 & ~w35595;
assign w35597 = ~w35590 & w35596;
assign w35598 = ~w35573 & ~w35586;
assign w35599 = w35567 & ~w35579;
assign w35600 = w35598 & w35599;
assign w35601 = ~w35573 & w35586;
assign w35602 = w35567 & w35579;
assign w35603 = w35601 & w35602;
assign w35604 = ~w35600 & ~w35603;
assign w35605 = w35573 & w35589;
assign w35606 = w35604 & ~w35605;
assign w35607 = w35597 & ~w35606;
assign w35608 = ~pi6315 & pi9040;
assign w35609 = pi6314 & ~pi9040;
assign w35610 = ~w35608 & ~w35609;
assign w35611 = pi1855 & ~w35610;
assign w35612 = ~pi1855 & w35610;
assign w35613 = ~w35611 & ~w35612;
assign w35614 = w35573 & ~w35586;
assign w35615 = w35602 & w35614;
assign w35616 = ~w35567 & ~w35579;
assign w35617 = ~w35602 & ~w35616;
assign w35618 = ~w35586 & ~w35596;
assign w35619 = ~w35617 & w35618;
assign w35620 = w35586 & ~w35596;
assign w35621 = ~w35573 & ~w35579;
assign w35622 = w35620 & w35621;
assign w35623 = w35579 & w35596;
assign w35624 = ~w35567 & ~w35573;
assign w35625 = w35623 & w35624;
assign w35626 = ~w35615 & ~w35622;
assign w35627 = ~w35625 & w35626;
assign w35628 = ~w35619 & w35627;
assign w35629 = w35613 & ~w35628;
assign w35630 = w35599 & w35620;
assign w35631 = ~w35567 & w35580;
assign w35632 = ~w35603 & ~w35631;
assign w35633 = w35598 & w35602;
assign w35634 = ~w35579 & ~w35586;
assign w35635 = w35601 & w35616;
assign w35636 = ~w35587 & ~w35635;
assign w35637 = ~w35633 & ~w35634;
assign w35638 = w35636 & w35637;
assign w35639 = w35596 & ~w35638;
assign w35640 = w35573 & w35586;
assign w35641 = ~w35579 & w35640;
assign w35642 = ~w35590 & ~w35641;
assign w35643 = ~w35596 & ~w35642;
assign w35644 = w35632 & ~w35643;
assign w35645 = ~w35639 & w35644;
assign w35646 = ~w35613 & ~w35645;
assign w35647 = ~w35588 & ~w35630;
assign w35648 = ~w35607 & w35647;
assign w35649 = ~w35629 & w35648;
assign w35650 = ~w35646 & w35649;
assign w35651 = pi1895 & w35650;
assign w35652 = ~pi1895 & ~w35650;
assign w35653 = ~w35651 & ~w35652;
assign w35654 = ~pi6295 & pi9040;
assign w35655 = ~pi6382 & ~pi9040;
assign w35656 = ~w35654 & ~w35655;
assign w35657 = pi1873 & ~w35656;
assign w35658 = ~pi1873 & w35656;
assign w35659 = ~w35657 & ~w35658;
assign w35660 = ~pi6287 & pi9040;
assign w35661 = ~pi6306 & ~pi9040;
assign w35662 = ~w35660 & ~w35661;
assign w35663 = pi1858 & ~w35662;
assign w35664 = ~pi1858 & w35662;
assign w35665 = ~w35663 & ~w35664;
assign w35666 = ~w35659 & ~w35665;
assign w35667 = ~pi6533 & pi9040;
assign w35668 = ~pi6282 & ~pi9040;
assign w35669 = ~w35667 & ~w35668;
assign w35670 = pi1881 & ~w35669;
assign w35671 = ~pi1881 & w35669;
assign w35672 = ~w35670 & ~w35671;
assign w35673 = ~w35666 & ~w35672;
assign w35674 = ~pi6367 & pi9040;
assign w35675 = ~pi6531 & ~pi9040;
assign w35676 = ~w35674 & ~w35675;
assign w35677 = pi1843 & ~w35676;
assign w35678 = ~pi1843 & w35676;
assign w35679 = ~w35677 & ~w35678;
assign w35680 = ~w35659 & w35679;
assign w35681 = ~w35665 & w35672;
assign w35682 = w35680 & w35681;
assign w35683 = ~w35673 & ~w35682;
assign w35684 = ~pi6306 & pi9040;
assign w35685 = ~pi6319 & ~pi9040;
assign w35686 = ~w35684 & ~w35685;
assign w35687 = pi1878 & ~w35686;
assign w35688 = ~pi1878 & w35686;
assign w35689 = ~w35687 & ~w35688;
assign w35690 = ~w35683 & w35689;
assign w35691 = ~w35672 & ~w35679;
assign w35692 = w35672 & w35679;
assign w35693 = ~w35691 & ~w35692;
assign w35694 = ~w35659 & w35665;
assign w35695 = ~w35693 & w35694;
assign w35696 = w35659 & w35689;
assign w35697 = w35665 & w35693;
assign w35698 = w35693 & w63905;
assign w35699 = ~w35659 & w35672;
assign w35700 = w35665 & ~w35699;
assign w35701 = ~w35681 & ~w35689;
assign w35702 = ~w35680 & w35701;
assign w35703 = w35672 & ~w35689;
assign w35704 = w35659 & w35703;
assign w35705 = w35665 & w35679;
assign w35706 = w35659 & w35705;
assign w35707 = ~w35704 & ~w35706;
assign w35708 = ~w35665 & ~w35679;
assign w35709 = ~w35659 & w35708;
assign w35710 = w35707 & ~w35709;
assign w35711 = ~w35665 & ~w35693;
assign w35712 = (~w35702 & ~w35710) | (~w35702 & w63906) | (~w35710 & w63906);
assign w35713 = (~w35698 & w35712) | (~w35698 & w66117) | (w35712 & w66117);
assign w35714 = ~pi6263 & pi9040;
assign w35715 = ~pi6533 & ~pi9040;
assign w35716 = ~w35714 & ~w35715;
assign w35717 = pi1874 & ~w35716;
assign w35718 = ~pi1874 & w35716;
assign w35719 = ~w35717 & ~w35718;
assign w35720 = ~w35713 & ~w35719;
assign w35721 = w35659 & ~w35679;
assign w35722 = ~w35665 & w35721;
assign w35723 = ~w35680 & ~w35721;
assign w35724 = ~w35672 & ~w35723;
assign w35725 = w35672 & w35723;
assign w35726 = ~w35724 & ~w35725;
assign w35727 = w35665 & ~w35726;
assign w35728 = (~w35722 & w35726) | (~w35722 & w66118) | (w35726 & w66118);
assign w35729 = ~w35689 & ~w35728;
assign w35730 = ~w35672 & w35689;
assign w35731 = w35679 & w35730;
assign w35732 = ~w35679 & w35699;
assign w35733 = ~w35731 & ~w35732;
assign w35734 = ~w35665 & ~w35733;
assign w35735 = w35680 & w35689;
assign w35736 = w35691 & w35696;
assign w35737 = ~w35735 & ~w35736;
assign w35738 = ~w35708 & ~w35737;
assign w35739 = ~w35659 & ~w35672;
assign w35740 = ~w35708 & w35739;
assign w35741 = ~w35704 & ~w35740;
assign w35742 = ~w35734 & w35741;
assign w35743 = ~w35738 & w35742;
assign w35744 = (w35719 & ~w35742) | (w35719 & w63907) | (~w35742 & w63907);
assign w35745 = ~w35665 & w35689;
assign w35746 = w35699 & w35745;
assign w35747 = (~w35746 & ~w35690) | (~w35746 & w66119) | (~w35690 & w66119);
assign w35748 = ~w35744 & w35747;
assign w35749 = ~w35729 & w35748;
assign w35750 = (~pi1897 & ~w35749) | (~pi1897 & w66120) | (~w35749 & w66120);
assign w35751 = w35749 & w66121;
assign w35752 = ~w35750 & ~w35751;
assign w35753 = ~pi6290 & pi9040;
assign w35754 = ~pi6395 & ~pi9040;
assign w35755 = ~w35753 & ~w35754;
assign w35756 = pi1880 & ~w35755;
assign w35757 = ~pi1880 & w35755;
assign w35758 = ~w35756 & ~w35757;
assign w35759 = ~pi6261 & pi9040;
assign w35760 = ~pi6288 & ~pi9040;
assign w35761 = ~w35759 & ~w35760;
assign w35762 = pi1864 & ~w35761;
assign w35763 = ~pi1864 & w35761;
assign w35764 = ~w35762 & ~w35763;
assign w35765 = ~w35758 & w35764;
assign w35766 = ~pi6271 & pi9040;
assign w35767 = ~pi6375 & ~pi9040;
assign w35768 = ~w35766 & ~w35767;
assign w35769 = pi1862 & ~w35768;
assign w35770 = ~pi1862 & w35768;
assign w35771 = ~w35769 & ~w35770;
assign w35772 = ~pi6278 & pi9040;
assign w35773 = ~pi6270 & ~pi9040;
assign w35774 = ~w35772 & ~w35773;
assign w35775 = pi1861 & ~w35774;
assign w35776 = ~pi1861 & w35774;
assign w35777 = ~w35775 & ~w35776;
assign w35778 = ~w35771 & ~w35777;
assign w35779 = ~pi6260 & pi9040;
assign w35780 = ~pi6466 & ~pi9040;
assign w35781 = ~w35779 & ~w35780;
assign w35782 = pi1885 & ~w35781;
assign w35783 = ~pi1885 & w35781;
assign w35784 = ~w35782 & ~w35783;
assign w35785 = w35778 & w35784;
assign w35786 = ~w35765 & w35785;
assign w35787 = w35764 & ~w35771;
assign w35788 = ~w35777 & ~w35784;
assign w35789 = w35777 & w35784;
assign w35790 = ~w35788 & ~w35789;
assign w35791 = ~w35787 & ~w35790;
assign w35792 = ~w35764 & w35771;
assign w35793 = ~w35787 & ~w35792;
assign w35794 = w35790 & ~w35793;
assign w35795 = w35771 & w35777;
assign w35796 = w35794 & ~w35795;
assign w35797 = ~w35791 & ~w35796;
assign w35798 = (~w35758 & w35796) | (~w35758 & w63908) | (w35796 & w63908);
assign w35799 = ~w35764 & w35777;
assign w35800 = w35771 & ~w35784;
assign w35801 = ~w35764 & ~w35777;
assign w35802 = w35800 & w35801;
assign w35803 = ~w35799 & ~w35802;
assign w35804 = (w35796 & w66122) | (w35796 & w66123) | (w66122 & w66123);
assign w35805 = ~w35786 & ~w35804;
assign w35806 = ~pi6270 & pi9040;
assign w35807 = pi6315 & ~pi9040;
assign w35808 = ~w35806 & ~w35807;
assign w35809 = pi1857 & ~w35808;
assign w35810 = ~pi1857 & w35808;
assign w35811 = ~w35809 & ~w35810;
assign w35812 = ~w35805 & ~w35811;
assign w35813 = w35758 & ~w35802;
assign w35814 = w35764 & ~w35777;
assign w35815 = ~w35799 & ~w35814;
assign w35816 = w35800 & ~w35815;
assign w35817 = ~w35801 & ~w35816;
assign w35818 = w35813 & ~w35817;
assign w35819 = w35788 & w35793;
assign w35820 = ~w35764 & w35784;
assign w35821 = w35764 & ~w35784;
assign w35822 = ~w35820 & ~w35821;
assign w35823 = w35777 & ~w35822;
assign w35824 = ~w35785 & ~w35823;
assign w35825 = (w35765 & w35823) | (w35765 & w66124) | (w35823 & w66124);
assign w35826 = ~w35778 & ~w35795;
assign w35827 = w35758 & w35784;
assign w35828 = ~w35799 & w35827;
assign w35829 = w35826 & w35828;
assign w35830 = ~w35819 & ~w35829;
assign w35831 = ~w35825 & w35830;
assign w35832 = w35811 & ~w35831;
assign w35833 = ~w35771 & w35784;
assign w35834 = w35758 & w35814;
assign w35835 = ~w35758 & w35777;
assign w35836 = w35764 & ~w35811;
assign w35837 = ~w35835 & ~w35836;
assign w35838 = ~w35800 & ~w35833;
assign w35839 = ~w35834 & w35838;
assign w35840 = ~w35837 & w35839;
assign w35841 = ~w35818 & ~w35840;
assign w35842 = ~w35832 & w35841;
assign w35843 = ~w35812 & w35842;
assign w35844 = pi1889 & ~w35843;
assign w35845 = ~pi1889 & w35843;
assign w35846 = ~w35844 & ~w35845;
assign w35847 = ~w35399 & ~w35539;
assign w35848 = ~w35402 & ~w35847;
assign w35849 = (w35378 & w35848) | (w35378 & w66125) | (w35848 & w66125);
assign w35850 = ~w35435 & ~w35849;
assign w35851 = ~w35414 & ~w35850;
assign w35852 = w35359 & w35381;
assign w35853 = (~w35852 & ~w35405) | (~w35852 & w66126) | (~w35405 & w66126);
assign w35854 = w35414 & ~w35853;
assign w35855 = (w35378 & w35534) | (w35378 & w66127) | (w35534 & w66127);
assign w35856 = ~w35365 & ~w35387;
assign w35857 = ~w35546 & ~w35856;
assign w35858 = w35414 & w35857;
assign w35859 = ~w35389 & ~w35532;
assign w35860 = w35542 & w35859;
assign w35861 = ~w35858 & ~w35860;
assign w35862 = ~w35426 & ~w35856;
assign w35863 = ~w35372 & ~w35862;
assign w35864 = ~w35552 & ~w35863;
assign w35865 = ~w35861 & w35864;
assign w35866 = ~w35378 & ~w35865;
assign w35867 = ~w35854 & ~w35855;
assign w35868 = ~w35851 & w35867;
assign w35869 = ~w35866 & w35868;
assign w35870 = ~pi1898 & w35869;
assign w35871 = pi1898 & ~w35869;
assign w35872 = ~w35870 & ~w35871;
assign w35873 = w35422 & ~w35857;
assign w35874 = ~w35366 & ~w35396;
assign w35875 = w35550 & ~w35874;
assign w35876 = (w35378 & w35426) | (w35378 & w66128) | (w35426 & w66128);
assign w35877 = w35365 & w35403;
assign w35878 = ~w35418 & ~w35877;
assign w35879 = ~w35378 & ~w35878;
assign w35880 = ~w35414 & w35428;
assign w35881 = w35547 & ~w35876;
assign w35882 = ~w35879 & w35881;
assign w35883 = w35880 & w35882;
assign w35884 = w35400 & ~w35877;
assign w35885 = ~w35435 & w35884;
assign w35886 = ~w35388 & ~w35399;
assign w35887 = w35539 & w35886;
assign w35888 = (~w35378 & ~w35404) | (~w35378 & w66129) | (~w35404 & w66129);
assign w35889 = ~w35887 & w35888;
assign w35890 = ~w35885 & ~w35889;
assign w35891 = (w35414 & w35431) | (w35414 & w66130) | (w35431 & w66130);
assign w35892 = ~w35890 & w35891;
assign w35893 = ~w35883 & ~w35892;
assign w35894 = ~w35873 & ~w35875;
assign w35895 = ~w35893 & w35894;
assign w35896 = pi1890 & ~w35895;
assign w35897 = ~pi1890 & w35895;
assign w35898 = ~w35896 & ~w35897;
assign w35899 = w35696 & ~w35743;
assign w35900 = w35659 & ~w35708;
assign w35901 = ~w35689 & ~w35900;
assign w35902 = ~w35693 & w35901;
assign w35903 = w35689 & w35725;
assign w35904 = w35697 & ~w35723;
assign w35905 = ~w35719 & ~w35902;
assign w35906 = ~w35903 & ~w35904;
assign w35907 = w35905 & w35906;
assign w35908 = ~w35673 & w35701;
assign w35909 = w35681 & w35721;
assign w35910 = w35719 & ~w35909;
assign w35911 = ~w35706 & ~w35908;
assign w35912 = w35910 & w35911;
assign w35913 = ~w35690 & w35912;
assign w35914 = ~w35907 & ~w35913;
assign w35915 = ~w35899 & ~w35914;
assign w35916 = ~pi1905 & w35915;
assign w35917 = pi1905 & ~w35915;
assign w35918 = ~w35916 & ~w35917;
assign w35919 = ~pi6382 & pi9040;
assign w35920 = ~pi6292 & ~pi9040;
assign w35921 = ~w35919 & ~w35920;
assign w35922 = pi1856 & ~w35921;
assign w35923 = ~pi1856 & w35921;
assign w35924 = ~w35922 & ~w35923;
assign w35925 = ~pi6309 & pi9040;
assign w35926 = ~pi6367 & ~pi9040;
assign w35927 = ~w35925 & ~w35926;
assign w35928 = pi1884 & ~w35927;
assign w35929 = ~pi1884 & w35927;
assign w35930 = ~w35928 & ~w35929;
assign w35931 = ~w35924 & w35930;
assign w35932 = ~pi6535 & pi9040;
assign w35933 = ~pi6263 & ~pi9040;
assign w35934 = ~w35932 & ~w35933;
assign w35935 = pi1860 & ~w35934;
assign w35936 = ~pi1860 & w35934;
assign w35937 = ~w35935 & ~w35936;
assign w35938 = ~pi6282 & pi9040;
assign w35939 = ~pi6401 & ~pi9040;
assign w35940 = ~w35938 & ~w35939;
assign w35941 = pi1872 & ~w35940;
assign w35942 = ~pi1872 & w35940;
assign w35943 = ~w35941 & ~w35942;
assign w35944 = ~w35937 & w35943;
assign w35945 = w35937 & ~w35943;
assign w35946 = ~w35944 & ~w35945;
assign w35947 = w35931 & w35946;
assign w35948 = ~pi6308 & pi9040;
assign w35949 = ~pi6309 & ~pi9040;
assign w35950 = ~w35948 & ~w35949;
assign w35951 = pi1875 & ~w35950;
assign w35952 = ~pi1875 & w35950;
assign w35953 = ~w35951 & ~w35952;
assign w35954 = w35947 & ~w35953;
assign w35955 = w35944 & w35953;
assign w35956 = w35930 & w35955;
assign w35957 = ~w35930 & w35953;
assign w35958 = w35937 & w35953;
assign w35959 = w35930 & ~w35958;
assign w35960 = w35945 & ~w35953;
assign w35961 = w35959 & ~w35960;
assign w35962 = w35924 & ~w35957;
assign w35963 = ~w35961 & w35962;
assign w35964 = w35930 & ~w35953;
assign w35965 = ~w35924 & ~w35937;
assign w35966 = w35964 & w35965;
assign w35967 = w35937 & w35943;
assign w35968 = ~w35924 & ~w35930;
assign w35969 = w35967 & w35968;
assign w35970 = ~pi6312 & pi9040;
assign w35971 = ~pi6284 & ~pi9040;
assign w35972 = ~w35970 & ~w35971;
assign w35973 = pi1882 & ~w35972;
assign w35974 = ~pi1882 & w35972;
assign w35975 = ~w35973 & ~w35974;
assign w35976 = ~w35937 & ~w35943;
assign w35977 = ~w35924 & ~w35953;
assign w35978 = w35976 & w35977;
assign w35979 = ~w35924 & w35955;
assign w35980 = ~w35975 & ~w35978;
assign w35981 = ~w35979 & w35980;
assign w35982 = ~w35966 & ~w35969;
assign w35983 = ~w35956 & w35982;
assign w35984 = ~w35963 & w35983;
assign w35985 = w35981 & w35984;
assign w35986 = w35924 & w35953;
assign w35987 = w35946 & w35986;
assign w35988 = ~w35937 & ~w35953;
assign w35989 = w35943 & w35988;
assign w35990 = w35968 & w35989;
assign w35991 = w35931 & w35958;
assign w35992 = w35924 & w35930;
assign w35993 = w35988 & w35992;
assign w35994 = ~w35958 & ~w35988;
assign w35995 = ~w35930 & ~w35943;
assign w35996 = w35994 & w35995;
assign w35997 = w35975 & ~w35991;
assign w35998 = ~w35993 & w35997;
assign w35999 = ~w35987 & ~w35990;
assign w36000 = ~w35996 & w35999;
assign w36001 = w35998 & w36000;
assign w36002 = ~w35985 & ~w36001;
assign w36003 = ~w35943 & w35991;
assign w36004 = w35976 & w35986;
assign w36005 = ~w35930 & w36004;
assign w36006 = ~w36003 & ~w36005;
assign w36007 = ~w35954 & w36006;
assign w36008 = ~w36002 & w36007;
assign w36009 = ~pi1892 & w36008;
assign w36010 = pi1892 & ~w36008;
assign w36011 = ~w36009 & ~w36010;
assign w36012 = ~pi6272 & pi9040;
assign w36013 = ~pi6281 & ~pi9040;
assign w36014 = ~w36012 & ~w36013;
assign w36015 = pi1868 & ~w36014;
assign w36016 = ~pi1868 & w36014;
assign w36017 = ~w36015 & ~w36016;
assign w36018 = ~pi6289 & pi9040;
assign w36019 = ~pi6312 & ~pi9040;
assign w36020 = ~w36018 & ~w36019;
assign w36021 = pi1843 & ~w36020;
assign w36022 = ~pi1843 & w36020;
assign w36023 = ~w36021 & ~w36022;
assign w36024 = ~pi6285 & pi9040;
assign w36025 = ~pi6374 & ~pi9040;
assign w36026 = ~w36024 & ~w36025;
assign w36027 = pi1869 & ~w36026;
assign w36028 = ~pi1869 & w36026;
assign w36029 = ~w36027 & ~w36028;
assign w36030 = ~w36023 & w36029;
assign w36031 = w36023 & ~w36029;
assign w36032 = ~w36030 & ~w36031;
assign w36033 = ~pi6268 & pi9040;
assign w36034 = ~pi6535 & ~pi9040;
assign w36035 = ~w36033 & ~w36034;
assign w36036 = pi1874 & ~w36035;
assign w36037 = ~pi1874 & w36035;
assign w36038 = ~w36036 & ~w36037;
assign w36039 = w36029 & w36038;
assign w36040 = ~w36032 & ~w36039;
assign w36041 = ~pi6292 & pi9040;
assign w36042 = ~pi6289 & ~pi9040;
assign w36043 = ~w36041 & ~w36042;
assign w36044 = pi1886 & ~w36043;
assign w36045 = ~pi1886 & w36043;
assign w36046 = ~w36044 & ~w36045;
assign w36047 = w36040 & ~w36046;
assign w36048 = ~pi6281 & pi9040;
assign w36049 = ~pi6307 & ~pi9040;
assign w36050 = ~w36048 & ~w36049;
assign w36051 = pi1877 & ~w36050;
assign w36052 = ~pi1877 & w36050;
assign w36053 = ~w36051 & ~w36052;
assign w36054 = w36023 & w36053;
assign w36055 = ~w36038 & w36046;
assign w36056 = w36054 & ~w36055;
assign w36057 = ~w36029 & ~w36038;
assign w36058 = ~w36023 & ~w36053;
assign w36059 = w36057 & w36058;
assign w36060 = ~w36056 & ~w36059;
assign w36061 = w36029 & ~w36038;
assign w36062 = w36053 & ~w36061;
assign w36063 = w36029 & ~w36046;
assign w36064 = ~w36058 & w36063;
assign w36065 = ~w36062 & ~w36064;
assign w36066 = w36032 & w63909;
assign w36067 = ~w36065 & ~w36066;
assign w36068 = ~w36046 & w36057;
assign w36069 = w36039 & w36046;
assign w36070 = ~w36068 & ~w36069;
assign w36071 = w36067 & ~w36070;
assign w36072 = w36067 & w66131;
assign w36073 = w36030 & w36038;
assign w36074 = ~w36053 & ~w36073;
assign w36075 = w36038 & w36046;
assign w36076 = ~w36030 & ~w36075;
assign w36077 = w36074 & ~w36076;
assign w36078 = ~w36047 & ~w36077;
assign w36079 = ~w36072 & w36078;
assign w36080 = ~w36017 & ~w36079;
assign w36081 = w36023 & ~w36046;
assign w36082 = ~w36057 & w36081;
assign w36083 = ~w36023 & w36046;
assign w36084 = w36057 & w36083;
assign w36085 = ~w36082 & ~w36084;
assign w36086 = w36062 & ~w36085;
assign w36087 = w36023 & w36061;
assign w36088 = ~w36063 & ~w36087;
assign w36089 = ~w36064 & ~w36088;
assign w36090 = ~w36038 & ~w36054;
assign w36091 = w36017 & ~w36090;
assign w36092 = w36089 & ~w36091;
assign w36093 = w36032 & w66132;
assign w36094 = ~w36057 & ~w36073;
assign w36095 = w36046 & ~w36053;
assign w36096 = ~w36094 & w36095;
assign w36097 = w36060 & ~w36093;
assign w36098 = ~w36096 & w36097;
assign w36099 = w36017 & ~w36098;
assign w36100 = ~w36086 & ~w36092;
assign w36101 = ~w36099 & w36100;
assign w36102 = ~w36080 & w36101;
assign w36103 = pi1910 & w36102;
assign w36104 = ~pi1910 & ~w36102;
assign w36105 = ~w36103 & ~w36104;
assign w36106 = w35924 & ~w35930;
assign w36107 = w35945 & w36106;
assign w36108 = w35924 & w35960;
assign w36109 = ~w35943 & w35953;
assign w36110 = ~w35964 & ~w36109;
assign w36111 = w35937 & ~w36110;
assign w36112 = ~w36108 & w36111;
assign w36113 = w35976 & w35992;
assign w36114 = ~w36107 & ~w36113;
assign w36115 = ~w35990 & w36114;
assign w36116 = w35981 & w36115;
assign w36117 = ~w36112 & w36116;
assign w36118 = ~w35964 & ~w35986;
assign w36119 = ~w36108 & ~w36118;
assign w36120 = w35959 & ~w36119;
assign w36121 = w35960 & w35968;
assign w36122 = w35975 & ~w36121;
assign w36123 = w35924 & w35943;
assign w36124 = ~w35994 & w36123;
assign w36125 = ~w35969 & ~w36005;
assign w36126 = ~w36124 & w36125;
assign w36127 = w36122 & w36126;
assign w36128 = ~w36120 & w36127;
assign w36129 = ~w35978 & ~w36124;
assign w36130 = ~w35930 & ~w36129;
assign w36131 = ~w35956 & ~w36003;
assign w36132 = ~w36130 & w36131;
assign w36133 = (w36132 & w36128) | (w36132 & w66133) | (w36128 & w66133);
assign w36134 = ~pi1899 & w36133;
assign w36135 = pi1899 & ~w36133;
assign w36136 = ~w36134 & ~w36135;
assign w36137 = ~w35977 & ~w35989;
assign w36138 = ~w35930 & ~w36137;
assign w36139 = w35924 & ~w35967;
assign w36140 = ~w35976 & ~w36139;
assign w36141 = w35930 & w35953;
assign w36142 = w36140 & w36141;
assign w36143 = ~w35975 & ~w36138;
assign w36144 = ~w36142 & w36143;
assign w36145 = ~w35924 & w35943;
assign w36146 = w35958 & w36145;
assign w36147 = w36106 & ~w36109;
assign w36148 = w35946 & w36147;
assign w36149 = w35965 & ~w36110;
assign w36150 = w35944 & ~w36118;
assign w36151 = w35975 & ~w36146;
assign w36152 = ~w36148 & w36151;
assign w36153 = ~w36149 & ~w36150;
assign w36154 = w36152 & w36153;
assign w36155 = ~w36144 & ~w36154;
assign w36156 = ~w36107 & ~w36149;
assign w36157 = w35957 & ~w36156;
assign w36158 = ~w35960 & ~w36004;
assign w36159 = ~w35992 & w36122;
assign w36160 = ~w36158 & ~w36159;
assign w36161 = ~w36157 & ~w36160;
assign w36162 = ~w36155 & w36161;
assign w36163 = pi1894 & ~w36162;
assign w36164 = ~pi1894 & w36162;
assign w36165 = ~w36163 & ~w36164;
assign w36166 = w36031 & w36075;
assign w36167 = w36030 & w36055;
assign w36168 = ~w36166 & ~w36167;
assign w36169 = ~w36029 & w36083;
assign w36170 = ~w36017 & ~w36087;
assign w36171 = ~w36169 & w36170;
assign w36172 = w36094 & w36171;
assign w36173 = ~w36084 & w36168;
assign w36174 = ~w36172 & w36173;
assign w36175 = ~w36053 & ~w36174;
assign w36176 = ~w36068 & ~w36087;
assign w36177 = w36053 & ~w36176;
assign w36178 = ~w36062 & w36176;
assign w36179 = ~w36032 & w36075;
assign w36180 = ~w36084 & ~w36179;
assign w36181 = ~w36178 & w36180;
assign w36182 = ~w36046 & w36073;
assign w36183 = w36017 & ~w36167;
assign w36184 = ~w36182 & w36183;
assign w36185 = (w36184 & ~w36181) | (w36184 & w66134) | (~w36181 & w66134);
assign w36186 = ~w36017 & ~w36177;
assign w36187 = w36180 & w36186;
assign w36188 = ~w36185 & ~w36187;
assign w36189 = ~w36175 & ~w36188;
assign w36190 = ~pi1896 & w36189;
assign w36191 = pi1896 & ~w36189;
assign w36192 = ~w36190 & ~w36191;
assign w36193 = w35567 & w35622;
assign w36194 = w35567 & w35573;
assign w36195 = w35634 & w36194;
assign w36196 = ~w35633 & ~w36195;
assign w36197 = ~w35632 & ~w35640;
assign w36198 = w35613 & ~w35636;
assign w36199 = w36196 & ~w36197;
assign w36200 = (w35596 & ~w36199) | (w35596 & w66135) | (~w36199 & w66135);
assign w36201 = ~w35596 & w36196;
assign w36202 = ~w35614 & ~w35641;
assign w36203 = w36201 & ~w36202;
assign w36204 = ~w35590 & w35604;
assign w36205 = ~w36203 & w36204;
assign w36206 = w35613 & ~w36205;
assign w36207 = w35589 & w35621;
assign w36208 = ~w35641 & ~w36207;
assign w36209 = w35596 & ~w36208;
assign w36210 = ~w35567 & w35620;
assign w36211 = w36196 & ~w36210;
assign w36212 = ~w36209 & w36211;
assign w36213 = (~w36193 & w36212) | (~w36193 & w66136) | (w36212 & w66136);
assign w36214 = ~w36200 & w36213;
assign w36215 = ~w36206 & w36214;
assign w36216 = pi1901 & ~w36215;
assign w36217 = ~pi1901 & w36215;
assign w36218 = ~w36216 & ~w36217;
assign w36219 = ~pi6368 & pi9040;
assign w36220 = ~pi6295 & ~pi9040;
assign w36221 = ~w36219 & ~w36220;
assign w36222 = pi1854 & ~w36221;
assign w36223 = ~pi1854 & w36221;
assign w36224 = ~w36222 & ~w36223;
assign w36225 = ~pi6401 & pi9040;
assign w36226 = ~pi6280 & ~pi9040;
assign w36227 = ~w36225 & ~w36226;
assign w36228 = pi1871 & ~w36227;
assign w36229 = ~pi1871 & w36227;
assign w36230 = ~w36228 & ~w36229;
assign w36231 = ~pi6374 & pi9040;
assign w36232 = ~pi6313 & ~pi9040;
assign w36233 = ~w36231 & ~w36232;
assign w36234 = pi1868 & ~w36233;
assign w36235 = ~pi1868 & w36233;
assign w36236 = ~w36234 & ~w36235;
assign w36237 = w36230 & w36236;
assign w36238 = ~pi6307 & pi9040;
assign w36239 = ~pi6368 & ~pi9040;
assign w36240 = ~w36238 & ~w36239;
assign w36241 = pi1869 & ~w36240;
assign w36242 = ~pi1869 & w36240;
assign w36243 = ~w36241 & ~w36242;
assign w36244 = w36237 & ~w36243;
assign w36245 = ~w36224 & ~w36244;
assign w36246 = ~pi6313 & pi9040;
assign w36247 = ~pi6272 & ~pi9040;
assign w36248 = ~w36246 & ~w36247;
assign w36249 = pi1875 & ~w36248;
assign w36250 = ~pi1875 & w36248;
assign w36251 = ~w36249 & ~w36250;
assign w36252 = w36230 & ~w36251;
assign w36253 = w36236 & ~w36243;
assign w36254 = ~w36236 & w36243;
assign w36255 = ~w36253 & ~w36254;
assign w36256 = w36252 & w36255;
assign w36257 = w36224 & ~w36256;
assign w36258 = ~w36245 & ~w36257;
assign w36259 = ~pi6284 & pi9040;
assign w36260 = ~pi6287 & ~pi9040;
assign w36261 = ~w36259 & ~w36260;
assign w36262 = pi1860 & ~w36261;
assign w36263 = ~pi1860 & w36261;
assign w36264 = ~w36262 & ~w36263;
assign w36265 = w36251 & ~w36255;
assign w36266 = w36236 & ~w36251;
assign w36267 = w36243 & w36266;
assign w36268 = (w36224 & w36265) | (w36224 & w66137) | (w36265 & w66137);
assign w36269 = ~w36252 & ~w36266;
assign w36270 = ~w36265 & w36269;
assign w36271 = ~w36224 & w36270;
assign w36272 = ~w36230 & ~w36243;
assign w36273 = ~w36236 & w36251;
assign w36274 = ~w36266 & ~w36273;
assign w36275 = w36272 & w36274;
assign w36276 = w36274 & w66138;
assign w36277 = ~w36264 & ~w36276;
assign w36278 = ~w36268 & w36277;
assign w36279 = ~w36271 & w36278;
assign w36280 = w36266 & w36272;
assign w36281 = ~w36230 & w36251;
assign w36282 = w36224 & ~w36230;
assign w36283 = ~w36255 & w36282;
assign w36284 = ~w36281 & ~w36283;
assign w36285 = w36270 & ~w36284;
assign w36286 = ~w36224 & ~w36237;
assign w36287 = ~w36269 & w36286;
assign w36288 = w36230 & w36243;
assign w36289 = w36273 & w36288;
assign w36290 = w36264 & ~w36280;
assign w36291 = ~w36289 & w36290;
assign w36292 = ~w36287 & w36291;
assign w36293 = ~w36285 & w36292;
assign w36294 = ~w36279 & ~w36293;
assign w36295 = ~w36258 & ~w36294;
assign w36296 = ~pi1918 & w36295;
assign w36297 = pi1918 & ~w36295;
assign w36298 = ~w36296 & ~w36297;
assign w36299 = w35765 & w35816;
assign w36300 = ~w35790 & ~w35821;
assign w36301 = w35813 & w36300;
assign w36302 = ~w35794 & w35811;
assign w36303 = ~w36299 & w36302;
assign w36304 = ~w36301 & w36303;
assign w36305 = ~w35758 & w35815;
assign w36306 = ~w35784 & w35826;
assign w36307 = ~w35764 & w36306;
assign w36308 = w35797 & ~w35824;
assign w36309 = w35771 & w35784;
assign w36310 = ~w35834 & ~w36309;
assign w36311 = ~w35827 & ~w36310;
assign w36312 = w35814 & w36309;
assign w36313 = ~w35811 & ~w36312;
assign w36314 = ~w36305 & w36313;
assign w36315 = ~w36307 & w36314;
assign w36316 = ~w36311 & w36315;
assign w36317 = ~w36308 & w36316;
assign w36318 = ~w36304 & ~w36317;
assign w36319 = pi1893 & w36318;
assign w36320 = ~pi1893 & ~w36318;
assign w36321 = ~w36319 & ~w36320;
assign w36322 = w36031 & ~w36038;
assign w36323 = w36168 & ~w36322;
assign w36324 = ~w36093 & w36323;
assign w36325 = w36323 & w66139;
assign w36326 = ~w36053 & ~w36324;
assign w36327 = ~w36017 & ~w36325;
assign w36328 = ~w36326 & w36327;
assign w36329 = w36074 & ~w36169;
assign w36330 = w36053 & w36067;
assign w36331 = ~w36329 & ~w36330;
assign w36332 = (w36081 & ~w36323) | (w36081 & w66140) | (~w36323 & w66140);
assign w36333 = w36017 & ~w36166;
assign w36334 = ~w36089 & w36333;
assign w36335 = ~w36332 & w36334;
assign w36336 = ~w36331 & w36335;
assign w36337 = ~w36328 & ~w36336;
assign w36338 = pi1921 & w36337;
assign w36339 = ~pi1921 & ~w36337;
assign w36340 = ~w36338 & ~w36339;
assign w36341 = w35601 & w35617;
assign w36342 = ~w35623 & w35640;
assign w36343 = ~w35617 & w36342;
assign w36344 = ~w36341 & ~w36343;
assign w36345 = ~w35580 & ~w35621;
assign w36346 = w35586 & ~w35602;
assign w36347 = w36345 & ~w36346;
assign w36348 = ~w35596 & ~w36347;
assign w36349 = ~w36347 & w66141;
assign w36350 = ~w35634 & ~w36194;
assign w36351 = ~w35614 & ~w36350;
assign w36352 = w35597 & ~w36351;
assign w36353 = ~w35598 & ~w35621;
assign w36354 = w36352 & w36353;
assign w36355 = w36344 & ~w36349;
assign w36356 = ~w36354 & w36355;
assign w36357 = ~w35613 & ~w36356;
assign w36358 = w35579 & w35601;
assign w36359 = ~w35567 & w36358;
assign w36360 = w35596 & ~w35600;
assign w36361 = ~w36359 & w36360;
assign w36362 = ~w36201 & ~w36361;
assign w36363 = w35586 & w36344;
assign w36364 = w36348 & ~w36363;
assign w36365 = w35613 & ~w36352;
assign w36366 = (~w36362 & w36364) | (~w36362 & w66142) | (w36364 & w66142);
assign w36367 = ~w36357 & w36366;
assign w36368 = pi1911 & ~w36367;
assign w36369 = ~pi1911 & w36367;
assign w36370 = ~w36368 & ~w36369;
assign w36371 = w35719 & w35728;
assign w36372 = w35705 & w35730;
assign w36373 = w35707 & w66143;
assign w36374 = ~w35719 & ~w36373;
assign w36375 = w35703 & w35705;
assign w36376 = ~w35736 & ~w36375;
assign w36377 = ~w36374 & w36376;
assign w36378 = ~w36371 & ~w36377;
assign w36379 = w35672 & w35698;
assign w36380 = (w35701 & w35724) | (w35701 & w63910) | (w35724 & w63910);
assign w36381 = ~w35692 & w35723;
assign w36382 = w35723 & w66144;
assign w36383 = ~w35683 & ~w35724;
assign w36384 = ~w36382 & w36383;
assign w36385 = ~w36379 & ~w36380;
assign w36386 = ~w36384 & w36385;
assign w36387 = w35719 & ~w36386;
assign w36388 = ~w35673 & ~w35741;
assign w36389 = w35901 & w36388;
assign w36390 = ~w35746 & ~w36389;
assign w36391 = ~w36387 & w36390;
assign w36392 = w36391 & w66145;
assign w36393 = (~pi1913 & ~w36391) | (~pi1913 & w66146) | (~w36391 & w66146);
assign w36394 = ~w36392 & ~w36393;
assign w36395 = w36252 & w36264;
assign w36396 = w36243 & ~w36251;
assign w36397 = w36230 & ~w36236;
assign w36398 = ~w36396 & ~w36397;
assign w36399 = ~w36274 & ~w36398;
assign w36400 = ~w36275 & ~w36399;
assign w36401 = ~w36224 & ~w36264;
assign w36402 = ~w36400 & w36401;
assign w36403 = (~w36400 & w66147) | (~w36400 & w66148) | (w66147 & w66148);
assign w36404 = ~w36243 & w36251;
assign w36405 = (w36224 & w36399) | (w36224 & w63912) | (w36399 & w63912);
assign w36406 = ~w36243 & ~w36266;
assign w36407 = ~w36224 & w36398;
assign w36408 = ~w36406 & w36407;
assign w36409 = ~w36405 & ~w36408;
assign w36410 = w36264 & ~w36409;
assign w36411 = ~w36252 & ~w36281;
assign w36412 = w36224 & w36406;
assign w36413 = w36411 & w36412;
assign w36414 = w36272 & ~w36274;
assign w36415 = ~w36405 & w36414;
assign w36416 = ~w36272 & w36274;
assign w36417 = ~w36288 & w36416;
assign w36418 = ~w36256 & ~w36283;
assign w36419 = w36243 & ~w36418;
assign w36420 = ~w36417 & ~w36419;
assign w36421 = (~w36264 & ~w36420) | (~w36264 & w66149) | (~w36420 & w66149);
assign w36422 = ~w36403 & ~w36413;
assign w36423 = ~w36410 & w36422;
assign w36424 = ~w36421 & w36423;
assign w36425 = pi1916 & ~w36424;
assign w36426 = ~pi1916 & w36424;
assign w36427 = ~w36425 & ~w36426;
assign w36428 = w35707 & w35719;
assign w36429 = w35681 & w35900;
assign w36430 = ~w35695 & ~w36429;
assign w36431 = ~w36382 & w36430;
assign w36432 = ~w36428 & ~w36431;
assign w36433 = ~w35719 & w35737;
assign w36434 = ~w36379 & w36433;
assign w36435 = w35745 & w36381;
assign w36436 = w35910 & ~w36435;
assign w36437 = ~w35727 & w36436;
assign w36438 = ~w36434 & ~w36437;
assign w36439 = ~w36432 & ~w36438;
assign w36440 = ~pi1917 & w36439;
assign w36441 = pi1917 & ~w36439;
assign w36442 = ~w36440 & ~w36441;
assign w36443 = ~w36274 & w36283;
assign w36444 = ~w36224 & w36416;
assign w36445 = w36236 & ~w36244;
assign w36446 = w36400 & ~w36445;
assign w36447 = ~w36230 & w36243;
assign w36448 = w36224 & ~w36447;
assign w36449 = (w36448 & ~w36400) | (w36448 & w66150) | (~w36400 & w66150);
assign w36450 = ~w36415 & ~w36444;
assign w36451 = (w36264 & ~w36450) | (w36264 & w66151) | (~w36450 & w66151);
assign w36452 = ~w36245 & ~w36264;
assign w36453 = ~w36444 & w36452;
assign w36454 = w36446 & w36453;
assign w36455 = w36288 & w36407;
assign w36456 = ~w36443 & ~w36455;
assign w36457 = ~w36402 & w36456;
assign w36458 = ~w36454 & w36457;
assign w36459 = ~w36451 & w36458;
assign w36460 = pi1908 & ~w36459;
assign w36461 = ~pi1908 & w36459;
assign w36462 = ~w36460 & ~w36461;
assign w36463 = w35957 & ~w36140;
assign w36464 = w35964 & ~w35965;
assign w36465 = ~w36145 & w36464;
assign w36466 = ~w36463 & ~w36465;
assign w36467 = w35975 & ~w36466;
assign w36468 = ~w35979 & ~w36124;
assign w36469 = w35930 & ~w36468;
assign w36470 = ~w35989 & ~w36146;
assign w36471 = ~w35968 & ~w35975;
assign w36472 = ~w36470 & ~w36471;
assign w36473 = w35947 & ~w35958;
assign w36474 = w35937 & ~w36145;
assign w36475 = w36118 & w36474;
assign w36476 = ~w35987 & ~w36475;
assign w36477 = ~w36473 & w36476;
assign w36478 = ~w35975 & ~w36477;
assign w36479 = ~w36469 & ~w36472;
assign w36480 = ~w36467 & w36479;
assign w36481 = ~w36478 & w36480;
assign w36482 = ~pi1912 & ~w36481;
assign w36483 = pi1912 & w36481;
assign w36484 = ~w36482 & ~w36483;
assign w36485 = ~w35822 & w35795;
assign w36486 = ~w36312 & ~w36485;
assign w36487 = w35784 & ~w35792;
assign w36488 = ~w36306 & ~w36487;
assign w36489 = (~w35758 & w36488) | (~w35758 & w66152) | (w36488 & w66152);
assign w36490 = ~w35771 & w35822;
assign w36491 = w35822 & w66153;
assign w36492 = w35758 & w36491;
assign w36493 = w36486 & ~w36492;
assign w36494 = ~w36489 & w36493;
assign w36495 = w35811 & ~w36494;
assign w36496 = ~w35811 & ~w36490;
assign w36497 = w36486 & w36496;
assign w36498 = w35813 & ~w36497;
assign w36499 = ~w35802 & ~w36491;
assign w36500 = ~w35811 & ~w36499;
assign w36501 = ~w35758 & w36486;
assign w36502 = ~w36500 & w36501;
assign w36503 = ~w36498 & ~w36502;
assign w36504 = ~w36495 & ~w36503;
assign w36505 = ~pi1904 & w36504;
assign w36506 = pi1904 & ~w36504;
assign w36507 = ~w36505 & ~w36506;
assign w36508 = w36243 & w36252;
assign w36509 = ~w36289 & ~w36508;
assign w36510 = ~w36251 & w36254;
assign w36511 = w36286 & ~w36510;
assign w36512 = ~w36236 & ~w36411;
assign w36513 = w36224 & ~w36280;
assign w36514 = ~w36512 & w36513;
assign w36515 = (w36509 & w36514) | (w36509 & w66154) | (w36514 & w66154);
assign w36516 = w36264 & ~w36515;
assign w36517 = (w36286 & w36408) | (w36286 & w66155) | (w36408 & w66155);
assign w36518 = ~w36243 & ~w36400;
assign w36519 = ~w36517 & ~w36518;
assign w36520 = ~w36264 & ~w36519;
assign w36521 = ~w36237 & ~w36396;
assign w36522 = w36224 & ~w36521;
assign w36523 = ~w36508 & ~w36522;
assign w36524 = ~w36264 & w36509;
assign w36525 = w36224 & ~w36404;
assign w36526 = ~w36524 & w36525;
assign w36527 = ~w36523 & ~w36526;
assign w36528 = ~w36516 & ~w36527;
assign w36529 = ~w36520 & w36528;
assign w36530 = pi1909 & ~w36529;
assign w36531 = ~pi1909 & w36529;
assign w36532 = ~w36530 & ~w36531;
assign w36533 = w35459 & ~w35472;
assign w36534 = (w35446 & ~w35459) | (w35446 & w63913) | (~w35459 & w63913);
assign w36535 = ~w35501 & w36534;
assign w36536 = w35459 & w35478;
assign w36537 = (~w35446 & ~w35489) | (~w35446 & w36541) | (~w35489 & w36541);
assign w36538 = ~w36536 & w36537;
assign w36539 = ~w36535 & ~w36538;
assign w36540 = ~w35465 & w36533;
assign w36541 = ~w35446 & w35458;
assign w36542 = w35488 & w35515;
assign w36543 = ~w35473 & ~w36542;
assign w36544 = ~w35481 & w36543;
assign w36545 = ~w35452 & w35465;
assign w36546 = w35472 & ~w36541;
assign w36547 = ~w36545 & w36546;
assign w36548 = w36544 & w36547;
assign w36549 = ~w36539 & ~w36540;
assign w36550 = ~w36548 & w36549;
assign w36551 = w35508 & ~w36550;
assign w36552 = ~w35514 & w66156;
assign w36553 = w35446 & ~w35452;
assign w36554 = w35477 & w36553;
assign w36555 = ~w35479 & w35483;
assign w36556 = ~w36544 & ~w36553;
assign w36557 = ~w35475 & ~w35494;
assign w36558 = w35446 & w35465;
assign w36559 = ~w36557 & w36558;
assign w36560 = ~w36555 & ~w36559;
assign w36561 = ~w36556 & w36560;
assign w36562 = ~w35508 & ~w36561;
assign w36563 = ~w36552 & ~w36554;
assign w36564 = ~w36551 & w36563;
assign w36565 = (pi1902 & ~w36564) | (pi1902 & w66157) | (~w36564 & w66157);
assign w36566 = w36564 & w66158;
assign w36567 = ~w36565 & ~w36566;
assign w36568 = w35483 & w35498;
assign w36569 = ~w35496 & ~w35501;
assign w36570 = w35508 & ~w36569;
assign w36571 = ~w35482 & ~w36570;
assign w36572 = ~w35446 & ~w36571;
assign w36573 = ~w35465 & ~w35476;
assign w36574 = w35452 & ~w36573;
assign w36575 = w35497 & w36574;
assign w36576 = ~w35513 & w36555;
assign w36577 = w35509 & ~w36533;
assign w36578 = ~w36575 & ~w36576;
assign w36579 = w36577 & w36578;
assign w36580 = w35458 & w35472;
assign w36581 = w36534 & ~w36580;
assign w36582 = ~w35494 & w36581;
assign w36583 = ~w36541 & ~w36581;
assign w36584 = w35478 & ~w36583;
assign w36585 = ~w35508 & w36543;
assign w36586 = ~w36582 & w36585;
assign w36587 = ~w36584 & w36586;
assign w36588 = ~w36579 & ~w36587;
assign w36589 = ~w35491 & ~w36568;
assign w36590 = ~w36572 & w36589;
assign w36591 = ~w36588 & w36590;
assign w36592 = pi1915 & ~w36591;
assign w36593 = ~pi1915 & w36591;
assign w36594 = ~w36592 & ~w36593;
assign w36595 = w35795 & w35820;
assign w36596 = ~w35800 & ~w35814;
assign w36597 = ~w35793 & w36596;
assign w36598 = w35813 & ~w35819;
assign w36599 = ~w36597 & w36598;
assign w36600 = ~w35798 & ~w36599;
assign w36601 = w35811 & ~w36595;
assign w36602 = ~w36600 & w36601;
assign w36603 = ~w35789 & ~w35827;
assign w36604 = ~w36597 & ~w36603;
assign w36605 = ~w35785 & w36305;
assign w36606 = ~w35811 & ~w35816;
assign w36607 = ~w36604 & w36606;
assign w36608 = ~w36605 & w36607;
assign w36609 = ~w36602 & ~w36608;
assign w36610 = ~pi1903 & w36609;
assign w36611 = pi1903 & ~w36609;
assign w36612 = ~w36610 & ~w36611;
assign w36613 = w35599 & ~w35601;
assign w36614 = (w35596 & ~w35589) | (w35596 & w66159) | (~w35589 & w66159);
assign w36615 = ~w36358 & w36614;
assign w36616 = ~w35596 & ~w35598;
assign w36617 = ~w36194 & w36616;
assign w36618 = ~w35641 & w36617;
assign w36619 = ~w36615 & ~w36618;
assign w36620 = w35613 & ~w36613;
assign w36621 = ~w36619 & w36620;
assign w36622 = ~w35621 & ~w36194;
assign w36623 = w36615 & w36622;
assign w36624 = ~w35623 & ~w36345;
assign w36625 = w35638 & w36624;
assign w36626 = ~w35588 & ~w35613;
assign w36627 = ~w36623 & w36626;
assign w36628 = ~w36625 & w36627;
assign w36629 = ~w36621 & ~w36628;
assign w36630 = ~w36208 & ~w36350;
assign w36631 = ~w35596 & ~w36359;
assign w36632 = ~w36630 & w36631;
assign w36633 = w35596 & ~w35635;
assign w36634 = ~w36195 & w36633;
assign w36635 = ~w36632 & ~w36634;
assign w36636 = ~w36629 & ~w36635;
assign w36637 = ~pi1930 & w36636;
assign w36638 = pi1930 & ~w36636;
assign w36639 = ~w36637 & ~w36638;
assign w36640 = w36039 & w36054;
assign w36641 = ~w36081 & ~w36083;
assign w36642 = w36090 & w36641;
assign w36643 = ~w36179 & ~w36640;
assign w36644 = w36643 & w66160;
assign w36645 = ~w36017 & ~w36644;
assign w36646 = ~w36053 & w36087;
assign w36647 = ~w36040 & w36181;
assign w36648 = w36040 & ~w36053;
assign w36649 = w36017 & ~w36069;
assign w36650 = ~w36648 & w36649;
assign w36651 = ~w36647 & w36650;
assign w36652 = ~w36071 & ~w36646;
assign w36653 = ~w36645 & w36652;
assign w36654 = ~w36651 & w36653;
assign w36655 = pi1931 & ~w36654;
assign w36656 = ~pi1931 & w36654;
assign w36657 = ~w36655 & ~w36656;
assign w36658 = ~w35466 & ~w36574;
assign w36659 = w35492 & w36658;
assign w36660 = ~w35508 & ~w36658;
assign w36661 = ~w35502 & ~w36540;
assign w36662 = ~w36660 & w36661;
assign w36663 = w35446 & ~w36662;
assign w36664 = w35452 & ~w36580;
assign w36665 = w35479 & w36664;
assign w36666 = w35475 & w36541;
assign w36667 = w35515 & w36553;
assign w36668 = ~w36536 & ~w36666;
assign w36669 = ~w36667 & w36668;
assign w36670 = ~w36665 & w36669;
assign w36671 = w35508 & ~w36670;
assign w36672 = w35472 & w36542;
assign w36673 = ~w35508 & w36545;
assign w36674 = ~w35498 & w36673;
assign w36675 = ~w36672 & ~w36674;
assign w36676 = ~w36659 & w36675;
assign w36677 = ~w36671 & w36676;
assign w36678 = ~w36663 & w36677;
assign w36679 = pi1914 & ~w36678;
assign w36680 = ~pi1914 & w36678;
assign w36681 = ~w36679 & ~w36680;
assign w36682 = ~pi6527 & pi9040;
assign w36683 = ~pi6695 & ~pi9040;
assign w36684 = ~w36682 & ~w36683;
assign w36685 = pi1920 & ~w36684;
assign w36686 = ~pi1920 & w36684;
assign w36687 = ~w36685 & ~w36686;
assign w36688 = ~pi6526 & pi9040;
assign w36689 = ~pi6609 & ~pi9040;
assign w36690 = ~w36688 & ~w36689;
assign w36691 = pi1925 & ~w36690;
assign w36692 = ~pi1925 & w36690;
assign w36693 = ~w36691 & ~w36692;
assign w36694 = ~pi6600 & pi9040;
assign w36695 = ~pi6528 & ~pi9040;
assign w36696 = ~w36694 & ~w36695;
assign w36697 = pi1943 & ~w36696;
assign w36698 = ~pi1943 & w36696;
assign w36699 = ~w36697 & ~w36698;
assign w36700 = ~pi6629 & pi9040;
assign w36701 = ~pi6530 & ~pi9040;
assign w36702 = ~w36700 & ~w36701;
assign w36703 = pi1940 & ~w36702;
assign w36704 = ~pi1940 & w36702;
assign w36705 = ~w36703 & ~w36704;
assign w36706 = ~w36687 & w36705;
assign w36707 = ~pi6525 & pi9040;
assign w36708 = ~pi6540 & ~pi9040;
assign w36709 = ~w36707 & ~w36708;
assign w36710 = pi1928 & ~w36709;
assign w36711 = ~pi1928 & w36709;
assign w36712 = ~w36710 & ~w36711;
assign w36713 = w36706 & w36712;
assign w36714 = w36706 & w36721;
assign w36715 = ~w36699 & ~w36705;
assign w36716 = w36712 & w36715;
assign w36717 = ~w36714 & ~w36716;
assign w36718 = ~w36693 & ~w36717;
assign w36719 = ~w36717 & w66161;
assign w36720 = ~w36687 & ~w36705;
assign w36721 = w36699 & w36712;
assign w36722 = w36720 & w36721;
assign w36723 = ~w36699 & ~w36712;
assign w36724 = w36687 & w36705;
assign w36725 = ~w36720 & ~w36724;
assign w36726 = w36723 & ~w36725;
assign w36727 = w36699 & ~w36712;
assign w36728 = w36706 & w36727;
assign w36729 = ~w36722 & ~w36728;
assign w36730 = ~w36726 & w36729;
assign w36731 = w36693 & ~w36730;
assign w36732 = ~w36693 & w36713;
assign w36733 = w36687 & ~w36699;
assign w36734 = ~w36705 & w36712;
assign w36735 = ~w36733 & w36734;
assign w36736 = ~w36721 & w36724;
assign w36737 = ~w36735 & ~w36736;
assign w36738 = ~w36687 & w36693;
assign w36739 = w36693 & ~w36723;
assign w36740 = ~w36738 & ~w36739;
assign w36741 = w36737 & ~w36740;
assign w36742 = w36724 & w36727;
assign w36743 = ~w36693 & ~w36742;
assign w36744 = ~w36712 & w36720;
assign w36745 = w36743 & ~w36744;
assign w36746 = ~w36741 & ~w36745;
assign w36747 = ~pi6693 & pi9040;
assign w36748 = ~pi6525 & ~pi9040;
assign w36749 = ~w36747 & ~w36748;
assign w36750 = pi1938 & ~w36749;
assign w36751 = ~pi1938 & w36749;
assign w36752 = ~w36750 & ~w36751;
assign w36753 = ~w36732 & w36752;
assign w36754 = ~w36746 & w36753;
assign w36755 = w36687 & w36699;
assign w36756 = w36705 & w36723;
assign w36757 = ~w36756 & w66162;
assign w36758 = ~w36693 & ~w36757;
assign w36759 = ~w36699 & w36705;
assign w36760 = w36738 & w36759;
assign w36761 = (~w36760 & ~w36737) | (~w36760 & w66163) | (~w36737 & w66163);
assign w36762 = w36712 & ~w36761;
assign w36763 = w36727 & w36738;
assign w36764 = ~w36752 & ~w36763;
assign w36765 = ~w36758 & w36764;
assign w36766 = ~w36762 & w36765;
assign w36767 = ~w36754 & ~w36766;
assign w36768 = ~w36719 & ~w36731;
assign w36769 = ~w36767 & w36768;
assign w36770 = pi1954 & w36769;
assign w36771 = ~pi1954 & ~w36769;
assign w36772 = ~w36770 & ~w36771;
assign w36773 = ~pi6528 & pi9040;
assign w36774 = ~pi6532 & ~pi9040;
assign w36775 = ~w36773 & ~w36774;
assign w36776 = pi1923 & ~w36775;
assign w36777 = ~pi1923 & w36775;
assign w36778 = ~w36776 & ~w36777;
assign w36779 = ~pi6609 & pi9040;
assign w36780 = ~pi6527 & ~pi9040;
assign w36781 = ~w36779 & ~w36780;
assign w36782 = pi1920 & ~w36781;
assign w36783 = ~pi1920 & w36781;
assign w36784 = ~w36782 & ~w36783;
assign w36785 = ~w36778 & ~w36784;
assign w36786 = ~pi6543 & pi9040;
assign w36787 = ~pi6492 & ~pi9040;
assign w36788 = ~w36786 & ~w36787;
assign w36789 = pi1939 & ~w36788;
assign w36790 = ~pi1939 & w36788;
assign w36791 = ~w36789 & ~w36790;
assign w36792 = ~pi6530 & pi9040;
assign w36793 = ~pi6625 & ~pi9040;
assign w36794 = ~w36792 & ~w36793;
assign w36795 = pi1924 & ~w36794;
assign w36796 = ~pi1924 & w36794;
assign w36797 = ~w36795 & ~w36796;
assign w36798 = ~w36791 & w36797;
assign w36799 = w36785 & w36798;
assign w36800 = ~pi6625 & pi9040;
assign w36801 = ~pi6626 & ~pi9040;
assign w36802 = ~w36800 & ~w36801;
assign w36803 = pi1933 & ~w36802;
assign w36804 = ~pi1933 & w36802;
assign w36805 = ~w36803 & ~w36804;
assign w36806 = ~w36799 & w36805;
assign w36807 = w36778 & w36784;
assign w36808 = w36798 & ~w36807;
assign w36809 = ~w36785 & ~w36808;
assign w36810 = w36806 & ~w36809;
assign w36811 = w36791 & ~w36797;
assign w36812 = ~w36798 & ~w36811;
assign w36813 = ~w36778 & w36805;
assign w36814 = w36784 & ~w36813;
assign w36815 = w36812 & w36814;
assign w36816 = w36778 & ~w36784;
assign w36817 = ~w36799 & ~w36816;
assign w36818 = ~w36778 & w36784;
assign w36819 = w36791 & w36797;
assign w36820 = w36818 & w36819;
assign w36821 = ~w36805 & ~w36820;
assign w36822 = ~w36791 & w36816;
assign w36823 = w36821 & ~w36822;
assign w36824 = ~w36817 & w36823;
assign w36825 = ~w36785 & ~w36813;
assign w36826 = w36811 & ~w36825;
assign w36827 = ~pi6523 & pi9040;
assign w36828 = ~pi6497 & ~pi9040;
assign w36829 = ~w36827 & ~w36828;
assign w36830 = pi1928 & ~w36829;
assign w36831 = ~pi1928 & w36829;
assign w36832 = ~w36830 & ~w36831;
assign w36833 = ~w36815 & ~w36832;
assign w36834 = ~w36826 & w36833;
assign w36835 = ~w36824 & w36834;
assign w36836 = ~w36778 & ~w36797;
assign w36837 = w36778 & w36797;
assign w36838 = ~w36836 & ~w36837;
assign w36839 = w36791 & w36805;
assign w36840 = ~w36816 & w36839;
assign w36841 = w36838 & w36840;
assign w36842 = w36784 & ~w36791;
assign w36843 = ~w36784 & w36791;
assign w36844 = ~w36842 & ~w36843;
assign w36845 = ~w36797 & w36844;
assign w36846 = w36844 & w63914;
assign w36847 = w36798 & w36818;
assign w36848 = w36778 & ~w36791;
assign w36849 = w36811 & w36818;
assign w36850 = ~w36848 & ~w36849;
assign w36851 = w36823 & ~w36850;
assign w36852 = w36832 & ~w36847;
assign w36853 = ~w36841 & w36852;
assign w36854 = ~w36846 & w36853;
assign w36855 = ~w36851 & w36854;
assign w36856 = ~w36835 & ~w36855;
assign w36857 = w36778 & ~w36805;
assign w36858 = w36812 & w36857;
assign w36859 = ~w36810 & ~w36858;
assign w36860 = ~w36856 & w36859;
assign w36861 = pi1959 & ~w36860;
assign w36862 = ~pi1959 & w36860;
assign w36863 = ~w36861 & ~w36862;
assign w36864 = ~pi6512 & pi9040;
assign w36865 = ~pi6622 & ~pi9040;
assign w36866 = ~w36864 & ~w36865;
assign w36867 = pi1927 & ~w36866;
assign w36868 = ~pi1927 & w36866;
assign w36869 = ~w36867 & ~w36868;
assign w36870 = ~pi6623 & pi9040;
assign w36871 = ~pi6517 & ~pi9040;
assign w36872 = ~w36870 & ~w36871;
assign w36873 = pi1938 & ~w36872;
assign w36874 = ~pi1938 & w36872;
assign w36875 = ~w36873 & ~w36874;
assign w36876 = ~pi6608 & pi9040;
assign w36877 = ~pi6520 & ~pi9040;
assign w36878 = ~w36876 & ~w36877;
assign w36879 = pi1950 & ~w36878;
assign w36880 = ~pi1950 & w36878;
assign w36881 = ~w36879 & ~w36880;
assign w36882 = w36875 & ~w36881;
assign w36883 = ~pi6546 & pi9040;
assign w36884 = ~pi6524 & ~pi9040;
assign w36885 = ~w36883 & ~w36884;
assign w36886 = pi1941 & ~w36885;
assign w36887 = ~pi1941 & w36885;
assign w36888 = ~w36886 & ~w36887;
assign w36889 = w36882 & w36888;
assign w36890 = ~pi6539 & pi9040;
assign w36891 = ~pi6513 & ~pi9040;
assign w36892 = ~w36890 & ~w36891;
assign w36893 = pi1900 & ~w36892;
assign w36894 = ~pi1900 & w36892;
assign w36895 = ~w36893 & ~w36894;
assign w36896 = ~w36888 & ~w36895;
assign w36897 = ~pi6489 & pi9040;
assign w36898 = ~pi6621 & ~pi9040;
assign w36899 = ~w36897 & ~w36898;
assign w36900 = pi1943 & ~w36899;
assign w36901 = ~pi1943 & w36899;
assign w36902 = ~w36900 & ~w36901;
assign w36903 = w36896 & ~w36902;
assign w36904 = w36888 & w36895;
assign w36905 = ~w36882 & ~w36904;
assign w36906 = w36902 & ~w36905;
assign w36907 = ~w36875 & ~w36881;
assign w36908 = w36875 & w36881;
assign w36909 = ~w36875 & ~w36895;
assign w36910 = w36902 & w36909;
assign w36911 = ~w36904 & ~w36910;
assign w36912 = ~w36907 & ~w36908;
assign w36913 = ~w36911 & w36912;
assign w36914 = ~w36903 & ~w36906;
assign w36915 = ~w36913 & w36914;
assign w36916 = w36889 & w36915;
assign w36917 = w36895 & ~w36902;
assign w36918 = ~w36910 & ~w36917;
assign w36919 = w36875 & w36902;
assign w36920 = ~w36881 & ~w36919;
assign w36921 = w36918 & w36920;
assign w36922 = w36875 & w36895;
assign w36923 = ~w36909 & ~w36922;
assign w36924 = w36888 & w36902;
assign w36925 = ~w36923 & ~w36924;
assign w36926 = ~w36888 & ~w36902;
assign w36927 = ~w36896 & ~w36926;
assign w36928 = w36925 & w36927;
assign w36929 = ~w36921 & ~w36928;
assign w36930 = (~w36888 & ~w36929) | (~w36888 & w63412) | (~w36929 & w63412);
assign w36931 = ~w36896 & ~w36904;
assign w36932 = ~w36875 & w36881;
assign w36933 = w36931 & w36932;
assign w36934 = w36896 & w63915;
assign w36935 = ~w36875 & ~w36902;
assign w36936 = ~w36896 & w36935;
assign w36937 = w36881 & ~w36917;
assign w36938 = ~w36920 & ~w36937;
assign w36939 = ~w36933 & ~w36936;
assign w36940 = ~w36934 & ~w36938;
assign w36941 = w36939 & w36940;
assign w36942 = ~w36908 & ~w36941;
assign w36943 = w36930 & ~w36942;
assign w36944 = ~w36919 & ~w36935;
assign w36945 = ~w36895 & ~w36944;
assign w36946 = w36895 & w36944;
assign w36947 = ~w36945 & ~w36946;
assign w36948 = ~w36947 & w63916;
assign w36949 = ~w36916 & ~w36948;
assign w36950 = ~w36943 & w36949;
assign w36951 = w36869 & ~w36941;
assign w36952 = ~w36881 & w36904;
assign w36953 = ~w36944 & w36952;
assign w36954 = w36908 & w36926;
assign w36955 = ~w36881 & w36902;
assign w36956 = w36896 & w36955;
assign w36957 = ~w36954 & ~w36956;
assign w36958 = ~w36953 & w36957;
assign w36959 = ~w36951 & w36958;
assign w36960 = (w36950 & w66164) | (w36950 & w66165) | (w66164 & w66165);
assign w36961 = (~w36950 & w66166) | (~w36950 & w66167) | (w66166 & w66167);
assign w36962 = ~w36960 & ~w36961;
assign w36963 = ~pi6486 & pi9040;
assign w36964 = ~pi6518 & ~pi9040;
assign w36965 = ~w36963 & ~w36964;
assign w36966 = pi1926 & ~w36965;
assign w36967 = ~pi1926 & w36965;
assign w36968 = ~w36966 & ~w36967;
assign w36969 = ~pi6493 & pi9040;
assign w36970 = ~pi6515 & ~pi9040;
assign w36971 = ~w36969 & ~w36970;
assign w36972 = pi1923 & ~w36971;
assign w36973 = ~pi1923 & w36971;
assign w36974 = ~w36972 & ~w36973;
assign w36975 = w36968 & w36974;
assign w36976 = ~pi6497 & pi9040;
assign w36977 = ~pi6488 & ~pi9040;
assign w36978 = ~w36976 & ~w36977;
assign w36979 = pi1906 & ~w36978;
assign w36980 = ~pi1906 & w36978;
assign w36981 = ~w36979 & ~w36980;
assign w36982 = w36975 & w36981;
assign w36983 = ~pi6488 & pi9040;
assign w36984 = ~pi6693 & ~pi9040;
assign w36985 = ~w36983 & ~w36984;
assign w36986 = pi1932 & ~w36985;
assign w36987 = ~pi1932 & w36985;
assign w36988 = ~w36986 & ~w36987;
assign w36989 = ~w36981 & w36988;
assign w36990 = ~w36968 & ~w36974;
assign w36991 = ~w36989 & w36990;
assign w36992 = ~w36982 & ~w36991;
assign w36993 = ~pi6626 & pi9040;
assign w36994 = ~pi6523 & ~pi9040;
assign w36995 = ~w36993 & ~w36994;
assign w36996 = pi1944 & ~w36995;
assign w36997 = ~pi1944 & w36995;
assign w36998 = ~w36996 & ~w36997;
assign w36999 = ~w36981 & ~w36998;
assign w37000 = ~w36992 & w36999;
assign w37001 = ~pi6492 & pi9040;
assign w37002 = ~pi6629 & ~pi9040;
assign w37003 = ~w37001 & ~w37002;
assign w37004 = pi1939 & ~w37003;
assign w37005 = ~pi1939 & w37003;
assign w37006 = ~w37004 & ~w37005;
assign w37007 = w36968 & ~w36988;
assign w37008 = ~w36974 & w37007;
assign w37009 = w37007 & w63918;
assign w37010 = w36968 & ~w36989;
assign w37011 = w36988 & w36990;
assign w37012 = ~w37010 & ~w37011;
assign w37013 = ~w37009 & ~w37012;
assign w37014 = ~w36974 & w36989;
assign w37015 = ~w36968 & ~w36988;
assign w37016 = w36974 & w37015;
assign w37017 = w37015 & w63919;
assign w37018 = ~w36998 & w37007;
assign w37019 = ~w37014 & ~w37018;
assign w37020 = ~w37017 & w37019;
assign w37021 = ~w37013 & ~w37020;
assign w37022 = w36968 & ~w36981;
assign w37023 = w36981 & ~w37007;
assign w37024 = (w36998 & w37023) | (w36998 & w66168) | (w37023 & w66168);
assign w37025 = w36981 & w36988;
assign w37026 = ~w37022 & ~w37025;
assign w37027 = ~w37010 & ~w37026;
assign w37028 = ~w36998 & ~w37027;
assign w37029 = ~w37024 & ~w37028;
assign w37030 = w36982 & ~w36988;
assign w37031 = ~w37021 & ~w37030;
assign w37032 = (~w37006 & ~w37031) | (~w37006 & w63920) | (~w37031 & w63920);
assign w37033 = w37021 & w37029;
assign w37034 = ~w36968 & w37014;
assign w37035 = ~w36982 & ~w37034;
assign w37036 = w36998 & ~w37035;
assign w37037 = w36975 & w36988;
assign w37038 = ~w36968 & w36988;
assign w37039 = (w36998 & ~w37038) | (w36998 & w66169) | (~w37038 & w66169);
assign w37040 = ~w37009 & ~w37037;
assign w37041 = w37039 & w37040;
assign w37042 = w37006 & ~w37041;
assign w37043 = ~w37036 & ~w37042;
assign w37044 = w36968 & ~w36974;
assign w37045 = ~w37015 & ~w37044;
assign w37046 = w36981 & ~w37045;
assign w37047 = ~w36981 & ~w36990;
assign w37048 = w37045 & w37047;
assign w37049 = ~w37037 & w37048;
assign w37050 = ~w36998 & ~w37046;
assign w37051 = ~w37049 & w37050;
assign w37052 = ~w37043 & ~w37051;
assign w37053 = ~w37000 & ~w37033;
assign w37054 = ~w37032 & w37053;
assign w37055 = (pi1953 & ~w37054) | (pi1953 & w66170) | (~w37054 & w66170);
assign w37056 = w37054 & w66171;
assign w37057 = ~w37055 & ~w37056;
assign w37058 = ~pi6718 & pi9040;
assign w37059 = ~pi6522 & ~pi9040;
assign w37060 = ~w37058 & ~w37059;
assign w37061 = pi1945 & ~w37060;
assign w37062 = ~pi1945 & w37060;
assign w37063 = ~w37061 & ~w37062;
assign w37064 = ~pi6606 & pi9040;
assign w37065 = ~pi6608 & ~pi9040;
assign w37066 = ~w37064 & ~w37065;
assign w37067 = pi1949 & ~w37066;
assign w37068 = ~pi1949 & w37066;
assign w37069 = ~w37067 & ~w37068;
assign w37070 = w37063 & ~w37069;
assign w37071 = ~pi6509 & pi9040;
assign w37072 = ~pi6529 & ~pi9040;
assign w37073 = ~w37071 & ~w37072;
assign w37074 = pi1935 & ~w37073;
assign w37075 = ~pi1935 & w37073;
assign w37076 = ~w37074 & ~w37075;
assign w37077 = ~pi6729 & pi9040;
assign w37078 = ~pi6539 & ~pi9040;
assign w37079 = ~w37077 & ~w37078;
assign w37080 = pi1922 & ~w37079;
assign w37081 = ~pi1922 & w37079;
assign w37082 = ~w37080 & ~w37081;
assign w37083 = ~w37076 & ~w37082;
assign w37084 = ~pi6490 & pi9040;
assign w37085 = ~pi6729 & ~pi9040;
assign w37086 = ~w37084 & ~w37085;
assign w37087 = pi1942 & ~w37086;
assign w37088 = ~pi1942 & w37086;
assign w37089 = ~w37087 & ~w37088;
assign w37090 = w37083 & ~w37089;
assign w37091 = ~w37069 & w37082;
assign w37092 = ~w37076 & w37089;
assign w37093 = w37091 & w37092;
assign w37094 = ~w37090 & ~w37093;
assign w37095 = ~pi6520 & pi9040;
assign w37096 = ~pi6509 & ~pi9040;
assign w37097 = ~w37095 & ~w37096;
assign w37098 = pi1948 & ~w37097;
assign w37099 = ~pi1948 & w37097;
assign w37100 = ~w37098 & ~w37099;
assign w37101 = w37083 & ~w37100;
assign w37102 = w37094 & ~w37101;
assign w37103 = w37070 & ~w37102;
assign w37104 = w37076 & ~w37089;
assign w37105 = ~w37070 & ~w37104;
assign w37106 = w37069 & ~w37082;
assign w37107 = ~w37091 & ~w37106;
assign w37108 = w37089 & w37107;
assign w37109 = w37063 & w37094;
assign w37110 = w37105 & ~w37108;
assign w37111 = w37109 & w37110;
assign w37112 = w37076 & w37082;
assign w37113 = w37063 & w37069;
assign w37114 = ~w37089 & w37091;
assign w37115 = ~w37113 & ~w37114;
assign w37116 = (w37112 & w37114) | (w37112 & w63921) | (w37114 & w63921);
assign w37117 = ~w37089 & ~w37107;
assign w37118 = w37083 & w37108;
assign w37119 = ~w37117 & ~w37118;
assign w37120 = w37083 & w37119;
assign w37121 = w37104 & w37106;
assign w37122 = ~w37076 & w37082;
assign w37123 = ~w37089 & w37122;
assign w37124 = w37069 & w37076;
assign w37125 = ~w37083 & ~w37124;
assign w37126 = ~w37123 & w37125;
assign w37127 = ~w37121 & ~w37126;
assign w37128 = ~w37063 & ~w37127;
assign w37129 = ~w37100 & ~w37116;
assign w37130 = ~w37111 & w37129;
assign w37131 = ~w37128 & w37130;
assign w37132 = ~w37120 & w37131;
assign w37133 = ~w37063 & ~w37119;
assign w37134 = w37089 & w37112;
assign w37135 = w37069 & ~w37134;
assign w37136 = w37069 & w37082;
assign w37137 = w37076 & ~w37082;
assign w37138 = w37063 & w37137;
assign w37139 = ~w37136 & ~w37138;
assign w37140 = ~w37135 & ~w37139;
assign w37141 = w37113 & w37122;
assign w37142 = w37100 & ~w37121;
assign w37143 = ~w37141 & w37142;
assign w37144 = ~w37140 & w37143;
assign w37145 = (w37132 & w66172) | (w37132 & w66173) | (w66172 & w66173);
assign w37146 = (~w37132 & w66174) | (~w37132 & w66175) | (w66174 & w66175);
assign w37147 = ~w37145 & ~w37146;
assign w37148 = w36920 & w36925;
assign w37149 = w36908 & w36947;
assign w37150 = w36888 & w36923;
assign w37151 = ~w36944 & w37150;
assign w37152 = ~w37148 & ~w37151;
assign w37153 = ~w37149 & w37152;
assign w37154 = ~w36869 & ~w37153;
assign w37155 = w36869 & ~w36909;
assign w37156 = ~w36931 & w37155;
assign w37157 = ~w36933 & ~w37156;
assign w37158 = w36902 & ~w37157;
assign w37159 = w36907 & w36926;
assign w37160 = w36875 & ~w36926;
assign w37161 = ~w36922 & w36926;
assign w37162 = w36881 & ~w37160;
assign w37163 = ~w37161 & w37162;
assign w37164 = ~w36889 & ~w37159;
assign w37165 = ~w37163 & w37164;
assign w37166 = w36869 & ~w37165;
assign w37167 = ~w37158 & ~w37166;
assign w37168 = ~w37154 & w37167;
assign w37169 = pi1965 & w37168;
assign w37170 = ~pi1965 & ~w37168;
assign w37171 = ~w37169 & ~w37170;
assign w37172 = ~pi6524 & pi9040;
assign w37173 = ~pi6489 & ~pi9040;
assign w37174 = ~w37172 & ~w37173;
assign w37175 = pi1900 & ~w37174;
assign w37176 = ~pi1900 & w37174;
assign w37177 = ~w37175 & ~w37176;
assign w37178 = ~pi6517 & pi9040;
assign w37179 = ~pi6718 & ~pi9040;
assign w37180 = ~w37178 & ~w37179;
assign w37181 = pi1927 & ~w37180;
assign w37182 = ~pi1927 & w37180;
assign w37183 = ~w37181 & ~w37182;
assign w37184 = w37177 & ~w37183;
assign w37185 = ~pi6534 & pi9040;
assign w37186 = ~pi6490 & ~pi9040;
assign w37187 = ~w37185 & ~w37186;
assign w37188 = pi1947 & ~w37187;
assign w37189 = ~pi1947 & w37187;
assign w37190 = ~w37188 & ~w37189;
assign w37191 = ~w37183 & w37190;
assign w37192 = ~w37177 & ~w37191;
assign w37193 = ~pi6511 & pi9040;
assign w37194 = ~pi6620 & ~pi9040;
assign w37195 = ~w37193 & ~w37194;
assign w37196 = pi1946 & ~w37195;
assign w37197 = ~pi1946 & w37195;
assign w37198 = ~w37196 & ~w37197;
assign w37199 = ~w37177 & ~w37190;
assign w37200 = w37183 & w37199;
assign w37201 = w37199 & w37232;
assign w37202 = w37192 & ~w37201;
assign w37203 = ~pi6496 & pi9040;
assign w37204 = ~pi6534 & ~pi9040;
assign w37205 = ~w37203 & ~w37204;
assign w37206 = pi1937 & ~w37205;
assign w37207 = ~pi1937 & w37205;
assign w37208 = ~w37206 & ~w37207;
assign w37209 = ~w37202 & ~w37208;
assign w37210 = ~w37183 & w37198;
assign w37211 = (~w37210 & w37202) | (~w37210 & w66176) | (w37202 & w66176);
assign w37212 = ~w37184 & ~w37211;
assign w37213 = w37177 & w37198;
assign w37214 = w37183 & ~w37190;
assign w37215 = w37213 & w37214;
assign w37216 = ~w37212 & ~w37215;
assign w37217 = ~pi6621 & pi9040;
assign w37218 = ~pi6516 & ~pi9040;
assign w37219 = ~w37217 & ~w37218;
assign w37220 = pi1934 & ~w37219;
assign w37221 = ~pi1934 & w37219;
assign w37222 = ~w37220 & ~w37221;
assign w37223 = ~w37216 & ~w37222;
assign w37224 = w37183 & w37190;
assign w37225 = w37177 & w37222;
assign w37226 = w37224 & w37225;
assign w37227 = w37184 & ~w37190;
assign w37228 = w37184 & w63923;
assign w37229 = w37222 & ~w37228;
assign w37230 = ~w37200 & ~w37227;
assign w37231 = w37229 & ~w37230;
assign w37232 = w37183 & ~w37198;
assign w37233 = ~w37177 & w37224;
assign w37234 = (~w37222 & ~w37224) | (~w37222 & w63924) | (~w37224 & w63924);
assign w37235 = w37232 & ~w37234;
assign w37236 = ~w37183 & ~w37190;
assign w37237 = ~w37198 & w37236;
assign w37238 = w37177 & w37190;
assign w37239 = ~w37183 & w37238;
assign w37240 = ~w37237 & ~w37239;
assign w37241 = ~w37222 & ~w37240;
assign w37242 = ~w37177 & w37210;
assign w37243 = w37210 & w66177;
assign w37244 = w37208 & ~w37226;
assign w37245 = ~w37243 & w37244;
assign w37246 = ~w37235 & w37245;
assign w37247 = w37246 & w66178;
assign w37248 = w37198 & w37224;
assign w37249 = ~w37177 & w37248;
assign w37250 = ~w37208 & ~w37215;
assign w37251 = ~w37249 & w37250;
assign w37252 = w37222 & ~w37240;
assign w37253 = ~w37190 & w37242;
assign w37254 = w37251 & ~w37253;
assign w37255 = ~w37252 & w37254;
assign w37256 = ~w37247 & ~w37255;
assign w37257 = ~w37223 & ~w37256;
assign w37258 = ~pi1961 & w37257;
assign w37259 = pi1961 & ~w37257;
assign w37260 = ~w37258 & ~w37259;
assign w37261 = ~w37177 & ~w37222;
assign w37262 = w37190 & ~w37198;
assign w37263 = w37261 & w37262;
assign w37264 = w37191 & w37213;
assign w37265 = ~w37263 & ~w37264;
assign w37266 = ~w37183 & ~w37225;
assign w37267 = ~w37265 & w37266;
assign w37268 = w37236 & w37261;
assign w37269 = w37183 & ~w37233;
assign w37270 = ~w37191 & ~w37222;
assign w37271 = w37198 & w37270;
assign w37272 = ~w37269 & w37271;
assign w37273 = w37177 & w37232;
assign w37274 = w37232 & w37238;
assign w37275 = ~w37201 & ~w37225;
assign w37276 = ~w37210 & ~w37275;
assign w37277 = w37208 & ~w37268;
assign w37278 = ~w37274 & w37277;
assign w37279 = ~w37272 & w37278;
assign w37280 = ~w37276 & w37279;
assign w37281 = ~w37208 & w37265;
assign w37282 = ~w37249 & ~w37271;
assign w37283 = ~w37272 & ~w37282;
assign w37284 = w37198 & ~w37261;
assign w37285 = ~w37192 & ~w37238;
assign w37286 = ~w37284 & w37285;
assign w37287 = w37281 & ~w37286;
assign w37288 = ~w37283 & w37287;
assign w37289 = ~w37280 & ~w37288;
assign w37290 = ~w37191 & w37222;
assign w37291 = ~w37242 & ~w37273;
assign w37292 = w37290 & ~w37291;
assign w37293 = ~w37267 & ~w37292;
assign w37294 = ~w37289 & w37293;
assign w37295 = pi1969 & w37294;
assign w37296 = ~pi1969 & ~w37294;
assign w37297 = ~w37295 & ~w37296;
assign w37298 = (w36805 & ~w36807) | (w36805 & w63925) | (~w36807 & w63925);
assign w37299 = w36838 & w36842;
assign w37300 = ~w37298 & w37299;
assign w37301 = w36805 & w36846;
assign w37302 = w36785 & w36819;
assign w37303 = ~w36849 & ~w37302;
assign w37304 = ~w37300 & w37303;
assign w37305 = ~w37301 & w37304;
assign w37306 = w36844 & w66179;
assign w37307 = w36805 & ~w37306;
assign w37308 = ~w36778 & ~w36812;
assign w37309 = ~w36785 & w36844;
assign w37310 = ~w37308 & ~w37309;
assign w37311 = w36778 & w36798;
assign w37312 = ~w36805 & ~w37311;
assign w37313 = ~w37310 & w37312;
assign w37314 = ~w37307 & ~w37313;
assign w37315 = w37304 & w63926;
assign w37316 = ~w37314 & w37315;
assign w37317 = w36837 & ~w36844;
assign w37318 = ~w36820 & ~w37317;
assign w37319 = (w36848 & ~w37318) | (w36848 & w66180) | (~w37318 & w66180);
assign w37320 = ~w36816 & ~w36818;
assign w37321 = ~w36819 & ~w37320;
assign w37322 = ~w36805 & ~w37321;
assign w37323 = ~w36832 & ~w37322;
assign w37324 = ~w37319 & w37323;
assign w37325 = ~w37316 & w37324;
assign w37326 = ~w36808 & ~w36839;
assign w37327 = w36778 & ~w37326;
assign w37328 = w36832 & ~w37327;
assign w37329 = w37305 & w37328;
assign w37330 = ~w37325 & w66181;
assign w37331 = (~pi1955 & w37325) | (~pi1955 & w66182) | (w37325 & w66182);
assign w37332 = ~w37330 & ~w37331;
assign w37333 = ~pi6536 & pi9040;
assign w37334 = ~pi6486 & ~pi9040;
assign w37335 = ~w37333 & ~w37334;
assign w37336 = pi1948 & ~w37335;
assign w37337 = ~pi1948 & w37335;
assign w37338 = ~w37336 & ~w37337;
assign w37339 = ~pi6628 & pi9040;
assign w37340 = ~pi6536 & ~pi9040;
assign w37341 = ~w37339 & ~w37340;
assign w37342 = pi1935 & ~w37341;
assign w37343 = ~pi1935 & w37341;
assign w37344 = ~w37342 & ~w37343;
assign w37345 = w37338 & w37344;
assign w37346 = ~pi6695 & pi9040;
assign w37347 = ~pi6493 & ~pi9040;
assign w37348 = ~w37346 & ~w37347;
assign w37349 = pi1951 & ~w37348;
assign w37350 = ~pi1951 & w37348;
assign w37351 = ~w37349 & ~w37350;
assign w37352 = ~pi6521 & pi9040;
assign w37353 = ~pi6543 & ~pi9040;
assign w37354 = ~w37352 & ~w37353;
assign w37355 = pi1932 & ~w37354;
assign w37356 = ~pi1932 & w37354;
assign w37357 = ~w37355 & ~w37356;
assign w37358 = ~w37351 & w37357;
assign w37359 = w37345 & w37358;
assign w37360 = w37351 & ~w37357;
assign w37361 = w37345 & w37360;
assign w37362 = ~w37344 & ~w37357;
assign w37363 = ~w37338 & w37351;
assign w37364 = w37362 & w37363;
assign w37365 = ~w37361 & ~w37364;
assign w37366 = ~w37338 & ~w37351;
assign w37367 = w37344 & w37366;
assign w37368 = ~pi6515 & pi9040;
assign w37369 = ~pi6607 & ~pi9040;
assign w37370 = ~w37368 & ~w37369;
assign w37371 = pi1936 & ~w37370;
assign w37372 = ~pi1936 & w37370;
assign w37373 = ~w37371 & ~w37372;
assign w37374 = (w37373 & ~w37366) | (w37373 & w66183) | (~w37366 & w66183);
assign w37375 = ~w37365 & w37374;
assign w37376 = w37338 & ~w37373;
assign w37377 = w37351 & w37376;
assign w37378 = ~w37345 & ~w37357;
assign w37379 = w37357 & ~w37366;
assign w37380 = w37373 & ~w37378;
assign w37381 = ~w37379 & w37380;
assign w37382 = ~w37377 & ~w37381;
assign w37383 = ~w37344 & ~w37382;
assign w37384 = w37338 & w37357;
assign w37385 = ~w37338 & ~w37357;
assign w37386 = ~w37384 & ~w37385;
assign w37387 = w37373 & ~w37386;
assign w37388 = w37344 & w37363;
assign w37389 = ~w37387 & w37388;
assign w37390 = w37344 & w37373;
assign w37391 = ~w37351 & ~w37357;
assign w37392 = w37390 & w37391;
assign w37393 = ~w37344 & ~w37363;
assign w37394 = ~w37373 & ~w37384;
assign w37395 = w37393 & w37394;
assign w37396 = ~pi6518 & pi9040;
assign w37397 = ~pi6526 & ~pi9040;
assign w37398 = ~w37396 & ~w37397;
assign w37399 = pi1926 & ~w37398;
assign w37400 = ~pi1926 & w37398;
assign w37401 = ~w37399 & ~w37400;
assign w37402 = ~w37392 & ~w37401;
assign w37403 = ~w37395 & w37402;
assign w37404 = ~w37389 & w37403;
assign w37405 = ~w37344 & w37384;
assign w37406 = ~w37367 & ~w37405;
assign w37407 = ~w37373 & ~w37406;
assign w37408 = w37338 & ~w37351;
assign w37409 = w37362 & w37408;
assign w37410 = w37344 & w37384;
assign w37411 = ~w37409 & ~w37410;
assign w37412 = w37373 & ~w37411;
assign w37413 = w37344 & w37358;
assign w37414 = w37344 & ~w37360;
assign w37415 = ~w37338 & w37373;
assign w37416 = ~w37414 & w37415;
assign w37417 = ~w37361 & w37401;
assign w37418 = ~w37413 & w37417;
assign w37419 = ~w37416 & w37418;
assign w37420 = ~w37407 & ~w37412;
assign w37421 = w37419 & w37420;
assign w37422 = ~w37404 & ~w37421;
assign w37423 = ~w37359 & ~w37375;
assign w37424 = ~w37383 & w37423;
assign w37425 = ~w37422 & w37424;
assign w37426 = pi1967 & ~w37425;
assign w37427 = ~pi1967 & w37425;
assign w37428 = ~w37426 & ~w37427;
assign w37429 = w37063 & w37104;
assign w37430 = ~w37107 & w37429;
assign w37431 = w37092 & w37136;
assign w37432 = ~w37063 & w37134;
assign w37433 = w37069 & ~w37092;
assign w37434 = w37105 & ~w37433;
assign w37435 = ~w37063 & ~w37069;
assign w37436 = w37104 & ~w37435;
assign w37437 = ~w37082 & ~w37436;
assign w37438 = ~w37434 & w37437;
assign w37439 = ~w37431 & ~w37432;
assign w37440 = ~w37438 & w37439;
assign w37441 = w37100 & w37440;
assign w37442 = ~w37100 & ~w37121;
assign w37443 = w37082 & ~w37104;
assign w37444 = w37433 & ~w37443;
assign w37445 = ~w37115 & ~w37444;
assign w37446 = w37442 & ~w37445;
assign w37447 = ~w37441 & ~w37446;
assign w37448 = ~w37063 & w37444;
assign w37449 = ~w37137 & w37448;
assign w37450 = ~w37100 & ~w37104;
assign w37451 = ~w37112 & w37450;
assign w37452 = ~w37123 & ~w37451;
assign w37453 = w37435 & ~w37452;
assign w37454 = ~w37430 & ~w37449;
assign w37455 = ~w37453 & w37454;
assign w37456 = ~w37447 & w37455;
assign w37457 = pi1956 & ~w37456;
assign w37458 = ~pi1956 & w37456;
assign w37459 = ~w37457 & ~w37458;
assign w37460 = w36991 & ~w37046;
assign w37461 = ~w37008 & ~w37037;
assign w37462 = ~w37460 & w37461;
assign w37463 = w36998 & ~w37006;
assign w37464 = (w37463 & w37460) | (w37463 & w66184) | (w37460 & w66184);
assign w37465 = w36999 & w37044;
assign w37466 = (w36974 & w37023) | (w36974 & w63927) | (w37023 & w63927);
assign w37467 = w37015 & ~w37466;
assign w37468 = w37462 & w37467;
assign w37469 = w37025 & w37044;
assign w37470 = ~w37034 & ~w37469;
assign w37471 = w36974 & w37038;
assign w37472 = w37470 & ~w37471;
assign w37473 = ~w36992 & ~w36998;
assign w37474 = ~w37030 & ~w37465;
assign w37475 = ~w37473 & w37474;
assign w37476 = ~w37468 & w37475;
assign w37477 = (w37006 & ~w37476) | (w37006 & w63928) | (~w37476 & w63928);
assign w37478 = w36981 & ~w37006;
assign w37479 = w37016 & w37478;
assign w37480 = w36974 & ~w36999;
assign w37481 = w36989 & w37480;
assign w37482 = ~w37048 & w37470;
assign w37483 = ~w36998 & ~w37006;
assign w37484 = ~w37482 & w37483;
assign w37485 = ~w37009 & ~w37479;
assign w37486 = ~w37481 & w37485;
assign w37487 = ~w37464 & w37486;
assign w37488 = ~w37484 & w37487;
assign w37489 = (pi1957 & w37477) | (pi1957 & w66185) | (w37477 & w66185);
assign w37490 = ~w37477 & w66186;
assign w37491 = ~w37489 & ~w37490;
assign w37492 = ~w36947 & w66187;
assign w37493 = (w36881 & w36910) | (w36881 & w63929) | (w36910 & w63929);
assign w37494 = ~w36946 & w37493;
assign w37495 = ~w36903 & ~w37160;
assign w37496 = ~w36921 & w37495;
assign w37497 = ~w37494 & w37496;
assign w37498 = ~w36916 & ~w37497;
assign w37499 = (w36869 & ~w37498) | (w36869 & w63930) | (~w37498 & w63930);
assign w37500 = ~w36869 & ~w36915;
assign w37501 = w36888 & ~w36953;
assign w37502 = w36913 & ~w37501;
assign w37503 = w36957 & ~w37159;
assign w37504 = ~w36941 & ~w37503;
assign w37505 = ~w37500 & ~w37502;
assign w37506 = ~w37504 & w37505;
assign w37507 = ~w37499 & w37506;
assign w37508 = ~pi1970 & w37507;
assign w37509 = pi1970 & ~w37507;
assign w37510 = ~w37508 & ~w37509;
assign w37511 = w37344 & w37357;
assign w37512 = w37394 & w37511;
assign w37513 = (w37357 & w37407) | (w37357 & w63931) | (w37407 & w63931);
assign w37514 = ~w37338 & ~w37362;
assign w37515 = ~w37511 & w37514;
assign w37516 = w37514 & w66188;
assign w37517 = w37338 & ~w37357;
assign w37518 = ~w37358 & ~w37517;
assign w37519 = ~w37514 & w37518;
assign w37520 = w37374 & ~w37519;
assign w37521 = ~w37519 & w66189;
assign w37522 = w37516 & w37521;
assign w37523 = (~w37401 & ~w37366) | (~w37401 & w63932) | (~w37366 & w63932);
assign w37524 = w37365 & w37523;
assign w37525 = ~w37512 & w37524;
assign w37526 = ~w37412 & w37525;
assign w37527 = ~w37513 & w37526;
assign w37528 = ~w37351 & w37376;
assign w37529 = w37387 & w37393;
assign w37530 = w37401 & ~w37528;
assign w37531 = ~w37516 & w37530;
assign w37532 = ~w37529 & w37531;
assign w37533 = w37362 & w37377;
assign w37534 = w37390 & ~w37391;
assign w37535 = ~w37379 & w37534;
assign w37536 = ~w37533 & ~w37535;
assign w37537 = (w37527 & w66190) | (w37527 & w66191) | (w66190 & w66191);
assign w37538 = pi1966 & w37537;
assign w37539 = ~pi1966 & ~w37537;
assign w37540 = ~w37538 & ~w37539;
assign w37541 = ~w37492 & ~w37493;
assign w37542 = ~w36869 & ~w37541;
assign w37543 = w36869 & ~w36906;
assign w37544 = ~w36929 & ~w37543;
assign w37545 = (w36869 & w36947) | (w36869 & w66192) | (w36947 & w66192);
assign w37546 = ~w36930 & w37545;
assign w37547 = ~w37544 & ~w37546;
assign w37548 = (pi1963 & ~w37547) | (pi1963 & w66193) | (~w37547 & w66193);
assign w37549 = w37547 & w66194;
assign w37550 = ~w37548 & ~w37549;
assign w37551 = w37090 & w37435;
assign w37552 = w37107 & w63934;
assign w37553 = ~w37113 & ~w37429;
assign w37554 = w37139 & ~w37553;
assign w37555 = ~w37552 & ~w37554;
assign w37556 = w37122 & ~w37433;
assign w37557 = (~w37063 & w37556) | (~w37063 & w63935) | (w37556 & w63935);
assign w37558 = w37555 & ~w37557;
assign w37559 = w37440 & w37558;
assign w37560 = (~w37100 & w37559) | (~w37100 & w63936) | (w37559 & w63936);
assign w37561 = (w37100 & ~w37555) | (w37100 & w66195) | (~w37555 & w66195);
assign w37562 = ~w37063 & w37552;
assign w37563 = ~w37111 & w66196;
assign w37564 = ~w37561 & w37563;
assign w37565 = ~w37560 & w66197;
assign w37566 = (pi1964 & w37560) | (pi1964 & w66198) | (w37560 & w66198);
assign w37567 = ~w37565 & ~w37566;
assign w37568 = ~w37373 & ~w37515;
assign w37569 = w37377 & w37511;
assign w37570 = w37408 & w37411;
assign w37571 = ~w37344 & w37351;
assign w37572 = w37517 & w37571;
assign w37573 = ~w37569 & ~w37572;
assign w37574 = ~w37570 & w37573;
assign w37575 = (w37568 & ~w37574) | (w37568 & w66199) | (~w37574 & w66199);
assign w37576 = ~w37401 & ~w37520;
assign w37577 = ~w37373 & w37516;
assign w37578 = w37345 & w37391;
assign w37579 = ~w37364 & ~w37578;
assign w37580 = w37373 & ~w37579;
assign w37581 = ~w37576 & w66200;
assign w37582 = ~w37575 & ~w37581;
assign w37583 = w37366 & w37568;
assign w37584 = ~w37521 & w37574;
assign w37585 = (w37401 & ~w37584) | (w37401 & w66201) | (~w37584 & w66201);
assign w37586 = ~w37582 & ~w37585;
assign w37587 = ~pi1968 & w37586;
assign w37588 = pi1968 & ~w37586;
assign w37589 = ~w37587 & ~w37588;
assign w37590 = w37433 & w37443;
assign w37591 = ~w37069 & w37112;
assign w37592 = ~w37063 & ~w37123;
assign w37593 = ~w37591 & w37592;
assign w37594 = ~w37109 & ~w37593;
assign w37595 = w37442 & ~w37590;
assign w37596 = ~w37594 & w37595;
assign w37597 = w37070 & w37094;
assign w37598 = w37100 & ~w37448;
assign w37599 = ~w37597 & w37598;
assign w37600 = ~w37596 & ~w37599;
assign w37601 = w37063 & w37089;
assign w37602 = ~w37555 & w37601;
assign w37603 = ~w37063 & ~w37076;
assign w37604 = ~w37100 & ~w37603;
assign w37605 = ~w37112 & ~w37604;
assign w37606 = w37108 & w37605;
assign w37607 = ~w37602 & ~w37606;
assign w37608 = ~w37600 & w37607;
assign w37609 = pi1973 & ~w37608;
assign w37610 = ~pi1973 & w37608;
assign w37611 = ~w37609 & ~w37610;
assign w37612 = w36975 & w36999;
assign w37613 = ~w37009 & ~w37612;
assign w37614 = (~w36998 & w36990) | (~w36998 & w66202) | (w36990 & w66202);
assign w37615 = ~w37011 & ~w37016;
assign w37616 = w37614 & ~w37615;
assign w37617 = (~w37006 & w37616) | (~w37006 & w66203) | (w37616 & w66203);
assign w37618 = (w37024 & ~w37476) | (w37024 & w63937) | (~w37476 & w63937);
assign w37619 = ~w37026 & w37480;
assign w37620 = w36999 & w37613;
assign w37621 = ~w37034 & ~w37619;
assign w37622 = ~w37620 & w37621;
assign w37623 = w37006 & ~w37622;
assign w37624 = (w37614 & ~w37461) | (w37614 & w66204) | (~w37461 & w66204);
assign w37625 = ~w36990 & w37463;
assign w37626 = ~w37008 & w37625;
assign w37627 = ~w37466 & w37626;
assign w37628 = ~w37624 & ~w37627;
assign w37629 = ~w37617 & w37628;
assign w37630 = ~w37623 & w37629;
assign w37631 = (pi1958 & w37618) | (pi1958 & w66205) | (w37618 & w66205);
assign w37632 = ~w37618 & w66206;
assign w37633 = ~w37631 & ~w37632;
assign w37634 = ~w37215 & ~w37274;
assign w37635 = w37230 & ~w37242;
assign w37636 = w37209 & ~w37635;
assign w37637 = w37634 & ~w37636;
assign w37638 = (~w37222 & w37636) | (~w37222 & w66207) | (w37636 & w66207);
assign w37639 = w37198 & w37199;
assign w37640 = w37234 & ~w37639;
assign w37641 = ~w37177 & ~w37198;
assign w37642 = ~w37191 & ~w37641;
assign w37643 = (w37222 & w37642) | (w37222 & w63938) | (w37642 & w63938);
assign w37644 = ~w37640 & ~w37643;
assign w37645 = ~w37228 & w37265;
assign w37646 = w37634 & w37645;
assign w37647 = (w37208 & ~w37646) | (w37208 & w63939) | (~w37646 & w63939);
assign w37648 = ~w37183 & w37262;
assign w37649 = w37281 & w37648;
assign w37650 = ~w37208 & w37290;
assign w37651 = w37637 & w37650;
assign w37652 = ~w37647 & ~w37649;
assign w37653 = ~w37638 & w37652;
assign w37654 = (pi1986 & ~w37653) | (pi1986 & w66208) | (~w37653 & w66208);
assign w37655 = w37653 & w66209;
assign w37656 = ~w37654 & ~w37655;
assign w37657 = ~w37039 & ~w37471;
assign w37658 = w37027 & ~w37657;
assign w37659 = w37020 & ~w37658;
assign w37660 = (w37006 & w37468) | (w37006 & w66210) | (w37468 & w66210);
assign w37661 = ~w36968 & w37483;
assign w37662 = w37615 & w37661;
assign w37663 = ~w37012 & w37463;
assign w37664 = ~w36988 & w37612;
assign w37665 = w37037 & w37478;
assign w37666 = ~w37664 & ~w37665;
assign w37667 = ~w37662 & w37666;
assign w37668 = ~w37663 & w37667;
assign w37669 = ~w37033 & w37668;
assign w37670 = ~w37660 & w37669;
assign w37671 = ~pi1962 & w37670;
assign w37672 = pi1962 & ~w37670;
assign w37673 = ~w37671 & ~w37672;
assign w37674 = (w37318 & w37313) | (w37318 & w66211) | (w37313 & w66211);
assign w37675 = w36832 & ~w37674;
assign w37676 = w37318 & w66212;
assign w37677 = w36806 & ~w37676;
assign w37678 = ~w36799 & ~w37306;
assign w37679 = ~w36832 & ~w37678;
assign w37680 = w36821 & ~w37317;
assign w37681 = ~w37679 & w37680;
assign w37682 = ~w37677 & ~w37681;
assign w37683 = ~w37675 & ~w37682;
assign w37684 = ~pi1971 & w37683;
assign w37685 = pi1971 & ~w37683;
assign w37686 = ~w37684 & ~w37685;
assign w37687 = (w37401 & w37363) | (w37401 & w66213) | (w37363 & w66213);
assign w37688 = w37518 & ~w37687;
assign w37689 = w37384 & w63932;
assign w37690 = ~w37578 & ~w37689;
assign w37691 = ~w37688 & w37690;
assign w37692 = ~w37373 & ~w37691;
assign w37693 = w37387 & ~w37519;
assign w37694 = ~w37359 & ~w37572;
assign w37695 = ~w37512 & w37694;
assign w37696 = ~w37693 & w37695;
assign w37697 = w37401 & ~w37696;
assign w37698 = w37373 & w37409;
assign w37699 = ~w37517 & w37571;
assign w37700 = ~w37381 & ~w37699;
assign w37701 = ~w37401 & ~w37700;
assign w37702 = ~w37522 & ~w37698;
assign w37703 = ~w37692 & ~w37697;
assign w37704 = w37703 & w66214;
assign w37705 = pi1980 & ~w37704;
assign w37706 = ~pi1980 & w37704;
assign w37707 = ~w37705 & ~w37706;
assign w37708 = w36693 & w36744;
assign w37709 = ~w36752 & ~w37708;
assign w37710 = ~w36699 & ~w36738;
assign w37711 = w36744 & ~w37710;
assign w37712 = w36687 & w36727;
assign w37713 = ~w36713 & ~w37712;
assign w37714 = ~w36726 & w37713;
assign w37715 = w36759 & w37714;
assign w37716 = (w36687 & w36756) | (w36687 & w63940) | (w36756 & w63940);
assign w37717 = w36693 & ~w36715;
assign w37718 = ~w36706 & w37717;
assign w37719 = ~w37716 & w37718;
assign w37720 = ~w36718 & ~w37711;
assign w37721 = ~w37715 & ~w37719;
assign w37722 = (~w37709 & ~w37721) | (~w37709 & w63941) | (~w37721 & w63941);
assign w37723 = w36712 & w36733;
assign w37724 = ~w36713 & ~w37723;
assign w37725 = w36693 & ~w37724;
assign w37726 = w36706 & w63942;
assign w37727 = ~w36742 & ~w37726;
assign w37728 = ~w36693 & ~w36712;
assign w37729 = w36699 & w36705;
assign w37730 = ~w36733 & ~w37729;
assign w37731 = w37728 & ~w37730;
assign w37732 = ~w36726 & ~w37731;
assign w37733 = ~w37725 & w37732;
assign w37734 = (~w36752 & ~w37733) | (~w36752 & w66215) | (~w37733 & w66215);
assign w37735 = ~w36687 & w36712;
assign w37736 = ~w37717 & w37735;
assign w37737 = w36687 & w36693;
assign w37738 = w37714 & w37737;
assign w37739 = (~w36752 & w37738) | (~w36752 & w63943) | (w37738 & w63943);
assign w37740 = w37714 & w66216;
assign w37741 = ~w36744 & ~w37712;
assign w37742 = (~w36693 & ~w37741) | (~w36693 & w63944) | (~w37741 & w63944);
assign w37743 = w36699 & w36720;
assign w37744 = w37727 & ~w37743;
assign w37745 = ~w37742 & w37744;
assign w37746 = ~w37740 & w37745;
assign w37747 = ~w36705 & w36721;
assign w37748 = (w37747 & w37746) | (w37747 & w63945) | (w37746 & w63945);
assign w37749 = ~w37722 & ~w37734;
assign w37750 = (pi1984 & ~w37749) | (pi1984 & w66217) | (~w37749 & w66217);
assign w37751 = w37749 & w66218;
assign w37752 = ~w37750 & ~w37751;
assign w37753 = ~w36730 & w36758;
assign w37754 = (w36752 & w37740) | (w36752 & w63946) | (w37740 & w63946);
assign w37755 = w36733 & w37728;
assign w37756 = (w37729 & w36742) | (w37729 & w66219) | (w36742 & w66219);
assign w37757 = ~w36739 & w66220;
assign w37758 = ~w37756 & ~w37757;
assign w37759 = w36687 & w36715;
assign w37760 = ~w37743 & ~w37759;
assign w37761 = w37758 & w37760;
assign w37762 = ~w36728 & ~w37755;
assign w37763 = ~w37761 & w37762;
assign w37764 = ~w36752 & ~w37763;
assign w37765 = ~w36719 & ~w36760;
assign w37766 = ~w37753 & w37765;
assign w37767 = ~w37754 & w37766;
assign w37768 = w37767 & w66221;
assign w37769 = (pi1996 & ~w37767) | (pi1996 & w66222) | (~w37767 & w66222);
assign w37770 = ~w37768 & ~w37769;
assign w37771 = w36805 & ~w36847;
assign w37772 = w36807 & w36811;
assign w37773 = w37312 & ~w37772;
assign w37774 = ~w37771 & ~w37773;
assign w37775 = w36816 & w36819;
assign w37776 = w36836 & ~w36844;
assign w37777 = w36823 & ~w37776;
assign w37778 = ~w36784 & ~w36811;
assign w37779 = ~w36848 & w37778;
assign w37780 = w37298 & ~w37779;
assign w37781 = w36832 & ~w37775;
assign w37782 = (w37781 & w37777) | (w37781 & w66223) | (w37777 & w66223);
assign w37783 = w37320 & ~w37776;
assign w37784 = ~w37776 & w63947;
assign w37785 = w36778 & ~w36842;
assign w37786 = w37318 & w63948;
assign w37787 = ~w37779 & w66224;
assign w37788 = ~w37783 & w37787;
assign w37789 = ~w36832 & ~w36847;
assign w37790 = ~w37784 & w37789;
assign w37791 = ~w37786 & w37790;
assign w37792 = ~w37788 & w37791;
assign w37793 = (~w37774 & w37792) | (~w37774 & w66225) | (w37792 & w66225);
assign w37794 = ~pi1976 & w37793;
assign w37795 = pi1976 & ~w37793;
assign w37796 = ~w37794 & ~w37795;
assign w37797 = ~pi6516 & pi9040;
assign w37798 = ~pi6487 & ~pi9040;
assign w37799 = ~w37797 & ~w37798;
assign w37800 = pi1937 & ~w37799;
assign w37801 = ~pi1937 & w37799;
assign w37802 = ~w37800 & ~w37801;
assign w37803 = ~pi6519 & pi9040;
assign w37804 = ~pi6605 & ~pi9040;
assign w37805 = ~w37803 & ~w37804;
assign w37806 = pi1949 & ~w37805;
assign w37807 = ~pi1949 & w37805;
assign w37808 = ~w37806 & ~w37807;
assign w37809 = ~w37802 & w37808;
assign w37810 = ~pi6529 & pi9040;
assign w37811 = ~pi6519 & ~pi9040;
assign w37812 = ~w37810 & ~w37811;
assign w37813 = pi1947 & ~w37812;
assign w37814 = ~pi1947 & w37812;
assign w37815 = ~w37813 & ~w37814;
assign w37816 = ~pi6487 & pi9040;
assign w37817 = ~pi6512 & ~pi9040;
assign w37818 = ~w37816 & ~w37817;
assign w37819 = pi1929 & ~w37818;
assign w37820 = ~pi1929 & w37818;
assign w37821 = ~w37819 & ~w37820;
assign w37822 = w37815 & w37821;
assign w37823 = ~pi6510 & pi9040;
assign w37824 = ~pi6511 & ~pi9040;
assign w37825 = ~w37823 & ~w37824;
assign w37826 = pi1922 & ~w37825;
assign w37827 = ~pi1922 & w37825;
assign w37828 = ~w37826 & ~w37827;
assign w37829 = w37822 & w37828;
assign w37830 = w37809 & w37829;
assign w37831 = ~w37802 & ~w37808;
assign w37832 = ~w37802 & w37815;
assign w37833 = w37802 & ~w37815;
assign w37834 = w37808 & ~w37833;
assign w37835 = ~w37832 & w37834;
assign w37836 = ~w37831 & ~w37835;
assign w37837 = ~pi6620 & pi9040;
assign w37838 = ~pi6496 & ~pi9040;
assign w37839 = ~w37837 & ~w37838;
assign w37840 = pi1919 & ~w37839;
assign w37841 = ~pi1919 & w37839;
assign w37842 = ~w37840 & ~w37841;
assign w37843 = ~w37836 & ~w37842;
assign w37844 = w37832 & w37842;
assign w37845 = (~w37808 & w37844) | (~w37808 & w66226) | (w37844 & w66226);
assign w37846 = ~w37835 & ~w37845;
assign w37847 = ~w37802 & ~w37815;
assign w37848 = ~w37842 & ~w37847;
assign w37849 = w37846 & ~w37848;
assign w37850 = ~w37843 & ~w37849;
assign w37851 = w37821 & w37831;
assign w37852 = ~w37828 & ~w37851;
assign w37853 = ~w37850 & w37852;
assign w37854 = ~w37821 & w37828;
assign w37855 = ~w37846 & w37854;
assign w37856 = w37821 & w37833;
assign w37857 = (w37842 & ~w37833) | (w37842 & w63949) | (~w37833 & w63949);
assign w37858 = w37821 & w37857;
assign w37859 = ~w37815 & ~w37821;
assign w37860 = ~w37822 & ~w37859;
assign w37861 = w37802 & ~w37808;
assign w37862 = ~w37809 & ~w37861;
assign w37863 = w37860 & w37862;
assign w37864 = ~w37808 & w37822;
assign w37865 = w37822 & w37861;
assign w37866 = ~w37863 & ~w37865;
assign w37867 = w37858 & ~w37866;
assign w37868 = ~w37821 & w37861;
assign w37869 = ~w37851 & ~w37868;
assign w37870 = w37828 & ~w37842;
assign w37871 = ~w37869 & w37870;
assign w37872 = ~w37842 & w37856;
assign w37873 = ~w37830 & ~w37872;
assign w37874 = ~w37871 & w37873;
assign w37875 = ~w37867 & w37874;
assign w37876 = ~w37855 & w37875;
assign w37877 = ~w37853 & w37876;
assign w37878 = pi1987 & w37877;
assign w37879 = ~pi1987 & ~w37877;
assign w37880 = ~w37878 & ~w37879;
assign w37881 = w37229 & ~w37248;
assign w37882 = ~w37222 & ~w37239;
assign w37883 = ~w37881 & ~w37882;
assign w37884 = w37222 & w37285;
assign w37885 = ~w37200 & ~w37262;
assign w37886 = w37270 & ~w37885;
assign w37887 = w37208 & ~w37253;
assign w37888 = ~w37884 & w37887;
assign w37889 = ~w37886 & w37888;
assign w37890 = ~w37213 & ~w37641;
assign w37891 = ~w37199 & ~w37266;
assign w37892 = ~w37890 & ~w37891;
assign w37893 = ~w37226 & w37251;
assign w37894 = ~w37892 & w37893;
assign w37895 = ~w37889 & ~w37894;
assign w37896 = ~w37883 & ~w37895;
assign w37897 = ~pi1995 & w37896;
assign w37898 = pi1995 & ~w37896;
assign w37899 = ~w37897 & ~w37898;
assign w37900 = ~w36687 & ~w36739;
assign w37901 = w37758 & w37900;
assign w37902 = ~w36714 & ~w37716;
assign w37903 = ~w37901 & w37902;
assign w37904 = w36752 & ~w37903;
assign w37905 = w36693 & w36727;
assign w37906 = ~w36725 & w37905;
assign w37907 = w36743 & ~w37714;
assign w37908 = ~w37906 & ~w37907;
assign w37909 = ~w37739 & w37908;
assign w37910 = ~w37904 & w37909;
assign w37911 = pi1994 & w37910;
assign w37912 = ~pi1994 & ~w37910;
assign w37913 = ~w37911 & ~w37912;
assign w37914 = w37802 & w37821;
assign w37915 = ~w37808 & w37815;
assign w37916 = ~w37914 & ~w37915;
assign w37917 = ~w37842 & ~w37916;
assign w37918 = w37834 & w37917;
assign w37919 = w37857 & w66227;
assign w37920 = w37859 & w37861;
assign w37921 = ~w37919 & ~w37920;
assign w37922 = w37809 & ~w37821;
assign w37923 = ~w37851 & ~w37922;
assign w37924 = w37857 & w37923;
assign w37925 = w37859 & w37862;
assign w37926 = w37809 & w37821;
assign w37927 = w37815 & w37861;
assign w37928 = ~w37926 & ~w37927;
assign w37929 = (~w37842 & ~w37862) | (~w37842 & w63413) | (~w37862 & w63413);
assign w37930 = w37928 & w37929;
assign w37931 = ~w37924 & ~w37930;
assign w37932 = ~w37848 & w37859;
assign w37933 = (~w37931 & w66228) | (~w37931 & w66229) | (w66228 & w66229);
assign w37934 = w37845 & w37921;
assign w37935 = ~w37931 & ~w37934;
assign w37936 = ~w37828 & ~w37935;
assign w37937 = ~w37821 & w37844;
assign w37938 = ~w37920 & ~w37937;
assign w37939 = ~w37864 & ~w37916;
assign w37940 = ~w37848 & ~w37939;
assign w37941 = ~w37938 & w37940;
assign w37942 = ~w37859 & w37870;
assign w37943 = w37862 & w37942;
assign w37944 = ~w37918 & ~w37943;
assign w37945 = ~w37941 & w37944;
assign w37946 = ~w37933 & w37945;
assign w37947 = ~w37936 & w37946;
assign w37948 = pi1979 & ~w37947;
assign w37949 = ~pi1979 & w37947;
assign w37950 = ~w37948 & ~w37949;
assign w37951 = w37829 & w37831;
assign w37952 = w37809 & ~w37842;
assign w37953 = ~w37860 & w37952;
assign w37954 = w37866 & ~w37953;
assign w37955 = (~w37828 & ~w37954) | (~w37828 & w66230) | (~w37954 & w66230);
assign w37956 = w37847 & w37923;
assign w37957 = w37808 & ~w37815;
assign w37958 = w37928 & ~w37957;
assign w37959 = w37828 & ~w37958;
assign w37960 = w37914 & w37957;
assign w37961 = ~w37956 & ~w37960;
assign w37962 = ~w37959 & w37961;
assign w37963 = w37842 & ~w37962;
assign w37964 = ~w37831 & w37870;
assign w37965 = w37958 & w37964;
assign w37966 = ~w37951 & ~w37965;
assign w37967 = ~w37955 & w37966;
assign w37968 = ~w37963 & w37967;
assign w37969 = pi1977 & w37968;
assign w37970 = ~pi1977 & ~w37968;
assign w37971 = ~w37969 & ~w37970;
assign w37972 = w37829 & ~w37939;
assign w37973 = (w37828 & ~w37923) | (w37828 & w64441) | (~w37923 & w64441);
assign w37974 = ~w37960 & ~w37973;
assign w37975 = w37842 & ~w37974;
assign w37976 = ~w37917 & ~w37940;
assign w37977 = ~w37925 & ~w37956;
assign w37978 = ~w37976 & w37977;
assign w37979 = ~w37828 & ~w37978;
assign w37980 = ~w37828 & ~w37864;
assign w37981 = ~w37868 & w37917;
assign w37982 = ~w37980 & w37981;
assign w37983 = ~w37972 & ~w37982;
assign w37984 = ~w37975 & w37983;
assign w37985 = ~w37979 & w37984;
assign w37986 = pi1988 & ~w37985;
assign w37987 = ~pi1988 & w37985;
assign w37988 = ~w37986 & ~w37987;
assign w37989 = ~pi6720 & pi9040;
assign w37990 = ~pi6759 & ~pi9040;
assign w37991 = ~w37989 & ~w37990;
assign w37992 = pi1985 & ~w37991;
assign w37993 = ~pi1985 & w37991;
assign w37994 = ~w37992 & ~w37993;
assign w37995 = ~pi6724 & pi9040;
assign w37996 = ~pi6779 & ~pi9040;
assign w37997 = ~w37995 & ~w37996;
assign w37998 = pi1972 & ~w37997;
assign w37999 = ~pi1972 & w37997;
assign w38000 = ~w37998 & ~w37999;
assign w38001 = ~pi6742 & pi9040;
assign w38002 = ~pi6775 & ~pi9040;
assign w38003 = ~w38001 & ~w38002;
assign w38004 = pi2008 & ~w38003;
assign w38005 = ~pi2008 & w38003;
assign w38006 = ~w38004 & ~w38005;
assign w38007 = ~pi6758 & pi9040;
assign w38008 = ~pi6725 & ~pi9040;
assign w38009 = ~w38007 & ~w38008;
assign w38010 = pi2003 & ~w38009;
assign w38011 = ~pi2003 & w38009;
assign w38012 = ~w38010 & ~w38011;
assign w38013 = ~w38006 & ~w38012;
assign w38014 = ~pi6767 & pi9040;
assign w38015 = ~pi6761 & ~pi9040;
assign w38016 = ~w38014 & ~w38015;
assign w38017 = pi1991 & ~w38016;
assign w38018 = ~pi1991 & w38016;
assign w38019 = ~w38017 & ~w38018;
assign w38020 = w38013 & w38019;
assign w38021 = w38013 & w66231;
assign w38022 = ~w37994 & w38021;
assign w38023 = ~w38006 & w38019;
assign w38024 = w38000 & ~w38012;
assign w38025 = ~w38023 & ~w38024;
assign w38026 = w38000 & ~w38019;
assign w38027 = w38006 & w38026;
assign w38028 = ~w38000 & w38012;
assign w38029 = ~w38027 & ~w38028;
assign w38030 = ~w38025 & ~w38029;
assign w38031 = ~w38000 & ~w38019;
assign w38032 = w38006 & ~w38012;
assign w38033 = ~w38000 & w38019;
assign w38034 = ~w38026 & ~w38033;
assign w38035 = w38032 & w38034;
assign w38036 = ~w38006 & w38031;
assign w38037 = w38031 & w66232;
assign w38038 = ~w38035 & ~w38037;
assign w38039 = ~w38035 & w66233;
assign w38040 = ~w38030 & ~w38039;
assign w38041 = w37994 & ~w38040;
assign w38042 = ~w37994 & w38012;
assign w38043 = w38012 & w38019;
assign w38044 = ~w38042 & ~w38043;
assign w38045 = (~w38023 & w38044) | (~w38023 & w66234) | (w38044 & w66234);
assign w38046 = w37994 & ~w38025;
assign w38047 = ~w38021 & w38046;
assign w38048 = ~w37994 & ~w38019;
assign w38049 = w38032 & w38048;
assign w38050 = ~w38012 & ~w38019;
assign w38051 = w38034 & ~w38050;
assign w38052 = w38006 & w38033;
assign w38053 = ~w38012 & w38052;
assign w38054 = ~w38051 & ~w38053;
assign w38055 = w37994 & ~w38000;
assign w38056 = ~w38054 & w38055;
assign w38057 = ~pi6759 & pi9040;
assign w38058 = ~pi6742 & ~pi9040;
assign w38059 = ~w38057 & ~w38058;
assign w38060 = pi2013 & ~w38059;
assign w38061 = ~pi2013 & w38059;
assign w38062 = ~w38060 & ~w38061;
assign w38063 = ~w38049 & ~w38062;
assign w38064 = (w38063 & w38047) | (w38063 & w66235) | (w38047 & w66235);
assign w38065 = ~w38056 & w38064;
assign w38066 = w38006 & w38012;
assign w38067 = w38026 & w38066;
assign w38068 = w38062 & ~w38067;
assign w38069 = ~w38036 & ~w38052;
assign w38070 = ~w37994 & ~w38069;
assign w38071 = ~w38047 & w38068;
assign w38072 = ~w38070 & w38071;
assign w38073 = ~w38065 & ~w38072;
assign w38074 = ~w38022 & ~w38041;
assign w38075 = ~w38073 & w38074;
assign w38076 = ~pi2019 & w38075;
assign w38077 = pi2019 & ~w38075;
assign w38078 = ~w38076 & ~w38077;
assign w38079 = ~pi6773 & pi9040;
assign w38080 = ~pi6762 & ~pi9040;
assign w38081 = ~w38079 & ~w38080;
assign w38082 = pi2006 & ~w38081;
assign w38083 = ~pi2006 & w38081;
assign w38084 = ~w38082 & ~w38083;
assign w38085 = ~pi6761 & pi9040;
assign w38086 = ~pi6758 & ~pi9040;
assign w38087 = ~w38085 & ~w38086;
assign w38088 = pi1975 & ~w38087;
assign w38089 = ~pi1975 & w38087;
assign w38090 = ~w38088 & ~w38089;
assign w38091 = ~w38084 & w38090;
assign w38092 = w38084 & ~w38090;
assign w38093 = ~w38091 & ~w38092;
assign w38094 = ~pi6757 & pi9040;
assign w38095 = ~pi6724 & ~pi9040;
assign w38096 = ~w38094 & ~w38095;
assign w38097 = pi1999 & ~w38096;
assign w38098 = ~pi1999 & w38096;
assign w38099 = ~w38097 & ~w38098;
assign w38100 = ~pi6827 & pi9040;
assign w38101 = ~pi6757 & ~pi9040;
assign w38102 = ~w38100 & ~w38101;
assign w38103 = pi2009 & ~w38102;
assign w38104 = ~pi2009 & w38102;
assign w38105 = ~w38103 & ~w38104;
assign w38106 = w38099 & ~w38105;
assign w38107 = w38093 & w38106;
assign w38108 = ~pi6725 & pi9040;
assign w38109 = ~pi6767 & ~pi9040;
assign w38110 = ~w38108 & ~w38109;
assign w38111 = pi1972 & ~w38110;
assign w38112 = ~pi1972 & w38110;
assign w38113 = ~w38111 & ~w38112;
assign w38114 = ~w38099 & ~w38113;
assign w38115 = ~w38084 & w38114;
assign w38116 = w38090 & w38115;
assign w38117 = w38105 & ~w38116;
assign w38118 = w38099 & w38113;
assign w38119 = ~w38114 & ~w38118;
assign w38120 = w38091 & w38119;
assign w38121 = ~w38114 & ~w38120;
assign w38122 = w38117 & ~w38121;
assign w38123 = ~w38105 & w38113;
assign w38124 = ~w38118 & ~w38123;
assign w38125 = w38093 & ~w38124;
assign w38126 = ~w38093 & ~w38099;
assign w38127 = ~w38105 & ~w38119;
assign w38128 = w38092 & w38114;
assign w38129 = w38127 & ~w38128;
assign w38130 = w38084 & ~w38113;
assign w38131 = ~w38084 & w38113;
assign w38132 = ~w38130 & ~w38131;
assign w38133 = ~w38114 & w38132;
assign w38134 = w38132 & w63414;
assign w38135 = w38105 & ~w38134;
assign w38136 = ~w38126 & ~w38133;
assign w38137 = w38091 & w38099;
assign w38138 = ~w38105 & ~w38137;
assign w38139 = ~w38136 & w38138;
assign w38140 = (~w38129 & w38139) | (~w38129 & w63415) | (w38139 & w63415);
assign w38141 = w38106 & w38130;
assign w38142 = ~pi6778 & pi9040;
assign w38143 = ~pi6821 & ~pi9040;
assign w38144 = ~w38142 & ~w38143;
assign w38145 = pi1991 & ~w38144;
assign w38146 = ~pi1991 & w38144;
assign w38147 = ~w38145 & ~w38146;
assign w38148 = ~w38128 & ~w38147;
assign w38149 = ~w38125 & ~w38141;
assign w38150 = w38148 & w38149;
assign w38151 = (w38150 & w38140) | (w38150 & w63951) | (w38140 & w63951);
assign w38152 = ~w38099 & w38113;
assign w38153 = w38092 & w38152;
assign w38154 = w38099 & ~w38132;
assign w38155 = ~w38153 & ~w38154;
assign w38156 = w38123 & ~w38155;
assign w38157 = w38114 & w66236;
assign w38158 = w38090 & ~w38099;
assign w38159 = w38131 & w38158;
assign w38160 = ~w38157 & ~w38159;
assign w38161 = ~w38090 & w38118;
assign w38162 = ~w38158 & ~w38161;
assign w38163 = w38084 & w38105;
assign w38164 = ~w38162 & w38163;
assign w38165 = w38147 & w38160;
assign w38166 = ~w38164 & w38165;
assign w38167 = ~w38156 & w38166;
assign w38168 = ~w38107 & ~w38122;
assign w38169 = (w38168 & w38151) | (w38168 & w66237) | (w38151 & w66237);
assign w38170 = pi2028 & w38169;
assign w38171 = ~pi2028 & ~w38169;
assign w38172 = ~w38170 & ~w38171;
assign w38173 = ~pi6754 & pi9040;
assign w38174 = ~pi6773 & ~pi9040;
assign w38175 = ~w38173 & ~w38174;
assign w38176 = pi1982 & ~w38175;
assign w38177 = ~pi1982 & w38175;
assign w38178 = ~w38176 & ~w38177;
assign w38179 = ~pi6764 & pi9040;
assign w38180 = ~pi6744 & ~pi9040;
assign w38181 = ~w38179 & ~w38180;
assign w38182 = pi1999 & ~w38181;
assign w38183 = ~pi1999 & w38181;
assign w38184 = ~w38182 & ~w38183;
assign w38185 = w38178 & w38184;
assign w38186 = ~pi6855 & pi9040;
assign w38187 = ~pi6754 & ~pi9040;
assign w38188 = ~w38186 & ~w38187;
assign w38189 = pi1983 & ~w38188;
assign w38190 = ~pi1983 & w38188;
assign w38191 = ~w38189 & ~w38190;
assign w38192 = ~pi6733 & pi9040;
assign w38193 = ~pi6854 & ~pi9040;
assign w38194 = ~w38192 & ~w38193;
assign w38195 = pi2010 & ~w38194;
assign w38196 = ~pi2010 & w38194;
assign w38197 = ~w38195 & ~w38196;
assign w38198 = ~w38191 & ~w38197;
assign w38199 = ~w38178 & ~w38184;
assign w38200 = w38198 & ~w38199;
assign w38201 = ~w38185 & w38200;
assign w38202 = ~w38184 & w38191;
assign w38203 = ~pi6719 & pi9040;
assign w38204 = ~pi6753 & ~pi9040;
assign w38205 = ~w38203 & ~w38204;
assign w38206 = pi2002 & ~w38205;
assign w38207 = ~pi2002 & w38205;
assign w38208 = ~w38206 & ~w38207;
assign w38209 = ~w38178 & ~w38208;
assign w38210 = w38202 & w38209;
assign w38211 = ~w38201 & ~w38210;
assign w38212 = w38184 & w38208;
assign w38213 = w38198 & w38212;
assign w38214 = w38197 & w38199;
assign w38215 = ~w38213 & ~w38214;
assign w38216 = ~w38211 & ~w38215;
assign w38217 = w38184 & w38191;
assign w38218 = w38178 & w38217;
assign w38219 = w38178 & w38197;
assign w38220 = ~w38178 & w38191;
assign w38221 = w38178 & ~w38191;
assign w38222 = ~w38220 & ~w38221;
assign w38223 = ~w38219 & w38222;
assign w38224 = ~pi6854 & pi9040;
assign w38225 = ~pi6776 & ~pi9040;
assign w38226 = ~w38224 & ~w38225;
assign w38227 = pi2006 & ~w38226;
assign w38228 = ~pi2006 & w38226;
assign w38229 = ~w38227 & ~w38228;
assign w38230 = ~w38191 & w38199;
assign w38231 = w38199 & w63952;
assign w38232 = w38229 & ~w38231;
assign w38233 = w38223 & ~w38232;
assign w38234 = w38184 & ~w38197;
assign w38235 = ~w38184 & w38197;
assign w38236 = ~w38234 & ~w38235;
assign w38237 = w38191 & w38236;
assign w38238 = (~w38219 & ~w38236) | (~w38219 & w66238) | (~w38236 & w66238);
assign w38239 = ~w38198 & ~w38202;
assign w38240 = w38178 & ~w38239;
assign w38241 = (w38229 & w38239) | (w38229 & w66239) | (w38239 & w66239);
assign w38242 = ~w38238 & w38241;
assign w38243 = ~w38218 & ~w38233;
assign w38244 = (w38208 & ~w38243) | (w38208 & w66240) | (~w38243 & w66240);
assign w38245 = ~w38178 & w38197;
assign w38246 = ~w38184 & ~w38191;
assign w38247 = ~w38245 & w38246;
assign w38248 = ~w38218 & ~w38247;
assign w38249 = w38208 & ~w38245;
assign w38250 = ~w38234 & w38249;
assign w38251 = ~w38248 & ~w38250;
assign w38252 = ~w38178 & w38251;
assign w38253 = ~w38191 & ~w38208;
assign w38254 = w38236 & w66241;
assign w38255 = w38209 & w38217;
assign w38256 = ~w38197 & w38255;
assign w38257 = ~w38240 & ~w38256;
assign w38258 = (~w38208 & ~w38257) | (~w38208 & w66242) | (~w38257 & w66242);
assign w38259 = w38229 & ~w38258;
assign w38260 = w38197 & ~w38208;
assign w38261 = ~w38222 & w38260;
assign w38262 = (w38191 & w38245) | (w38191 & w66243) | (w38245 & w66243);
assign w38263 = w38199 & w38262;
assign w38264 = ~w38197 & w38218;
assign w38265 = ~w38213 & ~w38229;
assign w38266 = ~w38261 & w38265;
assign w38267 = ~w38264 & w38266;
assign w38268 = ~w38263 & w38267;
assign w38269 = ~w38259 & ~w38268;
assign w38270 = ~w38216 & ~w38252;
assign w38271 = ~w38244 & w38270;
assign w38272 = ~w38269 & w38271;
assign w38273 = pi2039 & ~w38272;
assign w38274 = ~pi2039 & w38272;
assign w38275 = ~w38273 & ~w38274;
assign w38276 = w38199 & w38237;
assign w38277 = w38212 & w38245;
assign w38278 = ~w38260 & w38262;
assign w38279 = ~w38201 & ~w38278;
assign w38280 = w38197 & w38208;
assign w38281 = w38248 & w38280;
assign w38282 = w38279 & w38281;
assign w38283 = ~w38201 & w66244;
assign w38284 = ~w38251 & w38283;
assign w38285 = ~w38282 & w38284;
assign w38286 = ~w38184 & ~w38260;
assign w38287 = w38240 & ~w38286;
assign w38288 = ~w38200 & w38247;
assign w38289 = ~w38237 & ~w38288;
assign w38290 = w38208 & ~w38289;
assign w38291 = w38209 & w38239;
assign w38292 = ~w38229 & ~w38291;
assign w38293 = ~w38287 & w38292;
assign w38294 = ~w38290 & w38293;
assign w38295 = ~w38285 & ~w38294;
assign w38296 = ~w38276 & ~w38277;
assign w38297 = ~w38295 & w38296;
assign w38298 = ~pi2023 & w38297;
assign w38299 = pi2023 & ~w38297;
assign w38300 = ~w38298 & ~w38299;
assign w38301 = w38090 & w38130;
assign w38302 = ~w38137 & ~w38301;
assign w38303 = ~w38154 & ~w38302;
assign w38304 = w38084 & w38090;
assign w38305 = w38105 & w38152;
assign w38306 = ~w38304 & ~w38305;
assign w38307 = ~w38129 & w38306;
assign w38308 = ~w38160 & w38307;
assign w38309 = ~w38091 & w38131;
assign w38310 = ~w38163 & ~w38309;
assign w38311 = w38099 & ~w38310;
assign w38312 = w38147 & ~w38153;
assign w38313 = ~w38303 & w38312;
assign w38314 = ~w38311 & w38313;
assign w38315 = ~w38308 & w38314;
assign w38316 = ~w38116 & ~w38134;
assign w38317 = ~w38084 & ~w38316;
assign w38318 = ~w38163 & ~w38306;
assign w38319 = ~w38132 & w66245;
assign w38320 = w38152 & w38304;
assign w38321 = ~w38319 & ~w38320;
assign w38322 = w38113 & ~w38321;
assign w38323 = ~w38127 & w38148;
assign w38324 = ~w38318 & w38323;
assign w38325 = ~w38317 & w38324;
assign w38326 = ~w38322 & w38325;
assign w38327 = ~w38315 & ~w38326;
assign w38328 = ~pi2040 & w38327;
assign w38329 = pi2040 & ~w38327;
assign w38330 = ~w38328 & ~w38329;
assign w38331 = ~pi6858 & pi9040;
assign w38332 = ~pi6719 & ~pi9040;
assign w38333 = ~w38331 & ~w38332;
assign w38334 = pi1992 & ~w38333;
assign w38335 = ~pi1992 & w38333;
assign w38336 = ~w38334 & ~w38335;
assign w38337 = ~pi6821 & pi9040;
assign w38338 = ~pi6764 & ~pi9040;
assign w38339 = ~w38337 & ~w38338;
assign w38340 = pi2010 & ~w38339;
assign w38341 = ~pi2010 & w38339;
assign w38342 = ~w38340 & ~w38341;
assign w38343 = w38336 & w38342;
assign w38344 = ~pi6744 & pi9040;
assign w38345 = ~pi6778 & ~pi9040;
assign w38346 = ~w38344 & ~w38345;
assign w38347 = pi2012 & ~w38346;
assign w38348 = ~pi2012 & w38346;
assign w38349 = ~w38347 & ~w38348;
assign w38350 = ~pi6941 & pi9040;
assign w38351 = ~pi6858 & ~pi9040;
assign w38352 = ~w38350 & ~w38351;
assign w38353 = pi2014 & ~w38352;
assign w38354 = ~pi2014 & w38352;
assign w38355 = ~w38353 & ~w38354;
assign w38356 = w38349 & ~w38355;
assign w38357 = w38343 & w38356;
assign w38358 = ~pi6770 & pi9040;
assign w38359 = ~pi6733 & ~pi9040;
assign w38360 = ~w38358 & ~w38359;
assign w38361 = pi1983 & ~w38360;
assign w38362 = ~pi1983 & w38360;
assign w38363 = ~w38361 & ~w38362;
assign w38364 = w38336 & ~w38355;
assign w38365 = ~pi6762 & pi9040;
assign w38366 = ~pi6855 & ~pi9040;
assign w38367 = ~w38365 & ~w38366;
assign w38368 = pi1981 & ~w38367;
assign w38369 = ~pi1981 & w38367;
assign w38370 = ~w38368 & ~w38369;
assign w38371 = ~w38343 & w38370;
assign w38372 = ~w38364 & w38371;
assign w38373 = ~w38349 & w38372;
assign w38374 = w38349 & w38355;
assign w38375 = w38336 & ~w38342;
assign w38376 = w38374 & w38375;
assign w38377 = w38342 & w38364;
assign w38378 = ~w38376 & ~w38377;
assign w38379 = w38343 & w38349;
assign w38380 = ~w38336 & ~w38342;
assign w38381 = w38356 & w38380;
assign w38382 = ~w38379 & ~w38381;
assign w38383 = w38370 & ~w38382;
assign w38384 = ~w38336 & w38342;
assign w38385 = w38349 & w38384;
assign w38386 = ~w38349 & ~w38355;
assign w38387 = w38336 & w38386;
assign w38388 = ~w38385 & ~w38387;
assign w38389 = ~w38370 & ~w38388;
assign w38390 = ~w38373 & w38378;
assign w38391 = ~w38383 & ~w38389;
assign w38392 = w38390 & w38391;
assign w38393 = w38363 & ~w38392;
assign w38394 = (w38370 & ~w38386) | (w38370 & w66246) | (~w38386 & w66246);
assign w38395 = w38342 & w38386;
assign w38396 = ~w38349 & w38355;
assign w38397 = w38380 & w38396;
assign w38398 = ~w38376 & ~w38397;
assign w38399 = ~w38395 & w38398;
assign w38400 = w38394 & ~w38399;
assign w38401 = w38336 & ~w38396;
assign w38402 = ~w38371 & w38401;
assign w38403 = ~w38342 & w38349;
assign w38404 = ~w38336 & ~w38386;
assign w38405 = ~w38403 & w38404;
assign w38406 = ~w38363 & ~w38405;
assign w38407 = ~w38374 & ~w38406;
assign w38408 = ~w38372 & ~w38402;
assign w38409 = ~w38407 & w38408;
assign w38410 = ~w38357 & ~w38400;
assign w38411 = ~w38409 & w38410;
assign w38412 = ~w38393 & w38411;
assign w38413 = pi2018 & w38412;
assign w38414 = ~pi2018 & ~w38412;
assign w38415 = ~w38413 & ~w38414;
assign w38416 = ~pi6715 & pi9040;
assign w38417 = ~pi6747 & ~pi9040;
assign w38418 = ~w38416 & ~w38417;
assign w38419 = pi1992 & ~w38418;
assign w38420 = ~pi1992 & w38418;
assign w38421 = ~w38419 & ~w38420;
assign w38422 = ~pi6857 & pi9040;
assign w38423 = ~pi6746 & ~pi9040;
assign w38424 = ~w38422 & ~w38423;
assign w38425 = pi2015 & ~w38424;
assign w38426 = ~pi2015 & w38424;
assign w38427 = ~w38425 & ~w38426;
assign w38428 = w38421 & w38427;
assign w38429 = ~pi6859 & pi9040;
assign w38430 = ~pi6780 & ~pi9040;
assign w38431 = ~w38429 & ~w38430;
assign w38432 = pi1990 & ~w38431;
assign w38433 = ~pi1990 & w38431;
assign w38434 = ~w38432 & ~w38433;
assign w38435 = w38421 & ~w38434;
assign w38436 = ~pi6782 & pi9040;
assign w38437 = ~pi6857 & ~pi9040;
assign w38438 = ~w38436 & ~w38437;
assign w38439 = pi2001 & ~w38438;
assign w38440 = ~pi2001 & w38438;
assign w38441 = ~w38439 & ~w38440;
assign w38442 = ~pi6752 & pi9040;
assign w38443 = ~pi6760 & ~pi9040;
assign w38444 = ~w38442 & ~w38443;
assign w38445 = pi2011 & ~w38444;
assign w38446 = ~pi2011 & w38444;
assign w38447 = ~w38445 & ~w38446;
assign w38448 = ~w38441 & w38447;
assign w38449 = w38435 & w38448;
assign w38450 = w38434 & ~w38447;
assign w38451 = ~w38441 & w38450;
assign w38452 = ~w38449 & ~w38451;
assign w38453 = w38428 & ~w38452;
assign w38454 = ~pi6746 & pi9040;
assign w38455 = ~pi6716 & ~pi9040;
assign w38456 = ~w38454 & ~w38455;
assign w38457 = pi2012 & ~w38456;
assign w38458 = ~pi2012 & w38456;
assign w38459 = ~w38457 & ~w38458;
assign w38460 = ~w38421 & ~w38434;
assign w38461 = ~w38447 & w38460;
assign w38462 = w38427 & w38461;
assign w38463 = ~w38427 & w38441;
assign w38464 = w38421 & w38434;
assign w38465 = w38463 & w38464;
assign w38466 = ~w38460 & ~w38464;
assign w38467 = ~w38427 & ~w38447;
assign w38468 = w38441 & ~w38450;
assign w38469 = ~w38467 & w38468;
assign w38470 = w38466 & w38469;
assign w38471 = w38461 & w38463;
assign w38472 = ~w38441 & ~w38450;
assign w38473 = ~w38428 & ~w38434;
assign w38474 = w38472 & ~w38473;
assign w38475 = w38447 & w38460;
assign w38476 = w38460 & w66247;
assign w38477 = ~w38441 & w38460;
assign w38478 = w38460 & w66248;
assign w38479 = ~w38476 & ~w38478;
assign w38480 = ~w38427 & ~w38441;
assign w38481 = w38464 & w38480;
assign w38482 = ~w38471 & ~w38481;
assign w38483 = ~w38474 & w38482;
assign w38484 = w38482 & w66249;
assign w38485 = ~w38449 & w38472;
assign w38486 = w38483 & w63953;
assign w38487 = ~w38462 & ~w38465;
assign w38488 = ~w38470 & w38487;
assign w38489 = (w38459 & w38486) | (w38459 & w66250) | (w38486 & w66250);
assign w38490 = w38427 & w38447;
assign w38491 = w38434 & w38490;
assign w38492 = ~w38467 & ~w38491;
assign w38493 = ~w38434 & w38441;
assign w38494 = w38421 & ~w38493;
assign w38495 = ~w38492 & ~w38494;
assign w38496 = ~w38435 & w38441;
assign w38497 = w38490 & w38496;
assign w38498 = w38452 & ~w38497;
assign w38499 = ~w38495 & w38498;
assign w38500 = w38448 & w38466;
assign w38501 = ~w38434 & w38447;
assign w38502 = ~w38450 & ~w38501;
assign w38503 = w38441 & w38502;
assign w38504 = w38502 & w66251;
assign w38505 = w38447 & w38504;
assign w38506 = ~w38500 & ~w38505;
assign w38507 = (w38421 & w38491) | (w38421 & w66252) | (w38491 & w66252);
assign w38508 = w38479 & ~w38507;
assign w38509 = w38480 & w38508;
assign w38510 = w38506 & w38509;
assign w38511 = (~w38453 & w38499) | (~w38453 & w66253) | (w38499 & w66253);
assign w38512 = ~w38510 & w38511;
assign w38513 = ~w38489 & w38512;
assign w38514 = pi2021 & ~w38513;
assign w38515 = ~pi2021 & w38513;
assign w38516 = ~w38514 & ~w38515;
assign w38517 = ~pi6741 & pi9040;
assign w38518 = ~pi6743 & ~pi9040;
assign w38519 = ~w38517 & ~w38518;
assign w38520 = pi2003 & ~w38519;
assign w38521 = ~pi2003 & w38519;
assign w38522 = ~w38520 & ~w38521;
assign w38523 = ~pi6750 & pi9040;
assign w38524 = ~pi6741 & ~pi9040;
assign w38525 = ~w38523 & ~w38524;
assign w38526 = pi2007 & ~w38525;
assign w38527 = ~pi2007 & w38525;
assign w38528 = ~w38526 & ~w38527;
assign w38529 = ~w38522 & w38528;
assign w38530 = ~pi6749 & pi9040;
assign w38531 = ~pi6752 & ~pi9040;
assign w38532 = ~w38530 & ~w38531;
assign w38533 = pi2013 & ~w38532;
assign w38534 = ~pi2013 & w38532;
assign w38535 = ~w38533 & ~w38534;
assign w38536 = ~pi6717 & pi9040;
assign w38537 = ~pi6772 & ~pi9040;
assign w38538 = ~w38536 & ~w38537;
assign w38539 = pi1998 & ~w38538;
assign w38540 = ~pi1998 & w38538;
assign w38541 = ~w38539 & ~w38540;
assign w38542 = w38535 & ~w38541;
assign w38543 = w38529 & w38542;
assign w38544 = w38522 & ~w38535;
assign w38545 = w38528 & ~w38535;
assign w38546 = ~pi6751 & pi9040;
assign w38547 = ~pi6756 & ~pi9040;
assign w38548 = ~w38546 & ~w38547;
assign w38549 = pi1974 & ~w38548;
assign w38550 = ~pi1974 & w38548;
assign w38551 = ~w38549 & ~w38550;
assign w38552 = ~w38545 & w38551;
assign w38553 = ~w38541 & ~w38551;
assign w38554 = w38541 & w38551;
assign w38555 = ~w38553 & ~w38554;
assign w38556 = ~w38552 & ~w38555;
assign w38557 = w38544 & w38556;
assign w38558 = ~w38522 & ~w38551;
assign w38559 = ~w38544 & ~w38558;
assign w38560 = w38522 & w38535;
assign w38561 = ~w38528 & w38560;
assign w38562 = ~w38522 & ~w38535;
assign w38563 = ~w38553 & w38562;
assign w38564 = ~w38561 & ~w38563;
assign w38565 = w38564 & w63954;
assign w38566 = ~w38557 & ~w38565;
assign w38567 = ~pi6771 & pi9040;
assign w38568 = ~pi6852 & ~pi9040;
assign w38569 = ~w38567 & ~w38568;
assign w38570 = pi1989 & ~w38569;
assign w38571 = ~pi1989 & w38569;
assign w38572 = ~w38570 & ~w38571;
assign w38573 = ~w38566 & ~w38572;
assign w38574 = ~w38522 & w38535;
assign w38575 = ~w38558 & ~w38574;
assign w38576 = ~w38555 & w38575;
assign w38577 = w38522 & w38551;
assign w38578 = ~w38558 & ~w38577;
assign w38579 = ~w38560 & ~w38578;
assign w38580 = w38576 & ~w38579;
assign w38581 = ~w38535 & w38541;
assign w38582 = ~w38542 & ~w38581;
assign w38583 = ~w38559 & ~w38572;
assign w38584 = w38582 & w38583;
assign w38585 = ~w38580 & ~w38584;
assign w38586 = w38541 & ~w38551;
assign w38587 = w38545 & w38586;
assign w38588 = ~w38551 & ~w38574;
assign w38589 = (~w38541 & w38545) | (~w38541 & w38553) | (w38545 & w38553);
assign w38590 = ~w38588 & w38589;
assign w38591 = w38529 & w38551;
assign w38592 = ~w38587 & ~w38591;
assign w38593 = w38564 & w38592;
assign w38594 = ~w38590 & w38593;
assign w38595 = w38572 & ~w38594;
assign w38596 = ~w38522 & w38587;
assign w38597 = ~w38543 & ~w38596;
assign w38598 = (w38597 & w38585) | (w38597 & w66254) | (w38585 & w66254);
assign w38599 = ~w38595 & w38598;
assign w38600 = ~w38573 & w38599;
assign w38601 = pi2038 & ~w38600;
assign w38602 = ~pi2038 & w38600;
assign w38603 = ~w38601 & ~w38602;
assign w38604 = ~w38427 & ~w38449;
assign w38605 = ~w38421 & ~w38441;
assign w38606 = w38502 & w38605;
assign w38607 = w38421 & ~w38447;
assign w38608 = ~w38605 & ~w38607;
assign w38609 = (w38427 & ~w38608) | (w38427 & w66255) | (~w38608 & w66255);
assign w38610 = ~w38606 & w38609;
assign w38611 = ~w38604 & ~w38610;
assign w38612 = w38450 & w66256;
assign w38613 = ~w38421 & w38434;
assign w38614 = w38463 & w38613;
assign w38615 = w38490 & w38493;
assign w38616 = ~w38459 & ~w38614;
assign w38617 = ~w38615 & w38616;
assign w38618 = ~w38462 & ~w38612;
assign w38619 = w38617 & w38618;
assign w38620 = w38508 & w38619;
assign w38621 = w38427 & w38466;
assign w38622 = w38502 & w38621;
assign w38623 = w38480 & ~w38502;
assign w38624 = ~w38449 & w38459;
assign w38625 = ~w38471 & w38624;
assign w38626 = ~w38623 & w38625;
assign w38627 = w38626 & w66257;
assign w38628 = ~w38620 & ~w38627;
assign w38629 = ~w38611 & ~w38628;
assign w38630 = ~pi2017 & w38629;
assign w38631 = pi2017 & ~w38629;
assign w38632 = ~w38630 & ~w38631;
assign w38633 = w38250 & w38289;
assign w38634 = ~w38191 & ~w38229;
assign w38635 = ~w38236 & w38634;
assign w38636 = ~w38237 & ~w38635;
assign w38637 = (~w38230 & w38636) | (~w38230 & w66258) | (w38636 & w66258);
assign w38638 = ~w38208 & ~w38637;
assign w38639 = w38202 & w38280;
assign w38640 = w38212 & w38223;
assign w38641 = ~w38229 & ~w38255;
assign w38642 = ~w38639 & w38641;
assign w38643 = ~w38276 & w38642;
assign w38644 = ~w38640 & w38643;
assign w38645 = w38185 & w38197;
assign w38646 = w38212 & w38220;
assign w38647 = w38209 & ~w38217;
assign w38648 = ~w38276 & w38647;
assign w38649 = ~w38645 & ~w38646;
assign w38650 = w38232 & w38649;
assign w38651 = ~w38648 & w38650;
assign w38652 = ~w38644 & ~w38651;
assign w38653 = ~w38633 & ~w38638;
assign w38654 = ~w38652 & w38653;
assign w38655 = pi2027 & ~w38654;
assign w38656 = ~pi2027 & w38654;
assign w38657 = ~w38655 & ~w38656;
assign w38658 = ~pi6716 & pi9040;
assign w38659 = ~pi6782 & ~pi9040;
assign w38660 = ~w38658 & ~w38659;
assign w38661 = pi2005 & ~w38660;
assign w38662 = ~pi2005 & w38660;
assign w38663 = ~w38661 & ~w38662;
assign w38664 = ~pi6777 & pi9040;
assign w38665 = ~pi6849 & ~pi9040;
assign w38666 = ~w38664 & ~w38665;
assign w38667 = pi2004 & ~w38666;
assign w38668 = ~pi2004 & w38666;
assign w38669 = ~w38667 & ~w38668;
assign w38670 = ~pi6768 & pi9040;
assign w38671 = ~pi6750 & ~pi9040;
assign w38672 = ~w38670 & ~w38671;
assign w38673 = pi1989 & ~w38672;
assign w38674 = ~pi1989 & w38672;
assign w38675 = ~w38673 & ~w38674;
assign w38676 = w38669 & ~w38675;
assign w38677 = ~pi6760 & pi9040;
assign w38678 = ~pi6728 & ~pi9040;
assign w38679 = ~w38677 & ~w38678;
assign w38680 = pi1974 & ~w38679;
assign w38681 = ~pi1974 & w38679;
assign w38682 = ~w38680 & ~w38681;
assign w38683 = w38676 & ~w38682;
assign w38684 = ~pi6743 & pi9040;
assign w38685 = ~pi6768 & ~pi9040;
assign w38686 = ~w38684 & ~w38685;
assign w38687 = pi1997 & ~w38686;
assign w38688 = ~pi1997 & w38686;
assign w38689 = ~w38687 & ~w38688;
assign w38690 = w38669 & ~w38689;
assign w38691 = w38675 & w38682;
assign w38692 = w38690 & w38691;
assign w38693 = ~w38683 & ~w38692;
assign w38694 = ~pi6728 & pi9040;
assign w38695 = ~pi6749 & ~pi9040;
assign w38696 = ~w38694 & ~w38695;
assign w38697 = pi2000 & ~w38696;
assign w38698 = ~pi2000 & w38696;
assign w38699 = ~w38697 & ~w38698;
assign w38700 = ~w38682 & w38689;
assign w38701 = w38675 & ~w38700;
assign w38702 = ~w38675 & w38689;
assign w38703 = ~w38682 & w38702;
assign w38704 = ~w38701 & ~w38703;
assign w38705 = ~w38682 & ~w38689;
assign w38706 = w38669 & w38705;
assign w38707 = ~w38699 & ~w38706;
assign w38708 = ~w38704 & w38707;
assign w38709 = w38693 & ~w38708;
assign w38710 = ~w38663 & ~w38709;
assign w38711 = w38675 & w38689;
assign w38712 = w38663 & w38682;
assign w38713 = w38711 & w38712;
assign w38714 = w38682 & ~w38689;
assign w38715 = ~w38675 & w38714;
assign w38716 = ~w38669 & w38715;
assign w38717 = w38663 & ~w38716;
assign w38718 = w38675 & w38705;
assign w38719 = ~w38715 & ~w38718;
assign w38720 = w38717 & ~w38719;
assign w38721 = ~w38675 & ~w38690;
assign w38722 = ~w38663 & ~w38700;
assign w38723 = ~w38683 & ~w38722;
assign w38724 = w38721 & ~w38723;
assign w38725 = ~w38669 & w38675;
assign w38726 = ~w38722 & w38725;
assign w38727 = w38699 & ~w38713;
assign w38728 = ~w38726 & w38727;
assign w38729 = ~w38724 & w38728;
assign w38730 = ~w38720 & w38729;
assign w38731 = w38669 & w38711;
assign w38732 = w38711 & w66259;
assign w38733 = ~w38692 & ~w38699;
assign w38734 = ~w38732 & w38733;
assign w38735 = w38683 & ~w38689;
assign w38736 = w38663 & ~w38700;
assign w38737 = w38721 & w38736;
assign w38738 = ~w38735 & ~w38737;
assign w38739 = w38734 & w38738;
assign w38740 = ~w38730 & ~w38739;
assign w38741 = ~w38710 & ~w38740;
assign w38742 = ~pi2022 & w38741;
assign w38743 = pi2022 & ~w38741;
assign w38744 = ~w38742 & ~w38743;
assign w38745 = w38491 & w38605;
assign w38746 = w38427 & ~w38612;
assign w38747 = (~w38459 & ~w38484) | (~w38459 & w63955) | (~w38484 & w63955);
assign w38748 = ~w38475 & w38746;
assign w38749 = ~w38448 & w38613;
assign w38750 = w38604 & ~w38749;
assign w38751 = ~w38748 & ~w38750;
assign w38752 = ~w38504 & ~w38751;
assign w38753 = w38459 & ~w38752;
assign w38754 = ~w38478 & ~w38504;
assign w38755 = ~w38427 & ~w38754;
assign w38756 = ~w38615 & ~w38745;
assign w38757 = ~w38755 & w38756;
assign w38758 = ~w38747 & w38757;
assign w38759 = ~w38753 & w38758;
assign w38760 = pi2024 & ~w38759;
assign w38761 = ~pi2024 & w38759;
assign w38762 = ~w38760 & ~w38761;
assign w38763 = w38000 & w38023;
assign w38764 = w38042 & w38763;
assign w38765 = w38024 & w38048;
assign w38766 = ~w38062 & ~w38765;
assign w38767 = w38012 & w38023;
assign w38768 = ~w38055 & w38767;
assign w38769 = w38031 & w38066;
assign w38770 = ~w37994 & w38769;
assign w38771 = w38019 & w38024;
assign w38772 = w38069 & ~w38771;
assign w38773 = w38013 & w38031;
assign w38774 = ~w37994 & ~w38773;
assign w38775 = ~w38772 & ~w38774;
assign w38776 = ~w38027 & ~w38053;
assign w38777 = w38766 & ~w38768;
assign w38778 = ~w38770 & w38777;
assign w38779 = w38776 & w38778;
assign w38780 = ~w38775 & w38779;
assign w38781 = ~w38006 & w38028;
assign w38782 = w38000 & ~w38050;
assign w38783 = ~w38023 & w38782;
assign w38784 = (w37994 & ~w38031) | (w37994 & w66260) | (~w38031 & w66260);
assign w38785 = ~w38781 & w38784;
assign w38786 = ~w38783 & w38785;
assign w38787 = w38033 & w38066;
assign w38788 = ~w37994 & ~w38020;
assign w38789 = ~w38787 & w38788;
assign w38790 = ~w38786 & ~w38789;
assign w38791 = w38038 & w38062;
assign w38792 = ~w38790 & w38791;
assign w38793 = (~w38764 & w38780) | (~w38764 & w66261) | (w38780 & w66261);
assign w38794 = pi2031 & w38793;
assign w38795 = ~pi2031 & ~w38793;
assign w38796 = ~w38794 & ~w38795;
assign w38797 = w37994 & ~w38013;
assign w38798 = ~w38055 & ~w38797;
assign w38799 = ~w38027 & w66262;
assign w38800 = ~w38798 & w38799;
assign w38801 = ~w38043 & w38782;
assign w38802 = (~w37994 & ~w38782) | (~w37994 & w66263) | (~w38782 & w66263);
assign w38803 = w38066 & w38802;
assign w38804 = w38766 & ~w38769;
assign w38805 = ~w38800 & w38804;
assign w38806 = ~w38803 & w38805;
assign w38807 = ~w38027 & ~w38055;
assign w38808 = ~w38801 & w38807;
assign w38809 = w37994 & ~w38808;
assign w38810 = ~w38036 & w38802;
assign w38811 = ~w38809 & ~w38810;
assign w38812 = ~w38053 & ~w38781;
assign w38813 = w38068 & w38812;
assign w38814 = ~w38811 & w38813;
assign w38815 = ~w37994 & w38030;
assign w38816 = w38032 & w38055;
assign w38817 = ~w38022 & ~w38816;
assign w38818 = ~w38815 & w38817;
assign w38819 = (w38818 & w38814) | (w38818 & w66264) | (w38814 & w66264);
assign w38820 = ~pi2044 & ~w38819;
assign w38821 = pi2044 & w38819;
assign w38822 = ~w38820 & ~w38821;
assign w38823 = (w38321 & w38139) | (w38321 & w66265) | (w38139 & w66265);
assign w38824 = w38147 & ~w38823;
assign w38825 = w38090 & ~w38152;
assign w38826 = w38132 & ~w38825;
assign w38827 = ~w38147 & ~w38826;
assign w38828 = ~w38319 & w38827;
assign w38829 = w38117 & ~w38828;
assign w38830 = ~w38147 & ~w38316;
assign w38831 = ~w38105 & w38321;
assign w38832 = ~w38830 & w38831;
assign w38833 = ~w38829 & ~w38832;
assign w38834 = ~w38824 & ~w38833;
assign w38835 = ~pi2051 & w38834;
assign w38836 = pi2051 & ~w38834;
assign w38837 = ~w38835 & ~w38836;
assign w38838 = w38544 & ~w38594;
assign w38839 = w38535 & ~w38578;
assign w38840 = ~w38575 & ~w38839;
assign w38841 = ~w38557 & ~w38840;
assign w38842 = ~w38528 & ~w38841;
assign w38843 = w38528 & w38839;
assign w38844 = ~w38581 & ~w38586;
assign w38845 = w38559 & ~w38844;
assign w38846 = ~w38572 & ~w38845;
assign w38847 = ~w38843 & w38846;
assign w38848 = ~w38842 & w38847;
assign w38849 = ~w38544 & w38582;
assign w38850 = w38582 & w66266;
assign w38851 = ~w38545 & ~w38591;
assign w38852 = ~w38849 & ~w38851;
assign w38853 = w38541 & w38577;
assign w38854 = w38572 & ~w38853;
assign w38855 = w38553 & w38560;
assign w38856 = w38854 & ~w38855;
assign w38857 = ~w38850 & w38856;
assign w38858 = ~w38852 & w38857;
assign w38859 = (~w38838 & w38848) | (~w38838 & w66267) | (w38848 & w66267);
assign w38860 = ~pi2047 & w38859;
assign w38861 = pi2047 & ~w38859;
assign w38862 = ~w38860 & ~w38861;
assign w38863 = ~w38191 & w38645;
assign w38864 = w38215 & w38229;
assign w38865 = ~w38863 & w38864;
assign w38866 = w38279 & w38865;
assign w38867 = w38197 & w38218;
assign w38868 = ~w38191 & ~w38235;
assign w38869 = w38208 & ~w38868;
assign w38870 = ~w38262 & w38869;
assign w38871 = (~w38229 & ~w38236) | (~w38229 & w66268) | (~w38236 & w66268);
assign w38872 = ~w38867 & w38871;
assign w38873 = ~w38870 & w38872;
assign w38874 = ~w38216 & w38873;
assign w38875 = ~w38866 & ~w38874;
assign w38876 = ~w38256 & ~w38875;
assign w38877 = ~pi2046 & w38876;
assign w38878 = pi2046 & ~w38876;
assign w38879 = ~w38877 & ~w38878;
assign w38880 = ~w38375 & ~w38384;
assign w38881 = w38396 & ~w38880;
assign w38882 = w38380 & w38386;
assign w38883 = ~w38385 & ~w38882;
assign w38884 = w38363 & ~w38883;
assign w38885 = ~w38356 & ~w38378;
assign w38886 = w38370 & ~w38881;
assign w38887 = ~w38884 & w38886;
assign w38888 = ~w38885 & w38887;
assign w38889 = ~w38356 & ~w38881;
assign w38890 = w38363 & ~w38889;
assign w38891 = ~w38336 & w38355;
assign w38892 = w38403 & w38891;
assign w38893 = ~w38370 & ~w38892;
assign w38894 = ~w38890 & w38893;
assign w38895 = ~w38888 & ~w38894;
assign w38896 = ~w38370 & ~w38881;
assign w38897 = w38384 & w38896;
assign w38898 = ~w38349 & ~w38370;
assign w38899 = w38343 & w38898;
assign w38900 = ~w38387 & ~w38899;
assign w38901 = w38398 & w38900;
assign w38902 = ~w38383 & w38901;
assign w38903 = ~w38897 & w38902;
assign w38904 = ~w38363 & ~w38903;
assign w38905 = ~w38895 & ~w38904;
assign w38906 = ~pi2020 & w38905;
assign w38907 = pi2020 & ~w38905;
assign w38908 = ~w38906 & ~w38907;
assign w38909 = w38105 & ~w38159;
assign w38910 = w38092 & w38118;
assign w38911 = w38138 & ~w38910;
assign w38912 = ~w38909 & ~w38911;
assign w38913 = ~w38092 & ~w38131;
assign w38914 = w38119 & w38913;
assign w38915 = ~w38090 & ~w38099;
assign w38916 = ~w38132 & w38915;
assign w38917 = ~w38105 & ~w38914;
assign w38918 = ~w38916 & w38917;
assign w38919 = ~w38161 & ~w38301;
assign w38920 = w38105 & ~w38115;
assign w38921 = w38919 & w38920;
assign w38922 = w38147 & ~w38921;
assign w38923 = ~w38918 & w38922;
assign w38924 = ~w38099 & ~w38105;
assign w38925 = w38084 & ~w38924;
assign w38926 = w38919 & w38925;
assign w38927 = ~w38120 & ~w38129;
assign w38928 = ~w38926 & w38927;
assign w38929 = ~w38147 & ~w38928;
assign w38930 = ~w38912 & ~w38923;
assign w38931 = ~w38929 & w38930;
assign w38932 = pi2041 & w38931;
assign w38933 = ~pi2041 & ~w38931;
assign w38934 = ~w38932 & ~w38933;
assign w38935 = ~pi6747 & pi9040;
assign w38936 = ~pi6859 & ~pi9040;
assign w38937 = ~w38935 & ~w38936;
assign w38938 = pi2000 & ~w38937;
assign w38939 = ~pi2000 & w38937;
assign w38940 = ~w38938 & ~w38939;
assign w38941 = ~pi6849 & pi9040;
assign w38942 = ~pi6771 & ~pi9040;
assign w38943 = ~w38941 & ~w38942;
assign w38944 = pi2011 & ~w38943;
assign w38945 = ~pi2011 & w38943;
assign w38946 = ~w38944 & ~w38945;
assign w38947 = ~w38940 & w38946;
assign w38948 = ~pi6748 & pi9040;
assign w38949 = ~pi6751 & ~pi9040;
assign w38950 = ~w38948 & ~w38949;
assign w38951 = pi1993 & ~w38950;
assign w38952 = ~pi1993 & w38950;
assign w38953 = ~w38951 & ~w38952;
assign w38954 = w38947 & w38953;
assign w38955 = ~pi6755 & pi9040;
assign w38956 = ~pi6748 & ~pi9040;
assign w38957 = ~w38955 & ~w38956;
assign w38958 = pi1997 & ~w38957;
assign w38959 = ~pi1997 & w38957;
assign w38960 = ~w38958 & ~w38959;
assign w38961 = ~w38953 & ~w38960;
assign w38962 = w38953 & w38960;
assign w38963 = ~w38961 & ~w38962;
assign w38964 = ~w38954 & w38963;
assign w38965 = w38940 & ~w38946;
assign w38966 = ~w38947 & ~w38965;
assign w38967 = ~pi6772 & pi9040;
assign w38968 = ~pi6723 & ~pi9040;
assign w38969 = ~w38967 & ~w38968;
assign w38970 = pi1978 & ~w38969;
assign w38971 = ~pi1978 & w38969;
assign w38972 = ~w38970 & ~w38971;
assign w38973 = ~w38940 & w38972;
assign w38974 = ~w38966 & ~w38973;
assign w38975 = w38964 & ~w38974;
assign w38976 = w38947 & w38975;
assign w38977 = ~pi6756 & pi9040;
assign w38978 = ~pi6755 & ~pi9040;
assign w38979 = ~w38977 & ~w38978;
assign w38980 = pi1990 & ~w38979;
assign w38981 = ~pi1990 & w38979;
assign w38982 = ~w38980 & ~w38981;
assign w38983 = w38961 & w38966;
assign w38984 = ~w38983 & w63956;
assign w38985 = w38966 & ~w38972;
assign w38986 = w38940 & w38953;
assign w38987 = ~w38960 & w38986;
assign w38988 = ~w38985 & w38987;
assign w38989 = ~w38946 & w38960;
assign w38990 = w38940 & w38989;
assign w38991 = ~w38954 & ~w38990;
assign w38992 = ~w38983 & w38991;
assign w38993 = ~w38972 & ~w38992;
assign w38994 = ~w38984 & ~w38988;
assign w38995 = ~w38993 & w38994;
assign w38996 = w38964 & ~w38985;
assign w38997 = w38982 & ~w38996;
assign w38998 = w38995 & w38997;
assign w38999 = ~w38946 & w38953;
assign w39000 = ~w38965 & ~w38999;
assign w39001 = ~w38986 & ~w39000;
assign w39002 = (~w38947 & w39000) | (~w38947 & w63957) | (w39000 & w63957);
assign w39003 = w38991 & ~w39002;
assign w39004 = ~w38972 & ~w38986;
assign w39005 = ~w38940 & ~w38946;
assign w39006 = w38960 & w39005;
assign w39007 = w39004 & ~w39006;
assign w39008 = (~w39007 & w39003) | (~w39007 & w66269) | (w39003 & w66269);
assign w39009 = ~w38940 & ~w38960;
assign w39010 = ~w38989 & ~w39009;
assign w39011 = ~w38963 & w39010;
assign w39012 = w39008 & w39011;
assign w39013 = (~w38976 & w38995) | (~w38976 & w66270) | (w38995 & w66270);
assign w39014 = ~w38998 & ~w39012;
assign w39015 = (pi2034 & ~w39014) | (pi2034 & w66271) | (~w39014 & w66271);
assign w39016 = w39014 & w66272;
assign w39017 = ~w39015 & ~w39016;
assign w39018 = ~w38946 & ~w38972;
assign w39019 = w38962 & w39018;
assign w39020 = w39004 & w39010;
assign w39021 = (~w38960 & w38983) | (~w38960 & w66273) | (w38983 & w66273);
assign w39022 = w38986 & ~w38989;
assign w39023 = ~w38953 & w38989;
assign w39024 = ~w39022 & ~w39023;
assign w39025 = w38972 & ~w39024;
assign w39026 = ~w39020 & ~w39025;
assign w39027 = (~w38982 & ~w39026) | (~w38982 & w66274) | (~w39026 & w66274);
assign w39028 = w38962 & ~w39022;
assign w39029 = ~w39008 & ~w39028;
assign w39030 = w38982 & ~w39029;
assign w39031 = w38960 & ~w38966;
assign w39032 = w38946 & ~w38960;
assign w39033 = w38940 & w39032;
assign w39034 = ~w39031 & ~w39033;
assign w39035 = (w38972 & w39031) | (w38972 & w66275) | (w39031 & w66275);
assign w39036 = w38987 & w39035;
assign w39037 = ~w39019 & ~w39036;
assign w39038 = ~w39027 & w39037;
assign w39039 = ~w39030 & w39038;
assign w39040 = pi2048 & ~w39039;
assign w39041 = ~pi2048 & w39039;
assign w39042 = ~w39040 & ~w39041;
assign w39043 = ~w38669 & ~w38682;
assign w39044 = ~w38689 & w39043;
assign w39045 = (w38663 & ~w39043) | (w38663 & w66276) | (~w39043 & w66276);
assign w39046 = ~w38700 & w38725;
assign w39047 = ~w38735 & ~w39046;
assign w39048 = w39045 & ~w39047;
assign w39049 = ~w38663 & ~w38702;
assign w39050 = ~w38702 & w66277;
assign w39051 = ~w38701 & w39050;
assign w39052 = ~w38663 & ~w38675;
assign w39053 = ~w38722 & ~w39052;
assign w39054 = ~w38663 & ~w38682;
assign w39055 = ~w38669 & w38689;
assign w39056 = w39054 & w39055;
assign w39057 = w38669 & w38702;
assign w39058 = w38702 & w39281;
assign w39059 = ~w39056 & ~w39058;
assign w39060 = ~w39053 & ~w39059;
assign w39061 = ~w38714 & w39046;
assign w39062 = w38705 & w39052;
assign w39063 = ~w38676 & w38712;
assign w39064 = w38699 & ~w39062;
assign w39065 = ~w39063 & w39064;
assign w39066 = w39065 & w66278;
assign w39067 = ~w39060 & w39066;
assign w39068 = ~w38706 & ~w39053;
assign w39069 = w39045 & ~w39057;
assign w39070 = ~w39068 & ~w39069;
assign w39071 = ~w38703 & ~w38714;
assign w39072 = ~w38690 & ~w39071;
assign w39073 = ~w39070 & w39072;
assign w39074 = ~w38732 & ~w39050;
assign w39075 = ~w39051 & ~w39074;
assign w39076 = ~w38699 & w39059;
assign w39077 = ~w39075 & w39076;
assign w39078 = ~w39073 & w39077;
assign w39079 = (~w39048 & w39078) | (~w39048 & w66279) | (w39078 & w66279);
assign w39080 = pi2029 & ~w39079;
assign w39081 = ~pi2029 & w39079;
assign w39082 = ~w39080 & ~w39081;
assign w39083 = ~w38374 & ~w38380;
assign w39084 = ~w38403 & ~w39083;
assign w39085 = w38394 & ~w39084;
assign w39086 = ~w38356 & ~w38880;
assign w39087 = ~w38357 & ~w38370;
assign w39088 = ~w38381 & ~w39086;
assign w39089 = w39087 & w39088;
assign w39090 = (~w38363 & w39089) | (~w38363 & w66280) | (w39089 & w66280);
assign w39091 = ~w38379 & ~w38386;
assign w39092 = w39088 & w66281;
assign w39093 = ~w38356 & ~w38892;
assign w39094 = w38382 & ~w39093;
assign w39095 = ~w38342 & ~w38401;
assign w39096 = w39085 & ~w39095;
assign w39097 = w38363 & ~w39094;
assign w39098 = ~w39096 & w39097;
assign w39099 = ~w39092 & w39098;
assign w39100 = w38364 & w38403;
assign w39101 = w38370 & ~w38397;
assign w39102 = ~w39100 & w39101;
assign w39103 = ~w38896 & ~w39102;
assign w39104 = (~w39103 & w39099) | (~w39103 & w66282) | (w39099 & w66282);
assign w39105 = ~pi2016 & w39104;
assign w39106 = pi2016 & ~w39104;
assign w39107 = ~w39105 & ~w39106;
assign w39108 = ~w38477 & w38609;
assign w39109 = ~w38427 & w38608;
assign w39110 = ~w38427 & ~w38434;
assign w39111 = ~w39109 & ~w39110;
assign w39112 = ~w39108 & w39111;
assign w39113 = w38506 & ~w39112;
assign w39114 = ~w38459 & ~w39113;
assign w39115 = ~w38451 & ~w38607;
assign w39116 = w38459 & ~w39115;
assign w39117 = ~w38476 & ~w38504;
assign w39118 = ~w39116 & w39117;
assign w39119 = w38427 & ~w39118;
assign w39120 = ~w38459 & ~w39109;
assign w39121 = ~w38464 & w38503;
assign w39122 = ~w39120 & w39121;
assign w39123 = w38447 & w38459;
assign w39124 = ~w38496 & w39123;
assign w39125 = ~w39111 & w39124;
assign w39126 = ~w39122 & ~w39125;
assign w39127 = ~w39119 & w39126;
assign w39128 = ~w39114 & w39127;
assign w39129 = pi2030 & ~w39128;
assign w39130 = ~pi2030 & w39128;
assign w39131 = ~w39129 & ~w39130;
assign w39132 = ~w38535 & w38578;
assign w39133 = ~w38839 & ~w39132;
assign w39134 = ~w38565 & ~w38852;
assign w39135 = w39133 & ~w39134;
assign w39136 = ~w38522 & w38556;
assign w39137 = ~w38561 & ~w38853;
assign w39138 = ~w39136 & w39137;
assign w39139 = ~w38528 & ~w39133;
assign w39140 = w39138 & w39139;
assign w39141 = ~w39135 & ~w39140;
assign w39142 = w38572 & ~w39141;
assign w39143 = w38572 & ~w38576;
assign w39144 = w38554 & w38850;
assign w39145 = w38528 & ~w38551;
assign w39146 = w38544 & w39145;
assign w39147 = ~w39144 & ~w39146;
assign w39148 = ~w39143 & ~w39147;
assign w39149 = w38542 & w38577;
assign w39150 = ~w38591 & ~w39149;
assign w39151 = ~w38541 & ~w38564;
assign w39152 = (~w38572 & w39136) | (~w38572 & w66283) | (w39136 & w66283);
assign w39153 = (~w38543 & ~w39151) | (~w38543 & w66284) | (~w39151 & w66284);
assign w39154 = ~w39152 & w39153;
assign w39155 = ~w39148 & w39154;
assign w39156 = ~w39142 & w66285;
assign w39157 = (~pi2050 & w39142) | (~pi2050 & w66286) | (w39142 & w66286);
assign w39158 = ~w39156 & ~w39157;
assign w39159 = w38033 & ~w38797;
assign w39160 = (w37994 & w38808) | (w37994 & w66287) | (w38808 & w66287);
assign w39161 = ~w39159 & ~w39160;
assign w39162 = ~w38062 & ~w39161;
assign w39163 = w38050 & ~w38807;
assign w39164 = ~w38763 & ~w38787;
assign w39165 = ~w38770 & w39164;
assign w39166 = ~w39163 & w39165;
assign w39167 = w38062 & ~w39166;
assign w39168 = ~w38013 & w38026;
assign w39169 = ~w38066 & w39168;
assign w39170 = ~w38052 & w38774;
assign w39171 = ~w39169 & w39170;
assign w39172 = w37994 & ~w38067;
assign w39173 = ~w38037 & w39172;
assign w39174 = ~w39171 & ~w39173;
assign w39175 = ~w39167 & ~w39174;
assign w39176 = ~w39162 & w39175;
assign w39177 = ~pi2063 & w39176;
assign w39178 = pi2063 & ~w39176;
assign w39179 = ~w39177 & ~w39178;
assign w39180 = ~w38963 & w38974;
assign w39181 = ~w38975 & ~w39180;
assign w39182 = ~w38982 & ~w39181;
assign w39183 = w38953 & w39032;
assign w39184 = w38991 & ~w39032;
assign w39185 = (w38982 & ~w38991) | (w38982 & w66288) | (~w38991 & w66288);
assign w39186 = w38961 & w39005;
assign w39187 = ~w39183 & ~w39186;
assign w39188 = ~w39185 & w39187;
assign w39189 = w38972 & ~w39188;
assign w39190 = ~w38972 & ~w39005;
assign w39191 = w39184 & w39190;
assign w39192 = w38962 & w39005;
assign w39193 = ~w39191 & ~w39192;
assign w39194 = w38982 & ~w39193;
assign w39195 = ~w39182 & ~w39189;
assign w39196 = ~w39194 & w39195;
assign w39197 = ~pi2042 & w39196;
assign w39198 = pi2042 & ~w39196;
assign w39199 = ~w39197 & ~w39198;
assign w39200 = w38541 & ~w39133;
assign w39201 = w38564 & w63958;
assign w39202 = ~w38578 & w66289;
assign w39203 = ~w39146 & w39150;
assign w39204 = ~w39202 & w39203;
assign w39205 = ~w39201 & w39204;
assign w39206 = w38589 & ~w39132;
assign w39207 = w39204 & w63959;
assign w39208 = (w38572 & w39207) | (w38572 & w66290) | (w39207 & w66290);
assign w39209 = w38541 & w38840;
assign w39210 = ~w38561 & w38854;
assign w39211 = (~w39210 & ~w39205) | (~w39210 & w66291) | (~w39205 & w66291);
assign w39212 = ~w39208 & ~w39211;
assign w39213 = ~pi2033 & w39212;
assign w39214 = pi2033 & ~w39212;
assign w39215 = ~w39213 & ~w39214;
assign w39216 = ~w39000 & w39004;
assign w39217 = w38960 & ~w39018;
assign w39218 = w38966 & ~w39217;
assign w39219 = ~w39031 & ~w39218;
assign w39220 = ~w38953 & w39219;
assign w39221 = w38954 & w38960;
assign w39222 = ~w39216 & ~w39221;
assign w39223 = (w38982 & w39220) | (w38982 & w66292) | (w39220 & w66292);
assign w39224 = ~w38982 & ~w39001;
assign w39225 = w39034 & w39224;
assign w39226 = (~w38972 & w39225) | (~w38972 & w66293) | (w39225 & w66293);
assign w39227 = ~w39035 & ~w39186;
assign w39228 = ~w38982 & ~w39227;
assign w39229 = w38972 & w38999;
assign w39230 = ~w39219 & w39229;
assign w39231 = ~w39223 & ~w39230;
assign w39232 = ~w39226 & ~w39228;
assign w39233 = w39231 & w39232;
assign w39234 = pi2026 & w39233;
assign w39235 = ~pi2026 & ~w39233;
assign w39236 = ~w39234 & ~w39235;
assign w39237 = ~w38715 & ~w39061;
assign w39238 = w38693 & w39237;
assign w39239 = ~w39049 & ~w39054;
assign w39240 = (w38691 & ~w39237) | (w38691 & w66294) | (~w39237 & w66294);
assign w39241 = ~w39057 & w39239;
assign w39242 = w39237 & w39241;
assign w39243 = ~w39240 & w39242;
assign w39244 = (~w38699 & w39238) | (~w38699 & w66295) | (w39238 & w66295);
assign w39245 = ~w39243 & w39244;
assign w39246 = w38699 & ~w38716;
assign w39247 = w39059 & w39246;
assign w39248 = ~w39070 & w39247;
assign w39249 = ~w39240 & w39248;
assign w39250 = ~w39245 & ~w39249;
assign w39251 = pi2035 & w39250;
assign w39252 = ~pi2035 & ~w39250;
assign w39253 = ~w39251 & ~w39252;
assign w39254 = ~w38356 & ~w38883;
assign w39255 = ~w39100 & ~w39254;
assign w39256 = ~w38370 & ~w39255;
assign w39257 = ~w38395 & ~w38403;
assign w39258 = (~w38891 & w38357) | (~w38891 & w66296) | (w38357 & w66296);
assign w39259 = w39257 & ~w39258;
assign w39260 = ~w38381 & ~w39259;
assign w39261 = w39085 & ~w39260;
assign w39262 = ~w38356 & ~w38375;
assign w39263 = w38370 & ~w38403;
assign w39264 = ~w39262 & w39263;
assign w39265 = ~w38357 & w38363;
assign w39266 = ~w38892 & ~w38899;
assign w39267 = w39265 & w39266;
assign w39268 = ~w39264 & w39267;
assign w39269 = ~w38380 & ~w39087;
assign w39270 = ~w39257 & w39269;
assign w39271 = ~w38363 & ~w39259;
assign w39272 = ~w39270 & w39271;
assign w39273 = ~w39268 & ~w39272;
assign w39274 = ~w39256 & ~w39261;
assign w39275 = ~w39273 & w39274;
assign w39276 = pi2025 & ~w39275;
assign w39277 = ~pi2025 & w39275;
assign w39278 = ~w39276 & ~w39277;
assign w39279 = w38717 & ~w38731;
assign w39280 = w39239 & ~w39279;
assign w39281 = w38669 & w38682;
assign w39282 = ~w39043 & ~w39281;
assign w39283 = ~w38675 & ~w38712;
assign w39284 = ~w39282 & w39283;
assign w39285 = ~w38713 & ~w39044;
assign w39286 = ~w39284 & w39285;
assign w39287 = w38734 & w39286;
assign w39288 = ~w38718 & ~w39055;
assign w39289 = w39049 & ~w39288;
assign w39290 = w38663 & ~w39071;
assign w39291 = w38699 & ~w38735;
assign w39292 = ~w39289 & w39291;
assign w39293 = ~w39290 & w39292;
assign w39294 = ~w39287 & ~w39293;
assign w39295 = ~w39280 & ~w39294;
assign w39296 = pi2057 & w39295;
assign w39297 = ~pi2057 & ~w39295;
assign w39298 = ~w39296 & ~w39297;
assign w39299 = ~pi6960 & pi9040;
assign w39300 = ~pi6975 & ~pi9040;
assign w39301 = ~w39299 & ~w39300;
assign w39302 = pi2043 & ~w39301;
assign w39303 = ~pi2043 & w39301;
assign w39304 = ~w39302 & ~w39303;
assign w39305 = ~pi6956 & pi9040;
assign w39306 = ~pi6946 & ~pi9040;
assign w39307 = ~w39305 & ~w39306;
assign w39308 = pi2065 & ~w39307;
assign w39309 = ~pi2065 & w39307;
assign w39310 = ~w39308 & ~w39309;
assign w39311 = ~w39304 & ~w39310;
assign w39312 = ~pi6979 & pi9040;
assign w39313 = ~pi6958 & ~pi9040;
assign w39314 = ~w39312 & ~w39313;
assign w39315 = pi2061 & ~w39314;
assign w39316 = ~pi2061 & w39314;
assign w39317 = ~w39315 & ~w39316;
assign w39318 = ~pi6958 & pi9040;
assign w39319 = ~pi7002 & ~pi9040;
assign w39320 = ~w39318 & ~w39319;
assign w39321 = pi2037 & ~w39320;
assign w39322 = ~pi2037 & w39320;
assign w39323 = ~w39321 & ~w39322;
assign w39324 = ~w39317 & w39323;
assign w39325 = w39317 & ~w39323;
assign w39326 = ~w39324 & ~w39325;
assign w39327 = w39311 & ~w39326;
assign w39328 = w39304 & ~w39323;
assign w39329 = w39304 & w39323;
assign w39330 = ~w39310 & w39317;
assign w39331 = w39329 & w39330;
assign w39332 = ~w39328 & ~w39331;
assign w39333 = ~pi7002 & pi9040;
assign w39334 = ~pi6980 & ~pi9040;
assign w39335 = ~w39333 & ~w39334;
assign w39336 = pi2076 & ~w39335;
assign w39337 = ~pi2076 & w39335;
assign w39338 = ~w39336 & ~w39337;
assign w39339 = ~w39317 & ~w39338;
assign w39340 = ~w39331 & ~w39339;
assign w39341 = ~w39332 & ~w39340;
assign w39342 = ~w39327 & ~w39341;
assign w39343 = w39310 & ~w39317;
assign w39344 = ~w39323 & w39343;
assign w39345 = w39343 & w39353;
assign w39346 = w39310 & w39323;
assign w39347 = ~w39304 & w39346;
assign w39348 = w39338 & ~w39347;
assign w39349 = w39310 & w39317;
assign w39350 = w39328 & w39349;
assign w39351 = ~w39345 & ~w39350;
assign w39352 = w39348 & w39351;
assign w39353 = ~w39304 & ~w39323;
assign w39354 = ~w39343 & w39353;
assign w39355 = w39317 & w39329;
assign w39356 = ~w39338 & ~w39354;
assign w39357 = ~w39355 & w39356;
assign w39358 = ~w39352 & ~w39357;
assign w39359 = w39342 & ~w39358;
assign w39360 = ~pi7084 & pi9040;
assign w39361 = ~pi6960 & ~pi9040;
assign w39362 = ~w39360 & ~w39361;
assign w39363 = pi2074 & ~w39362;
assign w39364 = ~pi2074 & w39362;
assign w39365 = ~w39363 & ~w39364;
assign w39366 = ~w39359 & w39365;
assign w39367 = ~w39310 & w39328;
assign w39368 = w39328 & w66297;
assign w39369 = w39338 & w39343;
assign w39370 = w39317 & ~w39365;
assign w39371 = w39311 & w39370;
assign w39372 = ~w39369 & ~w39371;
assign w39373 = w39323 & ~w39372;
assign w39374 = w39304 & w39346;
assign w39375 = (w39338 & ~w39346) | (w39338 & w39598) | (~w39346 & w39598);
assign w39376 = ~w39330 & w39354;
assign w39377 = ~w39367 & w39375;
assign w39378 = ~w39376 & w39377;
assign w39379 = ~w39311 & ~w39328;
assign w39380 = ~w39317 & w39379;
assign w39381 = ~w39338 & ~w39350;
assign w39382 = ~w39380 & w39381;
assign w39383 = ~w39365 & ~w39382;
assign w39384 = ~w39378 & w39383;
assign w39385 = ~w39368 & ~w39373;
assign w39386 = ~w39384 & w39385;
assign w39387 = ~w39366 & w39386;
assign w39388 = pi2153 & w39387;
assign w39389 = ~pi2153 & ~w39387;
assign w39390 = ~w39388 & ~w39389;
assign w39391 = ~pi7005 & pi9040;
assign w39392 = ~pi6973 & ~pi9040;
assign w39393 = ~w39391 & ~w39392;
assign w39394 = pi2055 & ~w39393;
assign w39395 = ~pi2055 & w39393;
assign w39396 = ~w39394 & ~w39395;
assign w39397 = ~pi7004 & pi9040;
assign w39398 = ~pi6993 & ~pi9040;
assign w39399 = ~w39397 & ~w39398;
assign w39400 = pi2075 & ~w39399;
assign w39401 = ~pi2075 & w39399;
assign w39402 = ~w39400 & ~w39401;
assign w39403 = w39396 & w39402;
assign w39404 = ~w39396 & ~w39402;
assign w39405 = ~w39403 & ~w39404;
assign w39406 = ~pi6980 & pi9040;
assign w39407 = ~pi7009 & ~pi9040;
assign w39408 = ~w39406 & ~w39407;
assign w39409 = pi2049 & ~w39408;
assign w39410 = ~pi2049 & w39408;
assign w39411 = ~w39409 & ~w39410;
assign w39412 = ~pi7083 & pi9040;
assign w39413 = ~pi6982 & ~pi9040;
assign w39414 = ~w39412 & ~w39413;
assign w39415 = pi2060 & ~w39414;
assign w39416 = ~pi2060 & w39414;
assign w39417 = ~w39415 & ~w39416;
assign w39418 = ~w39411 & w39417;
assign w39419 = w39405 & w39418;
assign w39420 = w39402 & w39417;
assign w39421 = w39411 & ~w39420;
assign w39422 = ~w39396 & w39411;
assign w39423 = w39417 & w39422;
assign w39424 = ~w39402 & w39418;
assign w39425 = ~w39423 & ~w39424;
assign w39426 = ~w39421 & ~w39425;
assign w39427 = w39396 & ~w39411;
assign w39428 = w39402 & w39427;
assign w39429 = w39427 & w40471;
assign w39430 = (~w39429 & w39425) | (~w39429 & w66298) | (w39425 & w66298);
assign w39431 = w39402 & w39422;
assign w39432 = ~w39411 & ~w39417;
assign w39433 = ~w39405 & w39432;
assign w39434 = ~w39431 & ~w39433;
assign w39435 = (~w39419 & ~w39430) | (~w39419 & w63416) | (~w39430 & w63416);
assign w39436 = ~pi6984 & pi9040;
assign w39437 = ~pi7084 & ~pi9040;
assign w39438 = ~w39436 & ~w39437;
assign w39439 = pi2066 & ~w39438;
assign w39440 = ~pi2066 & w39438;
assign w39441 = ~w39439 & ~w39440;
assign w39442 = (~w63416 & w66299) | (~w63416 & w66300) | (w66299 & w66300);
assign w39443 = ~w39402 & ~w39417;
assign w39444 = w39402 & w39418;
assign w39445 = w39396 & ~w39441;
assign w39446 = (w39445 & w39444) | (w39445 & w66301) | (w39444 & w66301);
assign w39447 = w39411 & w39446;
assign w39448 = w39441 & ~w39443;
assign w39449 = w39396 & ~w39402;
assign w39450 = ~w39411 & w39441;
assign w39451 = w39449 & ~w39450;
assign w39452 = ~w39448 & w39451;
assign w39453 = w39411 & ~w39417;
assign w39454 = ~w39449 & ~w39453;
assign w39455 = ~w39431 & w39454;
assign w39456 = w39441 & ~w39452;
assign w39457 = ~w39422 & ~w39427;
assign w39458 = (~w39432 & w39457) | (~w39432 & w63960) | (w39457 & w63960);
assign w39459 = (~w39441 & ~w39405) | (~w39441 & w63961) | (~w39405 & w63961);
assign w39460 = ~w39458 & w39459;
assign w39461 = w39404 & ~w39411;
assign w39462 = w39396 & w39453;
assign w39463 = ~w39423 & ~w39461;
assign w39464 = (~w39441 & ~w39463) | (~w39441 & w63962) | (~w39463 & w63962);
assign w39465 = ~w39460 & ~w39464;
assign w39466 = ~w39421 & ~w39465;
assign w39467 = ~pi6982 & pi9040;
assign w39468 = ~pi6978 & ~pi9040;
assign w39469 = ~w39467 & ~w39468;
assign w39470 = pi2077 & ~w39469;
assign w39471 = ~pi2077 & w39469;
assign w39472 = ~w39470 & ~w39471;
assign w39473 = (w39472 & ~w39456) | (w39472 & w66302) | (~w39456 & w66302);
assign w39474 = ~w39466 & w39473;
assign w39475 = ~w39418 & ~w39441;
assign w39476 = (~w39441 & w39444) | (~w39441 & w63417) | (w39444 & w63417);
assign w39477 = ~w39428 & ~w39462;
assign w39478 = ~w39476 & w39477;
assign w39479 = (~w39452 & ~w39478) | (~w39452 & w63963) | (~w39478 & w63963);
assign w39480 = (w39450 & w39458) | (w39450 & w66303) | (w39458 & w66303);
assign w39481 = w39403 & w39411;
assign w39482 = w39417 & w39481;
assign w39483 = ~w39472 & ~w39482;
assign w39484 = ~w39480 & w39483;
assign w39485 = w39479 & w39484;
assign w39486 = ~w39474 & ~w39485;
assign w39487 = ~w39442 & ~w39447;
assign w39488 = ~w39486 & w66304;
assign w39489 = (~pi2152 & w39486) | (~pi2152 & w66305) | (w39486 & w66305);
assign w39490 = ~w39488 & ~w39489;
assign w39491 = ~pi6945 & pi9040;
assign w39492 = ~pi7081 & ~pi9040;
assign w39493 = ~w39491 & ~w39492;
assign w39494 = pi2032 & ~w39493;
assign w39495 = ~pi2032 & w39493;
assign w39496 = ~w39494 & ~w39495;
assign w39497 = ~pi7012 & pi9040;
assign w39498 = ~pi6947 & ~pi9040;
assign w39499 = ~w39497 & ~w39498;
assign w39500 = pi2067 & ~w39499;
assign w39501 = ~pi2067 & w39499;
assign w39502 = ~w39500 & ~w39501;
assign w39503 = w39496 & w39502;
assign w39504 = ~pi7082 & pi9040;
assign w39505 = ~pi7006 & ~pi9040;
assign w39506 = ~w39504 & ~w39505;
assign w39507 = pi2071 & ~w39506;
assign w39508 = ~pi2071 & w39506;
assign w39509 = ~w39507 & ~w39508;
assign w39510 = ~w39502 & ~w39509;
assign w39511 = ~pi7008 & pi9040;
assign w39512 = ~pi6945 & ~pi9040;
assign w39513 = ~w39511 & ~w39512;
assign w39514 = pi2070 & ~w39513;
assign w39515 = ~pi2070 & w39513;
assign w39516 = ~w39514 & ~w39515;
assign w39517 = ~pi6968 & pi9040;
assign w39518 = ~pi6962 & ~pi9040;
assign w39519 = ~w39517 & ~w39518;
assign w39520 = pi2073 & ~w39519;
assign w39521 = ~pi2073 & w39519;
assign w39522 = ~w39520 & ~w39521;
assign w39523 = ~w39516 & ~w39522;
assign w39524 = ~w39510 & w39523;
assign w39525 = ~w39503 & w39524;
assign w39526 = ~pi6962 & pi9040;
assign w39527 = ~pi6990 & ~pi9040;
assign w39528 = ~w39526 & ~w39527;
assign w39529 = pi2069 & ~w39528;
assign w39530 = ~pi2069 & w39528;
assign w39531 = ~w39529 & ~w39530;
assign w39532 = ~w39496 & w39516;
assign w39533 = ~w39502 & w39522;
assign w39534 = ~w39532 & ~w39533;
assign w39535 = ~w39516 & w39522;
assign w39536 = ~w39496 & w39502;
assign w39537 = w39535 & ~w39536;
assign w39538 = w39516 & ~w39522;
assign w39539 = ~w39510 & w39538;
assign w39540 = ~w39537 & ~w39539;
assign w39541 = w39534 & ~w39540;
assign w39542 = ~w39496 & ~w39538;
assign w39543 = w39516 & w39522;
assign w39544 = w39496 & ~w39543;
assign w39545 = ~w39542 & ~w39544;
assign w39546 = ~w39509 & ~w39536;
assign w39547 = w39545 & w39546;
assign w39548 = ~w39525 & w39531;
assign w39549 = ~w39541 & w39548;
assign w39550 = ~w39547 & w39549;
assign w39551 = w39510 & ~w39545;
assign w39552 = ~w39496 & w39533;
assign w39553 = w39502 & w39509;
assign w39554 = ~w39536 & ~w39539;
assign w39555 = ~w39535 & ~w39554;
assign w39556 = w39553 & ~w39555;
assign w39557 = w39536 & w39538;
assign w39558 = ~w39531 & ~w39552;
assign w39559 = ~w39557 & w39558;
assign w39560 = ~w39551 & w39559;
assign w39561 = ~w39556 & w39560;
assign w39562 = ~w39550 & ~w39561;
assign w39563 = w39502 & ~w39522;
assign w39564 = ~w39533 & ~w39563;
assign w39565 = w39509 & ~w39564;
assign w39566 = w39532 & w39565;
assign w39567 = ~w39537 & ~w39557;
assign w39568 = ~w39509 & ~w39567;
assign w39569 = ~w39496 & w39535;
assign w39570 = (~w39509 & ~w39535) | (~w39509 & w66306) | (~w39535 & w66306);
assign w39571 = ~w39554 & w39570;
assign w39572 = ~w39568 & ~w39571;
assign w39573 = w39542 & ~w39572;
assign w39574 = ~w39566 & ~w39573;
assign w39575 = ~w39562 & w39574;
assign w39576 = pi2173 & ~w39575;
assign w39577 = ~pi2173 & w39575;
assign w39578 = ~w39576 & ~w39577;
assign w39579 = w39311 & ~w39323;
assign w39580 = w39339 & w39579;
assign w39581 = ~w39345 & ~w39355;
assign w39582 = w39338 & ~w39581;
assign w39583 = ~w39304 & w39349;
assign w39584 = ~w39368 & ~w39583;
assign w39585 = w39375 & w39584;
assign w39586 = w39365 & ~w39585;
assign w39587 = ~w39582 & ~w39586;
assign w39588 = w39304 & w39343;
assign w39589 = ~w39311 & ~w39588;
assign w39590 = w39324 & w39589;
assign w39591 = w39317 & ~w39379;
assign w39592 = ~w39338 & ~w39591;
assign w39593 = ~w39590 & w39592;
assign w39594 = ~w39587 & ~w39593;
assign w39595 = ~w39583 & ~w39588;
assign w39596 = ~w39338 & ~w39595;
assign w39597 = ~w39325 & ~w39349;
assign w39598 = ~w39304 & w39338;
assign w39599 = w39597 & w39598;
assign w39600 = ~w39596 & ~w39599;
assign w39601 = ~w39342 & ~w39600;
assign w39602 = w39330 & w39338;
assign w39603 = ~w39344 & ~w39602;
assign w39604 = w39304 & ~w39603;
assign w39605 = ~w39341 & ~w39604;
assign w39606 = w39600 & w39605;
assign w39607 = ~w39365 & ~w39606;
assign w39608 = ~w39580 & ~w39601;
assign w39609 = ~w39607 & w39608;
assign w39610 = w39609 & w66307;
assign w39611 = (~pi2169 & ~w39609) | (~pi2169 & w66308) | (~w39609 & w66308);
assign w39612 = ~w39610 & ~w39611;
assign w39613 = w39317 & w39347;
assign w39614 = w39338 & ~w39353;
assign w39615 = ~w39589 & w39614;
assign w39616 = ~w39327 & ~w39344;
assign w39617 = ~w39613 & w39616;
assign w39618 = (w39365 & ~w39617) | (w39365 & w66309) | (~w39617 & w66309);
assign w39619 = w39317 & w39346;
assign w39620 = ~w39347 & ~w39579;
assign w39621 = ~w39619 & w39620;
assign w39622 = (~w39375 & ~w39620) | (~w39375 & w66310) | (~w39620 & w66310);
assign w39623 = w39348 & w39589;
assign w39624 = ~w39622 & ~w39623;
assign w39625 = w39365 & ~w39624;
assign w39626 = w39304 & ~w39310;
assign w39627 = w39329 & w39339;
assign w39628 = ~w39365 & ~w39627;
assign w39629 = w39626 & ~w39628;
assign w39630 = w39624 & ~w39629;
assign w39631 = ~w39625 & ~w39630;
assign w39632 = ~w39601 & ~w39618;
assign w39633 = ~w39631 & w39632;
assign w39634 = pi2163 & ~w39633;
assign w39635 = ~pi2163 & w39633;
assign w39636 = ~w39634 & ~w39635;
assign w39637 = ~pi7009 & pi9040;
assign w39638 = ~pi6984 & ~pi9040;
assign w39639 = ~w39637 & ~w39638;
assign w39640 = pi2045 & ~w39639;
assign w39641 = ~pi2045 & w39639;
assign w39642 = ~w39640 & ~w39641;
assign w39643 = ~pi6966 & pi9040;
assign w39644 = ~pi7005 & ~pi9040;
assign w39645 = ~w39643 & ~w39644;
assign w39646 = pi2037 & ~w39645;
assign w39647 = ~pi2037 & w39645;
assign w39648 = ~w39646 & ~w39647;
assign w39649 = ~w39642 & ~w39648;
assign w39650 = ~pi6992 & pi9040;
assign w39651 = ~pi6988 & ~pi9040;
assign w39652 = ~w39650 & ~w39651;
assign w39653 = pi2074 & ~w39652;
assign w39654 = ~pi2074 & w39652;
assign w39655 = ~w39653 & ~w39654;
assign w39656 = ~pi6983 & pi9040;
assign w39657 = ~pi7004 & ~pi9040;
assign w39658 = ~w39656 & ~w39657;
assign w39659 = pi2049 & ~w39658;
assign w39660 = ~pi2049 & w39658;
assign w39661 = ~w39659 & ~w39660;
assign w39662 = ~w39655 & ~w39661;
assign w39663 = w39649 & w39662;
assign w39664 = ~pi6959 & pi9040;
assign w39665 = ~pi7003 & ~pi9040;
assign w39666 = ~w39664 & ~w39665;
assign w39667 = pi2055 & ~w39666;
assign w39668 = ~pi2055 & w39666;
assign w39669 = ~w39667 & ~w39668;
assign w39670 = w39642 & ~w39648;
assign w39671 = ~w39655 & w39661;
assign w39672 = w39670 & w39671;
assign w39673 = ~pi6953 & pi9040;
assign w39674 = ~pi6983 & ~pi9040;
assign w39675 = ~w39673 & ~w39674;
assign w39676 = pi2062 & ~w39675;
assign w39677 = ~pi2062 & w39675;
assign w39678 = ~w39676 & ~w39677;
assign w39679 = w39661 & ~w39678;
assign w39680 = w39648 & w39655;
assign w39681 = ~w39642 & w39655;
assign w39682 = ~w39648 & ~w39681;
assign w39683 = ~w39680 & ~w39682;
assign w39684 = w39679 & w39683;
assign w39685 = w39648 & w39661;
assign w39686 = ~w39642 & w39685;
assign w39687 = ~w39670 & ~w39686;
assign w39688 = w39655 & w39678;
assign w39689 = ~w39687 & w39688;
assign w39690 = ~w39663 & w39669;
assign w39691 = ~w39672 & w39690;
assign w39692 = ~w39684 & w39691;
assign w39693 = ~w39689 & w39692;
assign w39694 = w39642 & ~w39655;
assign w39695 = ~w39681 & ~w39694;
assign w39696 = ~w39648 & w39678;
assign w39697 = w39695 & ~w39696;
assign w39698 = w39695 & w66311;
assign w39699 = w39649 & w39655;
assign w39700 = ~w39679 & w39699;
assign w39701 = ~w39698 & ~w39700;
assign w39702 = ~w39661 & w39680;
assign w39703 = w39662 & w39670;
assign w39704 = ~w39702 & ~w39703;
assign w39705 = ~w39678 & ~w39704;
assign w39706 = ~w39669 & ~w39705;
assign w39707 = w39701 & w39706;
assign w39708 = ~w39693 & ~w39707;
assign w39709 = w39648 & ~w39678;
assign w39710 = w39695 & w39709;
assign w39711 = w39678 & ~w39703;
assign w39712 = ~w39648 & ~w39661;
assign w39713 = ~w39685 & ~w39712;
assign w39714 = w39694 & w39713;
assign w39715 = ~w39712 & ~w39714;
assign w39716 = w39711 & ~w39715;
assign w39717 = ~w39710 & ~w39716;
assign w39718 = ~w39708 & w39717;
assign w39719 = ~pi2197 & ~w39718;
assign w39720 = pi2197 & w39718;
assign w39721 = ~w39719 & ~w39720;
assign w39722 = w39496 & w39564;
assign w39723 = ~w39509 & ~w39516;
assign w39724 = w39722 & w39723;
assign w39725 = ~w39522 & w39724;
assign w39726 = w39502 & w39545;
assign w39727 = ~w39496 & ~w39509;
assign w39728 = w39509 & ~w39533;
assign w39729 = ~w39502 & w39516;
assign w39730 = ~w39535 & ~w39729;
assign w39731 = w39728 & ~w39730;
assign w39732 = (w39531 & w39564) | (w39531 & w66312) | (w39564 & w66312);
assign w39733 = ~w39731 & w39732;
assign w39734 = ~w39726 & w39733;
assign w39735 = ~w39725 & w39734;
assign w39736 = w39570 & ~w39730;
assign w39737 = ~w39496 & w39523;
assign w39738 = ~w39524 & ~w39737;
assign w39739 = ~w39536 & ~w39738;
assign w39740 = ~w39564 & w66313;
assign w39741 = ~w39552 & ~w39553;
assign w39742 = w39543 & ~w39741;
assign w39743 = ~w39531 & ~w39736;
assign w39744 = ~w39739 & ~w39740;
assign w39745 = w39744 & w66314;
assign w39746 = ~w39735 & ~w39745;
assign w39747 = ~w39502 & w39509;
assign w39748 = ~w39557 & ~w39747;
assign w39749 = (w39509 & w39552) | (w39509 & w66315) | (w39552 & w66315);
assign w39750 = w39728 & ~w39737;
assign w39751 = ~w39749 & ~w39750;
assign w39752 = ~w39748 & w39751;
assign w39753 = w39553 & w39569;
assign w39754 = ~w39752 & ~w39753;
assign w39755 = ~w39746 & w39754;
assign w39756 = pi2145 & ~w39755;
assign w39757 = ~pi2145 & w39755;
assign w39758 = ~w39756 & ~w39757;
assign w39759 = ~pi6974 & pi9040;
assign w39760 = ~pi7008 & ~pi9040;
assign w39761 = ~w39759 & ~w39760;
assign w39762 = pi2036 & ~w39761;
assign w39763 = ~pi2036 & w39761;
assign w39764 = ~w39762 & ~w39763;
assign w39765 = ~pi7068 & pi9040;
assign w39766 = ~pi6972 & ~pi9040;
assign w39767 = ~w39765 & ~w39766;
assign w39768 = pi2059 & ~w39767;
assign w39769 = ~pi2059 & w39767;
assign w39770 = ~w39768 & ~w39769;
assign w39771 = ~pi6948 & pi9040;
assign w39772 = ~pi7068 & ~pi9040;
assign w39773 = ~w39771 & ~w39772;
assign w39774 = pi2077 & ~w39773;
assign w39775 = ~pi2077 & w39773;
assign w39776 = ~w39774 & ~w39775;
assign w39777 = w39770 & ~w39776;
assign w39778 = ~pi7081 & pi9040;
assign w39779 = ~pi6952 & ~pi9040;
assign w39780 = ~w39778 & ~w39779;
assign w39781 = pi2052 & ~w39780;
assign w39782 = ~pi2052 & w39780;
assign w39783 = ~w39781 & ~w39782;
assign w39784 = w39777 & w39783;
assign w39785 = w39777 & w66316;
assign w39786 = ~pi7006 & pi9040;
assign w39787 = ~pi6948 & ~pi9040;
assign w39788 = ~w39786 & ~w39787;
assign w39789 = pi2060 & ~w39788;
assign w39790 = ~pi2060 & w39788;
assign w39791 = ~w39789 & ~w39790;
assign w39792 = w39785 & ~w39791;
assign w39793 = ~w39764 & w39791;
assign w39794 = ~w39770 & ~w39793;
assign w39795 = ~w39776 & ~w39791;
assign w39796 = w39764 & w39776;
assign w39797 = w39770 & ~w39796;
assign w39798 = ~w39795 & w39797;
assign w39799 = ~w39764 & ~w39776;
assign w39800 = ~w39796 & ~w39799;
assign w39801 = ~w39791 & ~w39800;
assign w39802 = ~w39800 & w66317;
assign w39803 = ~w39798 & ~w39802;
assign w39804 = ~w39794 & w39803;
assign w39805 = w39776 & w39791;
assign w39806 = w39764 & ~w39791;
assign w39807 = ~w39805 & ~w39806;
assign w39808 = ~pi6954 & pi9040;
assign w39809 = ~pi6986 & ~pi9040;
assign w39810 = ~w39808 & ~w39809;
assign w39811 = pi2058 & ~w39810;
assign w39812 = ~pi2058 & w39810;
assign w39813 = ~w39811 & ~w39812;
assign w39814 = ~w39770 & w39776;
assign w39815 = ~w39777 & ~w39813;
assign w39816 = ~w39814 & w39815;
assign w39817 = w39807 & w39816;
assign w39818 = ~w39804 & ~w39817;
assign w39819 = ~w39783 & ~w39818;
assign w39820 = ~w39783 & w39805;
assign w39821 = ~w39770 & w39799;
assign w39822 = w39795 & ~w39821;
assign w39823 = ~w39820 & ~w39822;
assign w39824 = w39783 & w39806;
assign w39825 = ~w39783 & ~w39814;
assign w39826 = ~w39805 & w39825;
assign w39827 = w39794 & w39800;
assign w39828 = ~w39826 & w39827;
assign w39829 = ~w39785 & ~w39824;
assign w39830 = w39823 & w39829;
assign w39831 = ~w39828 & w39830;
assign w39832 = (w39813 & ~w39830) | (w39813 & w66318) | (~w39830 & w66318);
assign w39833 = w39783 & w39791;
assign w39834 = w39764 & ~w39776;
assign w39835 = w39833 & w39834;
assign w39836 = ~w39821 & ~w39835;
assign w39837 = ~w39794 & ~w39836;
assign w39838 = w39764 & w39791;
assign w39839 = ~w39814 & ~w39838;
assign w39840 = ~w39794 & ~w39839;
assign w39841 = w39806 & w39814;
assign w39842 = w39776 & w39783;
assign w39843 = w39791 & w39842;
assign w39844 = ~w39841 & ~w39843;
assign w39845 = ~w39840 & ~w39844;
assign w39846 = ~w39837 & ~w39845;
assign w39847 = ~w39770 & ~w39791;
assign w39848 = w39842 & w39847;
assign w39849 = ~w39792 & ~w39848;
assign w39850 = (w39849 & w39846) | (w39849 & w66319) | (w39846 & w66319);
assign w39851 = ~w39832 & w39850;
assign w39852 = ~w39819 & w39851;
assign w39853 = pi2147 & ~w39852;
assign w39854 = ~pi2147 & w39852;
assign w39855 = ~w39853 & ~w39854;
assign w39856 = w39378 & ~w39597;
assign w39857 = (~w39338 & w39353) | (~w39338 & w66320) | (w39353 & w66320);
assign w39858 = w39317 & ~w39367;
assign w39859 = ~w39374 & w39858;
assign w39860 = w39857 & ~w39859;
assign w39861 = ~w39332 & w39378;
assign w39862 = w39324 & w39338;
assign w39863 = (w39621 & w66321) | (w39621 & w66322) | (w66321 & w66322);
assign w39864 = ~w39368 & w39628;
assign w39865 = ~w39861 & w39864;
assign w39866 = w39304 & w39862;
assign w39867 = w39339 & ~w39626;
assign w39868 = ~w39345 & ~w39867;
assign w39869 = ~w39329 & ~w39868;
assign w39870 = w39365 & ~w39619;
assign w39871 = ~w39866 & w39870;
assign w39872 = ~w39869 & w39871;
assign w39873 = (~w39872 & ~w39865) | (~w39872 & w66323) | (~w39865 & w66323);
assign w39874 = ~w39856 & ~w39860;
assign w39875 = ~w39873 & w39874;
assign w39876 = ~pi2150 & ~w39875;
assign w39877 = pi2150 & w39875;
assign w39878 = ~w39876 & ~w39877;
assign w39879 = w39655 & w39661;
assign w39880 = w39670 & w39879;
assign w39881 = ~w39669 & ~w39880;
assign w39882 = ~w39648 & ~w39678;
assign w39883 = ~w39678 & ~w39694;
assign w39884 = ~w39882 & ~w39883;
assign w39885 = w39671 & ~w39697;
assign w39886 = w39884 & w39885;
assign w39887 = ~w39695 & w39712;
assign w39888 = ~w39678 & ~w39713;
assign w39889 = w39672 & ~w39678;
assign w39890 = (w39678 & w39663) | (w39678 & w66324) | (w39663 & w66324);
assign w39891 = ~w39642 & w39661;
assign w39892 = w39683 & w39891;
assign w39893 = ~w39889 & ~w39890;
assign w39894 = ~w39892 & w39893;
assign w39895 = ~w39649 & w39697;
assign w39896 = w39894 & w39895;
assign w39897 = w39881 & ~w39887;
assign w39898 = ~w39888 & w39897;
assign w39899 = ~w39886 & w39898;
assign w39900 = ~w39896 & w39899;
assign w39901 = w39642 & ~w39661;
assign w39902 = w39704 & w39901;
assign w39903 = w39669 & ~w39902;
assign w39904 = w39894 & w39903;
assign w39905 = ~w39900 & ~w39904;
assign w39906 = pi2154 & w39905;
assign w39907 = ~pi2154 & ~w39905;
assign w39908 = ~w39906 & ~w39907;
assign w39909 = ~pi6967 & pi9040;
assign w39910 = ~pi6950 & ~pi9040;
assign w39911 = ~w39909 & ~w39910;
assign w39912 = pi2036 & ~w39911;
assign w39913 = ~pi2036 & w39911;
assign w39914 = ~w39912 & ~w39913;
assign w39915 = ~pi6990 & pi9040;
assign w39916 = ~pi7012 & ~pi9040;
assign w39917 = ~w39915 & ~w39916;
assign w39918 = pi2072 & ~w39917;
assign w39919 = ~pi2072 & w39917;
assign w39920 = ~w39918 & ~w39919;
assign w39921 = w39914 & ~w39920;
assign w39922 = ~pi6985 & pi9040;
assign w39923 = ~pi6967 & ~pi9040;
assign w39924 = ~w39922 & ~w39923;
assign w39925 = pi2058 & ~w39924;
assign w39926 = ~pi2058 & w39924;
assign w39927 = ~w39925 & ~w39926;
assign w39928 = w39921 & w39927;
assign w39929 = ~w39914 & ~w39927;
assign w39930 = ~w39928 & ~w39929;
assign w39931 = ~pi6951 & pi9040;
assign w39932 = ~pi6985 & ~pi9040;
assign w39933 = ~w39931 & ~w39932;
assign w39934 = pi2078 & ~w39933;
assign w39935 = ~pi2078 & w39933;
assign w39936 = ~w39934 & ~w39935;
assign w39937 = ~pi6994 & pi9040;
assign w39938 = ~pi6969 & ~pi9040;
assign w39939 = ~w39937 & ~w39938;
assign w39940 = pi2068 & ~w39939;
assign w39941 = ~pi2068 & w39939;
assign w39942 = ~w39940 & ~w39941;
assign w39943 = ~w39936 & w39942;
assign w39944 = ~w39930 & w39943;
assign w39945 = ~w39914 & w39920;
assign w39946 = w39927 & w39945;
assign w39947 = (~w39936 & ~w39945) | (~w39936 & w66325) | (~w39945 & w66325);
assign w39948 = w39927 & ~w39942;
assign w39949 = ~w39947 & w39948;
assign w39950 = ~w39927 & w39942;
assign w39951 = w39945 & w39950;
assign w39952 = w39920 & ~w39927;
assign w39953 = w39914 & w39952;
assign w39954 = ~w39920 & ~w39927;
assign w39955 = ~w39942 & w39954;
assign w39956 = ~w39953 & ~w39955;
assign w39957 = ~w39936 & ~w39956;
assign w39958 = ~pi6952 & pi9040;
assign w39959 = ~pi6996 & ~pi9040;
assign w39960 = ~w39958 & ~w39959;
assign w39961 = pi2056 & ~w39960;
assign w39962 = ~pi2056 & w39960;
assign w39963 = ~w39961 & ~w39962;
assign w39964 = ~w39921 & ~w39945;
assign w39965 = ~w39950 & ~w39964;
assign w39966 = w39936 & ~w39952;
assign w39967 = ~w39929 & w39966;
assign w39968 = ~w39965 & w39967;
assign w39969 = ~w39951 & w39963;
assign w39970 = ~w39949 & w39969;
assign w39971 = ~w39957 & ~w39968;
assign w39972 = w39970 & w39971;
assign w39973 = w39936 & ~w39956;
assign w39974 = w39921 & w66326;
assign w39975 = ~w39963 & ~w39974;
assign w39976 = ~w39914 & w39942;
assign w39977 = ~w39946 & ~w39954;
assign w39978 = w39976 & ~w39977;
assign w39979 = ~w39914 & ~w39920;
assign w39980 = w39942 & w39979;
assign w39981 = w39947 & ~w39980;
assign w39982 = ~w39927 & ~w39945;
assign w39983 = w39981 & ~w39982;
assign w39984 = ~w39973 & w39975;
assign w39985 = w39984 & w66327;
assign w39986 = ~w39972 & ~w39985;
assign w39987 = ~w39944 & ~w39986;
assign w39988 = pi2144 & w39987;
assign w39989 = ~pi2144 & ~w39987;
assign w39990 = ~w39988 & ~w39989;
assign w39991 = ~w39831 & w39833;
assign w39992 = ~w39776 & ~w39847;
assign w39993 = w39825 & ~w39992;
assign w39994 = ~w39841 & ~w39992;
assign w39995 = w39783 & ~w39994;
assign w39996 = w39813 & ~w39840;
assign w39997 = ~w39993 & w39996;
assign w39998 = ~w39995 & w39997;
assign w39999 = ~w39801 & ~w39821;
assign w40000 = ~w39783 & ~w39999;
assign w40001 = ~w39793 & ~w39806;
assign w40002 = w39842 & w40001;
assign w40003 = w39797 & ~w39807;
assign w40004 = ~w39813 & ~w40002;
assign w40005 = ~w40003 & w40004;
assign w40006 = ~w40000 & w40005;
assign w40007 = ~w39998 & ~w40006;
assign w40008 = ~w39991 & ~w40007;
assign w40009 = ~pi2146 & w40008;
assign w40010 = pi2146 & ~w40008;
assign w40011 = ~w40009 & ~w40010;
assign w40012 = w39522 & w39532;
assign w40013 = w39509 & ~w39534;
assign w40014 = ~w40012 & w40013;
assign w40015 = w39503 & w39523;
assign w40016 = w39532 & w66328;
assign w40017 = w39542 & w39564;
assign w40018 = ~w40015 & ~w40016;
assign w40019 = ~w40017 & w40018;
assign w40020 = ~w40014 & w40019;
assign w40021 = ~w39725 & w40020;
assign w40022 = ~w39531 & ~w40021;
assign w40023 = ~w39523 & ~w40012;
assign w40024 = w39565 & ~w40023;
assign w40025 = w39564 & w66329;
assign w40026 = ~w39568 & ~w40024;
assign w40027 = (w39531 & ~w40026) | (w39531 & w66330) | (~w40026 & w66330);
assign w40028 = ~w39737 & ~w40025;
assign w40029 = w39546 & ~w40028;
assign w40030 = ~w39740 & ~w39753;
assign w40031 = ~w40029 & w40030;
assign w40032 = ~w40027 & w40031;
assign w40033 = ~w40022 & w40032;
assign w40034 = ~pi2171 & w40033;
assign w40035 = pi2171 & ~w40033;
assign w40036 = ~w40034 & ~w40035;
assign w40037 = w39791 & w39800;
assign w40038 = ~w39801 & ~w40037;
assign w40039 = w39770 & w40038;
assign w40040 = w39833 & w39839;
assign w40041 = ~w39824 & ~w40040;
assign w40042 = ~w40040 & w63965;
assign w40043 = ~w39783 & ~w39805;
assign w40044 = w39814 & w39838;
assign w40045 = ~w40043 & ~w40044;
assign w40046 = w40042 & w40045;
assign w40047 = ~w40039 & ~w40046;
assign w40048 = w39813 & ~w40047;
assign w40049 = w40001 & ~w40045;
assign w40050 = w39802 & ~w39813;
assign w40051 = w40041 & ~w40049;
assign w40052 = ~w40050 & w40051;
assign w40053 = w39770 & w39838;
assign w40054 = ~w39820 & ~w40053;
assign w40055 = w39813 & w40054;
assign w40056 = ~w40052 & ~w40055;
assign w40057 = ~w40048 & ~w40056;
assign w40058 = ~pi2149 & w40057;
assign w40059 = pi2149 & ~w40057;
assign w40060 = ~w40058 & ~w40059;
assign w40061 = ~w39946 & w66331;
assign w40062 = w39920 & w39927;
assign w40063 = w39914 & w39936;
assign w40064 = ~w39976 & ~w40063;
assign w40065 = w40062 & ~w40064;
assign w40066 = w39954 & w66332;
assign w40067 = ~w40065 & ~w40066;
assign w40068 = w39950 & w39979;
assign w40069 = w39914 & w39948;
assign w40070 = w39936 & ~w40068;
assign w40071 = ~w40069 & w40070;
assign w40072 = ~w40067 & w40071;
assign w40073 = ~w39914 & w40072;
assign w40074 = ~w39964 & ~w40062;
assign w40075 = ~w39964 & w66333;
assign w40076 = ~w39914 & ~w39936;
assign w40077 = ~w39950 & ~w40076;
assign w40078 = w39920 & ~w40077;
assign w40079 = ~w40077 & w66334;
assign w40080 = ~w40061 & ~w40075;
assign w40081 = ~w40079 & w40080;
assign w40082 = (~w39963 & w40073) | (~w39963 & w66335) | (w40073 & w66335);
assign w40083 = w39954 & w40076;
assign w40084 = w39943 & ~w39977;
assign w40085 = ~w39950 & w40063;
assign w40086 = w39948 & w39964;
assign w40087 = ~w40083 & ~w40085;
assign w40088 = ~w40086 & w40087;
assign w40089 = ~w40084 & w40088;
assign w40090 = w39963 & ~w40089;
assign w40091 = ~w39927 & w40079;
assign w40092 = ~w39936 & ~w40091;
assign w40093 = ~w40071 & ~w40092;
assign w40094 = ~w40090 & ~w40093;
assign w40095 = ~w40082 & w40094;
assign w40096 = ~pi2155 & w40095;
assign w40097 = pi2155 & ~w40095;
assign w40098 = ~w40096 & ~w40097;
assign w40099 = ~pi6988 & pi9040;
assign w40100 = ~pi6961 & ~pi9040;
assign w40101 = ~w40099 & ~w40100;
assign w40102 = pi2069 & ~w40101;
assign w40103 = ~pi2069 & w40101;
assign w40104 = ~w40102 & ~w40103;
assign w40105 = ~pi6955 & pi9040;
assign w40106 = ~pi6966 & ~pi9040;
assign w40107 = ~w40105 & ~w40106;
assign w40108 = pi2070 & ~w40107;
assign w40109 = ~pi2070 & w40107;
assign w40110 = ~w40108 & ~w40109;
assign w40111 = w40104 & ~w40110;
assign w40112 = ~pi7003 & pi9040;
assign w40113 = ~pi6953 & ~pi9040;
assign w40114 = ~w40112 & ~w40113;
assign w40115 = pi2079 & ~w40114;
assign w40116 = ~pi2079 & w40114;
assign w40117 = ~w40115 & ~w40116;
assign w40118 = ~w40104 & ~w40117;
assign w40119 = ~w40111 & ~w40118;
assign w40120 = ~w40104 & w40110;
assign w40121 = ~w40117 & w40120;
assign w40122 = ~pi6946 & pi9040;
assign w40123 = ~pi6959 & ~pi9040;
assign w40124 = ~w40122 & ~w40123;
assign w40125 = pi2064 & ~w40124;
assign w40126 = ~pi2064 & w40124;
assign w40127 = ~w40125 & ~w40126;
assign w40128 = ~pi6975 & pi9040;
assign w40129 = ~pi6955 & ~pi9040;
assign w40130 = ~w40128 & ~w40129;
assign w40131 = pi2065 & ~w40130;
assign w40132 = ~pi2065 & w40130;
assign w40133 = ~w40131 & ~w40132;
assign w40134 = w40104 & w40133;
assign w40135 = ~w40110 & w40134;
assign w40136 = (~w40127 & ~w40120) | (~w40127 & w40162) | (~w40120 & w40162);
assign w40137 = ~w40135 & w40136;
assign w40138 = ~w40119 & w40137;
assign w40139 = ~w40111 & w40127;
assign w40140 = ~w40120 & ~w40139;
assign w40141 = w40110 & ~w40117;
assign w40142 = w40133 & w40141;
assign w40143 = ~w40110 & ~w40133;
assign w40144 = w40117 & ~w40133;
assign w40145 = ~w40104 & ~w40110;
assign w40146 = ~w40144 & ~w40145;
assign w40147 = ~w40143 & ~w40146;
assign w40148 = ~w40146 & w66336;
assign w40149 = w40110 & w40134;
assign w40150 = ~w40117 & w40143;
assign w40151 = ~w40149 & ~w40150;
assign w40152 = ~w40104 & ~w40146;
assign w40153 = w40127 & w40151;
assign w40154 = (~w40137 & ~w40153) | (~w40137 & w66337) | (~w40153 & w66337);
assign w40155 = ~pi6993 & pi9040;
assign w40156 = ~pi6992 & ~pi9040;
assign w40157 = ~w40155 & ~w40156;
assign w40158 = pi2043 & ~w40157;
assign w40159 = ~pi2043 & w40157;
assign w40160 = ~w40158 & ~w40159;
assign w40161 = (~w63966 & w66338) | (~w63966 & w66339) | (w66338 & w66339);
assign w40162 = w40117 & ~w40127;
assign w40163 = w40111 & w40162;
assign w40164 = w40134 & w40141;
assign w40165 = (w40160 & w40154) | (w40160 & w63967) | (w40154 & w63967);
assign w40166 = w40118 & w40133;
assign w40167 = ~w40144 & ~w40166;
assign w40168 = ~w40120 & w40139;
assign w40169 = ~w40167 & w40168;
assign w40170 = ~w40163 & ~w40164;
assign w40171 = ~w40169 & w40170;
assign w40172 = ~w40165 & w40171;
assign w40173 = ~w40161 & w40172;
assign w40174 = ~pi2156 & w40173;
assign w40175 = pi2156 & ~w40173;
assign w40176 = ~w40174 & ~w40175;
assign w40177 = ~w40104 & ~w40133;
assign w40178 = (w40127 & ~w40177) | (w40127 & w40191) | (~w40177 & w40191);
assign w40179 = ~w40151 & w40178;
assign w40180 = ~w40127 & w40133;
assign w40181 = w40120 & w40180;
assign w40182 = ~w40119 & w40180;
assign w40183 = ~w40110 & w40117;
assign w40184 = w40177 & w40183;
assign w40185 = ~w40121 & ~w40181;
assign w40186 = ~w40184 & w40185;
assign w40187 = ~w40182 & w40186;
assign w40188 = ~w40148 & ~w40179;
assign w40189 = w40187 & w40188;
assign w40190 = ~w40160 & ~w40189;
assign w40191 = w40110 & w40127;
assign w40192 = ~w40167 & w40191;
assign w40193 = w40104 & ~w40117;
assign w40194 = ~w40134 & ~w40141;
assign w40195 = ~w40193 & ~w40194;
assign w40196 = w40178 & ~w40195;
assign w40197 = ~w40143 & ~w40177;
assign w40198 = ~w40195 & w66340;
assign w40199 = w40183 & w40198;
assign w40200 = w40104 & ~w40133;
assign w40201 = w40183 & w40200;
assign w40202 = ~w40127 & w40201;
assign w40203 = w40118 & w40143;
assign w40204 = ~w40135 & ~w40203;
assign w40205 = w40127 & ~w40204;
assign w40206 = ~w40177 & ~w40183;
assign w40207 = w40147 & ~w40206;
assign w40208 = ~w40127 & w40193;
assign w40209 = ~w40205 & ~w40208;
assign w40210 = ~w40207 & w40209;
assign w40211 = w40160 & ~w40210;
assign w40212 = ~w40192 & ~w40202;
assign w40213 = ~w40199 & w40212;
assign w40214 = ~w40190 & w40213;
assign w40215 = w40214 & w66341;
assign w40216 = (pi2148 & ~w40214) | (pi2148 & w66342) | (~w40214 & w66342);
assign w40217 = ~w40215 & ~w40216;
assign w40218 = ~w40194 & ~w40206;
assign w40219 = ~w40127 & ~w40164;
assign w40220 = ~w40147 & w40219;
assign w40221 = w40143 & w40193;
assign w40222 = w40220 & ~w40221;
assign w40223 = ~w40160 & ~w40218;
assign w40224 = (w40223 & w40222) | (w40223 & w66343) | (w40222 & w66343);
assign w40225 = ~w40193 & ~w40201;
assign w40226 = w40151 & ~w40225;
assign w40227 = ~w40142 & ~w40203;
assign w40228 = w40220 & ~w40227;
assign w40229 = (w40160 & ~w40149) | (w40160 & w66344) | (~w40149 & w66344);
assign w40230 = ~w40226 & w40229;
assign w40231 = ~w40198 & w40230;
assign w40232 = ~w40228 & w40231;
assign w40233 = ~w40127 & w40207;
assign w40234 = w40141 & w40200;
assign w40235 = ~w40184 & ~w40234;
assign w40236 = w40127 & ~w40235;
assign w40237 = ~w40233 & ~w40236;
assign w40238 = (w40237 & w40232) | (w40237 & w66345) | (w40232 & w66345);
assign w40239 = pi2165 & w40238;
assign w40240 = ~pi2165 & ~w40238;
assign w40241 = ~w40239 & ~w40240;
assign w40242 = w39796 & w39825;
assign w40243 = w39799 & w39833;
assign w40244 = ~w40242 & ~w40243;
assign w40245 = w39764 & w39784;
assign w40246 = ~w39764 & w39847;
assign w40247 = w40054 & ~w40246;
assign w40248 = ~w40245 & w40247;
assign w40249 = (~w39813 & ~w40248) | (~w39813 & w66346) | (~w40248 & w66346);
assign w40250 = (~w40044 & w39822) | (~w40044 & w63968) | (w39822 & w63968);
assign w40251 = w40042 & w40250;
assign w40252 = w39803 & ~w40244;
assign w40253 = ~w39785 & ~w39845;
assign w40254 = ~w40038 & ~w40253;
assign w40255 = (~w39835 & ~w40038) | (~w39835 & w66347) | (~w40038 & w66347);
assign w40256 = (w39813 & w40254) | (w39813 & w66348) | (w40254 & w66348);
assign w40257 = ~w39848 & ~w40251;
assign w40258 = ~w40252 & w40257;
assign w40259 = ~w40249 & w40258;
assign w40260 = (pi2151 & ~w40259) | (pi2151 & w66349) | (~w40259 & w66349);
assign w40261 = w40259 & w66350;
assign w40262 = ~w40260 & ~w40261;
assign w40263 = w39516 & w39533;
assign w40264 = w39570 & ~w40263;
assign w40265 = w39751 & ~w40264;
assign w40266 = w39535 & w39536;
assign w40267 = ~w39726 & ~w40266;
assign w40268 = ~w40265 & w40267;
assign w40269 = ~w39531 & ~w40268;
assign w40270 = (w39750 & ~w40026) | (w39750 & w63969) | (~w40026 & w63969);
assign w40271 = ~w39543 & w39722;
assign w40272 = ~w39571 & ~w39749;
assign w40273 = (w39531 & ~w40272) | (w39531 & w66351) | (~w40272 & w66351);
assign w40274 = ~w39724 & ~w40270;
assign w40275 = ~w40273 & w40274;
assign w40276 = w40275 & w66352;
assign w40277 = (pi2161 & ~w40275) | (pi2161 & w66353) | (~w40275 & w66353);
assign w40278 = ~w40276 & ~w40277;
assign w40279 = ~pi6957 & pi9040;
assign w40280 = ~pi6968 & ~pi9040;
assign w40281 = ~w40279 & ~w40280;
assign w40282 = pi2072 & ~w40281;
assign w40283 = ~pi2072 & w40281;
assign w40284 = ~w40282 & ~w40283;
assign w40285 = ~pi6965 & pi9040;
assign w40286 = ~pi7082 & ~pi9040;
assign w40287 = ~w40285 & ~w40286;
assign w40288 = pi2056 & ~w40287;
assign w40289 = ~pi2056 & w40287;
assign w40290 = ~w40288 & ~w40289;
assign w40291 = ~w40284 & ~w40290;
assign w40292 = ~pi6969 & pi9040;
assign w40293 = ~pi6981 & ~pi9040;
assign w40294 = ~w40292 & ~w40293;
assign w40295 = pi2054 & ~w40294;
assign w40296 = ~pi2054 & w40294;
assign w40297 = ~w40295 & ~w40296;
assign w40298 = ~w40290 & ~w40297;
assign w40299 = ~pi6972 & pi9040;
assign w40300 = ~pi6974 & ~pi9040;
assign w40301 = ~w40299 & ~w40300;
assign w40302 = pi2067 & ~w40301;
assign w40303 = ~pi2067 & w40301;
assign w40304 = ~w40302 & ~w40303;
assign w40305 = ~pi6947 & pi9040;
assign w40306 = ~pi6954 & ~pi9040;
assign w40307 = ~w40305 & ~w40306;
assign w40308 = pi2053 & ~w40307;
assign w40309 = ~pi2053 & w40307;
assign w40310 = ~w40308 & ~w40309;
assign w40311 = (w40310 & ~w40298) | (w40310 & w66354) | (~w40298 & w66354);
assign w40312 = w40290 & w40297;
assign w40313 = ~w40284 & w40312;
assign w40314 = ~w40284 & ~w40297;
assign w40315 = ~w40290 & ~w40304;
assign w40316 = ~w40314 & w40315;
assign w40317 = ~w40313 & ~w40316;
assign w40318 = w40311 & w40317;
assign w40319 = w40291 & w40318;
assign w40320 = ~pi6986 & pi9040;
assign w40321 = ~pi6965 & ~pi9040;
assign w40322 = ~w40320 & ~w40321;
assign w40323 = pi2073 & ~w40322;
assign w40324 = ~pi2073 & w40322;
assign w40325 = ~w40323 & ~w40324;
assign w40326 = w40284 & w40297;
assign w40327 = ~w40314 & ~w40326;
assign w40328 = w40290 & w40304;
assign w40329 = ~w40315 & ~w40328;
assign w40330 = w40304 & w40310;
assign w40331 = w40329 & ~w40330;
assign w40332 = ~w40327 & ~w40331;
assign w40333 = ~w40311 & ~w40331;
assign w40334 = w40327 & w40329;
assign w40335 = ~w40333 & w40334;
assign w40336 = ~w40332 & ~w40335;
assign w40337 = ~w40325 & w40336;
assign w40338 = w40315 & w40325;
assign w40339 = w40326 & w40338;
assign w40340 = ~w40284 & w40304;
assign w40341 = ~w40284 & ~w40304;
assign w40342 = ~w40298 & ~w40341;
assign w40343 = w40329 & w40342;
assign w40344 = ~w40340 & ~w40343;
assign w40345 = w40310 & w40325;
assign w40346 = ~w40344 & w40345;
assign w40347 = w40313 & w40330;
assign w40348 = ~w40310 & w40325;
assign w40349 = ~w40315 & w40348;
assign w40350 = w40344 & w40349;
assign w40351 = ~w40339 & ~w40347;
assign w40352 = ~w40319 & w40351;
assign w40353 = ~w40346 & ~w40350;
assign w40354 = w40352 & w40353;
assign w40355 = ~w40337 & w40354;
assign w40356 = pi2195 & w40355;
assign w40357 = ~pi2195 & ~w40355;
assign w40358 = ~w40356 & ~w40357;
assign w40359 = ~w39662 & ~w39879;
assign w40360 = w39648 & w40359;
assign w40361 = w40359 & w66355;
assign w40362 = ~w39880 & ~w40361;
assign w40363 = ~w39642 & ~w40359;
assign w40364 = ~w40359 & w66356;
assign w40365 = w39678 & ~w40364;
assign w40366 = ~w39649 & ~w39901;
assign w40367 = w39695 & ~w40366;
assign w40368 = ~w39884 & ~w40360;
assign w40369 = ~w40367 & w40368;
assign w40370 = (w40362 & w40369) | (w40362 & w66357) | (w40369 & w66357);
assign w40371 = w39669 & ~w40370;
assign w40372 = w39881 & ~w40363;
assign w40373 = ~w40361 & w40372;
assign w40374 = w39711 & ~w40373;
assign w40375 = ~w39703 & ~w40364;
assign w40376 = ~w39669 & ~w40375;
assign w40377 = ~w39678 & w40362;
assign w40378 = ~w40376 & w40377;
assign w40379 = ~w40374 & ~w40378;
assign w40380 = ~w40371 & ~w40379;
assign w40381 = ~pi2201 & w40380;
assign w40382 = pi2201 & ~w40380;
assign w40383 = ~w40381 & ~w40382;
assign w40384 = ~w40291 & ~w40315;
assign w40385 = w40310 & w40384;
assign w40386 = ~w40297 & ~w40315;
assign w40387 = ~w40342 & w40386;
assign w40388 = w40385 & w40387;
assign w40389 = (w40314 & w40331) | (w40314 & w66358) | (w40331 & w66358);
assign w40390 = w40314 & ~w40329;
assign w40391 = ~w40343 & ~w40390;
assign w40392 = ~w40310 & w40391;
assign w40393 = w40391 & w63970;
assign w40394 = (w40325 & w40393) | (w40325 & w66359) | (w40393 & w66359);
assign w40395 = w40312 & w40341;
assign w40396 = (~w40395 & w40392) | (~w40395 & w66360) | (w40392 & w66360);
assign w40397 = ~w40325 & ~w40396;
assign w40398 = (~w40291 & w40329) | (~w40291 & w66361) | (w40329 & w66361);
assign w40399 = w40297 & w40315;
assign w40400 = ~w40310 & ~w40399;
assign w40401 = ~w40398 & w40400;
assign w40402 = w40326 & w40401;
assign w40403 = w40297 & w40345;
assign w40404 = w40317 & w40403;
assign w40405 = ~w40388 & ~w40404;
assign w40406 = ~w40402 & w40405;
assign w40407 = ~w40394 & w40406;
assign w40408 = ~w40397 & w40407;
assign w40409 = pi2186 & ~w40408;
assign w40410 = ~pi2186 & w40408;
assign w40411 = ~w40409 & ~w40410;
assign w40412 = w40127 & w40221;
assign w40413 = ~w40166 & ~w40200;
assign w40414 = ~w40183 & ~w40219;
assign w40415 = w40413 & ~w40414;
assign w40416 = w40139 & ~w40413;
assign w40417 = ~w40160 & ~w40416;
assign w40418 = ~w40415 & w40417;
assign w40419 = w40133 & ~w40193;
assign w40420 = ~w40200 & ~w40419;
assign w40421 = w40178 & w40420;
assign w40422 = w40160 & ~w40181;
assign w40423 = ~w40201 & w40422;
assign w40424 = ~w40164 & w40423;
assign w40425 = ~w40421 & w40424;
assign w40426 = ~w40418 & ~w40425;
assign w40427 = ~w40193 & ~w40204;
assign w40428 = ~w40234 & ~w40427;
assign w40429 = ~w40127 & ~w40428;
assign w40430 = ~w40199 & ~w40412;
assign w40431 = ~w40429 & w40430;
assign w40432 = ~w40426 & w40431;
assign w40433 = pi2179 & ~w40432;
assign w40434 = ~pi2179 & w40432;
assign w40435 = ~w40433 & ~w40434;
assign w40436 = w40284 & ~w40304;
assign w40437 = ~w40312 & ~w40436;
assign w40438 = ~w40291 & ~w40310;
assign w40439 = w40437 & w40438;
assign w40440 = ~w40284 & ~w40391;
assign w40441 = w40290 & ~w40436;
assign w40442 = w40297 & ~w40441;
assign w40443 = w40310 & ~w40437;
assign w40444 = ~w40442 & w40443;
assign w40445 = ~w40439 & ~w40444;
assign w40446 = ~w40440 & w40445;
assign w40447 = ~w40325 & ~w40446;
assign w40448 = ~w40387 & ~w40399;
assign w40449 = w40345 & ~w40448;
assign w40450 = ~w40304 & ~w40310;
assign w40451 = ~w40325 & ~w40450;
assign w40452 = w40326 & ~w40328;
assign w40453 = ~w40451 & w40452;
assign w40454 = w40348 & ~w40386;
assign w40455 = ~w40437 & w40454;
assign w40456 = ~w40347 & ~w40453;
assign w40457 = ~w40455 & w40456;
assign w40458 = ~w40449 & w40457;
assign w40459 = ~w40447 & w40458;
assign w40460 = pi2205 & ~w40459;
assign w40461 = ~pi2205 & w40459;
assign w40462 = ~w40460 & ~w40461;
assign w40463 = w39430 & ~w39464;
assign w40464 = ~w39419 & ~w39459;
assign w40465 = w39430 & w63971;
assign w40466 = ~w39418 & ~w39453;
assign w40467 = ~w39403 & ~w40466;
assign w40468 = ~w39420 & w39441;
assign w40469 = ~w40467 & w40468;
assign w40470 = ~w40465 & ~w40469;
assign w40471 = w39402 & ~w39417;
assign w40472 = w39450 & w40471;
assign w40473 = w39441 & w39458;
assign w40474 = w39411 & ~w39462;
assign w40475 = w40473 & w40474;
assign w40476 = (w39472 & ~w40463) | (w39472 & w63972) | (~w40463 & w63972);
assign w40477 = ~w39447 & ~w40472;
assign w40478 = (w40477 & w39435) | (w40477 & w66362) | (w39435 & w66362);
assign w40479 = ~w40476 & w40478;
assign w40480 = (pi2200 & ~w40479) | (pi2200 & w63973) | (~w40479 & w63973);
assign w40481 = w40479 & w63974;
assign w40482 = ~w40480 & ~w40481;
assign w40483 = ~w39445 & ~w39478;
assign w40484 = w39434 & ~w40483;
assign w40485 = ~w39472 & ~w40484;
assign w40486 = w39472 & ~w39475;
assign w40487 = ~w39441 & ~w40486;
assign w40488 = w39461 & ~w40487;
assign w40489 = w39417 & w39451;
assign w40490 = ~w40486 & w40489;
assign w40491 = w39457 & w40471;
assign w40492 = (w39441 & ~w39425) | (w39441 & w66363) | (~w39425 & w66363);
assign w40493 = ~w39446 & ~w40491;
assign w40494 = ~w40492 & w40493;
assign w40495 = w39472 & ~w40494;
assign w40496 = ~w40488 & ~w40490;
assign w40497 = ~w40495 & w40496;
assign w40498 = ~w40485 & w40497;
assign w40499 = pi2172 & ~w40498;
assign w40500 = ~pi2172 & w40498;
assign w40501 = ~w40499 & ~w40500;
assign w40502 = w39952 & w40077;
assign w40503 = w39921 & ~w39948;
assign w40504 = ~w40086 & ~w40503;
assign w40505 = w39966 & w40504;
assign w40506 = ~w40502 & ~w40505;
assign w40507 = ~w39963 & ~w40506;
assign w40508 = ~w40086 & w66364;
assign w40509 = ~w39936 & ~w40508;
assign w40510 = ~w39963 & ~w40509;
assign w40511 = ~w39965 & ~w40069;
assign w40512 = ~w40504 & ~w40511;
assign w40513 = w39963 & w39981;
assign w40514 = ~w39942 & w39979;
assign w40515 = w39936 & ~w40514;
assign w40516 = ~w40078 & w40515;
assign w40517 = ~w40513 & ~w40516;
assign w40518 = ~w40079 & ~w40512;
assign w40519 = ~w40517 & w40518;
assign w40520 = ~w40510 & ~w40519;
assign w40521 = ~w40520 & w66365;
assign w40522 = (~pi2157 & w40520) | (~pi2157 & w66366) | (w40520 & w66366);
assign w40523 = ~w40521 & ~w40522;
assign w40524 = w40310 & w40442;
assign w40525 = ~w40335 & w66367;
assign w40526 = ~w40310 & w40313;
assign w40527 = w40304 & w40452;
assign w40528 = ~w40340 & w40441;
assign w40529 = ~w40341 & ~w40384;
assign w40530 = ~w40438 & w40529;
assign w40531 = (~w40297 & w40530) | (~w40297 & w66368) | (w40530 & w66368);
assign w40532 = ~w40298 & ~w40312;
assign w40533 = w40450 & w40532;
assign w40534 = w40325 & ~w40527;
assign w40535 = ~w40533 & w40534;
assign w40536 = ~w40531 & w40535;
assign w40537 = w40385 & ~w40528;
assign w40538 = w40298 & w40341;
assign w40539 = ~w40325 & ~w40538;
assign w40540 = ~w40537 & w40539;
assign w40541 = ~w40401 & w40540;
assign w40542 = ~w40536 & ~w40541;
assign w40543 = ~w40525 & ~w40526;
assign w40544 = ~w40542 & w40543;
assign w40545 = pi2180 & ~w40544;
assign w40546 = ~pi2180 & w40544;
assign w40547 = ~w40545 & ~w40546;
assign w40548 = ~w39700 & w39888;
assign w40549 = ~w39714 & ~w40548;
assign w40550 = ~w39696 & ~w39709;
assign w40551 = ~w39695 & ~w40550;
assign w40552 = w39669 & ~w40551;
assign w40553 = w39662 & ~w40550;
assign w40554 = ~w39701 & w39882;
assign w40555 = ~w40553 & ~w40554;
assign w40556 = w39669 & ~w40555;
assign w40557 = ~w39686 & ~w39901;
assign w40558 = w40552 & ~w40557;
assign w40559 = w40549 & w40558;
assign w40560 = w39655 & ~w39669;
assign w40561 = ~w39882 & w40560;
assign w40562 = w40557 & w40561;
assign w40563 = (~w40562 & w40549) | (~w40562 & w66369) | (w40549 & w66369);
assign w40564 = ~w40559 & w40563;
assign w40565 = ~w40556 & w40564;
assign w40566 = pi2177 & ~w40565;
assign w40567 = ~pi2177 & w40565;
assign w40568 = ~w40566 & ~w40567;
assign w40569 = ~w39921 & w39948;
assign w40570 = ~w39980 & ~w40569;
assign w40571 = w39963 & ~w40570;
assign w40572 = ~w39953 & ~w40571;
assign w40573 = ~w39936 & ~w40572;
assign w40574 = w39936 & w40074;
assign w40575 = w39963 & ~w40068;
assign w40576 = ~w40574 & w40575;
assign w40577 = ~w39929 & ~w39950;
assign w40578 = w40064 & ~w40577;
assign w40579 = ~w40065 & ~w40514;
assign w40580 = ~w40578 & w40579;
assign w40581 = w39975 & w40580;
assign w40582 = ~w40576 & ~w40581;
assign w40583 = ~w40072 & ~w40573;
assign w40584 = ~w40582 & w40583;
assign w40585 = pi2188 & w40584;
assign w40586 = ~pi2188 & ~w40584;
assign w40587 = ~w40585 & ~w40586;
assign w40588 = w39427 & ~w39448;
assign w40589 = ~w40473 & ~w40588;
assign w40590 = ~w39472 & ~w40589;
assign w40591 = ~w39396 & w39441;
assign w40592 = w39444 & ~w40591;
assign w40593 = w39405 & w39421;
assign w40594 = ~w40592 & ~w40593;
assign w40595 = w39472 & ~w40594;
assign w40596 = w39432 & w39472;
assign w40597 = ~w39426 & ~w40596;
assign w40598 = w40591 & ~w40597;
assign w40599 = ~w39460 & ~w40595;
assign w40600 = ~w40598 & w40599;
assign w40601 = ~w40590 & w40600;
assign w40602 = ~pi2191 & w40601;
assign w40603 = pi2191 & ~w40601;
assign w40604 = ~w40602 & ~w40603;
assign w40605 = ~pi7202 & pi9040;
assign w40606 = ~pi7185 & ~pi9040;
assign w40607 = ~w40605 & ~w40606;
assign w40608 = pi2225 & ~w40607;
assign w40609 = ~pi2225 & w40607;
assign w40610 = ~w40608 & ~w40609;
assign w40611 = ~pi7190 & pi9040;
assign w40612 = ~pi7200 & ~pi9040;
assign w40613 = ~w40611 & ~w40612;
assign w40614 = pi2211 & ~w40613;
assign w40615 = ~pi2211 & w40613;
assign w40616 = ~w40614 & ~w40615;
assign w40617 = w40610 & w40616;
assign w40618 = ~pi7241 & pi9040;
assign w40619 = ~pi7240 & ~pi9040;
assign w40620 = ~w40618 & ~w40619;
assign w40621 = pi2208 & ~w40620;
assign w40622 = ~pi2208 & w40620;
assign w40623 = ~w40621 & ~w40622;
assign w40624 = w40617 & w40623;
assign w40625 = ~pi7196 & pi9040;
assign w40626 = ~pi7204 & ~pi9040;
assign w40627 = ~w40625 & ~w40626;
assign w40628 = pi2158 & ~w40627;
assign w40629 = ~pi2158 & w40627;
assign w40630 = ~w40628 & ~w40629;
assign w40631 = ~w40623 & ~w40630;
assign w40632 = w40610 & w40630;
assign w40633 = ~w40631 & ~w40632;
assign w40634 = ~w40623 & w40633;
assign w40635 = ~w40624 & ~w40634;
assign w40636 = w40623 & w40630;
assign w40637 = ~w40616 & ~w40636;
assign w40638 = ~pi7239 & pi9040;
assign w40639 = ~pi7237 & ~pi9040;
assign w40640 = ~w40638 & ~w40639;
assign w40641 = pi2189 & ~w40640;
assign w40642 = ~pi2189 & w40640;
assign w40643 = ~w40641 & ~w40642;
assign w40644 = ~w40637 & w40643;
assign w40645 = ~w40610 & ~w40616;
assign w40646 = w40623 & ~w40630;
assign w40647 = w40645 & w40646;
assign w40648 = w40616 & w40636;
assign w40649 = ~w40647 & ~w40648;
assign w40650 = w40633 & w40649;
assign w40651 = ~w40644 & ~w40650;
assign w40652 = w40635 & ~w40651;
assign w40653 = w40631 & w40645;
assign w40654 = ~w40634 & w66370;
assign w40655 = ~w40610 & w40616;
assign w40656 = w40636 & w40655;
assign w40657 = ~w40616 & w40623;
assign w40658 = ~w40655 & ~w40657;
assign w40659 = w40633 & w40658;
assign w40660 = w40616 & w40631;
assign w40661 = ~w40616 & w40632;
assign w40662 = ~w40643 & ~w40647;
assign w40663 = ~w40660 & ~w40661;
assign w40664 = w40662 & w40663;
assign w40665 = ~w40656 & ~w40659;
assign w40666 = w40664 & w40665;
assign w40667 = ~w40654 & w40666;
assign w40668 = ~w40652 & ~w40667;
assign w40669 = ~pi7244 & pi9040;
assign w40670 = ~pi7209 & ~pi9040;
assign w40671 = ~w40669 & ~w40670;
assign w40672 = pi2162 & ~w40671;
assign w40673 = ~pi2162 & w40671;
assign w40674 = ~w40672 & ~w40673;
assign w40675 = ~w40668 & w40674;
assign w40676 = ~w40616 & w40631;
assign w40677 = w40643 & ~w40676;
assign w40678 = w40635 & w40677;
assign w40679 = ~w40666 & ~w40674;
assign w40680 = ~w40678 & w40679;
assign w40681 = w40616 & ~w40623;
assign w40682 = ~w40657 & ~w40681;
assign w40683 = ~w40636 & ~w40655;
assign w40684 = ~w40682 & ~w40683;
assign w40685 = w40643 & w40684;
assign w40686 = w40616 & w40646;
assign w40687 = ~w40658 & ~w40686;
assign w40688 = ~w40643 & ~w40687;
assign w40689 = ~w40632 & ~w40657;
assign w40690 = w40610 & w40689;
assign w40691 = ~w40685 & ~w40690;
assign w40692 = ~w40688 & w40691;
assign w40693 = ~w40645 & w40677;
assign w40694 = ~w40664 & ~w40693;
assign w40695 = ~w40692 & w40694;
assign w40696 = ~w40680 & ~w40695;
assign w40697 = ~w40675 & w40696;
assign w40698 = pi2080 & w40697;
assign w40699 = ~pi2080 & ~w40697;
assign w40700 = ~w40698 & ~w40699;
assign w40701 = ~pi7237 & pi9040;
assign w40702 = ~pi7197 & ~pi9040;
assign w40703 = ~w40701 & ~w40702;
assign w40704 = pi2160 & ~w40703;
assign w40705 = ~pi2160 & w40703;
assign w40706 = ~w40704 & ~w40705;
assign w40707 = ~pi7186 & pi9040;
assign w40708 = ~pi7241 & ~pi9040;
assign w40709 = ~w40707 & ~w40708;
assign w40710 = pi2176 & ~w40709;
assign w40711 = ~pi2176 & w40709;
assign w40712 = ~w40710 & ~w40711;
assign w40713 = ~pi7213 & pi9040;
assign w40714 = ~pi7202 & ~pi9040;
assign w40715 = ~w40713 & ~w40714;
assign w40716 = pi2192 & ~w40715;
assign w40717 = ~pi2192 & w40715;
assign w40718 = ~w40716 & ~w40717;
assign w40719 = w40712 & ~w40718;
assign w40720 = ~pi7209 & pi9040;
assign w40721 = ~pi7189 & ~pi9040;
assign w40722 = ~w40720 & ~w40721;
assign w40723 = pi2159 & ~w40722;
assign w40724 = ~pi2159 & w40722;
assign w40725 = ~w40723 & ~w40724;
assign w40726 = ~pi7216 & pi9040;
assign w40727 = ~pi7223 & ~pi9040;
assign w40728 = ~w40726 & ~w40727;
assign w40729 = pi2238 & ~w40728;
assign w40730 = ~pi2238 & w40728;
assign w40731 = ~w40729 & ~w40730;
assign w40732 = w40725 & ~w40731;
assign w40733 = ~w40719 & w40732;
assign w40734 = w40719 & ~w40732;
assign w40735 = ~w40733 & ~w40734;
assign w40736 = w40706 & ~w40735;
assign w40737 = w40712 & w40725;
assign w40738 = w40718 & w40737;
assign w40739 = ~w40732 & ~w40738;
assign w40740 = ~w40736 & ~w40739;
assign w40741 = ~w40718 & w40731;
assign w40742 = ~w40725 & w40741;
assign w40743 = w40712 & w40718;
assign w40744 = ~w40706 & ~w40743;
assign w40745 = ~w40742 & w40744;
assign w40746 = ~w40712 & ~w40725;
assign w40747 = w40718 & w40746;
assign w40748 = (w40706 & ~w40746) | (w40706 & w41468) | (~w40746 & w41468);
assign w40749 = ~w40712 & w40725;
assign w40750 = w40731 & w40749;
assign w40751 = w40749 & w40741;
assign w40752 = w40748 & ~w40751;
assign w40753 = ~w40745 & ~w40752;
assign w40754 = ~pi7195 & pi9040;
assign w40755 = ~pi7225 & ~pi9040;
assign w40756 = ~w40754 & ~w40755;
assign w40757 = pi2221 & ~w40756;
assign w40758 = ~pi2221 & w40756;
assign w40759 = ~w40757 & ~w40758;
assign w40760 = (~w40759 & w40740) | (~w40759 & w66371) | (w40740 & w66371);
assign w40761 = ~w40731 & w40746;
assign w40762 = ~w40750 & ~w40761;
assign w40763 = ~w40706 & ~w40762;
assign w40764 = ~w40725 & w40743;
assign w40765 = w40743 & w66372;
assign w40766 = (~w40765 & w40735) | (~w40765 & w66373) | (w40735 & w66373);
assign w40767 = ~w40763 & w40766;
assign w40768 = w40759 & ~w40767;
assign w40769 = w40741 & w63975;
assign w40770 = ~w40712 & w40718;
assign w40771 = ~w40731 & w40770;
assign w40772 = ~w40769 & ~w40771;
assign w40773 = ~w40735 & ~w40772;
assign w40774 = w40718 & w40731;
assign w40775 = ~w40718 & ~w40731;
assign w40776 = ~w40774 & ~w40775;
assign w40777 = w40746 & ~w40776;
assign w40778 = (w40706 & w40773) | (w40706 & w66374) | (w40773 & w66374);
assign w40779 = w40744 & ~w40776;
assign w40780 = w40737 & w40779;
assign w40781 = ~w40760 & ~w40780;
assign w40782 = ~w40768 & ~w40778;
assign w40783 = w40781 & w40782;
assign w40784 = pi2093 & ~w40783;
assign w40785 = ~pi2093 & w40783;
assign w40786 = ~w40784 & ~w40785;
assign w40787 = w40610 & w40646;
assign w40788 = ~w40643 & w40787;
assign w40789 = w40617 & w40631;
assign w40790 = w40643 & ~w40789;
assign w40791 = (w40610 & w40684) | (w40610 & w66375) | (w40684 & w66375);
assign w40792 = ~w40660 & ~w40791;
assign w40793 = w40790 & ~w40792;
assign w40794 = w40630 & w40643;
assign w40795 = w40645 & w40794;
assign w40796 = ~w40610 & ~w40643;
assign w40797 = w40630 & w40681;
assign w40798 = ~w40796 & ~w40797;
assign w40799 = ~w40633 & ~w40798;
assign w40800 = ~w40636 & ~w40643;
assign w40801 = ~w40689 & w40800;
assign w40802 = ~w40674 & ~w40795;
assign w40803 = ~w40801 & w40802;
assign w40804 = ~w40799 & w40803;
assign w40805 = ~w40687 & w66376;
assign w40806 = w40630 & w40655;
assign w40807 = ~w40650 & w40798;
assign w40808 = ~w40688 & w40807;
assign w40809 = w40674 & ~w40806;
assign w40810 = ~w40805 & w40809;
assign w40811 = (~w40804 & w40808) | (~w40804 & w66377) | (w40808 & w66377);
assign w40812 = ~w40656 & ~w40788;
assign w40813 = ~w40793 & w40812;
assign w40814 = ~w40811 & w40813;
assign w40815 = pi2081 & ~w40814;
assign w40816 = ~pi2081 & w40814;
assign w40817 = ~w40815 & ~w40816;
assign w40818 = ~pi7187 & pi9040;
assign w40819 = ~pi7208 & ~pi9040;
assign w40820 = ~w40818 & ~w40819;
assign w40821 = pi2158 & ~w40820;
assign w40822 = ~pi2158 & w40820;
assign w40823 = ~w40821 & ~w40822;
assign w40824 = ~pi7242 & pi9040;
assign w40825 = ~pi7217 & ~pi9040;
assign w40826 = ~w40824 & ~w40825;
assign w40827 = pi2196 & ~w40826;
assign w40828 = ~pi2196 & w40826;
assign w40829 = ~w40827 & ~w40828;
assign w40830 = ~w40823 & ~w40829;
assign w40831 = ~pi7243 & pi9040;
assign w40832 = ~pi7219 & ~pi9040;
assign w40833 = ~w40831 & ~w40832;
assign w40834 = pi2199 & ~w40833;
assign w40835 = ~pi2199 & w40833;
assign w40836 = ~w40834 & ~w40835;
assign w40837 = ~pi7199 & pi9040;
assign w40838 = ~pi7215 & ~pi9040;
assign w40839 = ~w40837 & ~w40838;
assign w40840 = pi2182 & ~w40839;
assign w40841 = ~pi2182 & w40839;
assign w40842 = ~w40840 & ~w40841;
assign w40843 = ~w40836 & w40842;
assign w40844 = w40836 & ~w40842;
assign w40845 = ~w40843 & ~w40844;
assign w40846 = w40830 & w40845;
assign w40847 = ~w40823 & w40836;
assign w40848 = w40829 & w40847;
assign w40849 = w40847 & w66378;
assign w40850 = ~pi7188 & pi9040;
assign w40851 = ~pi7203 & ~pi9040;
assign w40852 = ~w40850 & ~w40851;
assign w40853 = pi2229 & ~w40852;
assign w40854 = ~pi2229 & w40852;
assign w40855 = ~w40853 & ~w40854;
assign w40856 = ~w40849 & w40855;
assign w40857 = ~w40846 & w40856;
assign w40858 = w40823 & ~w40836;
assign w40859 = ~w40829 & w40842;
assign w40860 = w40858 & w40859;
assign w40861 = ~w40855 & ~w40860;
assign w40862 = ~w40857 & ~w40861;
assign w40863 = w40823 & ~w40842;
assign w40864 = ~w40855 & ~w40863;
assign w40865 = ~w40848 & w40864;
assign w40866 = ~w40847 & ~w40858;
assign w40867 = w40845 & w40866;
assign w40868 = w40855 & ~w40867;
assign w40869 = ~w40865 & ~w40868;
assign w40870 = w40829 & w40842;
assign w40871 = ~w40823 & ~w40836;
assign w40872 = w40870 & w40871;
assign w40873 = ~w40829 & ~w40842;
assign w40874 = w40866 & w40873;
assign w40875 = ~w40836 & w40855;
assign w40876 = w40870 & w40875;
assign w40877 = ~pi7221 & pi9040;
assign w40878 = ~pi7210 & ~pi9040;
assign w40879 = ~w40877 & ~w40878;
assign w40880 = pi2208 & ~w40879;
assign w40881 = ~pi2208 & w40879;
assign w40882 = ~w40880 & ~w40881;
assign w40883 = ~w40872 & ~w40882;
assign w40884 = ~w40876 & w40883;
assign w40885 = ~w40874 & w40884;
assign w40886 = ~w40869 & w40885;
assign w40887 = w40823 & w40836;
assign w40888 = w40870 & w40887;
assign w40889 = w40882 & ~w40888;
assign w40890 = w40845 & w63976;
assign w40891 = w40865 & w40890;
assign w40892 = w40842 & w40855;
assign w40893 = w40847 & w40892;
assign w40894 = ~w40842 & ~w40855;
assign w40895 = w40858 & ~w40894;
assign w40896 = ~w40870 & w40895;
assign w40897 = ~w40829 & ~w40855;
assign w40898 = ~w40845 & w40897;
assign w40899 = w40889 & ~w40893;
assign w40900 = ~w40896 & ~w40898;
assign w40901 = w40899 & w40900;
assign w40902 = ~w40891 & w40901;
assign w40903 = ~w40886 & ~w40902;
assign w40904 = ~w40862 & ~w40903;
assign w40905 = ~pi2082 & w40904;
assign w40906 = pi2082 & ~w40904;
assign w40907 = ~w40905 & ~w40906;
assign w40908 = w40823 & ~w40829;
assign w40909 = w40844 & w40855;
assign w40910 = w40908 & w40909;
assign w40911 = w40829 & w40895;
assign w40912 = ~w40829 & w40871;
assign w40913 = ~w40848 & ~w40912;
assign w40914 = w40842 & ~w40913;
assign w40915 = ~w40836 & ~w40873;
assign w40916 = ~w40829 & w40836;
assign w40917 = w40823 & ~w40855;
assign w40918 = ~w40916 & w40917;
assign w40919 = ~w40915 & w40918;
assign w40920 = w40867 & w40875;
assign w40921 = ~w40911 & ~w40919;
assign w40922 = ~w40914 & w40921;
assign w40923 = ~w40920 & w40922;
assign w40924 = w40882 & ~w40923;
assign w40925 = w40829 & ~w40858;
assign w40926 = w40842 & ~w40847;
assign w40927 = ~w40925 & w40926;
assign w40928 = ~w40855 & w40927;
assign w40929 = (~w40860 & ~w40927) | (~w40860 & w66379) | (~w40927 & w66379);
assign w40930 = ~w40918 & ~w40929;
assign w40931 = ~w40842 & w40916;
assign w40932 = ~w40892 & ~w40931;
assign w40933 = ~w40927 & ~w40932;
assign w40934 = ~w40860 & ~w40933;
assign w40935 = ~w40882 & ~w40934;
assign w40936 = ~w40882 & ~w40887;
assign w40937 = ~w40916 & ~w40936;
assign w40938 = w40894 & ~w40908;
assign w40939 = ~w40937 & w40938;
assign w40940 = ~w40910 & ~w40939;
assign w40941 = ~w40930 & w40940;
assign w40942 = ~w40935 & w40941;
assign w40943 = ~w40924 & w40942;
assign w40944 = pi2099 & ~w40943;
assign w40945 = ~pi2099 & w40943;
assign w40946 = ~w40944 & ~w40945;
assign w40947 = ~pi7206 & pi9040;
assign w40948 = ~pi7244 & ~pi9040;
assign w40949 = ~w40947 & ~w40948;
assign w40950 = pi2184 & ~w40949;
assign w40951 = ~pi2184 & w40949;
assign w40952 = ~w40950 & ~w40951;
assign w40953 = ~pi7204 & pi9040;
assign w40954 = ~pi7216 & ~pi9040;
assign w40955 = ~w40953 & ~w40954;
assign w40956 = pi2243 & ~w40955;
assign w40957 = ~pi2243 & w40955;
assign w40958 = ~w40956 & ~w40957;
assign w40959 = w40952 & w40958;
assign w40960 = ~pi7185 & pi9040;
assign w40961 = ~pi7195 & ~pi9040;
assign w40962 = ~w40960 & ~w40961;
assign w40963 = pi2162 & ~w40962;
assign w40964 = ~pi2162 & w40962;
assign w40965 = ~w40963 & ~w40964;
assign w40966 = w40959 & w40965;
assign w40967 = ~pi7240 & pi9040;
assign w40968 = ~pi7192 & ~pi9040;
assign w40969 = ~w40967 & ~w40968;
assign w40970 = pi2211 & ~w40969;
assign w40971 = ~pi2211 & w40969;
assign w40972 = ~w40970 & ~w40971;
assign w40973 = ~w40958 & w40972;
assign w40974 = ~w40952 & ~w40965;
assign w40975 = ~w40973 & w40974;
assign w40976 = ~w40966 & ~w40975;
assign w40977 = ~pi7189 & pi9040;
assign w40978 = ~pi7184 & ~pi9040;
assign w40979 = ~w40977 & ~w40978;
assign w40980 = pi2168 & ~w40979;
assign w40981 = ~pi2168 & w40979;
assign w40982 = ~w40980 & ~w40981;
assign w40983 = ~w40976 & ~w40982;
assign w40984 = ~w40965 & ~w40972;
assign w40985 = ~w40952 & ~w40958;
assign w40986 = ~w40959 & w40984;
assign w40987 = ~w40985 & w40986;
assign w40988 = ~w40952 & w40965;
assign w40989 = ~w40958 & ~w40982;
assign w40990 = w40988 & w40989;
assign w40991 = w40965 & ~w40972;
assign w40992 = w40959 & w40991;
assign w40993 = ~w40990 & ~w40992;
assign w40994 = ~w40987 & w40993;
assign w40995 = w40952 & w40972;
assign w40996 = ~w40965 & w40995;
assign w40997 = w40972 & w40988;
assign w40998 = w40988 & w63977;
assign w40999 = w40972 & w40974;
assign w41000 = w40974 & w40973;
assign w41001 = ~w40996 & ~w40998;
assign w41002 = (w40982 & ~w41001) | (w40982 & w66380) | (~w41001 & w66380);
assign w41003 = w40994 & ~w41002;
assign w41004 = ~w40983 & w41003;
assign w41005 = ~pi7222 & pi9040;
assign w41006 = ~pi7213 & ~pi9040;
assign w41007 = ~w41005 & ~w41006;
assign w41008 = pi2224 & ~w41007;
assign w41009 = ~pi2224 & w41007;
assign w41010 = ~w41008 & ~w41009;
assign w41011 = ~w41004 & w41010;
assign w41012 = w40982 & ~w41010;
assign w41013 = w40958 & ~w40965;
assign w41014 = ~w40972 & ~w41013;
assign w41015 = w40972 & w41013;
assign w41016 = ~w41014 & ~w41015;
assign w41017 = ~w40952 & ~w41016;
assign w41018 = w40965 & w40995;
assign w41019 = ~w41017 & ~w41018;
assign w41020 = w41012 & ~w41019;
assign w41021 = w40959 & ~w41010;
assign w41022 = w40984 & w41021;
assign w41023 = w40952 & w40982;
assign w41024 = w40973 & w41023;
assign w41025 = ~w40982 & ~w41010;
assign w41026 = ~w40984 & ~w40988;
assign w41027 = ~w40958 & w41026;
assign w41028 = ~w40998 & ~w41027;
assign w41029 = w41025 & ~w41028;
assign w41030 = w40985 & w40991;
assign w41031 = ~w41024 & ~w41030;
assign w41032 = ~w41022 & w41031;
assign w41033 = ~w41029 & w41032;
assign w41034 = ~w41020 & w41033;
assign w41035 = ~w41011 & w41034;
assign w41036 = pi2091 & w41035;
assign w41037 = ~pi2091 & ~w41035;
assign w41038 = ~w41036 & ~w41037;
assign w41039 = (~w40674 & ~w40691) | (~w40674 & w66381) | (~w40691 & w66381);
assign w41040 = ~w40647 & w40790;
assign w41041 = ~w40653 & ~w40686;
assign w41042 = w40683 & ~w41041;
assign w41043 = w40636 & w40645;
assign w41044 = ~w40643 & ~w41043;
assign w41045 = ~w41042 & w41044;
assign w41046 = ~w41040 & ~w41045;
assign w41047 = ~w40643 & w40797;
assign w41048 = ~w40616 & w40787;
assign w41049 = ~w40617 & w40682;
assign w41050 = w40677 & w41049;
assign w41051 = ~w40656 & ~w41047;
assign w41052 = ~w41048 & w41051;
assign w41053 = ~w41050 & w41052;
assign w41054 = w40674 & ~w41053;
assign w41055 = ~w41039 & ~w41046;
assign w41056 = ~w41054 & w41055;
assign w41057 = ~pi2088 & w41056;
assign w41058 = pi2088 & ~w41056;
assign w41059 = ~w41057 & ~w41058;
assign w41060 = ~w40966 & ~w41000;
assign w41061 = w40982 & ~w41060;
assign w41062 = w40984 & w41023;
assign w41063 = w40965 & w40972;
assign w41064 = w40985 & w41063;
assign w41065 = ~w41062 & ~w41064;
assign w41066 = ~w40994 & ~w41065;
assign w41067 = ~w40952 & w40984;
assign w41068 = w40989 & w41067;
assign w41069 = ~w40958 & w40965;
assign w41070 = w40965 & w40982;
assign w41071 = w40952 & ~w41070;
assign w41072 = w41069 & w41071;
assign w41073 = ~w40972 & w41072;
assign w41074 = w40989 & ~w40996;
assign w41075 = w40958 & ~w40982;
assign w41076 = w41026 & w41075;
assign w41077 = ~w41074 & ~w41076;
assign w41078 = ~w41073 & ~w41077;
assign w41079 = w40982 & ~w41015;
assign w41080 = ~w41018 & ~w41030;
assign w41081 = w41079 & w41080;
assign w41082 = w41010 & ~w41081;
assign w41083 = ~w41078 & w41082;
assign w41084 = ~w41013 & ~w41069;
assign w41085 = ~w40972 & ~w41084;
assign w41086 = ~w41063 & w41084;
assign w41087 = w40982 & ~w41086;
assign w41088 = ~w40982 & w41084;
assign w41089 = ~w41085 & ~w41088;
assign w41090 = ~w41087 & w41089;
assign w41091 = w40993 & w41065;
assign w41092 = ~w41090 & w41091;
assign w41093 = ~w41010 & ~w41092;
assign w41094 = ~w41061 & ~w41068;
assign w41095 = ~w41066 & w41094;
assign w41096 = ~w41083 & w41095;
assign w41097 = ~w41093 & w41096;
assign w41098 = ~pi2104 & ~w41097;
assign w41099 = pi2104 & w41097;
assign w41100 = ~w41098 & ~w41099;
assign w41101 = ~w40829 & w40893;
assign w41102 = w40845 & w66382;
assign w41103 = (w40864 & w40933) | (w40864 & w66383) | (w40933 & w66383);
assign w41104 = w40871 & w40892;
assign w41105 = ~w40910 & ~w41104;
assign w41106 = ~w41102 & w41105;
assign w41107 = ~w41103 & w41106;
assign w41108 = w40882 & ~w41107;
assign w41109 = ~w40908 & w40909;
assign w41110 = ~w40836 & ~w40855;
assign w41111 = w40908 & ~w40909;
assign w41112 = w40859 & ~w40866;
assign w41113 = ~w41111 & ~w41112;
assign w41114 = ~w41110 & ~w41113;
assign w41115 = w40871 & w40873;
assign w41116 = ~w40872 & ~w41115;
assign w41117 = ~w41109 & w41116;
assign w41118 = ~w40891 & w41117;
assign w41119 = ~w41114 & w41118;
assign w41120 = ~w40882 & ~w41119;
assign w41121 = ~w41102 & ~w41115;
assign w41122 = ~w40855 & ~w41121;
assign w41123 = ~w40876 & ~w41101;
assign w41124 = ~w41122 & w41123;
assign w41125 = ~w41120 & w41124;
assign w41126 = w41125 & w66384;
assign w41127 = (~pi2085 & ~w41125) | (~pi2085 & w66385) | (~w41125 & w66385);
assign w41128 = ~w41126 & ~w41127;
assign w41129 = ~pi7219 & pi9040;
assign w41130 = ~pi7226 & ~pi9040;
assign w41131 = ~w41129 & ~w41130;
assign w41132 = pi2242 & ~w41131;
assign w41133 = ~pi2242 & w41131;
assign w41134 = ~w41132 & ~w41133;
assign w41135 = ~pi7193 & pi9040;
assign w41136 = ~pi7187 & ~pi9040;
assign w41137 = ~w41135 & ~w41136;
assign w41138 = pi2185 & ~w41137;
assign w41139 = ~pi2185 & w41137;
assign w41140 = ~w41138 & ~w41139;
assign w41141 = w41134 & w41140;
assign w41142 = ~pi7180 & pi9040;
assign w41143 = ~pi7198 & ~pi9040;
assign w41144 = ~w41142 & ~w41143;
assign w41145 = pi2164 & ~w41144;
assign w41146 = ~pi2164 & w41144;
assign w41147 = ~w41145 & ~w41146;
assign w41148 = ~pi7191 & pi9040;
assign w41149 = ~pi7242 & ~pi9040;
assign w41150 = ~w41148 & ~w41149;
assign w41151 = pi2174 & ~w41150;
assign w41152 = ~pi2174 & w41150;
assign w41153 = ~w41151 & ~w41152;
assign w41154 = ~w41147 & w41153;
assign w41155 = w41141 & w41154;
assign w41156 = w41134 & ~w41153;
assign w41157 = ~w41140 & ~w41147;
assign w41158 = w41156 & w41157;
assign w41159 = ~w41155 & ~w41158;
assign w41160 = ~pi7211 & pi9040;
assign w41161 = ~pi7188 & ~pi9040;
assign w41162 = ~w41160 & ~w41161;
assign w41163 = pi2178 & ~w41162;
assign w41164 = ~pi2178 & w41162;
assign w41165 = ~w41163 & ~w41164;
assign w41166 = w41134 & ~w41140;
assign w41167 = w41147 & ~w41153;
assign w41168 = w41166 & w41167;
assign w41169 = w41165 & ~w41168;
assign w41170 = w41140 & ~w41167;
assign w41171 = ~w41156 & w41170;
assign w41172 = ~w41140 & w41147;
assign w41173 = ~w41153 & w41172;
assign w41174 = ~w41171 & ~w41173;
assign w41175 = ~w41169 & ~w41174;
assign w41176 = w41159 & ~w41175;
assign w41177 = ~pi7215 & pi9040;
assign w41178 = ~pi7183 & ~pi9040;
assign w41179 = ~w41177 & ~w41178;
assign w41180 = pi2244 & ~w41179;
assign w41181 = ~pi2244 & w41179;
assign w41182 = ~w41180 & ~w41181;
assign w41183 = ~w41176 & ~w41182;
assign w41184 = w41153 & w41182;
assign w41185 = w41140 & w41147;
assign w41186 = w41184 & w41185;
assign w41187 = w41153 & w41157;
assign w41188 = ~w41134 & w41187;
assign w41189 = w41182 & ~w41188;
assign w41190 = ~w41147 & ~w41153;
assign w41191 = w41140 & w41190;
assign w41192 = ~w41187 & ~w41191;
assign w41193 = w41189 & ~w41192;
assign w41194 = ~w41167 & ~w41182;
assign w41195 = ~w41134 & w41140;
assign w41196 = ~w41194 & w41195;
assign w41197 = w41134 & ~w41147;
assign w41198 = ~w41140 & ~w41197;
assign w41199 = w41194 & w41198;
assign w41200 = w41169 & ~w41186;
assign w41201 = ~w41196 & ~w41199;
assign w41202 = w41200 & w41201;
assign w41203 = ~w41193 & w41202;
assign w41204 = ~w41167 & w41182;
assign w41205 = w41198 & w41204;
assign w41206 = w41141 & w41147;
assign w41207 = ~w41153 & w41206;
assign w41208 = w41159 & ~w41165;
assign w41209 = ~w41205 & ~w41207;
assign w41210 = w41208 & w41209;
assign w41211 = ~w41203 & ~w41210;
assign w41212 = ~w41183 & ~w41211;
assign w41213 = ~pi2086 & w41212;
assign w41214 = pi2086 & ~w41212;
assign w41215 = ~w41213 & ~w41214;
assign w41216 = ~w40643 & ~w41048;
assign w41217 = ~w40623 & w40806;
assign w41218 = ~w40649 & ~w40674;
assign w41219 = ~w40661 & w40790;
assign w41220 = ~w41217 & w41219;
assign w41221 = (~w41216 & ~w41220) | (~w41216 & w66386) | (~w41220 & w66386);
assign w41222 = w40623 & w40796;
assign w41223 = w40643 & ~w41041;
assign w41224 = ~w40623 & w40661;
assign w41225 = ~w40789 & ~w41222;
assign w41226 = ~w41224 & w41225;
assign w41227 = ~w41223 & w41226;
assign w41228 = w40674 & ~w41227;
assign w41229 = w40616 & ~w40789;
assign w41230 = w40800 & w41229;
assign w41231 = ~w40634 & ~w41230;
assign w41232 = ~w40791 & w41231;
assign w41233 = ~w40674 & ~w41232;
assign w41234 = ~w41221 & ~w41228;
assign w41235 = ~w41233 & w41234;
assign w41236 = ~pi2087 & w41235;
assign w41237 = pi2087 & ~w41235;
assign w41238 = ~w41236 & ~w41237;
assign w41239 = w41084 & w66387;
assign w41240 = ~w40997 & ~w41239;
assign w41241 = w41088 & w41240;
assign w41242 = ~w41003 & w41087;
assign w41243 = w40959 & w40972;
assign w41244 = ~w41030 & ~w41072;
assign w41245 = ~w41072 & w66388;
assign w41246 = w41027 & ~w41071;
assign w41247 = w41010 & ~w41243;
assign w41248 = ~w41246 & w41247;
assign w41249 = ~w41245 & w41248;
assign w41250 = (~w40982 & w41022) | (~w40982 & w66389) | (w41022 & w66389);
assign w41251 = ~w41010 & w41244;
assign w41252 = ~w41250 & w41251;
assign w41253 = ~w41249 & ~w41252;
assign w41254 = w41012 & ~w41240;
assign w41255 = ~w41241 & ~w41254;
assign w41256 = ~w41253 & w66390;
assign w41257 = pi2095 & w41256;
assign w41258 = ~pi2095 & ~w41256;
assign w41259 = ~w41257 & ~w41258;
assign w41260 = ~w41134 & w41153;
assign w41261 = w41140 & w41260;
assign w41262 = ~w41158 & ~w41261;
assign w41263 = w41182 & ~w41262;
assign w41264 = ~w41154 & ~w41173;
assign w41265 = ~w41153 & ~w41182;
assign w41266 = w41134 & ~w41265;
assign w41267 = ~w41264 & ~w41266;
assign w41268 = ~w41172 & ~w41182;
assign w41269 = w41134 & w41268;
assign w41270 = ~w41170 & w41269;
assign w41271 = ~w41207 & ~w41269;
assign w41272 = ~w41270 & ~w41271;
assign w41273 = ~w41165 & ~w41267;
assign w41274 = ~w41272 & w41273;
assign w41275 = ~w41134 & w41147;
assign w41276 = ~w41191 & ~w41275;
assign w41277 = w41171 & ~w41276;
assign w41278 = ~w41166 & w41184;
assign w41279 = w41157 & w41265;
assign w41280 = w41165 & ~w41278;
assign w41281 = ~w41279 & w41280;
assign w41282 = ~w41270 & w41281;
assign w41283 = ~w41277 & w41282;
assign w41284 = ~w41274 & ~w41283;
assign w41285 = ~w41166 & ~w41190;
assign w41286 = ~w41197 & ~w41285;
assign w41287 = w41265 & ~w41286;
assign w41288 = ~w41265 & w41286;
assign w41289 = ~w41287 & ~w41288;
assign w41290 = ~w41140 & ~w41184;
assign w41291 = w41165 & ~w41290;
assign w41292 = ~w41156 & ~w41260;
assign w41293 = w41147 & w41292;
assign w41294 = ~w41291 & w41293;
assign w41295 = ~w41289 & w41294;
assign w41296 = ~w41263 & ~w41295;
assign w41297 = ~w41284 & w41296;
assign w41298 = pi2084 & ~w41297;
assign w41299 = ~pi2084 & w41297;
assign w41300 = ~w41298 & ~w41299;
assign w41301 = w40889 & w40928;
assign w41302 = ~w40830 & w40864;
assign w41303 = w40856 & ~w40912;
assign w41304 = ~w41110 & ~w41302;
assign w41305 = ~w41303 & w41304;
assign w41306 = ~w40888 & ~w41112;
assign w41307 = ~w41305 & w41306;
assign w41308 = ~w40882 & ~w41307;
assign w41309 = ~w40864 & ~w40882;
assign w41310 = w40890 & ~w41309;
assign w41311 = ~w40863 & ~w40931;
assign w41312 = w40882 & ~w41311;
assign w41313 = ~w40872 & ~w41102;
assign w41314 = ~w41312 & w41313;
assign w41315 = w40855 & ~w41314;
assign w41316 = ~w41301 & ~w41310;
assign w41317 = ~w41315 & w41316;
assign w41318 = ~w41308 & w41317;
assign w41319 = pi2097 & ~w41318;
assign w41320 = ~pi2097 & w41318;
assign w41321 = ~w41319 & ~w41320;
assign w41322 = ~pi7184 & pi9040;
assign w41323 = ~pi7201 & ~pi9040;
assign w41324 = ~w41322 & ~w41323;
assign w41325 = pi2224 & ~w41324;
assign w41326 = ~pi2224 & w41324;
assign w41327 = ~w41325 & ~w41326;
assign w41328 = ~pi7192 & pi9040;
assign w41329 = ~pi7220 & ~pi9040;
assign w41330 = ~w41328 & ~w41329;
assign w41331 = pi2212 & ~w41330;
assign w41332 = ~pi2212 & w41330;
assign w41333 = ~w41331 & ~w41332;
assign w41334 = ~w41327 & w41333;
assign w41335 = ~pi7223 & pi9040;
assign w41336 = ~pi7206 & ~pi9040;
assign w41337 = ~w41335 & ~w41336;
assign w41338 = pi2184 & ~w41337;
assign w41339 = ~pi2184 & w41337;
assign w41340 = ~w41338 & ~w41339;
assign w41341 = ~pi7182 & pi9040;
assign w41342 = ~pi7196 & ~pi9040;
assign w41343 = ~w41341 & ~w41342;
assign w41344 = pi2176 & ~w41343;
assign w41345 = ~pi2176 & w41343;
assign w41346 = ~w41344 & ~w41345;
assign w41347 = ~w41340 & ~w41346;
assign w41348 = w41334 & w41347;
assign w41349 = ~pi7225 & pi9040;
assign w41350 = ~pi7190 & ~pi9040;
assign w41351 = ~w41349 & ~w41350;
assign w41352 = pi2218 & ~w41351;
assign w41353 = ~pi2218 & w41351;
assign w41354 = ~w41352 & ~w41353;
assign w41355 = ~w41348 & w41354;
assign w41356 = w41340 & w41346;
assign w41357 = ~w41347 & ~w41356;
assign w41358 = w41334 & w41357;
assign w41359 = ~w41347 & ~w41358;
assign w41360 = w41355 & ~w41359;
assign w41361 = ~w41327 & w41346;
assign w41362 = w41327 & ~w41346;
assign w41363 = ~w41361 & ~w41362;
assign w41364 = ~w41333 & w41363;
assign w41365 = w41363 & w66391;
assign w41366 = ~w41327 & w41340;
assign w41367 = ~w41333 & ~w41340;
assign w41368 = w41327 & w41367;
assign w41369 = w41346 & w41368;
assign w41370 = ~w41366 & ~w41369;
assign w41371 = w41357 & ~w41361;
assign w41372 = ~w41362 & ~w41367;
assign w41373 = (~w41354 & ~w41371) | (~w41354 & w63979) | (~w41371 & w63979);
assign w41374 = ~w41370 & w41373;
assign w41375 = w41327 & w41354;
assign w41376 = (~w41375 & ~w41357) | (~w41375 & w66392) | (~w41357 & w66392);
assign w41377 = w41333 & ~w41340;
assign w41378 = ~w41333 & w41356;
assign w41379 = ~w41377 & ~w41378;
assign w41380 = ~w41376 & ~w41379;
assign w41381 = ~pi7179 & pi9040;
assign w41382 = ~pi7222 & ~pi9040;
assign w41383 = ~w41381 & ~w41382;
assign w41384 = pi2159 & ~w41383;
assign w41385 = ~pi2159 & w41383;
assign w41386 = ~w41384 & ~w41385;
assign w41387 = ~w41365 & w41386;
assign w41388 = ~w41380 & w41387;
assign w41389 = ~w41374 & w41388;
assign w41390 = w41346 & ~w41354;
assign w41391 = w41368 & ~w41390;
assign w41392 = w41340 & w41362;
assign w41393 = ~w41348 & ~w41392;
assign w41394 = ~w41354 & ~w41393;
assign w41395 = ~w41386 & ~w41391;
assign w41396 = ~w41394 & w41395;
assign w41397 = ~w41389 & ~w41396;
assign w41398 = w41327 & ~w41333;
assign w41399 = w41340 & ~w41354;
assign w41400 = ~w41356 & ~w41390;
assign w41401 = ~w41386 & ~w41400;
assign w41402 = ~w41399 & ~w41401;
assign w41403 = ~w41334 & ~w41398;
assign w41404 = ~w41402 & w41403;
assign w41405 = ~w41360 & ~w41404;
assign w41406 = ~w41397 & w41405;
assign w41407 = pi2094 & ~w41406;
assign w41408 = ~pi2094 & w41406;
assign w41409 = ~w41407 & ~w41408;
assign w41410 = ~w40751 & ~w40765;
assign w41411 = w40712 & w40775;
assign w41412 = ~w40737 & ~w40747;
assign w41413 = (w40706 & ~w41412) | (w40706 & w66393) | (~w41412 & w66393);
assign w41414 = w40719 & w40725;
assign w41415 = ~w40764 & ~w41414;
assign w41416 = w40712 & w41415;
assign w41417 = w41413 & w41416;
assign w41418 = ~w40771 & w41410;
assign w41419 = ~w41417 & w41418;
assign w41420 = w40759 & ~w41419;
assign w41421 = ~w40719 & ~w40774;
assign w41422 = ~w40761 & w41415;
assign w41423 = ~w40748 & ~w41421;
assign w41424 = w41422 & w41423;
assign w41425 = w40706 & ~w40774;
assign w41426 = ~w41411 & w41425;
assign w41427 = w40772 & w41426;
assign w41428 = (~w40759 & w41424) | (~w40759 & w63980) | (w41424 & w63980);
assign w41429 = (w40759 & ~w41415) | (w40759 & w66394) | (~w41415 & w66394);
assign w41430 = ~w40773 & ~w41429;
assign w41431 = ~w40706 & ~w41430;
assign w41432 = w40706 & ~w40712;
assign w41433 = w40741 & w41432;
assign w41434 = ~w40780 & ~w41433;
assign w41435 = ~w41428 & w41434;
assign w41436 = ~w41431 & w41435;
assign w41437 = (pi2101 & ~w41436) | (pi2101 & w66395) | (~w41436 & w66395);
assign w41438 = w41436 & w66396;
assign w41439 = ~w41437 & ~w41438;
assign w41440 = w40952 & w41015;
assign w41441 = w40973 & ~w41071;
assign w41442 = ~w40982 & w40991;
assign w41443 = ~w41062 & ~w41442;
assign w41444 = ~w40987 & w41443;
assign w41445 = ~w41440 & ~w41441;
assign w41446 = w41444 & w41445;
assign w41447 = w41010 & ~w41446;
assign w41448 = w41021 & w41063;
assign w41449 = w40965 & ~w40973;
assign w41450 = ~w40999 & ~w41449;
assign w41451 = w41012 & ~w41450;
assign w41452 = ~w40996 & ~w41067;
assign w41453 = w41025 & ~w41452;
assign w41454 = ~w41073 & ~w41448;
assign w41455 = ~w41451 & ~w41453;
assign w41456 = w41454 & w41455;
assign w41457 = ~w41066 & w41456;
assign w41458 = ~w41447 & w41457;
assign w41459 = ~pi2090 & ~w41458;
assign w41460 = pi2090 & w41458;
assign w41461 = ~w41459 & ~w41460;
assign w41462 = w40732 & w40753;
assign w41463 = w40706 & w40761;
assign w41464 = ~w40759 & ~w41463;
assign w41465 = w40725 & w40779;
assign w41466 = w40731 & w40737;
assign w41467 = ~w40746 & ~w41466;
assign w41468 = w40706 & ~w40718;
assign w41469 = ~w40776 & ~w41468;
assign w41470 = ~w41467 & ~w41469;
assign w41471 = ~w40764 & ~w40771;
assign w41472 = (w40706 & ~w41471) | (w40706 & w66397) | (~w41471 & w66397);
assign w41473 = ~w41465 & ~w41470;
assign w41474 = (~w41464 & ~w41473) | (~w41464 & w66398) | (~w41473 & w66398);
assign w41475 = ~w40706 & ~w41421;
assign w41476 = ~w41421 & w66399;
assign w41477 = ~w40750 & ~w41414;
assign w41478 = w40706 & ~w41477;
assign w41479 = (~w40718 & w40773) | (~w40718 & w66400) | (w40773 & w66400);
assign w41480 = w40718 & w40732;
assign w41481 = ~w41432 & w41480;
assign w41482 = w41410 & ~w41481;
assign w41483 = ~w41476 & ~w41478;
assign w41484 = w41482 & w41483;
assign w41485 = (~w40759 & ~w41484) | (~w40759 & w66401) | (~w41484 & w66401);
assign w41486 = ~w41462 & ~w41474;
assign w41487 = ~w41485 & w41486;
assign w41488 = pi2098 & w41487;
assign w41489 = ~pi2098 & ~w41487;
assign w41490 = ~w41488 & ~w41489;
assign w41491 = ~pi7183 & pi9040;
assign w41492 = ~pi7207 & ~pi9040;
assign w41493 = ~w41491 & ~w41492;
assign w41494 = pi2174 & ~w41493;
assign w41495 = ~pi2174 & w41493;
assign w41496 = ~w41494 & ~w41495;
assign w41497 = ~pi7238 & pi9040;
assign w41498 = ~pi7243 & ~pi9040;
assign w41499 = ~w41497 & ~w41498;
assign w41500 = pi2192 & ~w41499;
assign w41501 = ~pi2192 & w41499;
assign w41502 = ~w41500 & ~w41501;
assign w41503 = ~pi7212 & pi9040;
assign w41504 = ~pi7180 & ~pi9040;
assign w41505 = ~w41503 & ~w41504;
assign w41506 = pi2183 & ~w41505;
assign w41507 = ~pi2183 & w41505;
assign w41508 = ~w41506 & ~w41507;
assign w41509 = ~w41502 & ~w41508;
assign w41510 = ~pi7226 & pi9040;
assign w41511 = ~pi7221 & ~pi9040;
assign w41512 = ~w41510 & ~w41511;
assign w41513 = pi2221 & ~w41512;
assign w41514 = ~pi2221 & w41512;
assign w41515 = ~w41513 & ~w41514;
assign w41516 = ~w41509 & ~w41515;
assign w41517 = ~w41508 & w41515;
assign w41518 = ~w41516 & ~w41517;
assign w41519 = w41496 & ~w41502;
assign w41520 = ~w41516 & ~w41519;
assign w41521 = ~w41518 & ~w41520;
assign w41522 = ~w41496 & w41502;
assign w41523 = ~w41519 & ~w41522;
assign w41524 = ~w41515 & ~w41523;
assign w41525 = ~w41496 & w41515;
assign w41526 = ~w41502 & w41508;
assign w41527 = w41525 & w41526;
assign w41528 = ~w41524 & ~w41527;
assign w41529 = ~pi7205 & pi9040;
assign w41530 = ~pi7181 & ~pi9040;
assign w41531 = ~w41529 & ~w41530;
assign w41532 = pi2215 & ~w41531;
assign w41533 = ~pi2215 & w41531;
assign w41534 = ~w41532 & ~w41533;
assign w41535 = ~w41519 & ~w41534;
assign w41536 = w41521 & ~w41535;
assign w41537 = w41536 & w66402;
assign w41538 = ~pi7208 & pi9040;
assign w41539 = ~pi7191 & ~pi9040;
assign w41540 = ~w41538 & ~w41539;
assign w41541 = pi2185 & ~w41540;
assign w41542 = ~pi2185 & w41540;
assign w41543 = ~w41541 & ~w41542;
assign w41544 = w41502 & w41534;
assign w41545 = w41496 & ~w41515;
assign w41546 = ~w41525 & ~w41545;
assign w41547 = w41508 & ~w41546;
assign w41548 = ~w41546 & w66403;
assign w41549 = w41515 & w41534;
assign w41550 = w41523 & ~w41549;
assign w41551 = ~w41508 & w41546;
assign w41552 = ~w41550 & w41551;
assign w41553 = (~w41543 & w41552) | (~w41543 & w66404) | (w41552 & w66404);
assign w41554 = ~w41508 & ~w41515;
assign w41555 = ~w41519 & w41554;
assign w41556 = ~w41527 & ~w41555;
assign w41557 = ~w41508 & w41522;
assign w41558 = w41515 & w41523;
assign w41559 = ~w41524 & ~w41558;
assign w41560 = w41496 & w41508;
assign w41561 = ~w41559 & w41560;
assign w41562 = (~w41557 & w41556) | (~w41557 & w66405) | (w41556 & w66405);
assign w41563 = (~w41534 & w41561) | (~w41534 & w66406) | (w41561 & w66406);
assign w41564 = w41509 & w41549;
assign w41565 = w41509 & w41525;
assign w41566 = ~w41508 & w41534;
assign w41567 = w41496 & w41566;
assign w41568 = ~w41526 & ~w41567;
assign w41569 = ~w41515 & ~w41568;
assign w41570 = w41515 & ~w41534;
assign w41571 = w41519 & ~w41570;
assign w41572 = ~w41496 & ~w41515;
assign w41573 = w41508 & w41534;
assign w41574 = w41572 & w41573;
assign w41575 = w41502 & w41570;
assign w41576 = ~w41565 & ~w41571;
assign w41577 = ~w41574 & ~w41575;
assign w41578 = w41576 & w41577;
assign w41579 = ~w41569 & w41578;
assign w41580 = w41543 & ~w41579;
assign w41581 = ~w41553 & ~w41564;
assign w41582 = ~w41580 & w41581;
assign w41583 = ~w41537 & ~w41563;
assign w41584 = w41582 & w41583;
assign w41585 = pi2092 & w41584;
assign w41586 = ~pi2092 & ~w41584;
assign w41587 = ~w41585 & ~w41586;
assign w41588 = w41154 & ~w41195;
assign w41589 = ~w41277 & w66407;
assign w41590 = ~w41182 & ~w41589;
assign w41591 = ~w41140 & ~w41265;
assign w41592 = w41275 & w41591;
assign w41593 = ~w41172 & w41182;
assign w41594 = ~w41277 & w66408;
assign w41595 = ~w41165 & ~w41592;
assign w41596 = ~w41594 & w41595;
assign w41597 = ~w41590 & w41596;
assign w41598 = ~w41166 & w41588;
assign w41599 = w41147 & w41261;
assign w41600 = w41165 & ~w41598;
assign w41601 = ~w41599 & w41600;
assign w41602 = w41289 & w41601;
assign w41603 = ~w41597 & ~w41602;
assign w41604 = pi2096 & w41603;
assign w41605 = ~pi2096 & ~w41603;
assign w41606 = ~w41604 & ~w41605;
assign w41607 = ~pi7207 & pi9040;
assign w41608 = ~pi7193 & ~pi9040;
assign w41609 = ~w41607 & ~w41608;
assign w41610 = pi2209 & ~w41609;
assign w41611 = ~pi2209 & w41609;
assign w41612 = ~w41610 & ~w41611;
assign w41613 = ~pi7227 & pi9040;
assign w41614 = ~pi7199 & ~pi9040;
assign w41615 = ~w41613 & ~w41614;
assign w41616 = pi2182 & ~w41615;
assign w41617 = ~pi2182 & w41615;
assign w41618 = ~w41616 & ~w41617;
assign w41619 = ~pi7203 & pi9040;
assign w41620 = ~pi7214 & ~pi9040;
assign w41621 = ~w41619 & ~w41620;
assign w41622 = pi2164 & ~w41621;
assign w41623 = ~pi2164 & w41621;
assign w41624 = ~w41622 & ~w41623;
assign w41625 = w41618 & ~w41624;
assign w41626 = ~pi7210 & pi9040;
assign w41627 = ~pi7212 & ~pi9040;
assign w41628 = ~w41626 & ~w41627;
assign w41629 = pi2210 & ~w41628;
assign w41630 = ~pi2210 & w41628;
assign w41631 = ~w41629 & ~w41630;
assign w41632 = ~pi7181 & pi9040;
assign w41633 = ~pi7245 & ~pi9040;
assign w41634 = ~w41632 & ~w41633;
assign w41635 = pi2178 & ~w41634;
assign w41636 = ~pi2178 & w41634;
assign w41637 = ~w41635 & ~w41636;
assign w41638 = ~w41618 & ~w41637;
assign w41639 = ~w41624 & ~w41631;
assign w41640 = w41638 & w41639;
assign w41641 = ~pi7217 & pi9040;
assign w41642 = ~pi7194 & ~pi9040;
assign w41643 = ~w41641 & ~w41642;
assign w41644 = pi2199 & ~w41643;
assign w41645 = ~pi2199 & w41643;
assign w41646 = ~w41644 & ~w41645;
assign w41647 = ~w41640 & ~w41646;
assign w41648 = ~w41631 & w41647;
assign w41649 = w41625 & ~w41648;
assign w41650 = ~w41631 & ~w41637;
assign w41651 = w41618 & w41650;
assign w41652 = w41618 & w41637;
assign w41653 = w41631 & ~w41637;
assign w41654 = ~w41618 & w41624;
assign w41655 = ~w41625 & ~w41638;
assign w41656 = ~w41653 & ~w41654;
assign w41657 = w41655 & w41656;
assign w41658 = ~w41652 & w41657;
assign w41659 = ~w41638 & ~w41652;
assign w41660 = ~w41639 & ~w41659;
assign w41661 = ~w41651 & ~w41660;
assign w41662 = ~w41658 & w41661;
assign w41663 = ~w41647 & w41662;
assign w41664 = (w41612 & w41663) | (w41612 & w66409) | (w41663 & w66409);
assign w41665 = w41624 & w41631;
assign w41666 = ~w41639 & ~w41665;
assign w41667 = ~w41659 & w41666;
assign w41668 = ~w41631 & w41637;
assign w41669 = w41612 & ~w41668;
assign w41670 = w41639 & w41659;
assign w41671 = ~w41669 & w41670;
assign w41672 = ~w41652 & w41665;
assign w41673 = ~w41618 & ~w41650;
assign w41674 = ~w41612 & ~w41673;
assign w41675 = w41672 & w41674;
assign w41676 = w41631 & w41637;
assign w41677 = w41654 & w41676;
assign w41678 = w41612 & w41624;
assign w41679 = w41650 & w41678;
assign w41680 = ~w41677 & ~w41679;
assign w41681 = ~w41667 & w41680;
assign w41682 = ~w41671 & w41681;
assign w41683 = ~w41675 & w41682;
assign w41684 = (~w41646 & ~w41682) | (~w41646 & w66410) | (~w41682 & w66410);
assign w41685 = ~w41612 & w41657;
assign w41686 = w41631 & w41638;
assign w41687 = w41624 & w41686;
assign w41688 = ~w41685 & ~w41687;
assign w41689 = w41646 & ~w41688;
assign w41690 = ~w41684 & ~w41689;
assign w41691 = ~w41664 & w41690;
assign w41692 = pi2105 & w41691;
assign w41693 = ~pi2105 & ~w41691;
assign w41694 = ~w41692 & ~w41693;
assign w41695 = ~w41654 & ~w41676;
assign w41696 = ~w41672 & ~w41695;
assign w41697 = w41612 & ~w41696;
assign w41698 = ~w41657 & w41697;
assign w41699 = ~w41612 & ~w41624;
assign w41700 = w41676 & w41699;
assign w41701 = w41624 & w41659;
assign w41702 = w41625 & w41637;
assign w41703 = ~w41701 & ~w41702;
assign w41704 = w41638 & ~w41678;
assign w41705 = ~w41631 & ~w41704;
assign w41706 = ~w41612 & ~w41618;
assign w41707 = w41659 & w66411;
assign w41708 = ~w41706 & ~w41707;
assign w41709 = ~w41650 & ~w41676;
assign w41710 = ~w41708 & w41709;
assign w41711 = (w41646 & ~w41703) | (w41646 & w66412) | (~w41703 & w66412);
assign w41712 = ~w41710 & w41711;
assign w41713 = (w41612 & w41701) | (w41612 & w66413) | (w41701 & w66413);
assign w41714 = w41674 & w41703;
assign w41715 = w41647 & ~w41713;
assign w41716 = ~w41714 & w41715;
assign w41717 = ~w41712 & ~w41716;
assign w41718 = (~w41700 & w41683) | (~w41700 & w66414) | (w41683 & w66414);
assign w41719 = ~w41717 & w41718;
assign w41720 = pi2125 & ~w41719;
assign w41721 = ~pi2125 & w41719;
assign w41722 = ~w41720 & ~w41721;
assign w41723 = w41544 & ~w41579;
assign w41724 = w41502 & ~w41554;
assign w41725 = ~w41534 & w41546;
assign w41726 = ~w41724 & w41725;
assign w41727 = ~w41523 & ~w41547;
assign w41728 = ~w41550 & ~w41727;
assign w41729 = ~w41543 & ~w41726;
assign w41730 = ~w41728 & w41729;
assign w41731 = w41502 & w41560;
assign w41732 = w41543 & ~w41731;
assign w41733 = w41517 & w41522;
assign w41734 = w41521 & w41534;
assign w41735 = w41518 & ~w41534;
assign w41736 = w41732 & ~w41733;
assign w41737 = ~w41735 & w41736;
assign w41738 = ~w41734 & w41737;
assign w41739 = ~w41730 & ~w41738;
assign w41740 = ~w41723 & ~w41739;
assign w41741 = ~pi2112 & w41740;
assign w41742 = pi2112 & ~w41740;
assign w41743 = ~w41741 & ~w41742;
assign w41744 = w40748 & ~w40765;
assign w41745 = ~w40725 & ~w40744;
assign w41746 = ~w41475 & w41745;
assign w41747 = ~w40731 & w40759;
assign w41748 = w40749 & ~w41747;
assign w41749 = ~w41746 & ~w41748;
assign w41750 = ~w41479 & w41749;
assign w41751 = ~w40778 & ~w41744;
assign w41752 = ~w41750 & w41751;
assign w41753 = w40746 & w41468;
assign w41754 = ~w40744 & ~w40749;
assign w41755 = w40774 & ~w41754;
assign w41756 = ~w40732 & ~w40742;
assign w41757 = w40712 & ~w41756;
assign w41758 = w40759 & ~w41753;
assign w41759 = ~w41755 & w41758;
assign w41760 = ~w41757 & w41759;
assign w41761 = w40749 & w40775;
assign w41762 = ~w40759 & ~w41761;
assign w41763 = ~w41413 & w41762;
assign w41764 = ~w41760 & ~w41763;
assign w41765 = ~w41752 & ~w41764;
assign w41766 = ~pi2103 & w41765;
assign w41767 = pi2103 & ~w41765;
assign w41768 = ~w41766 & ~w41767;
assign w41769 = w41508 & ~w41559;
assign w41770 = w41502 & ~w41545;
assign w41771 = ~w41519 & w41566;
assign w41772 = ~w41770 & w41771;
assign w41773 = ~w41733 & ~w41772;
assign w41774 = ~w41769 & w41773;
assign w41775 = w41543 & ~w41774;
assign w41776 = w41502 & ~w41517;
assign w41777 = ~w41509 & w41546;
assign w41778 = ~w41776 & w41777;
assign w41779 = w41544 & w41572;
assign w41780 = w41535 & ~w41770;
assign w41781 = ~w41523 & ~w41557;
assign w41782 = w41534 & ~w41543;
assign w41783 = w41781 & w41782;
assign w41784 = ~w41779 & ~w41780;
assign w41785 = ~w41778 & w41784;
assign w41786 = ~w41783 & w41785;
assign w41787 = ~w41575 & w41732;
assign w41788 = ~w41786 & ~w41787;
assign w41789 = ~w41775 & ~w41788;
assign w41790 = ~pi2113 & w41789;
assign w41791 = pi2113 & ~w41789;
assign w41792 = ~w41790 & ~w41791;
assign w41793 = w41327 & w41333;
assign w41794 = w41357 & w63981;
assign w41795 = w41354 & ~w41794;
assign w41796 = w41793 & ~w41795;
assign w41797 = ~w41363 & w41367;
assign w41798 = (~w41361 & w41363) | (~w41361 & w66415) | (w41363 & w66415);
assign w41799 = w41400 & ~w41798;
assign w41800 = w41361 & ~w41379;
assign w41801 = ~w41358 & w41366;
assign w41802 = ~w41800 & w41801;
assign w41803 = (~w41386 & w41355) | (~w41386 & w66416) | (w41355 & w66416);
assign w41804 = ~w41799 & w41803;
assign w41805 = ~w41802 & w41804;
assign w41806 = ~w41796 & w41805;
assign w41807 = w41354 & w41365;
assign w41808 = w41354 & ~w41378;
assign w41809 = w41800 & ~w41808;
assign w41810 = w41362 & w41377;
assign w41811 = w41340 & ~w41376;
assign w41812 = w41386 & ~w41810;
assign w41813 = ~w41369 & w41812;
assign w41814 = ~w41807 & w41813;
assign w41815 = ~w41809 & ~w41811;
assign w41816 = w41814 & w41815;
assign w41817 = ~w41806 & ~w41816;
assign w41818 = pi2119 & w41817;
assign w41819 = ~pi2119 & ~w41817;
assign w41820 = ~w41818 & ~w41819;
assign w41821 = w41658 & w41697;
assign w41822 = ~w41653 & w41666;
assign w41823 = ~w41651 & ~w41686;
assign w41824 = ~w41822 & w41823;
assign w41825 = (w41660 & w41824) | (w41660 & w66417) | (w41824 & w66417);
assign w41826 = ~w41646 & w41662;
assign w41827 = (~w41612 & w41826) | (~w41612 & w66418) | (w41826 & w66418);
assign w41828 = w41612 & w41824;
assign w41829 = (w41646 & w41828) | (w41646 & w63982) | (w41828 & w63982);
assign w41830 = w41669 & ~w41824;
assign w41831 = w41657 & w66419;
assign w41832 = (~w41646 & w41830) | (~w41646 & w66420) | (w41830 & w66420);
assign w41833 = ~w41821 & ~w41829;
assign w41834 = ~w41832 & w41833;
assign w41835 = (pi2127 & ~w41834) | (pi2127 & w66421) | (~w41834 & w66421);
assign w41836 = w41834 & w66422;
assign w41837 = ~w41835 & ~w41836;
assign w41838 = ~w41624 & w41662;
assign w41839 = ~w41612 & ~w41695;
assign w41840 = ~w41637 & w41699;
assign w41841 = ~w41839 & ~w41840;
assign w41842 = ~w41697 & w41841;
assign w41843 = (~w41646 & w41838) | (~w41646 & w66423) | (w41838 & w66423);
assign w41844 = w41665 & w41706;
assign w41845 = ~w41824 & w66424;
assign w41846 = ~w41670 & w41823;
assign w41847 = w41612 & ~w41846;
assign w41848 = ~w41695 & w66425;
assign w41849 = ~w41672 & ~w41848;
assign w41850 = (w41646 & w41847) | (w41646 & w66426) | (w41847 & w66426);
assign w41851 = ~w41844 & ~w41845;
assign w41852 = ~w41850 & w41851;
assign w41853 = ~w41843 & w41852;
assign w41854 = pi2116 & ~w41853;
assign w41855 = ~pi2116 & w41853;
assign w41856 = ~w41854 & ~w41855;
assign w41857 = (~w41548 & ~w41536) | (~w41548 & w66427) | (~w41536 & w66427);
assign w41858 = w41543 & ~w41857;
assign w41859 = ~w41547 & w66428;
assign w41860 = (w41543 & w41524) | (w41543 & w66429) | (w41524 & w66429);
assign w41861 = ~w41859 & ~w41860;
assign w41862 = ~w41534 & ~w41861;
assign w41863 = ~w41496 & w41509;
assign w41864 = w41545 & w41573;
assign w41865 = ~w41575 & ~w41731;
assign w41866 = ~w41863 & ~w41864;
assign w41867 = w41865 & w41866;
assign w41868 = w41560 & w41570;
assign w41869 = ~w41779 & ~w41868;
assign w41870 = w41543 & w41781;
assign w41871 = ~w41869 & ~w41870;
assign w41872 = (~w41564 & w41867) | (~w41564 & w66430) | (w41867 & w66430);
assign w41873 = ~w41871 & w41872;
assign w41874 = ~w41862 & w41873;
assign w41875 = ~w41858 & w41874;
assign w41876 = ~pi2131 & w41875;
assign w41877 = pi2131 & ~w41875;
assign w41878 = ~w41876 & ~w41877;
assign w41879 = w41361 & w41377;
assign w41880 = w41354 & ~w41879;
assign w41881 = (~w41354 & ~w41366) | (~w41354 & w66431) | (~w41366 & w66431);
assign w41882 = w41327 & w41378;
assign w41883 = w41881 & ~w41882;
assign w41884 = ~w41880 & ~w41883;
assign w41885 = w41333 & w41392;
assign w41886 = ~w41346 & ~w41398;
assign w41887 = ~w41366 & w41886;
assign w41888 = w41808 & ~w41887;
assign w41889 = w41373 & ~w41797;
assign w41890 = w41386 & ~w41885;
assign w41891 = (w41890 & w41889) | (w41890 & w66432) | (w41889 & w66432);
assign w41892 = w41346 & ~w41793;
assign w41893 = w41340 & ~w41886;
assign w41894 = ~w41892 & w41893;
assign w41895 = ~w41357 & ~w41368;
assign w41896 = ~w41354 & ~w41895;
assign w41897 = ~w41333 & w41362;
assign w41898 = ~w41794 & w66433;
assign w41899 = ~w41896 & ~w41898;
assign w41900 = ~w41358 & ~w41386;
assign w41901 = ~w41894 & w41900;
assign w41902 = ~w41899 & w41901;
assign w41903 = ~w41891 & ~w41902;
assign w41904 = ~w41884 & ~w41903;
assign w41905 = ~pi2121 & w41904;
assign w41906 = pi2121 & ~w41904;
assign w41907 = ~w41905 & ~w41906;
assign w41908 = w41340 & ~w41363;
assign w41909 = ~w41794 & ~w41908;
assign w41910 = w41333 & ~w41909;
assign w41911 = w41363 & w66434;
assign w41912 = w41354 & ~w41911;
assign w41913 = ~w41372 & ~w41398;
assign w41914 = w41881 & ~w41908;
assign w41915 = ~w41913 & w41914;
assign w41916 = ~w41912 & ~w41915;
assign w41917 = (w41386 & w41916) | (w41386 & w66435) | (w41916 & w66435);
assign w41918 = ~w41364 & ~w41386;
assign w41919 = (w41355 & w41910) | (w41355 & w66436) | (w41910 & w66436);
assign w41920 = ~w41348 & ~w41911;
assign w41921 = ~w41386 & ~w41920;
assign w41922 = (~w41354 & w41909) | (~w41354 & w66431) | (w41909 & w66431);
assign w41923 = ~w41921 & w41922;
assign w41924 = ~w41919 & ~w41923;
assign w41925 = ~w41917 & ~w41924;
assign w41926 = ~pi2130 & w41925;
assign w41927 = pi2130 & ~w41925;
assign w41928 = ~w41926 & ~w41927;
assign w41929 = w41182 & ~w41264;
assign w41930 = w41268 & ~w41276;
assign w41931 = ~w41158 & ~w41929;
assign w41932 = ~w41930 & w41931;
assign w41933 = w41165 & ~w41932;
assign w41934 = ~w41190 & ~w41290;
assign w41935 = w41292 & ~w41934;
assign w41936 = ~w41155 & ~w41186;
assign w41937 = ~w41207 & w41936;
assign w41938 = ~w41935 & w41937;
assign w41939 = ~w41165 & ~w41938;
assign w41940 = w41189 & ~w41206;
assign w41941 = ~w41265 & ~w41268;
assign w41942 = ~w41940 & w41941;
assign w41943 = ~w41939 & ~w41942;
assign w41944 = ~w41933 & w41943;
assign w41945 = ~pi2126 & w41944;
assign w41946 = pi2126 & ~w41944;
assign w41947 = ~w41945 & ~w41946;
assign w41948 = ~pi4312 & pi9040;
assign w41949 = ~pi4440 & ~pi9040;
assign w41950 = ~w41948 & ~w41949;
assign w41951 = pi2261 & ~w41950;
assign w41952 = ~pi2261 & w41950;
assign w41953 = ~w41951 & ~w41952;
assign w41954 = ~pi4585 & pi9040;
assign w41955 = ~pi4657 & ~pi9040;
assign w41956 = ~w41954 & ~w41955;
assign w41957 = pi2262 & ~w41956;
assign w41958 = ~pi2262 & w41956;
assign w41959 = ~w41957 & ~w41958;
assign w41960 = w41953 & ~w41959;
assign w41961 = ~pi4601 & pi9040;
assign w41962 = ~pi4474 & ~pi9040;
assign w41963 = ~w41961 & ~w41962;
assign w41964 = pi2206 & ~w41963;
assign w41965 = ~pi2206 & w41963;
assign w41966 = ~w41964 & ~w41965;
assign w41967 = ~w41960 & w41966;
assign w41968 = ~pi4395 & pi9040;
assign w41969 = ~pi4386 & ~pi9040;
assign w41970 = ~w41968 & ~w41969;
assign w41971 = pi2264 & ~w41970;
assign w41972 = ~pi2264 & w41970;
assign w41973 = ~w41971 & ~w41972;
assign w41974 = w41959 & ~w41973;
assign w41975 = ~w41966 & ~w41974;
assign w41976 = ~w41967 & ~w41975;
assign w41977 = ~w41953 & w41959;
assign w41978 = ~w41959 & w41973;
assign w41979 = ~w41977 & ~w41978;
assign w41980 = w41976 & w41979;
assign w41981 = ~pi4323 & pi9040;
assign w41982 = ~pi4537 & ~pi9040;
assign w41983 = ~w41981 & ~w41982;
assign w41984 = pi2247 & ~w41983;
assign w41985 = ~pi2247 & w41983;
assign w41986 = ~w41984 & ~w41985;
assign w41987 = w41980 & w41986;
assign w41988 = w41959 & w41973;
assign w41989 = ~w41966 & w41973;
assign w41990 = w41966 & ~w41973;
assign w41991 = ~w41989 & ~w41990;
assign w41992 = (w41986 & w41991) | (w41986 & w63983) | (w41991 & w63983);
assign w41993 = (w41991 & w66437) | (w41991 & w66438) | (w66437 & w66438);
assign w41994 = ~w41953 & w41966;
assign w41995 = w41988 & w41994;
assign w41996 = w41960 & w41991;
assign w41997 = w41991 & w63984;
assign w41998 = ~w41995 & ~w41997;
assign w41999 = ~w41993 & w41998;
assign w42000 = w41998 & w66439;
assign w42001 = ~w41973 & w41994;
assign w42002 = w41959 & w41989;
assign w42003 = ~w42001 & ~w42002;
assign w42004 = ~w41977 & ~w42003;
assign w42005 = ~w41953 & ~w41959;
assign w42006 = w41989 & w42005;
assign w42007 = ~w41995 & ~w42006;
assign w42008 = ~w41976 & w42007;
assign w42009 = w41986 & ~w42008;
assign w42010 = ~w42004 & ~w42009;
assign w42011 = ~w41994 & ~w42005;
assign w42012 = ~w41973 & ~w42011;
assign w42013 = ~w42009 & w63985;
assign w42014 = ~w41978 & ~w41986;
assign w42015 = ~w41974 & ~w41977;
assign w42016 = ~w42001 & ~w42015;
assign w42017 = w42014 & ~w42016;
assign w42018 = w42008 & w42017;
assign w42019 = (~w42018 & w42013) | (~w42018 & w66440) | (w42013 & w66440);
assign w42020 = ~w41959 & w41966;
assign w42021 = w41973 & w42020;
assign w42022 = (~w41986 & w42016) | (~w41986 & w66441) | (w42016 & w66441);
assign w42023 = ~w42019 & ~w42022;
assign w42024 = ~pi4757 & pi9040;
assign w42025 = ~pi4407 & ~pi9040;
assign w42026 = ~w42024 & ~w42025;
assign w42027 = pi2227 & ~w42026;
assign w42028 = ~pi2227 & w42026;
assign w42029 = ~w42027 & ~w42028;
assign w42030 = ~w42023 & w42029;
assign w42031 = w42010 & ~w42018;
assign w42032 = ~w42029 & ~w42031;
assign w42033 = ~w41986 & w41991;
assign w42034 = w41973 & w42029;
assign w42035 = ~w42033 & ~w42034;
assign w42036 = w41953 & ~w41966;
assign w42037 = ~w41994 & ~w42036;
assign w42038 = ~w41959 & ~w42037;
assign w42039 = ~w42035 & w42038;
assign w42040 = ~w41987 & ~w42039;
assign w42041 = ~w42032 & w42040;
assign w42042 = ~w42030 & w42041;
assign w42043 = ~w41973 & w41977;
assign w42044 = ~w42021 & ~w42043;
assign w42045 = ~w41986 & ~w42044;
assign w42046 = ~w41966 & w42045;
assign w42047 = w41966 & ~w42005;
assign w42048 = ~w41979 & w42047;
assign w42049 = w41986 & ~w42003;
assign w42050 = w41973 & ~w42005;
assign w42051 = ~w41967 & ~w41986;
assign w42052 = ~w42050 & w42051;
assign w42053 = w41966 & ~w41986;
assign w42054 = w41988 & w42053;
assign w42055 = ~w42048 & ~w42054;
assign w42056 = ~w42049 & w42055;
assign w42057 = ~w42052 & w42056;
assign w42058 = w42029 & ~w42057;
assign w42059 = w41960 & w41989;
assign w42060 = w41986 & w42059;
assign w42061 = w42005 & w42053;
assign w42062 = w42037 & ~w42050;
assign w42063 = ~w42051 & w42062;
assign w42064 = ~w42060 & ~w42061;
assign w42065 = ~w42063 & w42064;
assign w42066 = ~w42029 & ~w42065;
assign w42067 = w41999 & ~w42046;
assign w42068 = ~w42066 & w42067;
assign w42069 = ~w42058 & w42068;
assign w42070 = ~pi4501 & pi9040;
assign w42071 = ~pi4502 & ~pi9040;
assign w42072 = ~w42070 & ~w42071;
assign w42073 = pi2258 & ~w42072;
assign w42074 = ~pi2258 & w42072;
assign w42075 = ~w42073 & ~w42074;
assign w42076 = ~pi4803 & pi9040;
assign w42077 = ~pi4476 & ~pi9040;
assign w42078 = ~w42076 & ~w42077;
assign w42079 = pi2245 & ~w42078;
assign w42080 = ~pi2245 & w42078;
assign w42081 = ~w42079 & ~w42080;
assign w42082 = w42075 & w42081;
assign w42083 = ~pi4498 & pi9040;
assign w42084 = ~pi4822 & ~pi9040;
assign w42085 = ~w42083 & ~w42084;
assign w42086 = pi2206 & ~w42085;
assign w42087 = ~pi2206 & w42085;
assign w42088 = ~w42086 & ~w42087;
assign w42089 = ~w42082 & ~w42088;
assign w42090 = ~pi4656 & pi9040;
assign w42091 = ~pi4439 & ~pi9040;
assign w42092 = ~w42090 & ~w42091;
assign w42093 = pi2240 & ~w42092;
assign w42094 = ~pi2240 & w42092;
assign w42095 = ~w42093 & ~w42094;
assign w42096 = w42088 & w42095;
assign w42097 = w42075 & ~w42095;
assign w42098 = ~w42081 & w42088;
assign w42099 = w42097 & w42098;
assign w42100 = ~pi4387 & pi9040;
assign w42101 = ~pi4534 & ~pi9040;
assign w42102 = ~w42100 & ~w42101;
assign w42103 = pi2269 & ~w42102;
assign w42104 = ~pi2269 & w42102;
assign w42105 = ~w42103 & ~w42104;
assign w42106 = ~w42099 & ~w42105;
assign w42107 = ~w42096 & ~w42106;
assign w42108 = ~w42089 & w42107;
assign w42109 = ~w42075 & w42095;
assign w42110 = ~w42097 & ~w42109;
assign w42111 = ~w42081 & ~w42110;
assign w42112 = ~w42075 & ~w42088;
assign w42113 = ~w42081 & w42112;
assign w42114 = ~w42095 & w42113;
assign w42115 = w42105 & ~w42114;
assign w42116 = ~w42096 & ~w42112;
assign w42117 = ~w42111 & ~w42116;
assign w42118 = ~w42115 & w42117;
assign w42119 = ~w42108 & ~w42118;
assign w42120 = ~w42075 & w42081;
assign w42121 = ~w42088 & w42095;
assign w42122 = w42120 & w42121;
assign w42123 = w42119 & ~w42122;
assign w42124 = ~pi4496 & pi9040;
assign w42125 = ~pi4536 & ~pi9040;
assign w42126 = ~w42124 & ~w42125;
assign w42127 = pi2264 & ~w42126;
assign w42128 = ~pi2264 & w42126;
assign w42129 = ~w42127 & ~w42128;
assign w42130 = ~w42123 & ~w42129;
assign w42131 = w42098 & w42109;
assign w42132 = w42105 & ~w42131;
assign w42133 = w42075 & ~w42081;
assign w42134 = w42121 & w42133;
assign w42135 = ~w42105 & ~w42134;
assign w42136 = w42081 & ~w42088;
assign w42137 = w42097 & w42136;
assign w42138 = w42135 & ~w42137;
assign w42139 = ~w42114 & w42138;
assign w42140 = ~w42132 & ~w42139;
assign w42141 = ~w42120 & ~w42133;
assign w42142 = w42096 & w42141;
assign w42143 = ~w42075 & ~w42095;
assign w42144 = w42119 & w42143;
assign w42145 = w42105 & w42111;
assign w42146 = w42075 & w42095;
assign w42147 = ~w42088 & ~w42105;
assign w42148 = w42146 & w42147;
assign w42149 = ~w42142 & ~w42148;
assign w42150 = ~w42145 & w42149;
assign w42151 = ~w42144 & w42150;
assign w42152 = w42129 & ~w42151;
assign w42153 = ~w42130 & ~w42140;
assign w42154 = ~w42152 & w42153;
assign w42155 = ~pi4324 & pi9040;
assign w42156 = ~pi4803 & ~pi9040;
assign w42157 = ~w42155 & ~w42156;
assign w42158 = pi2230 & ~w42157;
assign w42159 = ~pi2230 & w42157;
assign w42160 = ~w42158 & ~w42159;
assign w42161 = ~pi4439 & pi9040;
assign w42162 = ~pi4500 & ~pi9040;
assign w42163 = ~w42161 & ~w42162;
assign w42164 = pi2270 & ~w42163;
assign w42165 = ~pi2270 & w42163;
assign w42166 = ~w42164 & ~w42165;
assign w42167 = w42160 & ~w42166;
assign w42168 = ~pi4764 & pi9040;
assign w42169 = ~pi4498 & ~pi9040;
assign w42170 = ~w42168 & ~w42169;
assign w42171 = pi2246 & ~w42170;
assign w42172 = ~pi2246 & w42170;
assign w42173 = ~w42171 & ~w42172;
assign w42174 = ~w42167 & ~w42173;
assign w42175 = ~pi4717 & pi9040;
assign w42176 = ~pi4387 & ~pi9040;
assign w42177 = ~w42175 & ~w42176;
assign w42178 = pi2234 & ~w42177;
assign w42179 = ~pi2234 & w42177;
assign w42180 = ~w42178 & ~w42179;
assign w42181 = ~w42174 & w42180;
assign w42182 = ~pi4502 & pi9040;
assign w42183 = ~pi4434 & ~pi9040;
assign w42184 = ~w42182 & ~w42183;
assign w42185 = pi2267 & ~w42184;
assign w42186 = ~pi2267 & w42184;
assign w42187 = ~w42185 & ~w42186;
assign w42188 = w42173 & w42187;
assign w42189 = ~pi4321 & pi9040;
assign w42190 = ~pi4443 & ~pi9040;
assign w42191 = ~w42189 & ~w42190;
assign w42192 = pi2217 & ~w42191;
assign w42193 = ~pi2217 & w42191;
assign w42194 = ~w42192 & ~w42193;
assign w42195 = w42160 & ~w42187;
assign w42196 = ~w42160 & w42187;
assign w42197 = ~w42195 & ~w42196;
assign w42198 = ~w42160 & ~w42166;
assign w42199 = ~w42188 & w42194;
assign w42200 = ~w42198 & w42199;
assign w42201 = w42197 & w42200;
assign w42202 = ~w42181 & w42201;
assign w42203 = ~w42160 & ~w42194;
assign w42204 = ~w42173 & w42187;
assign w42205 = w42203 & w42204;
assign w42206 = w42180 & ~w42205;
assign w42207 = ~w42160 & w42194;
assign w42208 = w42188 & w42207;
assign w42209 = ~w42205 & ~w42208;
assign w42210 = ~w42166 & ~w42206;
assign w42211 = ~w42209 & w42210;
assign w42212 = w42173 & ~w42187;
assign w42213 = w42167 & w42212;
assign w42214 = w42167 & ~w42204;
assign w42215 = w42173 & w42194;
assign w42216 = ~w42187 & w42215;
assign w42217 = w42160 & w42216;
assign w42218 = w42180 & ~w42217;
assign w42219 = ~w42173 & w42194;
assign w42220 = w42160 & w42219;
assign w42221 = w42166 & ~w42220;
assign w42222 = ~w42188 & ~w42207;
assign w42223 = ~w42160 & w42215;
assign w42224 = w42166 & ~w42223;
assign w42225 = ~w42222 & w42224;
assign w42226 = w42187 & w42221;
assign w42227 = ~w42225 & w42226;
assign w42228 = w42173 & w42203;
assign w42229 = w42160 & ~w42194;
assign w42230 = w42204 & w42229;
assign w42231 = ~w42166 & ~w42228;
assign w42232 = ~w42230 & w42231;
assign w42233 = ~w42188 & w42203;
assign w42234 = ~w42232 & w42233;
assign w42235 = ~w42214 & w42218;
assign w42236 = ~w42227 & w42235;
assign w42237 = ~w42234 & w42236;
assign w42238 = ~w42207 & ~w42229;
assign w42239 = ~w42215 & ~w42238;
assign w42240 = ~w42187 & w42239;
assign w42241 = ~w42180 & ~w42225;
assign w42242 = ~w42240 & w42241;
assign w42243 = ~w42237 & ~w42242;
assign w42244 = ~w42202 & ~w42213;
assign w42245 = ~w42211 & w42244;
assign w42246 = ~w42243 & w42245;
assign w42247 = w42081 & w42110;
assign w42248 = w42088 & w42247;
assign w42249 = w42115 & ~w42248;
assign w42250 = ~w42135 & ~w42249;
assign w42251 = ~w42082 & ~w42097;
assign w42252 = ~w42088 & ~w42251;
assign w42253 = w42132 & ~w42252;
assign w42254 = w42095 & w42112;
assign w42255 = w42106 & ~w42254;
assign w42256 = ~w42253 & ~w42255;
assign w42257 = ~w42248 & ~w42256;
assign w42258 = w42129 & ~w42257;
assign w42259 = w42097 & w42106;
assign w42260 = w42088 & w42105;
assign w42261 = ~w42095 & ~w42260;
assign w42262 = ~w42122 & ~w42133;
assign w42263 = ~w42261 & ~w42262;
assign w42264 = ~w42121 & ~w42260;
assign w42265 = w42081 & ~w42105;
assign w42266 = ~w42075 & ~w42265;
assign w42267 = w42264 & w42266;
assign w42268 = ~w42259 & ~w42267;
assign w42269 = ~w42263 & w42268;
assign w42270 = ~w42129 & ~w42269;
assign w42271 = w42109 & w42265;
assign w42272 = ~w42250 & ~w42271;
assign w42273 = ~w42258 & w42272;
assign w42274 = ~w42270 & w42273;
assign w42275 = w42188 & w42229;
assign w42276 = ~w42205 & ~w42275;
assign w42277 = w42204 & w42207;
assign w42278 = ~w42173 & ~w42207;
assign w42279 = ~w42188 & ~w42215;
assign w42280 = ~w42278 & w42279;
assign w42281 = ~w42160 & ~w42280;
assign w42282 = ~w42180 & ~w42278;
assign w42283 = ~w42281 & w42282;
assign w42284 = w42276 & ~w42277;
assign w42285 = ~w42283 & w42284;
assign w42286 = w42166 & ~w42285;
assign w42287 = w42167 & w42215;
assign w42288 = ~w42173 & ~w42187;
assign w42289 = ~w42194 & w42288;
assign w42290 = w42221 & ~w42289;
assign w42291 = ~w42232 & ~w42290;
assign w42292 = w42212 & ~w42224;
assign w42293 = w42180 & ~w42277;
assign w42294 = ~w42287 & w42293;
assign w42295 = ~w42292 & w42294;
assign w42296 = ~w42291 & w42295;
assign w42297 = ~w42220 & ~w42289;
assign w42298 = ~w42166 & ~w42297;
assign w42299 = ~w42180 & ~w42208;
assign w42300 = w42276 & w42299;
assign w42301 = ~w42298 & w42300;
assign w42302 = ~w42296 & ~w42301;
assign w42303 = ~w42286 & ~w42302;
assign w42304 = ~w41953 & w41973;
assign w42305 = w41986 & w42304;
assign w42306 = (w42051 & w42013) | (w42051 & w66442) | (w42013 & w66442);
assign w42307 = w42029 & ~w42305;
assign w42308 = ~w41980 & w42307;
assign w42309 = ~w42306 & w42308;
assign w42310 = w41959 & w41986;
assign w42311 = w41991 & ~w42043;
assign w42312 = w42310 & ~w42311;
assign w42313 = ~w41986 & w42006;
assign w42314 = ~w42001 & ~w42029;
assign w42315 = ~w42054 & w42314;
assign w42316 = ~w41996 & ~w42313;
assign w42317 = w42315 & w42316;
assign w42318 = ~w42312 & w42317;
assign w42319 = ~w42309 & ~w42318;
assign w42320 = ~w41978 & w42036;
assign w42321 = w42022 & w42320;
assign w42322 = ~w41960 & ~w42043;
assign w42323 = w42053 & ~w42322;
assign w42324 = ~w42060 & ~w42323;
assign w42325 = ~w42321 & w42324;
assign w42326 = ~w42319 & w42325;
assign w42327 = ~w41979 & ~w42002;
assign w42328 = w41986 & ~w42327;
assign w42329 = ~w42045 & ~w42320;
assign w42330 = ~w42328 & w42329;
assign w42331 = ~w42029 & ~w42330;
assign w42332 = ~w42020 & ~w42304;
assign w42333 = w42014 & ~w42332;
assign w42334 = w41990 & w42310;
assign w42335 = ~w41995 & ~w42059;
assign w42336 = ~w42334 & w42335;
assign w42337 = ~w42333 & w42336;
assign w42338 = w42029 & ~w42337;
assign w42339 = ~w42002 & ~w42005;
assign w42340 = w41992 & ~w42339;
assign w42341 = ~w42313 & ~w42340;
assign w42342 = ~w42321 & w42341;
assign w42343 = ~w42338 & w42342;
assign w42344 = ~w42331 & w42343;
assign w42345 = pi2331 & ~w42344;
assign w42346 = ~pi2331 & w42344;
assign w42347 = ~w42345 & ~w42346;
assign w42348 = ~pi4478 & pi9040;
assign w42349 = ~pi4395 & ~pi9040;
assign w42350 = ~w42348 & ~w42349;
assign w42351 = pi2233 & ~w42350;
assign w42352 = ~pi2233 & w42350;
assign w42353 = ~w42351 & ~w42352;
assign w42354 = ~pi4532 & pi9040;
assign w42355 = ~pi4312 & ~pi9040;
assign w42356 = ~w42354 & ~w42355;
assign w42357 = pi2254 & ~w42356;
assign w42358 = ~pi2254 & w42356;
assign w42359 = ~w42357 & ~w42358;
assign w42360 = w42353 & ~w42359;
assign w42361 = ~pi4546 & pi9040;
assign w42362 = ~pi4646 & ~pi9040;
assign w42363 = ~w42361 & ~w42362;
assign w42364 = pi2265 & ~w42363;
assign w42365 = ~pi2265 & w42363;
assign w42366 = ~w42364 & ~w42365;
assign w42367 = ~pi4407 & pi9040;
assign w42368 = ~pi4488 & ~pi9040;
assign w42369 = ~w42367 & ~w42368;
assign w42370 = pi2222 & ~w42369;
assign w42371 = ~pi2222 & w42369;
assign w42372 = ~w42370 & ~w42371;
assign w42373 = ~w42366 & w42372;
assign w42374 = ~pi4537 & pi9040;
assign w42375 = ~pi4390 & ~pi9040;
assign w42376 = ~w42374 & ~w42375;
assign w42377 = pi2198 & ~w42376;
assign w42378 = ~pi2198 & w42376;
assign w42379 = ~w42377 & ~w42378;
assign w42380 = w42373 & w42379;
assign w42381 = w42360 & w42380;
assign w42382 = ~pi4662 & pi9040;
assign w42383 = ~pi4706 & ~pi9040;
assign w42384 = ~w42382 & ~w42383;
assign w42385 = pi2271 & ~w42384;
assign w42386 = ~pi2271 & w42384;
assign w42387 = ~w42385 & ~w42386;
assign w42388 = w42359 & ~w42372;
assign w42389 = w42353 & w42366;
assign w42390 = w42388 & w42389;
assign w42391 = w42387 & ~w42390;
assign w42392 = ~w42360 & ~w42373;
assign w42393 = w42360 & w42372;
assign w42394 = w42360 & w42373;
assign w42395 = ~w42392 & ~w42394;
assign w42396 = ~w42379 & ~w42395;
assign w42397 = ~w42353 & ~w42372;
assign w42398 = ~w42366 & w42397;
assign w42399 = ~w42353 & w42372;
assign w42400 = w42366 & w42399;
assign w42401 = w42379 & ~w42400;
assign w42402 = ~w42398 & w42401;
assign w42403 = ~w42396 & ~w42402;
assign w42404 = w42391 & ~w42403;
assign w42405 = ~w42353 & ~w42379;
assign w42406 = w42399 & w42819;
assign w42407 = ~w42388 & ~w42406;
assign w42408 = w42405 & ~w42407;
assign w42409 = w42366 & w42372;
assign w42410 = ~w42379 & ~w42409;
assign w42411 = w42353 & w42359;
assign w42412 = ~w42410 & w42411;
assign w42413 = w42366 & ~w42372;
assign w42414 = ~w42373 & ~w42413;
assign w42415 = w42379 & ~w42414;
assign w42416 = ~w42388 & w42415;
assign w42417 = ~w42387 & ~w42394;
assign w42418 = ~w42412 & w42417;
assign w42419 = ~w42416 & w42418;
assign w42420 = ~w42408 & w42419;
assign w42421 = ~w42404 & ~w42420;
assign w42422 = ~w42353 & w42359;
assign w42423 = ~w42413 & ~w42422;
assign w42424 = ~w42392 & ~w42423;
assign w42425 = w42397 & w42913;
assign w42426 = ~w42424 & ~w42425;
assign w42427 = w42413 & w42422;
assign w42428 = w42426 & ~w42427;
assign w42429 = ~w42379 & ~w42428;
assign w42430 = ~w42381 & ~w42429;
assign w42431 = ~w42421 & w42430;
assign w42432 = ~pi2272 & w42431;
assign w42433 = pi2272 & ~w42431;
assign w42434 = ~w42432 & ~w42433;
assign w42435 = ~w42257 & w42265;
assign w42436 = ~w42096 & ~w42113;
assign w42437 = w42249 & ~w42436;
assign w42438 = ~w42095 & ~w42112;
assign w42439 = w42138 & w42438;
assign w42440 = ~w42437 & ~w42439;
assign w42441 = w42129 & w42440;
assign w42442 = w42075 & ~w42096;
assign w42443 = ~w42136 & w42442;
assign w42444 = w42105 & ~w42443;
assign w42445 = ~w42105 & ~w42113;
assign w42446 = ~w42137 & w42445;
assign w42447 = ~w42444 & ~w42446;
assign w42448 = ~w42129 & ~w42134;
assign w42449 = ~w42142 & w42448;
assign w42450 = ~w42447 & w42449;
assign w42451 = ~w42441 & ~w42450;
assign w42452 = ~w42129 & ~w42249;
assign w42453 = ~w42096 & w42247;
assign w42454 = ~w42452 & w42453;
assign w42455 = ~w42435 & ~w42454;
assign w42456 = ~w42451 & w42455;
assign w42457 = ~pi4386 & pi9040;
assign w42458 = ~pi4320 & ~pi9040;
assign w42459 = ~w42457 & ~w42458;
assign w42460 = pi2262 & ~w42459;
assign w42461 = ~pi2262 & w42459;
assign w42462 = ~w42460 & ~w42461;
assign w42463 = ~pi4720 & pi9040;
assign w42464 = ~pi4757 & ~pi9040;
assign w42465 = ~w42463 & ~w42464;
assign w42466 = pi2241 & ~w42465;
assign w42467 = ~pi2241 & w42465;
assign w42468 = ~w42466 & ~w42467;
assign w42469 = ~w42462 & w42468;
assign w42470 = w42462 & ~w42468;
assign w42471 = ~w42469 & ~w42470;
assign w42472 = ~pi4440 & pi9040;
assign w42473 = ~pi4662 & ~pi9040;
assign w42474 = ~w42472 & ~w42473;
assign w42475 = pi2227 & ~w42474;
assign w42476 = ~pi2227 & w42474;
assign w42477 = ~w42475 & ~w42476;
assign w42478 = ~pi4474 & pi9040;
assign w42479 = ~pi4546 & ~pi9040;
assign w42480 = ~w42478 & ~w42479;
assign w42481 = pi2268 & ~w42480;
assign w42482 = ~pi2268 & w42480;
assign w42483 = ~w42481 & ~w42482;
assign w42484 = w42477 & ~w42483;
assign w42485 = ~w42468 & w42484;
assign w42486 = w42462 & ~w42483;
assign w42487 = w42470 & w42477;
assign w42488 = ~w42486 & ~w42487;
assign w42489 = ~w42469 & w42488;
assign w42490 = ~pi4488 & pi9040;
assign w42491 = ~pi4596 & ~pi9040;
assign w42492 = ~w42490 & ~w42491;
assign w42493 = pi2216 & ~w42492;
assign w42494 = ~pi2216 & w42492;
assign w42495 = ~w42493 & ~w42494;
assign w42496 = ~w42489 & ~w42495;
assign w42497 = ~w42485 & ~w42496;
assign w42498 = w42471 & ~w42497;
assign w42499 = w42462 & w42468;
assign w42500 = ~w42477 & w42499;
assign w42501 = ~w42495 & ~w42500;
assign w42502 = ~w42477 & w42483;
assign w42503 = w42471 & ~w42502;
assign w42504 = w42501 & w42503;
assign w42505 = ~pi4597 & pi9040;
assign w42506 = ~pi4532 & ~pi9040;
assign w42507 = ~w42505 & ~w42506;
assign w42508 = pi2266 & ~w42507;
assign w42509 = ~pi2266 & w42507;
assign w42510 = ~w42508 & ~w42509;
assign w42511 = ~w42484 & ~w42488;
assign w42512 = w42468 & w42484;
assign w42513 = ~w42511 & ~w42512;
assign w42514 = w42495 & ~w42513;
assign w42515 = w42477 & ~w42486;
assign w42516 = w42470 & ~w42477;
assign w42517 = ~w42515 & ~w42516;
assign w42518 = ~w42495 & ~w42517;
assign w42519 = ~w42469 & ~w42518;
assign w42520 = w42502 & ~w42519;
assign w42521 = ~w42504 & ~w42510;
assign w42522 = ~w42514 & w42521;
assign w42523 = ~w42520 & w42522;
assign w42524 = w42485 & w42495;
assign w42525 = w42501 & ~w42511;
assign w42526 = w42468 & w42477;
assign w42527 = w42483 & w42526;
assign w42528 = ~w42468 & ~w42477;
assign w42529 = ~w42486 & w42528;
assign w42530 = w42495 & ~w42529;
assign w42531 = ~w42527 & w42530;
assign w42532 = ~w42525 & ~w42531;
assign w42533 = w42471 & w42502;
assign w42534 = ~w42484 & ~w42502;
assign w42535 = w42468 & w42534;
assign w42536 = ~w42533 & ~w42535;
assign w42537 = ~w42462 & ~w42536;
assign w42538 = w42510 & ~w42524;
assign w42539 = ~w42537 & w42538;
assign w42540 = ~w42532 & w42539;
assign w42541 = ~w42523 & ~w42540;
assign w42542 = ~w42498 & ~w42541;
assign w42543 = ~w42495 & w42512;
assign w42544 = w42468 & ~w42543;
assign w42545 = w42486 & ~w42544;
assign w42546 = w42469 & ~w42477;
assign w42547 = w42483 & w42495;
assign w42548 = w42546 & ~w42547;
assign w42549 = ~w42533 & ~w42548;
assign w42550 = ~w42545 & w42549;
assign w42551 = w42510 & ~w42550;
assign w42552 = w42469 & w42484;
assign w42553 = ~w42462 & w42477;
assign w42554 = w42510 & w42553;
assign w42555 = ~w42477 & ~w42510;
assign w42556 = w42471 & w42555;
assign w42557 = ~w42552 & ~w42554;
assign w42558 = ~w42556 & w42557;
assign w42559 = w42495 & ~w42558;
assign w42560 = w42483 & w42499;
assign w42561 = w42477 & w42560;
assign w42562 = ~w42518 & ~w42561;
assign w42563 = ~w42510 & ~w42562;
assign w42564 = ~w42483 & ~w42499;
assign w42565 = w42462 & w42495;
assign w42566 = ~w42534 & w42565;
assign w42567 = ~w42495 & w42546;
assign w42568 = ~w42566 & ~w42567;
assign w42569 = w42564 & ~w42568;
assign w42570 = ~w42559 & ~w42569;
assign w42571 = ~w42563 & w42570;
assign w42572 = ~w42551 & w42571;
assign w42573 = ~pi4729 & pi9040;
assign w42574 = ~pi4321 & ~pi9040;
assign w42575 = ~w42573 & ~w42574;
assign w42576 = pi2223 & ~w42575;
assign w42577 = ~pi2223 & w42575;
assign w42578 = ~w42576 & ~w42577;
assign w42579 = ~pi4434 & pi9040;
assign w42580 = ~pi4496 & ~pi9040;
assign w42581 = ~w42579 & ~w42580;
assign w42582 = pi2271 & ~w42581;
assign w42583 = ~pi2271 & w42581;
assign w42584 = ~w42582 & ~w42583;
assign w42585 = ~pi4500 & pi9040;
assign w42586 = ~pi4504 & ~pi9040;
assign w42587 = ~w42585 & ~w42586;
assign w42588 = pi2230 & ~w42587;
assign w42589 = ~pi2230 & w42587;
assign w42590 = ~w42588 & ~w42589;
assign w42591 = ~w42584 & ~w42590;
assign w42592 = w42584 & w42590;
assign w42593 = ~w42591 & ~w42592;
assign w42594 = ~pi4487 & pi9040;
assign w42595 = ~pi4501 & ~pi9040;
assign w42596 = ~w42594 & ~w42595;
assign w42597 = pi2254 & ~w42596;
assign w42598 = ~pi2254 & w42596;
assign w42599 = ~w42597 & ~w42598;
assign w42600 = ~w42578 & ~w42599;
assign w42601 = ~w42590 & w42600;
assign w42602 = w42584 & w42599;
assign w42603 = ~pi4445 & pi9040;
assign w42604 = ~pi4804 & ~pi9040;
assign w42605 = ~w42603 & ~w42604;
assign w42606 = pi2255 & ~w42605;
assign w42607 = ~pi2255 & w42605;
assign w42608 = ~w42606 & ~w42607;
assign w42609 = w42602 & ~w42608;
assign w42610 = w42578 & w42599;
assign w42611 = w42590 & w42610;
assign w42612 = ~w42609 & ~w42611;
assign w42613 = ~w42601 & w42612;
assign w42614 = w42612 & w63419;
assign w42615 = ~w42578 & ~w42614;
assign w42616 = w42599 & w42608;
assign w42617 = ~w42584 & ~w42599;
assign w42618 = ~w42602 & ~w42617;
assign w42619 = ~w42590 & w42618;
assign w42620 = w42590 & ~w42618;
assign w42621 = ~w42619 & ~w42620;
assign w42622 = w42578 & w42621;
assign w42623 = w42621 & w63420;
assign w42624 = ~w42584 & w42590;
assign w42625 = w42608 & w42624;
assign w42626 = (w42616 & w42623) | (w42616 & w63986) | (w42623 & w63986);
assign w42627 = (~w42623 & w66443) | (~w42623 & w66444) | (w66443 & w66444);
assign w42628 = ~w42615 & ~w42627;
assign w42629 = ~w42619 & ~w42625;
assign w42630 = ~w42601 & w42617;
assign w42631 = w42578 & w42608;
assign w42632 = w42591 & w42631;
assign w42633 = ~w42630 & ~w42632;
assign w42634 = (w42633 & ~w42615) | (w42633 & w63987) | (~w42615 & w63987);
assign w42635 = w42590 & ~w42599;
assign w42636 = w42608 & w42635;
assign w42637 = ~w42609 & ~w42636;
assign w42638 = w42634 & w42637;
assign w42639 = ~w42608 & ~w42610;
assign w42640 = ~w42602 & w42639;
assign w42641 = ~w42592 & w42640;
assign w42642 = w42634 & w66445;
assign w42643 = ~w42628 & ~w42642;
assign w42644 = ~pi4822 & pi9040;
assign w42645 = ~pi4324 & ~pi9040;
assign w42646 = ~w42644 & ~w42645;
assign w42647 = pi2246 & ~w42646;
assign w42648 = ~pi2246 & w42646;
assign w42649 = ~w42647 & ~w42648;
assign w42650 = ~w42643 & ~w42649;
assign w42651 = w42584 & w42608;
assign w42652 = w42600 & w42651;
assign w42653 = ~w42638 & w42649;
assign w42654 = ~w42599 & w42632;
assign w42655 = w42578 & ~w42608;
assign w42656 = w42620 & w42655;
assign w42657 = ~w42590 & w42599;
assign w42658 = w42639 & w42657;
assign w42659 = ~w42652 & ~w42654;
assign w42660 = ~w42658 & w42659;
assign w42661 = ~w42656 & w42660;
assign w42662 = ~w42653 & w42661;
assign w42663 = ~w42650 & w42662;
assign w42664 = ~pi4646 & pi9040;
assign w42665 = ~pi4720 & ~pi9040;
assign w42666 = ~w42664 & ~w42665;
assign w42667 = pi2241 & ~w42666;
assign w42668 = ~pi2241 & w42666;
assign w42669 = ~w42667 & ~w42668;
assign w42670 = ~pi4596 & pi9040;
assign w42671 = ~pi4389 & ~pi9040;
assign w42672 = ~w42670 & ~w42671;
assign w42673 = pi2266 & ~w42672;
assign w42674 = ~pi2266 & w42672;
assign w42675 = ~w42673 & ~w42674;
assign w42676 = ~w42669 & w42675;
assign w42677 = ~pi4320 & pi9040;
assign w42678 = ~pi4499 & ~pi9040;
assign w42679 = ~w42677 & ~w42678;
assign w42680 = pi2252 & ~w42679;
assign w42681 = ~pi2252 & w42679;
assign w42682 = ~w42680 & ~w42681;
assign w42683 = w42676 & w42682;
assign w42684 = ~pi4388 & pi9040;
assign w42685 = ~pi4601 & ~pi9040;
assign w42686 = ~w42684 & ~w42685;
assign w42687 = pi2233 & ~w42686;
assign w42688 = ~pi2233 & w42686;
assign w42689 = ~w42687 & ~w42688;
assign w42690 = w42669 & w42689;
assign w42691 = w42675 & ~w42682;
assign w42692 = w42690 & w42691;
assign w42693 = ~w42683 & ~w42692;
assign w42694 = ~pi4706 & pi9040;
assign w42695 = ~pi4585 & ~pi9040;
assign w42696 = ~w42694 & ~w42695;
assign w42697 = pi2263 & ~w42696;
assign w42698 = ~pi2263 & w42696;
assign w42699 = ~w42697 & ~w42698;
assign w42700 = ~w42693 & ~w42699;
assign w42701 = ~w42669 & ~w42689;
assign w42702 = ~w42675 & ~w42682;
assign w42703 = w42701 & w42702;
assign w42704 = ~w42675 & w42689;
assign w42705 = ~w42669 & ~w42682;
assign w42706 = ~w42690 & ~w42701;
assign w42707 = ~w42705 & w42706;
assign w42708 = w42704 & w42707;
assign w42709 = w42675 & ~w42689;
assign w42710 = ~w42704 & ~w42709;
assign w42711 = w42669 & ~w42710;
assign w42712 = w42676 & w42689;
assign w42713 = ~w42711 & ~w42712;
assign w42714 = w42699 & ~w42707;
assign w42715 = ~w42713 & w42714;
assign w42716 = ~w42700 & ~w42703;
assign w42717 = ~w42708 & w42716;
assign w42718 = ~w42715 & w42717;
assign w42719 = ~pi4423 & pi9040;
assign w42720 = pi4597 & ~pi9040;
assign w42721 = ~w42719 & ~w42720;
assign w42722 = pi2222 & ~w42721;
assign w42723 = ~pi2222 & w42721;
assign w42724 = ~w42722 & ~w42723;
assign w42725 = ~w42718 & ~w42724;
assign w42726 = ~w42689 & w42699;
assign w42727 = ~w42702 & w42726;
assign w42728 = w42699 & ~w42709;
assign w42729 = ~w42669 & ~w42728;
assign w42730 = ~w42675 & w42682;
assign w42731 = ~w42691 & ~w42730;
assign w42732 = w42689 & w42731;
assign w42733 = ~w42727 & ~w42729;
assign w42734 = ~w42732 & w42733;
assign w42735 = ~w42691 & w42729;
assign w42736 = w42669 & w42730;
assign w42737 = w42724 & ~w42736;
assign w42738 = ~w42735 & w42737;
assign w42739 = ~w42734 & w42738;
assign w42740 = w42669 & w42731;
assign w42741 = w42699 & ~w42740;
assign w42742 = ~w42699 & ~w42708;
assign w42743 = w42701 & ~w42730;
assign w42744 = ~w42689 & w42736;
assign w42745 = ~w42743 & ~w42744;
assign w42746 = w42742 & w42745;
assign w42747 = ~w42741 & ~w42746;
assign w42748 = ~w42739 & ~w42747;
assign w42749 = ~w42725 & w42748;
assign w42750 = w42503 & w42547;
assign w42751 = (~w42516 & ~w42536) | (~w42516 & w66446) | (~w42536 & w66446);
assign w42752 = w42496 & w42751;
assign w42753 = w42495 & ~w42751;
assign w42754 = ~w42462 & w42485;
assign w42755 = ~w42752 & ~w42754;
assign w42756 = ~w42753 & w42755;
assign w42757 = ~w42510 & ~w42756;
assign w42758 = ~w42484 & ~w42495;
assign w42759 = ~w42487 & ~w42533;
assign w42760 = w42758 & ~w42759;
assign w42761 = ~w42510 & ~w42528;
assign w42762 = ~w42495 & ~w42527;
assign w42763 = ~w42547 & ~w42762;
assign w42764 = ~w42470 & w42477;
assign w42765 = ~w42761 & ~w42764;
assign w42766 = w42763 & w42765;
assign w42767 = ~w42483 & w42516;
assign w42768 = ~w42543 & ~w42560;
assign w42769 = ~w42767 & w42768;
assign w42770 = w42510 & ~w42769;
assign w42771 = ~w42750 & ~w42760;
assign w42772 = ~w42766 & w42771;
assign w42773 = ~w42770 & w42772;
assign w42774 = ~w42757 & w42773;
assign w42775 = ~w42187 & w42219;
assign w42776 = ~w42221 & w42775;
assign w42777 = w42229 & w42292;
assign w42778 = w42187 & w42215;
assign w42779 = ~w42166 & ~w42778;
assign w42780 = ~w42281 & w42779;
assign w42781 = ~w42240 & w42280;
assign w42782 = ~w42212 & w42229;
assign w42783 = w42166 & ~w42782;
assign w42784 = ~w42217 & w42783;
assign w42785 = ~w42781 & w42784;
assign w42786 = ~w42780 & ~w42785;
assign w42787 = ~w42180 & ~w42776;
assign w42788 = ~w42777 & w42787;
assign w42789 = ~w42786 & w42788;
assign w42790 = ~w42194 & w42196;
assign w42791 = w42224 & ~w42790;
assign w42792 = ~w42195 & ~w42297;
assign w42793 = ~w42166 & ~w42792;
assign w42794 = ~w42781 & w42793;
assign w42795 = ~w42791 & ~w42794;
assign w42796 = ~w42204 & w42782;
assign w42797 = ~w42201 & ~w42796;
assign w42798 = w42218 & w42797;
assign w42799 = ~w42795 & w42798;
assign w42800 = ~w42789 & ~w42799;
assign w42801 = w42359 & w42415;
assign w42802 = ~w42393 & ~w42400;
assign w42803 = ~w42379 & ~w42802;
assign w42804 = w42353 & w42413;
assign w42805 = w42353 & w42373;
assign w42806 = w42359 & w42805;
assign w42807 = w42353 & w42379;
assign w42808 = ~w42359 & ~w42372;
assign w42809 = w42807 & w42808;
assign w42810 = ~w42804 & ~w42809;
assign w42811 = ~w42406 & w42810;
assign w42812 = ~w42425 & ~w42806;
assign w42813 = w42811 & w42812;
assign w42814 = ~w42801 & ~w42803;
assign w42815 = w42813 & w42814;
assign w42816 = ~w42387 & ~w42815;
assign w42817 = ~w42380 & ~w42400;
assign w42818 = w42815 & ~w42817;
assign w42819 = ~w42359 & w42366;
assign w42820 = ~w42399 & w42819;
assign w42821 = ~w42804 & w42820;
assign w42822 = ~w42366 & w42422;
assign w42823 = w42353 & ~w42373;
assign w42824 = ~w42808 & w42823;
assign w42825 = ~w42822 & ~w42824;
assign w42826 = ~w42379 & ~w42825;
assign w42827 = w42359 & w42398;
assign w42828 = ~w42821 & ~w42827;
assign w42829 = ~w42826 & w42828;
assign w42830 = ~w42818 & w42829;
assign w42831 = w42387 & ~w42830;
assign w42832 = ~w42398 & ~w42806;
assign w42833 = ~w42403 & ~w42832;
assign w42834 = ~w42816 & ~w42833;
assign w42835 = ~w42831 & w42834;
assign w42836 = ~w42131 & w42141;
assign w42837 = ~w42264 & w42836;
assign w42838 = w42143 & w42147;
assign w42839 = w42088 & w42120;
assign w42840 = ~w42107 & w42839;
assign w42841 = ~w42837 & ~w42838;
assign w42842 = ~w42840 & w42841;
assign w42843 = w42129 & ~w42842;
assign w42844 = ~w42121 & ~w42146;
assign w42845 = ~w42440 & ~w42844;
assign w42846 = w42106 & ~w42131;
assign w42847 = w42129 & ~w42133;
assign w42848 = w42088 & ~w42120;
assign w42849 = ~w42095 & ~w42847;
assign w42850 = ~w42848 & w42849;
assign w42851 = w42105 & ~w42850;
assign w42852 = ~w42846 & ~w42851;
assign w42853 = w42111 & ~w42121;
assign w42854 = w42265 & ~w42844;
assign w42855 = ~w42148 & ~w42854;
assign w42856 = ~w42853 & w42855;
assign w42857 = ~w42129 & ~w42856;
assign w42858 = ~w42852 & ~w42857;
assign w42859 = ~w42843 & w42858;
assign w42860 = ~w42845 & w42859;
assign w42861 = ~w42389 & ~w42405;
assign w42862 = w42359 & ~w42861;
assign w42863 = ~w42379 & ~w42390;
assign w42864 = w42360 & ~w42409;
assign w42865 = ~w42862 & ~w42864;
assign w42866 = w42863 & w42865;
assign w42867 = w42359 & w42379;
assign w42868 = w42409 & w42867;
assign w42869 = ~w42387 & ~w42427;
assign w42870 = ~w42809 & ~w42868;
assign w42871 = w42869 & w42870;
assign w42872 = ~w42866 & w42871;
assign w42873 = ~w42379 & ~w42399;
assign w42874 = w42353 & w42388;
assign w42875 = ~w42393 & ~w42398;
assign w42876 = ~w42874 & w42875;
assign w42877 = ~w42413 & w42873;
assign w42878 = w42876 & w42877;
assign w42879 = w42379 & ~w42876;
assign w42880 = w42391 & w66447;
assign w42881 = ~w42878 & w42880;
assign w42882 = ~w42879 & w42881;
assign w42883 = w42379 & w42424;
assign w42884 = w42405 & w42819;
assign w42885 = ~w42381 & ~w42884;
assign w42886 = ~w42883 & w42885;
assign w42887 = (w42886 & w42882) | (w42886 & w66448) | (w42882 & w66448);
assign w42888 = pi2288 & ~w42887;
assign w42889 = ~pi2288 & w42887;
assign w42890 = ~w42888 & ~w42889;
assign w42891 = w42462 & w42502;
assign w42892 = ~w42526 & ~w42564;
assign w42893 = ~w42891 & w42892;
assign w42894 = ~w42552 & ~w42893;
assign w42895 = w42495 & w42894;
assign w42896 = w42483 & ~w42553;
assign w42897 = w42758 & ~w42896;
assign w42898 = w42485 & ~w42518;
assign w42899 = w42568 & ~w42897;
assign w42900 = ~w42898 & w42899;
assign w42901 = w42894 & w42900;
assign w42902 = ~w42495 & ~w42901;
assign w42903 = w42510 & ~w42895;
assign w42904 = ~w42902 & w42903;
assign w42905 = ~w42763 & ~w42767;
assign w42906 = ~w42530 & ~w42905;
assign w42907 = ~w42462 & w42527;
assign w42908 = w42900 & ~w42907;
assign w42909 = ~w42510 & ~w42908;
assign w42910 = ~w42569 & ~w42906;
assign w42911 = ~w42909 & w42910;
assign w42912 = ~w42904 & w42911;
assign w42913 = ~w42359 & ~w42366;
assign w42914 = ~w42397 & w42913;
assign w42915 = ~w42807 & w42914;
assign w42916 = w42399 & ~w42863;
assign w42917 = ~w42372 & ~w42422;
assign w42918 = w42873 & ~w42917;
assign w42919 = ~w42915 & ~w42918;
assign w42920 = ~w42916 & w42919;
assign w42921 = ~w42387 & ~w42920;
assign w42922 = ~w42827 & w42863;
assign w42923 = ~w42366 & w42874;
assign w42924 = (~w42359 & w42424) | (~w42359 & w66449) | (w42424 & w66449);
assign w42925 = w42401 & ~w42923;
assign w42926 = ~w42924 & w42925;
assign w42927 = ~w42922 & ~w42926;
assign w42928 = w42808 & ~w42861;
assign w42929 = w42366 & w42422;
assign w42930 = ~w42408 & w42929;
assign w42931 = ~w42805 & ~w42928;
assign w42932 = ~w42930 & w42931;
assign w42933 = w42387 & ~w42932;
assign w42934 = ~w42921 & ~w42927;
assign w42935 = ~w42933 & w42934;
assign w42936 = ~pi2276 & w42935;
assign w42937 = pi2276 & ~w42935;
assign w42938 = ~w42936 & ~w42937;
assign w42939 = ~pi4504 & pi9040;
assign w42940 = ~pi4764 & ~pi9040;
assign w42941 = ~w42939 & ~w42940;
assign w42942 = pi2251 & ~w42941;
assign w42943 = ~pi2251 & w42941;
assign w42944 = ~w42942 & ~w42943;
assign w42945 = ~pi4804 & pi9040;
assign w42946 = ~pi4584 & ~pi9040;
assign w42947 = ~w42945 & ~w42946;
assign w42948 = pi2234 & ~w42947;
assign w42949 = ~pi2234 & w42947;
assign w42950 = ~w42948 & ~w42949;
assign w42951 = ~pi4313 & pi9040;
assign w42952 = ~pi4656 & ~pi9040;
assign w42953 = ~w42951 & ~w42952;
assign w42954 = pi2240 & ~w42953;
assign w42955 = ~pi2240 & w42953;
assign w42956 = ~w42954 & ~w42955;
assign w42957 = ~w42950 & ~w42956;
assign w42958 = ~pi4536 & pi9040;
assign w42959 = ~pi4729 & ~pi9040;
assign w42960 = ~w42958 & ~w42959;
assign w42961 = pi2253 & ~w42960;
assign w42962 = ~pi2253 & w42960;
assign w42963 = ~w42961 & ~w42962;
assign w42964 = ~pi4534 & pi9040;
assign w42965 = ~pi4503 & ~pi9040;
assign w42966 = ~w42964 & ~w42965;
assign w42967 = pi2217 & ~w42966;
assign w42968 = ~pi2217 & w42966;
assign w42969 = ~w42967 & ~w42968;
assign w42970 = ~w42963 & ~w42969;
assign w42971 = w42957 & w42970;
assign w42972 = ~w42956 & w42969;
assign w42973 = ~w42950 & w42963;
assign w42974 = ~w42972 & ~w42973;
assign w42975 = ~w42957 & ~w42974;
assign w42976 = ~pi4476 & pi9040;
assign w42977 = ~pi4645 & ~pi9040;
assign w42978 = ~w42976 & ~w42977;
assign w42979 = pi2258 & ~w42978;
assign w42980 = ~pi2258 & w42978;
assign w42981 = ~w42979 & ~w42980;
assign w42982 = w42975 & w42981;
assign w42983 = w42956 & ~w42969;
assign w42984 = ~w42963 & ~w42981;
assign w42985 = w42983 & ~w42984;
assign w42986 = ~w42971 & ~w42985;
assign w42987 = ~w42982 & w42986;
assign w42988 = w42944 & ~w42987;
assign w42989 = w42957 & w42969;
assign w42990 = w42963 & w42989;
assign w42991 = w42981 & ~w42990;
assign w42992 = w42944 & ~w42950;
assign w42993 = w42950 & w42956;
assign w42994 = ~w42957 & ~w42993;
assign w42995 = ~w42992 & w42994;
assign w42996 = w42963 & w42969;
assign w42997 = ~w42970 & ~w42996;
assign w42998 = w42995 & ~w42997;
assign w42999 = ~w42975 & w42997;
assign w43000 = ~w42995 & w42999;
assign w43001 = ~w42981 & ~w42998;
assign w43002 = ~w43000 & w43001;
assign w43003 = ~w42991 & ~w43002;
assign w43004 = ~w42944 & w42981;
assign w43005 = w42974 & w43004;
assign w43006 = w42987 & w43005;
assign w43007 = ~w42988 & ~w43006;
assign w43008 = ~w43003 & w43007;
assign w43009 = ~w42669 & ~w42702;
assign w43010 = ~w42675 & ~w42701;
assign w43011 = ~w42699 & ~w43009;
assign w43012 = ~w43010 & w43011;
assign w43013 = w42690 & w42702;
assign w43014 = w42705 & ~w42710;
assign w43015 = w42707 & w42710;
assign w43016 = ~w43014 & ~w43015;
assign w43017 = ~w42682 & ~w42704;
assign w43018 = (w43017 & w43015) | (w43017 & w66450) | (w43015 & w66450);
assign w43019 = w42682 & ~w42713;
assign w43020 = ~w43012 & w43019;
assign w43021 = w42704 & w42729;
assign w43022 = w42701 & w42730;
assign w43023 = ~w43021 & ~w43022;
assign w43024 = ~w43018 & w43023;
assign w43025 = ~w43020 & w43024;
assign w43026 = w43009 & w43025;
assign w43027 = ~w42724 & ~w43013;
assign w43028 = ~w42744 & w43027;
assign w43029 = ~w43012 & w43028;
assign w43030 = ~w43026 & w43029;
assign w43031 = w42699 & ~w42706;
assign w43032 = w42724 & ~w43031;
assign w43033 = w43025 & w43032;
assign w43034 = ~w43030 & ~w43033;
assign w43035 = w42616 & ~w42634;
assign w43036 = ~w42635 & ~w42657;
assign w43037 = w42651 & w43036;
assign w43038 = ~w42593 & w42640;
assign w43039 = w42578 & ~w43036;
assign w43040 = w42593 & w43039;
assign w43041 = ~w42649 & ~w43037;
assign w43042 = ~w43038 & w43041;
assign w43043 = ~w43040 & w43042;
assign w43044 = ~w42578 & w42584;
assign w43045 = ~w42657 & w43044;
assign w43046 = ~w42584 & ~w42600;
assign w43047 = w42608 & ~w43044;
assign w43048 = ~w43045 & ~w43046;
assign w43049 = ~w43047 & w43048;
assign w43050 = w42592 & w42600;
assign w43051 = ~w43046 & ~w43050;
assign w43052 = w42608 & ~w43051;
assign w43053 = ~w42611 & w42649;
assign w43054 = ~w43049 & w43053;
assign w43055 = ~w43052 & w43054;
assign w43056 = ~w43043 & ~w43055;
assign w43057 = ~w43035 & ~w43056;
assign w43058 = w42591 & w42616;
assign w43059 = ~w42592 & ~w42608;
assign w43060 = w42599 & w43044;
assign w43061 = ~w43059 & ~w43060;
assign w43062 = w43036 & ~w43061;
assign w43063 = ~w42636 & ~w43058;
assign w43064 = ~w43062 & w43063;
assign w43065 = ~w42623 & w43064;
assign w43066 = ~w42609 & w43053;
assign w43067 = ~w43065 & ~w43066;
assign w43068 = ~w43062 & w66451;
assign w43069 = ~w42578 & ~w43068;
assign w43070 = ~w42622 & w42649;
assign w43071 = ~w43069 & w43070;
assign w43072 = ~w43067 & ~w43071;
assign w43073 = ~pi2306 & w43072;
assign w43074 = pi2306 & ~w43072;
assign w43075 = ~w43073 & ~w43074;
assign w43076 = ~w42682 & w42709;
assign w43077 = w43031 & ~w43076;
assign w43078 = ~w42709 & w43017;
assign w43079 = ~w43019 & ~w43078;
assign w43080 = ~w42701 & ~w42702;
assign w43081 = w43079 & w43080;
assign w43082 = ~w43077 & ~w43081;
assign w43083 = w42724 & ~w43082;
assign w43084 = w42699 & ~w42736;
assign w43085 = ~w42692 & w43084;
assign w43086 = ~w42742 & ~w43085;
assign w43087 = ~w42699 & w42724;
assign w43088 = ~w42712 & ~w43076;
assign w43089 = w43087 & ~w43088;
assign w43090 = ~w42682 & w42690;
assign w43091 = ~w42701 & ~w42709;
assign w43092 = ~w42691 & ~w43091;
assign w43093 = ~w42699 & ~w43090;
assign w43094 = ~w43092 & w43093;
assign w43095 = ~w42705 & ~w42709;
assign w43096 = ~w42691 & ~w43095;
assign w43097 = w43084 & ~w43096;
assign w43098 = ~w42741 & ~w43097;
assign w43099 = w43016 & ~w43098;
assign w43100 = ~w42724 & ~w43094;
assign w43101 = ~w43099 & w43100;
assign w43102 = ~w43086 & ~w43089;
assign w43103 = ~w43101 & w43102;
assign w43104 = ~w43083 & w43103;
assign w43105 = w42160 & w42289;
assign w43106 = w42779 & ~w43105;
assign w43107 = ~w42221 & ~w43106;
assign w43108 = ~w42216 & ~w42228;
assign w43109 = w42166 & ~w43108;
assign w43110 = ~w42166 & w42239;
assign w43111 = w42206 & ~w43109;
assign w43112 = ~w43110 & w43111;
assign w43113 = ~w42174 & ~w42203;
assign w43114 = w42197 & ~w43113;
assign w43115 = ~w42275 & ~w42287;
assign w43116 = w42299 & w43115;
assign w43117 = ~w43114 & w43116;
assign w43118 = ~w43112 & ~w43117;
assign w43119 = ~w43107 & ~w43118;
assign w43120 = ~pi2321 & w43119;
assign w43121 = pi2321 & ~w43119;
assign w43122 = ~w43120 & ~w43121;
assign w43123 = ~w42944 & w42956;
assign w43124 = w42950 & w42963;
assign w43125 = ~w42969 & w43124;
assign w43126 = ~w43123 & w43125;
assign w43127 = w42956 & w43126;
assign w43128 = ~w42989 & ~w43124;
assign w43129 = ~w42944 & ~w43128;
assign w43130 = w42970 & ~w42994;
assign w43131 = ~w42975 & ~w43130;
assign w43132 = ~w42950 & w42956;
assign w43133 = w42970 & ~w43132;
assign w43134 = (~w43133 & ~w43131) | (~w43133 & w63421) | (~w43131 & w63421);
assign w43135 = ~w42972 & ~w43124;
assign w43136 = ~w42950 & ~w42969;
assign w43137 = w43135 & ~w43136;
assign w43138 = w43135 & w63422;
assign w43139 = ~w42969 & ~w43131;
assign w43140 = ~w42993 & w42996;
assign w43141 = w42944 & ~w43135;
assign w43142 = ~w43140 & w43141;
assign w43143 = ~w43138 & ~w43142;
assign w43144 = ~w43139 & w43143;
assign w43145 = (~w43129 & ~w43144) | (~w43129 & w63423) | (~w43144 & w63423);
assign w43146 = w42981 & ~w43145;
assign w43147 = ~w42950 & ~w42963;
assign w43148 = ~w42944 & ~w42956;
assign w43149 = ~w43147 & w43148;
assign w43150 = ~w42981 & ~w43149;
assign w43151 = w43140 & ~w43150;
assign w43152 = ~w43127 & ~w43151;
assign w43153 = (w43152 & w43144) | (w43152 & w66452) | (w43144 & w66452);
assign w43154 = (pi2297 & w43146) | (pi2297 & w66453) | (w43146 & w66453);
assign w43155 = ~w43146 & w66454;
assign w43156 = ~w43154 & ~w43155;
assign w43157 = (~w43126 & ~w43131) | (~w43126 & w63989) | (~w43131 & w63989);
assign w43158 = w42944 & w42963;
assign w43159 = (~w43131 & w66455) | (~w43131 & w66456) | (w66455 & w66456);
assign w43160 = (~w43131 & w66457) | (~w43131 & w66458) | (w66457 & w66458);
assign w43161 = ~w43159 & w43160;
assign w43162 = (~w42981 & w43131) | (~w42981 & w66459) | (w43131 & w66459);
assign w43163 = w43157 & w43162;
assign w43164 = ~w43161 & ~w43163;
assign w43165 = ~w42970 & w42994;
assign w43166 = w43004 & ~w43133;
assign w43167 = ~w43165 & w43166;
assign w43168 = w42950 & w42969;
assign w43169 = w42963 & w43123;
assign w43170 = w43168 & w43169;
assign w43171 = ~w43167 & ~w43170;
assign w43172 = (w43171 & w43145) | (w43171 & w63990) | (w43145 & w63990);
assign w43173 = (pi2289 & ~w43172) | (pi2289 & w66460) | (~w43172 & w66460);
assign w43174 = w43172 & w66461;
assign w43175 = ~w43173 & ~w43174;
assign w43176 = ~w43136 & ~w43168;
assign w43177 = ~w42956 & ~w43176;
assign w43178 = w42944 & ~w43177;
assign w43179 = ~w43125 & ~w43158;
assign w43180 = ~w43178 & ~w43179;
assign w43181 = ~w43124 & w43149;
assign w43182 = ~w42997 & w43132;
assign w43183 = ~w42950 & ~w43141;
assign w43184 = ~w42972 & ~w42983;
assign w43185 = w42950 & ~w43184;
assign w43186 = ~w42963 & ~w43185;
assign w43187 = ~w43183 & w43186;
assign w43188 = ~w43181 & ~w43182;
assign w43189 = ~w43187 & w43188;
assign w43190 = w42981 & ~w43189;
assign w43191 = w43123 & w43176;
assign w43192 = w42969 & w43132;
assign w43193 = w42944 & ~w42971;
assign w43194 = ~w43192 & w43193;
assign w43195 = ~w43185 & w43194;
assign w43196 = w43150 & ~w43191;
assign w43197 = ~w43195 & w43196;
assign w43198 = ~w43180 & ~w43197;
assign w43199 = ~w43190 & w43198;
assign w43200 = pi2281 & ~w43199;
assign w43201 = ~pi2281 & w43199;
assign w43202 = ~w43200 & ~w43201;
assign w43203 = ~w43036 & w66462;
assign w43204 = w42592 & w42655;
assign w43205 = ~w43058 & ~w43204;
assign w43206 = ~w43203 & ~w43205;
assign w43207 = ~w42630 & ~w42658;
assign w43208 = w43049 & ~w43207;
assign w43209 = w42578 & w42625;
assign w43210 = w42613 & ~w43209;
assign w43211 = ~w42649 & ~w43210;
assign w43212 = ~w43044 & w43059;
assign w43213 = ~w42621 & w43212;
assign w43214 = ~w42654 & ~w43050;
assign w43215 = ~w43213 & w43214;
assign w43216 = ~w42626 & w43215;
assign w43217 = w42649 & ~w43216;
assign w43218 = ~w42652 & ~w43206;
assign w43219 = ~w43208 & w43218;
assign w43220 = ~w43211 & w43219;
assign w43221 = ~w43217 & w66463;
assign w43222 = (pi2311 & w43217) | (pi2311 & w66464) | (w43217 & w66464);
assign w43223 = ~w43221 & ~w43222;
assign w43224 = ~w42699 & w43022;
assign w43225 = w43079 & w43087;
assign w43226 = ~w42711 & w43097;
assign w43227 = ~w42701 & w43078;
assign w43228 = ~w42699 & ~w43227;
assign w43229 = ~w42724 & ~w43226;
assign w43230 = ~w43228 & w43229;
assign w43231 = w43078 & w43097;
assign w43232 = ~w43022 & ~w43231;
assign w43233 = w42724 & ~w43232;
assign w43234 = w43019 & ~w43087;
assign w43235 = ~w43224 & ~w43234;
assign w43236 = ~w43225 & w43235;
assign w43237 = ~w43230 & ~w43233;
assign w43238 = w43236 & w43237;
assign w43239 = ~pi4873 & pi9040;
assign w43240 = ~pi4725 & ~pi9040;
assign w43241 = ~w43239 & ~w43240;
assign w43242 = pi2335 & ~w43241;
assign w43243 = ~pi2335 & w43241;
assign w43244 = ~w43242 & ~w43243;
assign w43245 = ~pi4658 & pi9040;
assign w43246 = ~pi4980 & ~pi9040;
assign w43247 = ~w43245 & ~w43246;
assign w43248 = pi2275 & ~w43247;
assign w43249 = ~pi2275 & w43247;
assign w43250 = ~w43248 & ~w43249;
assign w43251 = w43244 & w43250;
assign w43252 = ~pi4732 & pi9040;
assign w43253 = ~pi4756 & ~pi9040;
assign w43254 = ~w43252 & ~w43253;
assign w43255 = pi2312 & ~w43254;
assign w43256 = ~pi2312 & w43254;
assign w43257 = ~w43255 & ~w43256;
assign w43258 = w43250 & w43257;
assign w43259 = ~w43250 & ~w43257;
assign w43260 = ~w43258 & ~w43259;
assign w43261 = ~pi4756 & pi9040;
assign w43262 = ~pi4672 & ~pi9040;
assign w43263 = ~w43261 & ~w43262;
assign w43264 = pi2319 & ~w43263;
assign w43265 = ~pi2319 & w43263;
assign w43266 = ~w43264 & ~w43265;
assign w43267 = (~w43251 & w43260) | (~w43251 & w63991) | (w43260 & w63991);
assign w43268 = ~pi4722 & pi9040;
assign w43269 = ~pi4732 & ~pi9040;
assign w43270 = ~w43268 & ~w43269;
assign w43271 = pi2327 & ~w43270;
assign w43272 = ~pi2327 & w43270;
assign w43273 = ~w43271 & ~w43272;
assign w43274 = w43250 & w43273;
assign w43275 = ~w43267 & w66465;
assign w43276 = w43257 & ~w43273;
assign w43277 = ~w43251 & ~w43276;
assign w43278 = ~w43258 & ~w43266;
assign w43279 = ~w43277 & w43278;
assign w43280 = ~w43275 & ~w43279;
assign w43281 = ~w43257 & w43273;
assign w43282 = ~w43276 & ~w43281;
assign w43283 = w43244 & w43257;
assign w43284 = w43282 & ~w43283;
assign w43285 = ~w43250 & ~w43266;
assign w43286 = ~w43273 & w43285;
assign w43287 = w43284 & ~w43286;
assign w43288 = w43280 & ~w43287;
assign w43289 = ~pi4674 & pi9040;
assign w43290 = ~pi4969 & ~pi9040;
assign w43291 = ~w43289 & ~w43290;
assign w43292 = pi2324 & ~w43291;
assign w43293 = ~pi2324 & w43291;
assign w43294 = ~w43292 & ~w43293;
assign w43295 = ~w43288 & w43294;
assign w43296 = w43257 & ~w43266;
assign w43297 = ~w43257 & w43266;
assign w43298 = ~w43296 & ~w43297;
assign w43299 = ~w43250 & ~w43273;
assign w43300 = ~w43281 & ~w43299;
assign w43301 = ~w43294 & ~w43300;
assign w43302 = w43298 & w43301;
assign w43303 = w43250 & w43282;
assign w43304 = (~w43244 & w43302) | (~w43244 & w63993) | (w43302 & w63993);
assign w43305 = ~w43267 & w66466;
assign w43306 = ~w43266 & ~w43273;
assign w43307 = w43283 & w43306;
assign w43308 = (~w43244 & ~w43285) | (~w43244 & w66467) | (~w43285 & w66467);
assign w43309 = w43285 & w43308;
assign w43310 = w43244 & w43273;
assign w43311 = ~w43296 & w43310;
assign w43312 = w43260 & w43311;
assign w43313 = w43266 & ~w43312;
assign w43314 = (~w43266 & w43284) | (~w43266 & w66468) | (w43284 & w66468);
assign w43315 = ~w43294 & ~w43314;
assign w43316 = ~w43313 & w43315;
assign w43317 = ~w43307 & ~w43309;
assign w43318 = ~w43304 & w66469;
assign w43319 = ~w43316 & w43318;
assign w43320 = ~w43295 & w43319;
assign w43321 = pi2357 & ~w43320;
assign w43322 = ~pi2357 & w43320;
assign w43323 = ~w43321 & ~w43322;
assign w43324 = ~w43280 & w43281;
assign w43325 = ~w43274 & ~w43299;
assign w43326 = w43283 & ~w43325;
assign w43327 = ~w43258 & w43266;
assign w43328 = w43300 & w43327;
assign w43329 = w43273 & ~w43278;
assign w43330 = ~w43244 & ~w43260;
assign w43331 = ~w43329 & w43330;
assign w43332 = ~w43294 & ~w43326;
assign w43333 = ~w43328 & w43332;
assign w43334 = ~w43331 & w43333;
assign w43335 = w43285 & w43300;
assign w43336 = w43294 & ~w43335;
assign w43337 = ~w43257 & ~w43306;
assign w43338 = ~w43244 & ~w43296;
assign w43339 = ~w43337 & w43338;
assign w43340 = w43258 & w43306;
assign w43341 = ~w43337 & ~w43340;
assign w43342 = w43244 & ~w43341;
assign w43343 = w43266 & w43274;
assign w43344 = ~w43339 & ~w43343;
assign w43345 = w43336 & w43344;
assign w43346 = ~w43342 & w43345;
assign w43347 = ~w43334 & ~w43346;
assign w43348 = ~w43324 & ~w43347;
assign w43349 = ~pi2363 & w43348;
assign w43350 = pi2363 & ~w43348;
assign w43351 = ~w43349 & ~w43350;
assign w43352 = ~w43312 & ~w43340;
assign w43353 = ~w43305 & w43352;
assign w43354 = w43294 & ~w43353;
assign w43355 = ~w43250 & ~w43282;
assign w43356 = ~w43303 & ~w43355;
assign w43357 = ~w43314 & w43356;
assign w43358 = ~w43274 & w43308;
assign w43359 = ~w43315 & w43358;
assign w43360 = ~w43357 & w43359;
assign w43361 = w43250 & ~w43296;
assign w43362 = ~w43274 & ~w43311;
assign w43363 = ~w43361 & ~w43362;
assign w43364 = (~w43285 & w43300) | (~w43285 & w66470) | (w43300 & w66470);
assign w43365 = w43363 & ~w43364;
assign w43366 = w43251 & w43297;
assign w43367 = ~w43286 & ~w43343;
assign w43368 = ~w43366 & w43367;
assign w43369 = ~w43294 & ~w43368;
assign w43370 = ~w43294 & ~w43299;
assign w43371 = ~w43343 & ~w43370;
assign w43372 = ~w43244 & w43257;
assign w43373 = ~w43306 & w43372;
assign w43374 = (~w43307 & w43371) | (~w43307 & w66471) | (w43371 & w66471);
assign w43375 = ~w43365 & w43374;
assign w43376 = ~w43369 & w43375;
assign w43377 = ~w43354 & w43376;
assign w43378 = (pi2368 & ~w43377) | (pi2368 & w66472) | (~w43377 & w66472);
assign w43379 = w43377 & w66473;
assign w43380 = ~w43378 & ~w43379;
assign w43381 = w43244 & w43278;
assign w43382 = ~w43325 & w43381;
assign w43383 = w43266 & ~w43356;
assign w43384 = w43336 & ~w43382;
assign w43385 = ~w43383 & w43384;
assign w43386 = ~w43267 & ~w43273;
assign w43387 = ~w43294 & ~w43363;
assign w43388 = ~w43386 & w43387;
assign w43389 = ~w43385 & ~w43388;
assign w43390 = w43273 & ~w43298;
assign w43391 = ~w43301 & ~w43390;
assign w43392 = ~w43244 & ~w43325;
assign w43393 = ~w43391 & w43392;
assign w43394 = ~w43389 & ~w43393;
assign w43395 = ~pi2373 & w43394;
assign w43396 = pi2373 & ~w43394;
assign w43397 = ~w43395 & ~w43396;
assign w43398 = ~pi4719 & pi9040;
assign w43399 = ~pi4724 & ~pi9040;
assign w43400 = ~w43398 & ~w43399;
assign w43401 = pi2314 & ~w43400;
assign w43402 = ~pi2314 & w43400;
assign w43403 = ~w43401 & ~w43402;
assign w43404 = ~pi5054 & pi9040;
assign w43405 = ~pi4661 & ~pi9040;
assign w43406 = ~w43404 & ~w43405;
assign w43407 = pi2275 & ~w43406;
assign w43408 = ~pi2275 & w43406;
assign w43409 = ~w43407 & ~w43408;
assign w43410 = ~pi4871 & pi9040;
assign w43411 = ~pi4542 & ~pi9040;
assign w43412 = ~w43410 & ~w43411;
assign w43413 = pi2329 & ~w43412;
assign w43414 = ~pi2329 & w43412;
assign w43415 = ~w43413 & ~w43414;
assign w43416 = w43409 & ~w43415;
assign w43417 = ~pi4721 & pi9040;
assign w43418 = ~pi5054 & ~pi9040;
assign w43419 = ~w43417 & ~w43418;
assign w43420 = pi2324 & ~w43419;
assign w43421 = ~pi2324 & w43419;
assign w43422 = ~w43420 & ~w43421;
assign w43423 = w43403 & ~w43422;
assign w43424 = w43416 & ~w43423;
assign w43425 = w43403 & w43424;
assign w43426 = ~pi4867 & pi9040;
assign w43427 = ~pi4721 & ~pi9040;
assign w43428 = ~w43426 & ~w43427;
assign w43429 = pi2308 & ~w43428;
assign w43430 = ~pi2308 & w43428;
assign w43431 = ~w43429 & ~w43430;
assign w43432 = ~pi4725 & pi9040;
assign w43433 = ~pi4666 & ~pi9040;
assign w43434 = ~w43432 & ~w43433;
assign w43435 = pi2334 & ~w43434;
assign w43436 = ~pi2334 & w43434;
assign w43437 = ~w43435 & ~w43436;
assign w43438 = ~w43431 & ~w43437;
assign w43439 = w43415 & ~w43422;
assign w43440 = w43409 & w43439;
assign w43441 = ~w43403 & ~w43422;
assign w43442 = ~w43415 & w43441;
assign w43443 = ~w43440 & ~w43442;
assign w43444 = ~w43437 & w43443;
assign w43445 = ~w43438 & ~w43444;
assign w43446 = ~w43409 & w43415;
assign w43447 = w43422 & ~w43446;
assign w43448 = ~w43416 & ~w43447;
assign w43449 = ~w43403 & ~w43409;
assign w43450 = ~w43439 & ~w43449;
assign w43451 = w43448 & w43450;
assign w43452 = ~w43425 & ~w43451;
assign w43453 = ~w43445 & w43452;
assign w43454 = w43423 & w43446;
assign w43455 = ~w43424 & w43431;
assign w43456 = ~w43448 & w43455;
assign w43457 = ~w43431 & ~w43443;
assign w43458 = ~w43431 & ~w43446;
assign w43459 = ~w43403 & w43422;
assign w43460 = ~w43458 & w43459;
assign w43461 = w43437 & ~w43454;
assign w43462 = ~w43460 & w43461;
assign w43463 = ~w43456 & w43462;
assign w43464 = ~w43457 & w43463;
assign w43465 = ~w43453 & ~w43464;
assign w43466 = ~w43409 & ~w43415;
assign w43467 = w43459 & w43466;
assign w43468 = w43409 & w43422;
assign w43469 = ~w43467 & ~w43468;
assign w43470 = ~w43409 & w43439;
assign w43471 = w43469 & ~w43470;
assign w43472 = ~w43437 & ~w43471;
assign w43473 = ~w43409 & w43423;
assign w43474 = ~w43425 & ~w43473;
assign w43475 = ~w43472 & w43474;
assign w43476 = ~w43431 & ~w43475;
assign w43477 = ~w43465 & ~w43476;
assign w43478 = ~pi2349 & w43477;
assign w43479 = pi2349 & ~w43477;
assign w43480 = ~w43478 & ~w43479;
assign w43481 = ~w43403 & w43415;
assign w43482 = ~w43466 & ~w43481;
assign w43483 = w43422 & w43437;
assign w43484 = ~w43482 & w43483;
assign w43485 = ~w43469 & w43484;
assign w43486 = w43409 & ~w43423;
assign w43487 = ~w43437 & ~w43459;
assign w43488 = w43486 & ~w43487;
assign w43489 = w43423 & w43466;
assign w43490 = ~w43488 & ~w43489;
assign w43491 = w43431 & ~w43490;
assign w43492 = ~w43409 & ~w43431;
assign w43493 = w43481 & ~w43492;
assign w43494 = ~w43440 & ~w43481;
assign w43495 = ~w43493 & ~w43494;
assign w43496 = ~w43416 & ~w43470;
assign w43497 = (~w43403 & w43470) | (~w43403 & w66474) | (w43470 & w66474);
assign w43498 = w43415 & w43422;
assign w43499 = w43431 & ~w43481;
assign w43500 = w43498 & w43499;
assign w43501 = ~w43409 & w43500;
assign w43502 = ~w43495 & ~w43497;
assign w43503 = (~w43437 & ~w43502) | (~w43437 & w66475) | (~w43502 & w66475);
assign w43504 = ~w43447 & ~w43470;
assign w43505 = ~w43437 & ~w43504;
assign w43506 = w43437 & ~w43439;
assign w43507 = ~w43486 & w43506;
assign w43508 = (~w43447 & w43495) | (~w43447 & w66476) | (w43495 & w66476);
assign w43509 = ~w43505 & ~w43508;
assign w43510 = ~w43431 & ~w43459;
assign w43511 = ~w43509 & w43510;
assign w43512 = ~w43485 & ~w43491;
assign w43513 = ~w43503 & w43512;
assign w43514 = ~w43511 & w43513;
assign w43515 = pi2361 & ~w43514;
assign w43516 = ~pi2361 & w43514;
assign w43517 = ~w43515 & ~w43516;
assign w43518 = ~pi4659 & pi9040;
assign w43519 = ~pi4595 & ~pi9040;
assign w43520 = ~w43518 & ~w43519;
assign w43521 = pi2295 & ~w43520;
assign w43522 = ~pi2295 & w43520;
assign w43523 = ~w43521 & ~w43522;
assign w43524 = ~pi4542 & pi9040;
assign w43525 = ~pi4726 & ~pi9040;
assign w43526 = ~w43524 & ~w43525;
assign w43527 = pi2320 & ~w43526;
assign w43528 = ~pi2320 & w43526;
assign w43529 = ~w43527 & ~w43528;
assign w43530 = ~w43523 & w43529;
assign w43531 = w43523 & ~w43529;
assign w43532 = ~w43530 & ~w43531;
assign w43533 = ~pi4950 & pi9040;
assign w43534 = ~pi4722 & ~pi9040;
assign w43535 = ~w43533 & ~w43534;
assign w43536 = pi2304 & ~w43535;
assign w43537 = ~pi2304 & w43535;
assign w43538 = ~w43536 & ~w43537;
assign w43539 = ~pi4980 & pi9040;
assign w43540 = ~pi4540 & ~pi9040;
assign w43541 = ~w43539 & ~w43540;
assign w43542 = pi2326 & ~w43541;
assign w43543 = ~pi2326 & w43541;
assign w43544 = ~w43542 & ~w43543;
assign w43545 = ~w43523 & w43544;
assign w43546 = w43523 & ~w43544;
assign w43547 = ~w43545 & ~w43546;
assign w43548 = w43538 & w43547;
assign w43549 = ~pi4540 & pi9040;
assign w43550 = ~pi4873 & ~pi9040;
assign w43551 = ~w43549 & ~w43550;
assign w43552 = pi2333 & ~w43551;
assign w43553 = ~pi2333 & w43551;
assign w43554 = ~w43552 & ~w43553;
assign w43555 = ~w43544 & w43554;
assign w43556 = ~w43538 & w43555;
assign w43557 = w43555 & w66477;
assign w43558 = ~w43529 & ~w43538;
assign w43559 = w43531 & ~w43554;
assign w43560 = (w43544 & w43559) | (w43544 & w66478) | (w43559 & w66478);
assign w43561 = w43538 & w43554;
assign w43562 = w43530 & w43561;
assign w43563 = w43523 & w43538;
assign w43564 = w43529 & ~w43547;
assign w43565 = ~w43547 & w66479;
assign w43566 = w43563 & w43565;
assign w43567 = ~w43562 & ~w43566;
assign w43568 = ~pi4595 & pi9040;
assign w43569 = ~pi4871 & ~pi9040;
assign w43570 = ~w43568 & ~w43569;
assign w43571 = pi2313 & ~w43570;
assign w43572 = ~pi2313 & w43570;
assign w43573 = ~w43571 & ~w43572;
assign w43574 = ~w43523 & ~w43544;
assign w43575 = ~w43554 & w43574;
assign w43576 = w43574 & w66480;
assign w43577 = w43529 & w43554;
assign w43578 = w43574 & w43577;
assign w43579 = ~w43573 & ~w43578;
assign w43580 = ~w43576 & w43579;
assign w43581 = (~w43557 & ~w43548) | (~w43557 & w66481) | (~w43548 & w66481);
assign w43582 = ~w43560 & w43580;
assign w43583 = w43581 & w43582;
assign w43584 = w43567 & w43583;
assign w43585 = w43532 & w43556;
assign w43586 = ~w43523 & w43585;
assign w43587 = ~w43558 & ~w43577;
assign w43588 = w43545 & w43587;
assign w43589 = ~w43547 & w63994;
assign w43590 = ~w43538 & ~w43554;
assign w43591 = ~w43532 & w43590;
assign w43592 = ~w43588 & ~w43591;
assign w43593 = ~w43586 & w43592;
assign w43594 = w43523 & w43544;
assign w43595 = w43577 & w43594;
assign w43596 = w43573 & ~w43595;
assign w43597 = w43593 & w66482;
assign w43598 = w43531 & w43555;
assign w43599 = w43538 & ~w43598;
assign w43600 = ~w43575 & w43599;
assign w43601 = w43529 & ~w43545;
assign w43602 = w43587 & ~w43601;
assign w43603 = ~w43600 & w43602;
assign w43604 = (~w43603 & w43584) | (~w43603 & w66483) | (w43584 & w66483);
assign w43605 = ~pi2343 & w43604;
assign w43606 = pi2343 & ~w43604;
assign w43607 = ~w43605 & ~w43606;
assign w43608 = ~pi4594 & pi9040;
assign w43609 = ~pi4670 & ~pi9040;
assign w43610 = ~w43608 & ~w43609;
assign w43611 = pi2312 & ~w43610;
assign w43612 = ~pi2312 & w43610;
assign w43613 = ~w43611 & ~w43612;
assign w43614 = ~pi4975 & pi9040;
assign w43615 = ~pi4830 & ~pi9040;
assign w43616 = ~w43614 & ~w43615;
assign w43617 = pi2305 & ~w43616;
assign w43618 = ~pi2305 & w43616;
assign w43619 = ~w43617 & ~w43618;
assign w43620 = ~pi4592 & pi9040;
assign w43621 = ~pi4599 & ~pi9040;
assign w43622 = ~w43620 & ~w43621;
assign w43623 = pi2316 & ~w43622;
assign w43624 = ~pi2316 & w43622;
assign w43625 = ~w43623 & ~w43624;
assign w43626 = w43619 & w43625;
assign w43627 = ~pi4668 & pi9040;
assign w43628 = ~pi4955 & ~pi9040;
assign w43629 = ~w43627 & ~w43628;
assign w43630 = pi2322 & ~w43629;
assign w43631 = ~pi2322 & w43629;
assign w43632 = ~w43630 & ~w43631;
assign w43633 = ~pi4723 & pi9040;
assign w43634 = ~pi4594 & ~pi9040;
assign w43635 = ~w43633 & ~w43634;
assign w43636 = pi2327 & ~w43635;
assign w43637 = ~pi2327 & w43635;
assign w43638 = ~w43636 & ~w43637;
assign w43639 = w43632 & w43638;
assign w43640 = ~w43632 & w43638;
assign w43641 = ~w43625 & w43640;
assign w43642 = ~w43639 & ~w43641;
assign w43643 = ~w43632 & ~w43638;
assign w43644 = w43625 & w43643;
assign w43645 = w43642 & ~w43644;
assign w43646 = (w43626 & ~w43642) | (w43626 & w66484) | (~w43642 & w66484);
assign w43647 = ~w43619 & w43632;
assign w43648 = w43619 & ~w43632;
assign w43649 = ~w43647 & ~w43648;
assign w43650 = ~w43639 & ~w43649;
assign w43651 = ~pi4541 & pi9040;
assign w43652 = ~pi4664 & ~pi9040;
assign w43653 = ~w43651 & ~w43652;
assign w43654 = pi2298 & ~w43653;
assign w43655 = ~pi2298 & w43653;
assign w43656 = ~w43654 & ~w43655;
assign w43657 = ~w43625 & ~w43656;
assign w43658 = ~w43638 & ~w43656;
assign w43659 = ~w43657 & ~w43658;
assign w43660 = ~w43650 & ~w43659;
assign w43661 = ~w43625 & w43632;
assign w43662 = ~w43638 & w43661;
assign w43663 = w43661 & w66485;
assign w43664 = ~w43619 & ~w43625;
assign w43665 = w43638 & w43664;
assign w43666 = w43656 & ~w43665;
assign w43667 = ~w43663 & w43666;
assign w43668 = ~w43660 & ~w43667;
assign w43669 = ~w43613 & ~w43646;
assign w43670 = ~w43668 & w43669;
assign w43671 = ~w43619 & w43625;
assign w43672 = w43639 & w43671;
assign w43673 = w43613 & ~w43672;
assign w43674 = w43649 & w43657;
assign w43675 = w43673 & ~w43674;
assign w43676 = w43625 & ~w43638;
assign w43677 = ~w43648 & ~w43676;
assign w43678 = w43648 & w43676;
assign w43679 = w43656 & ~w43677;
assign w43680 = ~w43678 & w43679;
assign w43681 = w43675 & ~w43680;
assign w43682 = ~w43670 & ~w43681;
assign w43683 = ~w43656 & ~w43678;
assign w43684 = ~w43626 & ~w43643;
assign w43685 = ~w43677 & w43684;
assign w43686 = w43656 & ~w43685;
assign w43687 = w43619 & ~w43656;
assign w43688 = ~w43664 & ~w43687;
assign w43689 = w43639 & ~w43688;
assign w43690 = w43686 & ~w43689;
assign w43691 = ~w43638 & w43664;
assign w43692 = w43664 & w43643;
assign w43693 = w43690 & ~w43692;
assign w43694 = ~w43683 & ~w43693;
assign w43695 = ~w43682 & ~w43694;
assign w43696 = pi2341 & w43695;
assign w43697 = ~pi2341 & ~w43695;
assign w43698 = ~w43696 & ~w43697;
assign w43699 = ~pi4860 & pi9040;
assign w43700 = ~pi4663 & ~pi9040;
assign w43701 = ~w43699 & ~w43700;
assign w43702 = pi2328 & ~w43701;
assign w43703 = ~pi2328 & w43701;
assign w43704 = ~w43702 & ~w43703;
assign w43705 = ~pi4823 & pi9040;
assign w43706 = ~pi4860 & ~pi9040;
assign w43707 = ~w43705 & ~w43706;
assign w43708 = pi2291 & ~w43707;
assign w43709 = ~pi2291 & w43707;
assign w43710 = ~w43708 & ~w43709;
assign w43711 = ~w43704 & ~w43710;
assign w43712 = ~pi4543 & pi9040;
assign w43713 = ~pi4872 & ~pi9040;
assign w43714 = ~w43712 & ~w43713;
assign w43715 = pi2310 & ~w43714;
assign w43716 = ~pi2310 & w43714;
assign w43717 = ~w43715 & ~w43716;
assign w43718 = ~pi4600 & pi9040;
assign w43719 = ~pi4728 & ~pi9040;
assign w43720 = ~w43718 & ~w43719;
assign w43721 = pi2296 & ~w43720;
assign w43722 = ~pi2296 & w43720;
assign w43723 = ~w43721 & ~w43722;
assign w43724 = w43717 & ~w43723;
assign w43725 = w43711 & w43724;
assign w43726 = ~w43710 & w43723;
assign w43727 = ~pi4663 & pi9040;
assign w43728 = ~pi4592 & ~pi9040;
assign w43729 = ~w43727 & ~w43728;
assign w43730 = pi2323 & ~w43729;
assign w43731 = ~pi2323 & w43729;
assign w43732 = ~w43730 & ~w43731;
assign w43733 = w43704 & w43732;
assign w43734 = w43726 & w43733;
assign w43735 = w43710 & ~w43732;
assign w43736 = ~w43704 & w43723;
assign w43737 = w43717 & w43736;
assign w43738 = w43735 & w43737;
assign w43739 = ~pi4664 & pi9040;
assign w43740 = ~pi4543 & ~pi9040;
assign w43741 = ~w43739 & ~w43740;
assign w43742 = pi2315 & ~w43741;
assign w43743 = ~pi2315 & w43741;
assign w43744 = ~w43742 & ~w43743;
assign w43745 = ~w43710 & ~w43732;
assign w43746 = ~w43717 & w43723;
assign w43747 = w43704 & w43717;
assign w43748 = ~w43746 & ~w43747;
assign w43749 = w43745 & ~w43748;
assign w43750 = ~w43717 & ~w43723;
assign w43751 = w43704 & w43710;
assign w43752 = w43750 & w43751;
assign w43753 = ~w43704 & ~w43726;
assign w43754 = ~w43717 & ~w43753;
assign w43755 = w43704 & ~w43723;
assign w43756 = ~w43736 & ~w43755;
assign w43757 = w43717 & ~w43756;
assign w43758 = ~w43711 & ~w43751;
assign w43759 = w43750 & w43758;
assign w43760 = w43732 & ~w43754;
assign w43761 = ~w43757 & ~w43759;
assign w43762 = w43760 & w43761;
assign w43763 = ~w43744 & ~w43752;
assign w43764 = ~w43738 & w43763;
assign w43765 = ~w43749 & w43764;
assign w43766 = ~w43762 & w43765;
assign w43767 = ~w43710 & w43717;
assign w43768 = w43710 & ~w43724;
assign w43769 = ~w43768 & w63424;
assign w43770 = ~w43704 & w43745;
assign w43771 = (w43717 & w43769) | (w43717 & w63995) | (w43769 & w63995);
assign w43772 = ~w43759 & ~w43771;
assign w43773 = w43704 & w43746;
assign w43774 = w43710 & w43746;
assign w43775 = w43717 & w43726;
assign w43776 = ~w43774 & ~w43775;
assign w43777 = (~w43773 & ~w43776) | (~w43773 & w63996) | (~w43776 & w63996);
assign w43778 = w43732 & ~w43777;
assign w43779 = w43772 & ~w43778;
assign w43780 = w43717 & ~w43751;
assign w43781 = (~w43732 & w43751) | (~w43732 & w66486) | (w43751 & w66486);
assign w43782 = ~w43754 & w43781;
assign w43783 = w43744 & ~w43782;
assign w43784 = w43779 & w43783;
assign w43785 = ~w43725 & ~w43734;
assign w43786 = (w43785 & w43784) | (w43785 & w66487) | (w43784 & w66487);
assign w43787 = pi2336 & ~w43786;
assign w43788 = ~pi2336 & w43786;
assign w43789 = ~w43787 & ~w43788;
assign w43790 = ~pi4667 & pi9040;
assign w43791 = ~pi4538 & ~pi9040;
assign w43792 = ~w43790 & ~w43791;
assign w43793 = pi2313 & ~w43792;
assign w43794 = ~pi2313 & w43792;
assign w43795 = ~w43793 & ~w43794;
assign w43796 = ~pi4727 & pi9040;
assign w43797 = ~pi4864 & ~pi9040;
assign w43798 = ~w43796 & ~w43797;
assign w43799 = pi2330 & ~w43798;
assign w43800 = ~pi2330 & w43798;
assign w43801 = ~w43799 & ~w43800;
assign w43802 = w43795 & w43801;
assign w43803 = ~pi4872 & pi9040;
assign w43804 = ~pi4598 & ~pi9040;
assign w43805 = ~w43803 & ~w43804;
assign w43806 = pi2296 & ~w43805;
assign w43807 = ~pi2296 & w43805;
assign w43808 = ~w43806 & ~w43807;
assign w43809 = w43802 & w43808;
assign w43810 = ~pi4728 & pi9040;
assign w43811 = ~pi4514 & ~pi9040;
assign w43812 = ~w43810 & ~w43811;
assign w43813 = pi2332 & ~w43812;
assign w43814 = ~pi2332 & w43812;
assign w43815 = ~w43813 & ~w43814;
assign w43816 = (w43815 & ~w43802) | (w43815 & w43913) | (~w43802 & w43913);
assign w43817 = ~pi4598 & pi9040;
assign w43818 = ~pi4763 & ~pi9040;
assign w43819 = ~w43817 & ~w43818;
assign w43820 = pi2326 & ~w43819;
assign w43821 = ~pi2326 & w43819;
assign w43822 = ~w43820 & ~w43821;
assign w43823 = ~w43808 & ~w43822;
assign w43824 = w43808 & w43822;
assign w43825 = ~w43823 & ~w43824;
assign w43826 = w43801 & w43825;
assign w43827 = w43816 & w43826;
assign w43828 = ~w43801 & w43808;
assign w43829 = ~w43795 & w43828;
assign w43830 = w43815 & ~w43829;
assign w43831 = ~w43795 & ~w43822;
assign w43832 = w43815 & ~w43831;
assign w43833 = w43802 & w43823;
assign w43834 = ~w43832 & ~w43833;
assign w43835 = ~w43830 & ~w43834;
assign w43836 = ~pi4955 & pi9040;
assign w43837 = ~pi4660 & ~pi9040;
assign w43838 = ~w43836 & ~w43837;
assign w43839 = pi2310 & ~w43838;
assign w43840 = ~pi2310 & w43838;
assign w43841 = ~w43839 & ~w43840;
assign w43842 = w43795 & ~w43801;
assign w43843 = ~w43815 & w43842;
assign w43844 = w43795 & ~w43808;
assign w43845 = ~w43822 & ~w43844;
assign w43846 = ~w43795 & w43801;
assign w43847 = w43845 & ~w43846;
assign w43848 = w43830 & w43847;
assign w43849 = ~w43795 & w43826;
assign w43850 = w43841 & ~w43843;
assign w43851 = ~w43848 & w43850;
assign w43852 = ~w43849 & w43851;
assign w43853 = ~w43844 & w63997;
assign w43854 = ~w43815 & w43853;
assign w43855 = ~w43801 & w43822;
assign w43856 = ~w43795 & w43855;
assign w43857 = ~w43854 & ~w43856;
assign w43858 = w43795 & w43815;
assign w43859 = ~w43802 & ~w43808;
assign w43860 = ~w43855 & w43859;
assign w43861 = w43859 & w66488;
assign w43862 = w43822 & w43844;
assign w43863 = ~w43808 & w43831;
assign w43864 = ~w43862 & ~w43863;
assign w43865 = w43801 & ~w43864;
assign w43866 = (~w43841 & w43864) | (~w43841 & w66489) | (w43864 & w66489);
assign w43867 = ~w43824 & ~w43829;
assign w43868 = ~w43795 & ~w43815;
assign w43869 = ~w43858 & ~w43868;
assign w43870 = ~w43867 & ~w43869;
assign w43871 = ~w43861 & ~w43870;
assign w43872 = w43871 & w66490;
assign w43873 = ~w43852 & ~w43872;
assign w43874 = ~w43827 & ~w43835;
assign w43875 = ~w43873 & w43874;
assign w43876 = pi2340 & w43875;
assign w43877 = ~pi2340 & ~w43875;
assign w43878 = ~w43876 & ~w43877;
assign w43879 = ~w43441 & ~w43492;
assign w43880 = w43450 & ~w43879;
assign w43881 = ~w43450 & w43499;
assign w43882 = w43468 & w43481;
assign w43883 = ~w43425 & ~w43882;
assign w43884 = ~w43880 & ~w43881;
assign w43885 = w43883 & w43884;
assign w43886 = ~w43495 & w43885;
assign w43887 = w43437 & ~w43886;
assign w43888 = w43416 & ~w43459;
assign w43889 = ~w43454 & ~w43467;
assign w43890 = ~w43882 & ~w43888;
assign w43891 = w43889 & w43890;
assign w43892 = w43438 & ~w43891;
assign w43893 = w43487 & w43493;
assign w43894 = w43431 & ~w43437;
assign w43895 = ~w43439 & w43894;
assign w43896 = w43891 & w43895;
assign w43897 = ~w43892 & ~w43893;
assign w43898 = ~w43896 & w43897;
assign w43899 = ~w43887 & w43898;
assign w43900 = pi2375 & ~w43899;
assign w43901 = ~pi2375 & w43899;
assign w43902 = ~w43900 & ~w43901;
assign w43903 = ~w43815 & ~w43857;
assign w43904 = (~w43828 & w43864) | (~w43828 & w66491) | (w43864 & w66491);
assign w43905 = w43822 & ~w43904;
assign w43906 = ~w43903 & ~w43905;
assign w43907 = w43841 & ~w43906;
assign w43908 = w43822 & ~w43846;
assign w43909 = (~w43841 & w43844) | (~w43841 & w66492) | (w43844 & w66492);
assign w43910 = ~w43802 & ~w43909;
assign w43911 = ~w43815 & ~w43908;
assign w43912 = ~w43910 & w43911;
assign w43913 = ~w43808 & w43815;
assign w43914 = w43855 & w43913;
assign w43915 = ~w43801 & ~w43815;
assign w43916 = w43831 & w43915;
assign w43917 = ~w43914 & ~w43916;
assign w43918 = w43824 & w43846;
assign w43919 = (~w43841 & ~w43917) | (~w43841 & w66493) | (~w43917 & w66493);
assign w43920 = ~w43801 & w43864;
assign w43921 = w43795 & w43824;
assign w43922 = ~w43831 & ~w43921;
assign w43923 = w43917 & ~w43922;
assign w43924 = w43920 & w43923;
assign w43925 = ~w43860 & w43922;
assign w43926 = ~w43865 & w43925;
assign w43927 = w43815 & ~w43866;
assign w43928 = ~w43926 & w43927;
assign w43929 = ~w43912 & ~w43919;
assign w43930 = ~w43924 & w43929;
assign w43931 = ~w43928 & w43930;
assign w43932 = ~w43907 & w43931;
assign w43933 = pi2348 & ~w43932;
assign w43934 = ~pi2348 & w43932;
assign w43935 = ~w43933 & ~w43934;
assign w43936 = w43825 & w43842;
assign w43937 = w43801 & w43845;
assign w43938 = ~w43936 & ~w43937;
assign w43939 = w43913 & ~w43938;
assign w43940 = w43816 & ~w43856;
assign w43941 = ~w43863 & w43940;
assign w43942 = ~w43825 & ~w43842;
assign w43943 = ~w43936 & ~w43942;
assign w43944 = ~w43815 & ~w43943;
assign w43945 = (~w43841 & w43944) | (~w43841 & w66494) | (w43944 & w66494);
assign w43946 = ~w43854 & ~w43915;
assign w43947 = w43942 & ~w43946;
assign w43948 = ~w43815 & ~w43853;
assign w43949 = w43809 & w43948;
assign w43950 = ~w43823 & ~w43940;
assign w43951 = ~w43860 & ~w43950;
assign w43952 = (w43841 & ~w43825) | (w43841 & w66495) | (~w43825 & w66495);
assign w43953 = ~w43949 & w43952;
assign w43954 = ~w43947 & w43953;
assign w43955 = ~w43951 & w43954;
assign w43956 = ~w43815 & w43849;
assign w43957 = ~w43939 & ~w43956;
assign w43958 = (w43957 & w43955) | (w43957 & w66496) | (w43955 & w66496);
assign w43959 = pi2353 & w43958;
assign w43960 = ~pi2353 & ~w43958;
assign w43961 = ~w43959 & ~w43960;
assign w43962 = (w43732 & w43768) | (w43732 & w66497) | (w43768 & w66497);
assign w43963 = ~w43779 & w43962;
assign w43964 = ~w43717 & ~w43770;
assign w43965 = w43717 & ~w43735;
assign w43966 = ~w43757 & ~w43965;
assign w43967 = ~w43964 & w43966;
assign w43968 = w43733 & w43767;
assign w43969 = ~w43758 & ~w43767;
assign w43970 = ~w43758 & w66498;
assign w43971 = w43745 & w43747;
assign w43972 = ~w43725 & ~w43971;
assign w43973 = w43745 & w43972;
assign w43974 = w43744 & ~w43968;
assign w43975 = ~w43970 & w43974;
assign w43976 = ~w43973 & w43975;
assign w43977 = ~w43736 & ~w43752;
assign w43978 = w43781 & ~w43977;
assign w43979 = (w43732 & w43769) | (w43732 & w66499) | (w43769 & w66499);
assign w43980 = ~w43744 & w43972;
assign w43981 = ~w43978 & w43980;
assign w43982 = ~w43979 & w43981;
assign w43983 = (~w43967 & w43982) | (~w43967 & w66500) | (w43982 & w66500);
assign w43984 = ~w43963 & w43983;
assign w43985 = pi2337 & ~w43984;
assign w43986 = ~pi2337 & w43984;
assign w43987 = ~w43985 & ~w43986;
assign w43988 = ~w43723 & w43971;
assign w43989 = w43746 & w43751;
assign w43990 = w43733 & w43750;
assign w43991 = w43711 & w43723;
assign w43992 = ~w43990 & ~w43991;
assign w43993 = (w43732 & ~w43726) | (w43732 & w66501) | (~w43726 & w66501);
assign w43994 = ~w43724 & ~w43732;
assign w43995 = ~w43993 & ~w43994;
assign w43996 = ~w43759 & ~w43989;
assign w43997 = w43996 & w66502;
assign w43998 = w43744 & ~w43997;
assign w43999 = ~w43746 & ~w43992;
assign w44000 = ~w43772 & w43999;
assign w44001 = ~w43717 & ~w43736;
assign w44002 = w43993 & ~w44001;
assign w44003 = (w43732 & ~w43747) | (w43732 & w63998) | (~w43747 & w63998);
assign w44004 = w43756 & ~w43780;
assign w44005 = ~w44003 & w44004;
assign w44006 = ~w44002 & ~w44005;
assign w44007 = (~w43744 & w44005) | (~w43744 & w66503) | (w44005 & w66503);
assign w44008 = ~w43988 & ~w44007;
assign w44009 = ~w43998 & w44008;
assign w44010 = ~w44000 & w44009;
assign w44011 = pi2339 & ~w44010;
assign w44012 = ~pi2339 & w44010;
assign w44013 = ~w44011 & ~w44012;
assign w44014 = ~w43732 & w43776;
assign w44015 = ~w43962 & ~w44014;
assign w44016 = (~w43744 & w43992) | (~w43744 & w66504) | (w43992 & w66504);
assign w44017 = ~w44015 & w66505;
assign w44018 = w43735 & ~w43748;
assign w44019 = ~w43725 & ~w43774;
assign w44020 = w44003 & w44019;
assign w44021 = w43745 & ~w43773;
assign w44022 = ~w43988 & w44021;
assign w44023 = ~w44018 & ~w44020;
assign w44024 = (w43744 & ~w44023) | (w43744 & w63999) | (~w44023 & w63999);
assign w44025 = ~w44000 & w44024;
assign w44026 = ~w43735 & w43969;
assign w44027 = ~w44006 & w44026;
assign w44028 = (~w44027 & w44025) | (~w44027 & w66506) | (w44025 & w66506);
assign w44029 = pi2338 & w44028;
assign w44030 = ~pi2338 & ~w44028;
assign w44031 = ~w44029 & ~w44030;
assign w44032 = w43561 & w43601;
assign w44033 = w43545 & w43558;
assign w44034 = ~w43554 & ~w44033;
assign w44035 = w43554 & ~w43594;
assign w44036 = (~w43538 & w43594) | (~w43538 & w43590) | (w43594 & w43590);
assign w44037 = ~w43564 & ~w43588;
assign w44038 = (~w44034 & ~w44037) | (~w44034 & w63425) | (~w44037 & w63425);
assign w44039 = w43558 & ~w43594;
assign w44040 = (~w44038 & w66507) | (~w44038 & w66508) | (w66507 & w66508);
assign w44041 = ~w43529 & ~w43546;
assign w44042 = w43590 & ~w44041;
assign w44043 = ~w43564 & w44042;
assign w44044 = w43538 & w43544;
assign w44045 = w43573 & ~w44044;
assign w44046 = (w43593 & w64001) | (w43593 & w64002) | (w64001 & w64002);
assign w44047 = ~w44045 & ~w44046;
assign w44048 = ~w43574 & ~w44038;
assign w44049 = ~w43587 & ~w44038;
assign w44050 = (w43573 & w44038) | (w43573 & w64003) | (w44038 & w64003);
assign w44051 = ~w44049 & w44050;
assign w44052 = ~w44040 & ~w44043;
assign w44053 = ~w44047 & ~w44051;
assign w44054 = w44053 & w66509;
assign w44055 = (~pi2345 & ~w44053) | (~pi2345 & w66510) | (~w44053 & w66510);
assign w44056 = ~w44054 & ~w44055;
assign w44057 = w43544 & w43554;
assign w44058 = w43532 & w44057;
assign w44059 = ~w43547 & w43590;
assign w44060 = w43547 & w63427;
assign w44061 = ~w44059 & ~w44060;
assign w44062 = ~w43532 & ~w44061;
assign w44063 = ~w43557 & ~w44058;
assign w44064 = ~w44062 & w44063;
assign w44065 = ~w44062 & w66511;
assign w44066 = w44048 & w44064;
assign w44067 = w43580 & ~w43586;
assign w44068 = ~w44066 & w44067;
assign w44069 = ~w43576 & ~w44058;
assign w44070 = ~w43538 & ~w44069;
assign w44071 = w43567 & ~w44070;
assign w44072 = (~w44068 & w66512) | (~w44068 & w66513) | (w66512 & w66513);
assign w44073 = (w44068 & w66514) | (w44068 & w66515) | (w66514 & w66515);
assign w44074 = ~w44072 & ~w44073;
assign w44075 = w43561 & ~w44064;
assign w44076 = w43532 & w44035;
assign w44077 = ~w43538 & ~w43546;
assign w44078 = (w44077 & w43564) | (w44077 & w66516) | (w43564 & w66516);
assign w44079 = ~w43529 & ~w43574;
assign w44080 = w43599 & w44079;
assign w44081 = w43573 & ~w44076;
assign w44082 = ~w44080 & w44081;
assign w44083 = ~w44078 & w44082;
assign w44084 = ~w43531 & w44077;
assign w44085 = ~w43557 & ~w44084;
assign w44086 = ~w43600 & w44085;
assign w44087 = ~w43573 & ~w43595;
assign w44088 = ~w43565 & w44087;
assign w44089 = ~w44086 & w44088;
assign w44090 = ~w44083 & ~w44089;
assign w44091 = ~w43585 & ~w44090;
assign w44092 = (pi2362 & ~w44091) | (pi2362 & w66517) | (~w44091 & w66517);
assign w44093 = w44091 & w66518;
assign w44094 = ~w44092 & ~w44093;
assign w44095 = w43826 & w66519;
assign w44096 = w43830 & ~w43862;
assign w44097 = ~w43828 & ~w43844;
assign w44098 = w43948 & ~w44097;
assign w44099 = ~w44096 & ~w44098;
assign w44100 = ~w43937 & ~w44099;
assign w44101 = ~w43841 & ~w44100;
assign w44102 = ~w43920 & ~w43946;
assign w44103 = ~w43824 & w43834;
assign w44104 = w43808 & ~w43842;
assign w44105 = ~w43844 & ~w44104;
assign w44106 = ~w43833 & ~w43868;
assign w44107 = ~w44105 & w44106;
assign w44108 = w43841 & ~w44103;
assign w44109 = ~w44107 & w44108;
assign w44110 = ~w43861 & ~w44095;
assign w44111 = ~w44102 & w44110;
assign w44112 = ~w44109 & w44111;
assign w44113 = ~w44101 & w44112;
assign w44114 = pi2359 & ~w44113;
assign w44115 = ~pi2359 & w44113;
assign w44116 = ~w44114 & ~w44115;
assign w44117 = ~pi4763 & pi9040;
assign w44118 = ~pi4975 & ~pi9040;
assign w44119 = ~w44117 & ~w44118;
assign w44120 = pi2328 & ~w44119;
assign w44121 = ~pi2328 & w44119;
assign w44122 = ~w44120 & ~w44121;
assign w44123 = ~pi4599 & pi9040;
assign w44124 = ~pi4541 & ~pi9040;
assign w44125 = ~w44123 & ~w44124;
assign w44126 = pi2301 & ~w44125;
assign w44127 = ~pi2301 & w44125;
assign w44128 = ~w44126 & ~w44127;
assign w44129 = w44122 & w44128;
assign w44130 = ~pi4864 & pi9040;
assign w44131 = ~pi4858 & ~pi9040;
assign w44132 = ~w44130 & ~w44131;
assign w44133 = pi2307 & ~w44132;
assign w44134 = ~pi2307 & w44132;
assign w44135 = ~w44133 & ~w44134;
assign w44136 = ~w44122 & w44135;
assign w44137 = ~w44129 & ~w44136;
assign w44138 = ~pi4858 & pi9040;
assign w44139 = ~pi4668 & ~pi9040;
assign w44140 = ~w44138 & ~w44139;
assign w44141 = pi2316 & ~w44140;
assign w44142 = ~pi2316 & w44140;
assign w44143 = ~w44141 & ~w44142;
assign w44144 = ~pi4660 & pi9040;
assign w44145 = ~pi4667 & ~pi9040;
assign w44146 = ~w44144 & ~w44145;
assign w44147 = pi2315 & ~w44146;
assign w44148 = ~pi2315 & w44146;
assign w44149 = ~w44147 & ~w44148;
assign w44150 = w44143 & ~w44149;
assign w44151 = ~w44122 & ~w44128;
assign w44152 = w44150 & ~w44151;
assign w44153 = w44137 & w44152;
assign w44154 = ~w44143 & w44149;
assign w44155 = ~w44150 & ~w44154;
assign w44156 = ~w44128 & w44155;
assign w44157 = ~w44122 & w44149;
assign w44158 = w44143 & w44157;
assign w44159 = ~w44151 & ~w44158;
assign w44160 = ~w44156 & ~w44159;
assign w44161 = ~w44122 & ~w44143;
assign w44162 = ~w44128 & ~w44149;
assign w44163 = ~w44161 & ~w44162;
assign w44164 = ~w44143 & ~w44149;
assign w44165 = ~w44122 & w44128;
assign w44166 = w44164 & w44165;
assign w44167 = w44155 & w64005;
assign w44168 = ~w44166 & ~w44167;
assign w44169 = (~w44163 & w44167) | (~w44163 & w66520) | (w44167 & w66520);
assign w44170 = ~w44137 & w44150;
assign w44171 = (~w44170 & ~w44160) | (~w44170 & w64006) | (~w44160 & w64006);
assign w44172 = ~w44169 & w44171;
assign w44173 = w44171 & w66521;
assign w44174 = w44129 & w44164;
assign w44175 = ~w44157 & ~w44174;
assign w44176 = ~w44160 & ~w44175;
assign w44177 = ~pi4514 & pi9040;
assign w44178 = ~pi4727 & ~pi9040;
assign w44179 = ~w44177 & ~w44178;
assign w44180 = pi2305 & ~w44179;
assign w44181 = ~pi2305 & w44179;
assign w44182 = ~w44180 & ~w44181;
assign w44183 = ~w44153 & w44182;
assign w44184 = ~w44176 & w44183;
assign w44185 = ~w44173 & w44184;
assign w44186 = w44122 & w44143;
assign w44187 = ~w44161 & ~w44186;
assign w44188 = ~w44135 & ~w44187;
assign w44189 = w44128 & w44149;
assign w44190 = ~w44135 & w44189;
assign w44191 = ~w44182 & ~w44190;
assign w44192 = ~w44188 & w44191;
assign w44193 = w44172 & w44192;
assign w44194 = ~w44185 & ~w44193;
assign w44195 = ~pi2344 & w44194;
assign w44196 = pi2344 & ~w44194;
assign w44197 = ~w44195 & ~w44196;
assign w44198 = w43403 & w43409;
assign w44199 = ~w43449 & ~w44198;
assign w44200 = w43423 & w43431;
assign w44201 = ~w43498 & ~w44199;
assign w44202 = ~w44200 & w44201;
assign w44203 = ~w43449 & w43498;
assign w44204 = ~w43458 & w44203;
assign w44205 = ~w44202 & ~w44204;
assign w44206 = ~w43437 & ~w44205;
assign w44207 = ~w43440 & ~w43484;
assign w44208 = ~w43431 & ~w44207;
assign w44209 = w43437 & w43489;
assign w44210 = w43431 & ~w43496;
assign w44211 = ~w43444 & w44210;
assign w44212 = ~w43500 & ~w44209;
assign w44213 = ~w44208 & w44212;
assign w44214 = ~w44211 & w44213;
assign w44215 = ~w44206 & w44214;
assign w44216 = ~pi2382 & ~w44215;
assign w44217 = pi2382 & w44215;
assign w44218 = ~w44216 & ~w44217;
assign w44219 = w43640 & w43687;
assign w44220 = ~w43692 & ~w44219;
assign w44221 = w43664 & w43640;
assign w44222 = w44220 & ~w44221;
assign w44223 = ~w43657 & ~w44222;
assign w44224 = ~w43661 & ~w43676;
assign w44225 = ~w43656 & ~w43662;
assign w44226 = w43619 & ~w44224;
assign w44227 = ~w44225 & w44226;
assign w44228 = w43632 & w43671;
assign w44229 = w43658 & w43671;
assign w44230 = ~w43613 & ~w44229;
assign w44231 = ~w43649 & w66522;
assign w44232 = w43619 & ~w43625;
assign w44233 = ~w43657 & ~w44232;
assign w44234 = w43639 & ~w44233;
assign w44235 = ~w44231 & ~w44234;
assign w44236 = ~w43626 & ~w43665;
assign w44237 = w43638 & ~w44236;
assign w44238 = ~w44235 & w44237;
assign w44239 = ~w44228 & w44230;
assign w44240 = w44220 & w44239;
assign w44241 = ~w44227 & w44240;
assign w44242 = ~w44238 & w44241;
assign w44243 = w43613 & ~w44221;
assign w44244 = w43626 & ~w43638;
assign w44245 = ~w43691 & ~w44244;
assign w44246 = w43632 & ~w44245;
assign w44247 = (~w43643 & w44233) | (~w43643 & w66523) | (w44233 & w66523);
assign w44248 = w43687 & ~w44247;
assign w44249 = ~w43643 & w43656;
assign w44250 = ~w43661 & w44249;
assign w44251 = ~w44231 & w44250;
assign w44252 = w44243 & ~w44246;
assign w44253 = w44252 & w66524;
assign w44254 = (~w44223 & w44242) | (~w44223 & w66525) | (w44242 & w66525);
assign w44255 = ~pi2351 & w44254;
assign w44256 = pi2351 & ~w44254;
assign w44257 = ~w44255 & ~w44256;
assign w44258 = w43683 & ~w43685;
assign w44259 = w43656 & ~w43662;
assign w44260 = ~w44258 & ~w44259;
assign w44261 = ~w43619 & w44224;
assign w44262 = ~w44261 & w66526;
assign w44263 = w43690 & w44262;
assign w44264 = (~w43656 & w44261) | (~w43656 & w66527) | (w44261 & w66527);
assign w44265 = ~w43641 & ~w43663;
assign w44266 = w43673 & w44265;
assign w44267 = ~w44264 & w44266;
assign w44268 = ~w44263 & w44267;
assign w44269 = w43645 & w43686;
assign w44270 = ~w43689 & w44230;
assign w44271 = ~w44269 & w44270;
assign w44272 = (~w44260 & w44268) | (~w44260 & w66528) | (w44268 & w66528);
assign w44273 = ~pi2374 & w44272;
assign w44274 = pi2374 & ~w44272;
assign w44275 = ~w44273 & ~w44274;
assign w44276 = ~pi4669 & pi9040;
assign w44277 = ~pi4950 & ~pi9040;
assign w44278 = ~w44276 & ~w44277;
assign w44279 = pi2334 & ~w44278;
assign w44280 = ~pi2334 & w44278;
assign w44281 = ~w44279 & ~w44280;
assign w44282 = ~pi4672 & pi9040;
assign w44283 = ~pi4658 & ~pi9040;
assign w44284 = ~w44282 & ~w44283;
assign w44285 = pi2320 & ~w44284;
assign w44286 = ~pi2320 & w44284;
assign w44287 = ~w44285 & ~w44286;
assign w44288 = ~w44281 & ~w44287;
assign w44289 = ~pi4614 & pi9040;
assign w44290 = ~pi4659 & ~pi9040;
assign w44291 = ~w44289 & ~w44290;
assign w44292 = pi2329 & ~w44291;
assign w44293 = ~pi2329 & w44291;
assign w44294 = ~w44292 & ~w44293;
assign w44295 = ~pi4724 & pi9040;
assign w44296 = ~pi4544 & ~pi9040;
assign w44297 = ~w44295 & ~w44296;
assign w44298 = pi2325 & ~w44297;
assign w44299 = ~pi2325 & w44297;
assign w44300 = ~w44298 & ~w44299;
assign w44301 = ~w44294 & ~w44300;
assign w44302 = w44288 & w44301;
assign w44303 = ~pi4726 & pi9040;
assign w44304 = ~pi4674 & ~pi9040;
assign w44305 = ~w44303 & ~w44304;
assign w44306 = pi2318 & ~w44305;
assign w44307 = ~pi2318 & w44305;
assign w44308 = ~w44306 & ~w44307;
assign w44309 = w44281 & ~w44294;
assign w44310 = ~w44281 & w44294;
assign w44311 = ~w44309 & ~w44310;
assign w44312 = w44287 & ~w44311;
assign w44313 = w44281 & ~w44287;
assign w44314 = ~w44287 & w44300;
assign w44315 = ~w44313 & ~w44314;
assign w44316 = ~w44308 & w44315;
assign w44317 = ~w44312 & w44316;
assign w44318 = ~w44287 & w44294;
assign w44319 = w44287 & ~w44294;
assign w44320 = ~w44318 & ~w44319;
assign w44321 = w44281 & w44320;
assign w44322 = ~w44287 & ~w44308;
assign w44323 = ~w44281 & ~w44322;
assign w44324 = ~w44320 & w44323;
assign w44325 = ~w44321 & ~w44324;
assign w44326 = ~w44288 & w44308;
assign w44327 = w44325 & w44326;
assign w44328 = ~pi4969 & pi9040;
assign w44329 = ~pi4669 & ~pi9040;
assign w44330 = ~w44328 & ~w44329;
assign w44331 = pi2295 & ~w44330;
assign w44332 = ~pi2295 & w44330;
assign w44333 = ~w44331 & ~w44332;
assign w44334 = ~w44302 & ~w44333;
assign w44335 = ~w44317 & w44334;
assign w44336 = ~w44327 & w44335;
assign w44337 = ~w44281 & w44287;
assign w44338 = w44294 & w44300;
assign w44339 = w44337 & w44338;
assign w44340 = ~w44300 & ~w44325;
assign w44341 = w44281 & w44300;
assign w44342 = ~w44308 & ~w44341;
assign w44343 = ~w44315 & w44342;
assign w44344 = w44333 & ~w44339;
assign w44345 = ~w44343 & w44344;
assign w44346 = ~w44340 & w44345;
assign w44347 = ~w44336 & ~w44346;
assign w44348 = (w44308 & ~w44311) | (w44308 & w66529) | (~w44311 & w66529);
assign w44349 = w44300 & w44309;
assign w44350 = ~w44308 & ~w44349;
assign w44351 = ~w44348 & ~w44350;
assign w44352 = ~w44347 & ~w44351;
assign w44353 = ~pi2372 & w44352;
assign w44354 = pi2372 & ~w44352;
assign w44355 = ~w44353 & ~w44354;
assign w44356 = ~w44318 & ~w44341;
assign w44357 = w44348 & ~w44356;
assign w44358 = w44319 & w44357;
assign w44359 = w44287 & ~w44300;
assign w44360 = w44315 & ~w44359;
assign w44361 = (~w44281 & ~w44315) | (~w44281 & w64007) | (~w44315 & w64007);
assign w44362 = ~w44281 & ~w44359;
assign w44363 = w44320 & ~w44362;
assign w44364 = ~w44308 & w44363;
assign w44365 = ~w44319 & w44326;
assign w44366 = w44356 & ~w44365;
assign w44367 = ~w44357 & ~w44366;
assign w44368 = (~w44333 & w44364) | (~w44333 & w66530) | (w44364 & w66530);
assign w44369 = ~w44367 & w44368;
assign w44370 = ~w44322 & ~w44333;
assign w44371 = w44338 & ~w44370;
assign w44372 = ~w44363 & w44371;
assign w44373 = ~w44311 & ~w44356;
assign w44374 = w44342 & ~w44373;
assign w44375 = w44308 & ~w44361;
assign w44376 = ~w44308 & w44337;
assign w44377 = ~w44313 & ~w44376;
assign w44378 = (w44301 & w44376) | (w44301 & w66531) | (w44376 & w66531);
assign w44379 = w44375 & ~w44378;
assign w44380 = w44333 & ~w44374;
assign w44381 = ~w44379 & w44380;
assign w44382 = ~w44358 & ~w44372;
assign w44383 = ~w44369 & w44382;
assign w44384 = ~w44381 & w44383;
assign w44385 = ~pi2358 & ~w44384;
assign w44386 = pi2358 & w44384;
assign w44387 = ~w44385 & ~w44386;
assign w44388 = w44317 & w44338;
assign w44389 = ~w44361 & ~w44373;
assign w44390 = (~w44308 & ~w44320) | (~w44308 & w66532) | (~w44320 & w66532);
assign w44391 = ~w44389 & ~w44390;
assign w44392 = w44389 & w44390;
assign w44393 = ~w44391 & ~w44392;
assign w44394 = ~w44333 & ~w44393;
assign w44395 = ~w44300 & w44308;
assign w44396 = w44310 & w44395;
assign w44397 = ~w44378 & ~w44396;
assign w44398 = w44326 & ~w44397;
assign w44399 = ~w44301 & ~w44337;
assign w44400 = ~w44338 & w44399;
assign w44401 = w44375 & ~w44400;
assign w44402 = ~w44308 & ~w44313;
assign w44403 = w44399 & w44402;
assign w44404 = ~w44378 & ~w44403;
assign w44405 = ~w44401 & w44404;
assign w44406 = w44333 & ~w44405;
assign w44407 = ~w44388 & ~w44398;
assign w44408 = ~w44394 & w44407;
assign w44409 = (pi2356 & ~w44408) | (pi2356 & w66533) | (~w44408 & w66533);
assign w44410 = w44408 & w66534;
assign w44411 = ~w44409 & ~w44410;
assign w44412 = w44310 & w44314;
assign w44413 = w44326 & ~w44363;
assign w44414 = (~w44412 & ~w44363) | (~w44412 & w66535) | (~w44363 & w66535);
assign w44415 = ~w44413 & w44414;
assign w44416 = w44333 & ~w44415;
assign w44417 = w44338 & ~w44377;
assign w44418 = ~w44313 & w44400;
assign w44419 = ~w44417 & ~w44418;
assign w44420 = w44397 & w44419;
assign w44421 = ~w44333 & ~w44420;
assign w44422 = ~w44294 & w44308;
assign w44423 = w44360 & w44422;
assign w44424 = ~w44416 & ~w44423;
assign w44425 = ~w44421 & w44424;
assign w44426 = ~pi2369 & w44425;
assign w44427 = pi2369 & ~w44425;
assign w44428 = ~w44426 & ~w44427;
assign w44429 = w44150 & w44165;
assign w44430 = w44161 & w44162;
assign w44431 = ~w44429 & ~w44430;
assign w44432 = (~w44143 & w44174) | (~w44143 & w66536) | (w44174 & w66536);
assign w44433 = w44431 & ~w44432;
assign w44434 = w44135 & ~w44433;
assign w44435 = ~w44128 & w44154;
assign w44436 = ~w44166 & ~w44435;
assign w44437 = ~w44135 & ~w44436;
assign w44438 = w44135 & w44149;
assign w44439 = w44151 & w44438;
assign w44440 = ~w44437 & ~w44439;
assign w44441 = ~w44182 & ~w44440;
assign w44442 = ~w44162 & ~w44189;
assign w44443 = w44122 & ~w44135;
assign w44444 = w44143 & ~w44182;
assign w44445 = ~w44443 & ~w44444;
assign w44446 = ~w44136 & ~w44442;
assign w44447 = ~w44445 & w44446;
assign w44448 = ~w44150 & ~w44158;
assign w44449 = ~w44160 & w66537;
assign w44450 = ~w44128 & w44186;
assign w44451 = ~w44165 & ~w44450;
assign w44452 = w44438 & ~w44451;
assign w44453 = w44431 & ~w44452;
assign w44454 = ~w44449 & w44453;
assign w44455 = w44182 & ~w44454;
assign w44456 = ~w44434 & ~w44447;
assign w44457 = ~w44441 & w44456;
assign w44458 = ~w44455 & w44457;
assign w44459 = pi2342 & w44458;
assign w44460 = ~pi2342 & ~w44458;
assign w44461 = ~w44459 & ~w44460;
assign w44462 = w43613 & ~w44235;
assign w44463 = w43613 & w43691;
assign w44464 = ~w43644 & w44236;
assign w44465 = ~w44243 & ~w44464;
assign w44466 = ~w43672 & ~w44463;
assign w44467 = ~w44465 & w44466;
assign w44468 = w43656 & ~w44467;
assign w44469 = w44232 & ~w44249;
assign w44470 = ~w43675 & w44469;
assign w44471 = ~w44228 & ~w44261;
assign w44472 = w43642 & ~w43656;
assign w44473 = ~w44471 & w44472;
assign w44474 = ~w44470 & ~w44473;
assign w44475 = ~w44462 & w44474;
assign w44476 = ~w44468 & w44475;
assign w44477 = pi2378 & ~w44476;
assign w44478 = ~pi2378 & w44476;
assign w44479 = ~w44477 & ~w44478;
assign w44480 = w44122 & ~w44155;
assign w44481 = (w44128 & w44480) | (w44128 & w63330) | (w44480 & w63330);
assign w44482 = w44135 & ~w44167;
assign w44483 = w44128 & w44154;
assign w44484 = w44129 & ~w44149;
assign w44485 = ~w44135 & ~w44484;
assign w44486 = ~w44149 & w44151;
assign w44487 = ~w44483 & ~w44486;
assign w44488 = ~w44480 & w44487;
assign w44489 = w44485 & w44488;
assign w44490 = (~w44481 & w44489) | (~w44481 & w66538) | (w44489 & w66538);
assign w44491 = w44182 & ~w44490;
assign w44492 = ~w44168 & ~w44182;
assign w44493 = ~w44135 & ~w44481;
assign w44494 = ~w44492 & w44493;
assign w44495 = ~w44481 & w66539;
assign w44496 = w44135 & ~w44166;
assign w44497 = ~w44495 & w44496;
assign w44498 = ~w44494 & ~w44497;
assign w44499 = ~w44491 & ~w44498;
assign w44500 = ~pi2347 & w44499;
assign w44501 = pi2347 & ~w44499;
assign w44502 = ~w44500 & ~w44501;
assign w44503 = ~w44481 & w63428;
assign w44504 = ~w44158 & ~w44435;
assign w44505 = w44135 & ~w44504;
assign w44506 = w44188 & ~w44435;
assign w44507 = ~w44505 & ~w44506;
assign w44508 = ~w44503 & w44507;
assign w44509 = w44483 & w44508;
assign w44510 = ~w44136 & ~w44443;
assign w44511 = w44164 & ~w44510;
assign w44512 = w44135 & ~w44450;
assign w44513 = (~w44512 & w44160) | (~w44512 & w64008) | (w44160 & w64008);
assign w44514 = (w44182 & w44509) | (w44182 & w64009) | (w44509 & w64009);
assign w44515 = w44149 & w44450;
assign w44516 = w44485 & ~w44515;
assign w44517 = w44135 & ~w44429;
assign w44518 = ~w44516 & ~w44517;
assign w44519 = (~w44518 & w44508) | (~w44518 & w66540) | (w44508 & w66540);
assign w44520 = ~w44514 & w66541;
assign w44521 = (pi2354 & w44514) | (pi2354 & w66542) | (w44514 & w66542);
assign w44522 = ~w44520 & ~w44521;
assign w44523 = ~pi4857 & pi9040;
assign w44524 = ~pi4828 & ~pi9040;
assign w44525 = ~w44523 & ~w44524;
assign w44526 = pi2384 & ~w44525;
assign w44527 = ~pi2384 & w44525;
assign w44528 = ~w44526 & ~w44527;
assign w44529 = ~pi5111 & pi9040;
assign w44530 = ~pi4856 & ~pi9040;
assign w44531 = ~w44529 & ~w44530;
assign w44532 = pi2381 & ~w44531;
assign w44533 = ~pi2381 & w44531;
assign w44534 = ~w44532 & ~w44533;
assign w44535 = ~pi4828 & pi9040;
assign w44536 = ~pi4863 & ~pi9040;
assign w44537 = ~w44535 & ~w44536;
assign w44538 = pi2388 & ~w44537;
assign w44539 = ~pi2388 & w44537;
assign w44540 = ~w44538 & ~w44539;
assign w44541 = w44534 & ~w44540;
assign w44542 = ~pi4752 & pi9040;
assign w44543 = ~pi4857 & ~pi9040;
assign w44544 = ~w44542 & ~w44543;
assign w44545 = pi2392 & ~w44544;
assign w44546 = ~pi2392 & w44544;
assign w44547 = ~w44545 & ~w44546;
assign w44548 = w44541 & ~w44547;
assign w44549 = ~pi4800 & pi9040;
assign w44550 = ~pi5087 & ~pi9040;
assign w44551 = ~w44549 & ~w44550;
assign w44552 = pi2390 & ~w44551;
assign w44553 = ~pi2390 & w44551;
assign w44554 = ~w44552 & ~w44553;
assign w44555 = w44540 & ~w44554;
assign w44556 = ~pi4941 & pi9040;
assign w44557 = ~pi4968 & ~pi9040;
assign w44558 = ~w44556 & ~w44557;
assign w44559 = pi2346 & ~w44558;
assign w44560 = ~pi2346 & w44558;
assign w44561 = ~w44559 & ~w44560;
assign w44562 = w44534 & ~w44561;
assign w44563 = w44555 & w44562;
assign w44564 = ~w44534 & ~w44561;
assign w44565 = w44554 & w44564;
assign w44566 = ~w44563 & ~w44565;
assign w44567 = w44547 & ~w44566;
assign w44568 = ~w44534 & w44540;
assign w44569 = ~w44554 & ~w44568;
assign w44570 = w44554 & ~w44561;
assign w44571 = ~w44547 & ~w44570;
assign w44572 = ~w44569 & w44571;
assign w44573 = ~w44540 & ~w44554;
assign w44574 = w44540 & w44554;
assign w44575 = ~w44573 & ~w44574;
assign w44576 = w44534 & w44561;
assign w44577 = ~w44575 & w44576;
assign w44578 = ~w44548 & ~w44572;
assign w44579 = ~w44577 & w44578;
assign w44580 = (~w44528 & ~w44579) | (~w44528 & w66543) | (~w44579 & w66543);
assign w44581 = w44561 & w44568;
assign w44582 = ~w44540 & w44570;
assign w44583 = ~w44581 & ~w44582;
assign w44584 = ~w44534 & ~w44554;
assign w44585 = ~w44541 & ~w44584;
assign w44586 = (~w44585 & ~w44583) | (~w44585 & w66544) | (~w44583 & w66544);
assign w44587 = w44564 & ~w44575;
assign w44588 = ~w44586 & ~w44587;
assign w44589 = w44573 & w44576;
assign w44590 = ~w44547 & ~w44589;
assign w44591 = ~w44588 & ~w44590;
assign w44592 = ~w44541 & ~w44568;
assign w44593 = ~w44561 & w44592;
assign w44594 = w44568 & w66545;
assign w44595 = ~w44593 & ~w44594;
assign w44596 = ~w44593 & w66546;
assign w44597 = ~w44554 & w44561;
assign w44598 = ~w44541 & ~w44597;
assign w44599 = ~w44581 & w44598;
assign w44600 = ~w44589 & ~w44599;
assign w44601 = w44547 & ~w44600;
assign w44602 = w44528 & ~w44596;
assign w44603 = ~w44601 & w44602;
assign w44604 = ~w44580 & ~w44591;
assign w44605 = ~w44603 & w44604;
assign w44606 = pi2408 & ~w44605;
assign w44607 = ~pi2408 & w44605;
assign w44608 = ~w44606 & ~w44607;
assign w44609 = ~pi4856 & pi9040;
assign w44610 = ~pi4800 & ~pi9040;
assign w44611 = ~w44609 & ~w44610;
assign w44612 = pi2366 & ~w44611;
assign w44613 = ~pi2366 & w44611;
assign w44614 = ~w44612 & ~w44613;
assign w44615 = ~pi5210 & pi9040;
assign w44616 = ~pi4819 & ~pi9040;
assign w44617 = ~w44615 & ~w44616;
assign w44618 = pi2383 & ~w44617;
assign w44619 = ~pi2383 & w44617;
assign w44620 = ~w44618 & ~w44619;
assign w44621 = ~w44614 & w44620;
assign w44622 = ~pi4751 & pi9040;
assign w44623 = ~pi5052 & ~pi9040;
assign w44624 = ~w44622 & ~w44623;
assign w44625 = pi2391 & ~w44624;
assign w44626 = ~pi2391 & w44624;
assign w44627 = ~w44625 & ~w44626;
assign w44628 = ~pi5052 & pi9040;
assign w44629 = ~pi4941 & ~pi9040;
assign w44630 = ~w44628 & ~w44629;
assign w44631 = pi2377 & ~w44630;
assign w44632 = ~pi2377 & w44630;
assign w44633 = ~w44631 & ~w44632;
assign w44634 = w44627 & ~w44633;
assign w44635 = ~w44614 & ~w44633;
assign w44636 = ~pi5087 & pi9040;
assign w44637 = ~pi5111 & ~pi9040;
assign w44638 = ~w44636 & ~w44637;
assign w44639 = pi2346 & ~w44638;
assign w44640 = ~pi2346 & w44638;
assign w44641 = ~w44639 & ~w44640;
assign w44642 = ~w44620 & ~w44641;
assign w44643 = w44620 & w44641;
assign w44644 = ~w44642 & ~w44643;
assign w44645 = w44635 & w44644;
assign w44646 = ~w44634 & ~w44645;
assign w44647 = w44621 & ~w44646;
assign w44648 = w44614 & ~w44620;
assign w44649 = ~w44633 & w44648;
assign w44650 = w44620 & w44633;
assign w44651 = ~w44649 & ~w44650;
assign w44652 = ~w44627 & ~w44641;
assign w44653 = (w44652 & w44649) | (w44652 & w66547) | (w44649 & w66547);
assign w44654 = ~w44621 & ~w44648;
assign w44655 = ~w44634 & w44654;
assign w44656 = w44641 & w44655;
assign w44657 = ~pi4759 & pi9040;
assign w44658 = ~pi4826 & ~pi9040;
assign w44659 = ~w44657 & ~w44658;
assign w44660 = pi2381 & ~w44659;
assign w44661 = ~pi2381 & w44659;
assign w44662 = ~w44660 & ~w44661;
assign w44663 = ~w44653 & ~w44662;
assign w44664 = ~w44656 & w44663;
assign w44665 = ~w44647 & w44664;
assign w44666 = w44635 & w44642;
assign w44667 = w44662 & ~w44666;
assign w44668 = w44641 & w44649;
assign w44669 = w44633 & w44642;
assign w44670 = ~w44633 & w44641;
assign w44671 = w44614 & w44620;
assign w44672 = w44670 & w44671;
assign w44673 = ~w44669 & ~w44672;
assign w44674 = ~w44645 & w44673;
assign w44675 = ~w44649 & w64010;
assign w44676 = w44674 & w64011;
assign w44677 = w44633 & ~w44641;
assign w44678 = ~w44670 & ~w44677;
assign w44679 = ~w44627 & w44678;
assign w44680 = ~w44641 & w44671;
assign w44681 = ~w44614 & w44633;
assign w44682 = w44641 & w44681;
assign w44683 = ~w44680 & ~w44682;
assign w44684 = ~w44679 & ~w44683;
assign w44685 = (~w44655 & w44684) | (~w44655 & w66548) | (w44684 & w66548);
assign w44686 = w44667 & ~w44668;
assign w44687 = ~w44676 & w44686;
assign w44688 = ~w44685 & w44687;
assign w44689 = ~w44665 & ~w44688;
assign w44690 = ~w44627 & ~w44654;
assign w44691 = ~w44627 & ~w44633;
assign w44692 = w44627 & ~w44668;
assign w44693 = ~w44643 & ~w44669;
assign w44694 = (~w44614 & w44669) | (~w44614 & w64012) | (w44669 & w64012);
assign w44695 = ~w44641 & w44651;
assign w44696 = ~w44694 & w44695;
assign w44697 = w44692 & ~w44696;
assign w44698 = ~w44690 & ~w44691;
assign w44699 = ~w44697 & w44698;
assign w44700 = ~w44689 & w66549;
assign w44701 = (pi2425 & w44689) | (pi2425 & w66550) | (w44689 & w66550);
assign w44702 = ~w44700 & ~w44701;
assign w44703 = ~w44627 & w44662;
assign w44704 = ~w44650 & w44667;
assign w44705 = ~w44703 & ~w44704;
assign w44706 = w44648 & ~w44678;
assign w44707 = ~w44634 & w44706;
assign w44708 = w44614 & w44633;
assign w44709 = w44644 & w44708;
assign w44710 = (~w44680 & ~w44674) | (~w44680 & w66551) | (~w44674 & w66551);
assign w44711 = ~w44709 & ~w44710;
assign w44712 = ~w44705 & ~w44707;
assign w44713 = ~w44711 & w44712;
assign w44714 = ~w44620 & ~w44691;
assign w44715 = ~w44708 & w44714;
assign w44716 = ~w44678 & ~w44715;
assign w44717 = ~w44654 & ~w44681;
assign w44718 = w44627 & w44678;
assign w44719 = ~w44717 & w44718;
assign w44720 = ~w44716 & ~w44719;
assign w44721 = w44627 & ~w44670;
assign w44722 = w44671 & ~w44721;
assign w44723 = ~w44662 & ~w44722;
assign w44724 = ~w44720 & w44723;
assign w44725 = ~w44713 & ~w44724;
assign w44726 = pi2420 & w44725;
assign w44727 = ~pi2420 & ~w44725;
assign w44728 = ~w44726 & ~w44727;
assign w44729 = w44541 & w44572;
assign w44730 = w44547 & ~w44576;
assign w44731 = w44554 & ~w44592;
assign w44732 = ~w44730 & w44731;
assign w44733 = ~w44554 & w44593;
assign w44734 = ~w44547 & w44561;
assign w44735 = w44584 & w44734;
assign w44736 = w44540 & ~w44561;
assign w44737 = ~w44597 & ~w44736;
assign w44738 = w44534 & w44547;
assign w44739 = ~w44737 & w44738;
assign w44740 = ~w44581 & ~w44735;
assign w44741 = ~w44739 & w44740;
assign w44742 = ~w44732 & w44741;
assign w44743 = (~w44528 & ~w44742) | (~w44528 & w66552) | (~w44742 & w66552);
assign w44744 = ~w44540 & w44564;
assign w44745 = w44547 & w44744;
assign w44746 = ~w44528 & ~w44745;
assign w44747 = w44547 & ~w44573;
assign w44748 = ~w44736 & w44747;
assign w44749 = w44561 & ~w44574;
assign w44750 = ~w44592 & w44749;
assign w44751 = w44748 & ~w44750;
assign w44752 = ~w44571 & w44744;
assign w44753 = ~w44564 & ~w44576;
assign w44754 = w44555 & ~w44753;
assign w44755 = w44534 & ~w44547;
assign w44756 = w44562 & w44574;
assign w44757 = ~w44573 & ~w44756;
assign w44758 = w44755 & ~w44757;
assign w44759 = ~w44752 & ~w44754;
assign w44760 = ~w44751 & w44759;
assign w44761 = ~w44758 & w44760;
assign w44762 = ~w44746 & ~w44761;
assign w44763 = ~w44729 & ~w44743;
assign w44764 = ~w44762 & w44763;
assign w44765 = pi2431 & ~w44764;
assign w44766 = ~pi2431 & w44764;
assign w44767 = ~w44765 & ~w44766;
assign w44768 = ~pi4829 & pi9040;
assign w44769 = ~pi4953 & ~pi9040;
assign w44770 = ~w44768 & ~w44769;
assign w44771 = pi2390 & ~w44770;
assign w44772 = ~pi2390 & w44770;
assign w44773 = ~w44771 & ~w44772;
assign w44774 = ~pi4825 & pi9040;
assign w44775 = ~pi5095 & ~pi9040;
assign w44776 = ~w44774 & ~w44775;
assign w44777 = pi2389 & ~w44776;
assign w44778 = ~pi2389 & w44776;
assign w44779 = ~w44777 & ~w44778;
assign w44780 = ~w44773 & ~w44779;
assign w44781 = ~pi5211 & pi9040;
assign w44782 = ~pi4829 & ~pi9040;
assign w44783 = ~w44781 & ~w44782;
assign w44784 = pi2387 & ~w44783;
assign w44785 = ~pi2387 & w44783;
assign w44786 = ~w44784 & ~w44785;
assign w44787 = ~pi4827 & pi9040;
assign w44788 = ~pi4750 & ~pi9040;
assign w44789 = ~w44787 & ~w44788;
assign w44790 = pi2384 & ~w44789;
assign w44791 = ~pi2384 & w44789;
assign w44792 = ~w44790 & ~w44791;
assign w44793 = w44786 & w44792;
assign w44794 = w44780 & w44793;
assign w44795 = ~pi4758 & pi9040;
assign w44796 = ~pi5295 & ~pi9040;
assign w44797 = ~w44795 & ~w44796;
assign w44798 = pi2364 & ~w44797;
assign w44799 = ~pi2364 & w44797;
assign w44800 = ~w44798 & ~w44799;
assign w44801 = w44792 & w44800;
assign w44802 = ~w44792 & ~w44800;
assign w44803 = ~w44801 & ~w44802;
assign w44804 = ~w44779 & ~w44800;
assign w44805 = w44773 & w44792;
assign w44806 = w44804 & w44805;
assign w44807 = w44803 & ~w44806;
assign w44808 = w44773 & w44786;
assign w44809 = w44807 & w44808;
assign w44810 = w44807 & w66553;
assign w44811 = ~pi4865 & pi9040;
assign w44812 = ~pi4978 & ~pi9040;
assign w44813 = ~w44811 & ~w44812;
assign w44814 = pi2360 & ~w44813;
assign w44815 = ~pi2360 & w44813;
assign w44816 = ~w44814 & ~w44815;
assign w44817 = ~w44779 & w44786;
assign w44818 = ~w44780 & ~w44817;
assign w44819 = w44773 & w44804;
assign w44820 = ~w44792 & w44819;
assign w44821 = (~w44816 & w44818) | (~w44816 & w66554) | (w44818 & w66554);
assign w44822 = ~w44820 & w44821;
assign w44823 = ~w44810 & w44822;
assign w44824 = ~w44773 & ~w44792;
assign w44825 = ~w44773 & ~w44800;
assign w44826 = w44773 & w44800;
assign w44827 = ~w44825 & ~w44826;
assign w44828 = w44786 & ~w44805;
assign w44829 = w44827 & w44828;
assign w44830 = (~w44804 & w44829) | (~w44804 & w64013) | (w44829 & w64013);
assign w44831 = ~w44779 & ~w44786;
assign w44832 = w44824 & w44831;
assign w44833 = ~w44818 & ~w44832;
assign w44834 = w44807 & w44833;
assign w44835 = ~w44830 & ~w44834;
assign w44836 = ~w44786 & w44805;
assign w44837 = w44816 & ~w44836;
assign w44838 = w44835 & w44837;
assign w44839 = w44779 & ~w44792;
assign w44840 = w44786 & w44839;
assign w44841 = w44825 & w44840;
assign w44842 = ~w44779 & ~w44792;
assign w44843 = w44803 & w44827;
assign w44844 = w44779 & w44792;
assign w44845 = w44825 & w44844;
assign w44846 = (~w44845 & w44843) | (~w44845 & w64014) | (w44843 & w64014);
assign w44847 = ~w44773 & ~w44803;
assign w44848 = (w44779 & ~w44803) | (w44779 & w66555) | (~w44803 & w66555);
assign w44849 = ~w44847 & w44848;
assign w44850 = w44800 & w44849;
assign w44851 = (~w44819 & w44846) | (~w44819 & w66556) | (w44846 & w66556);
assign w44852 = ~w44850 & w44851;
assign w44853 = ~w44786 & ~w44852;
assign w44854 = ~w44794 & ~w44841;
assign w44855 = (w44854 & w44838) | (w44854 & w66557) | (w44838 & w66557);
assign w44856 = ~w44853 & w44855;
assign w44857 = pi2402 & ~w44856;
assign w44858 = ~pi2402 & w44856;
assign w44859 = ~w44857 & ~w44858;
assign w44860 = ~pi4951 & pi9040;
assign w44861 = ~pi4862 & ~pi9040;
assign w44862 = ~w44860 & ~w44861;
assign w44863 = pi2386 & ~w44862;
assign w44864 = ~pi2386 & w44862;
assign w44865 = ~w44863 & ~w44864;
assign w44866 = ~pi4866 & pi9040;
assign w44867 = ~pi4977 & ~pi9040;
assign w44868 = ~w44866 & ~w44867;
assign w44869 = pi2367 & ~w44868;
assign w44870 = ~pi2367 & w44868;
assign w44871 = ~w44869 & ~w44870;
assign w44872 = w44865 & ~w44871;
assign w44873 = ~pi5114 & pi9040;
assign w44874 = ~pi4870 & ~pi9040;
assign w44875 = ~w44873 & ~w44874;
assign w44876 = pi2396 & ~w44875;
assign w44877 = ~pi2396 & w44875;
assign w44878 = ~w44876 & ~w44877;
assign w44879 = ~pi4869 & pi9040;
assign w44880 = ~pi5114 & ~pi9040;
assign w44881 = ~w44879 & ~w44880;
assign w44882 = pi2379 & ~w44881;
assign w44883 = ~pi2379 & w44881;
assign w44884 = ~w44882 & ~w44883;
assign w44885 = w44871 & w44884;
assign w44886 = w44865 & ~w44885;
assign w44887 = ~w44871 & ~w44884;
assign w44888 = ~w44886 & ~w44887;
assign w44889 = ~pi4750 & pi9040;
assign w44890 = ~pi5277 & ~pi9040;
assign w44891 = ~w44889 & ~w44890;
assign w44892 = pi2398 & ~w44891;
assign w44893 = ~pi2398 & w44891;
assign w44894 = ~w44892 & ~w44893;
assign w44895 = ~w44878 & w44894;
assign w44896 = ~w44888 & w44895;
assign w44897 = ~w44872 & w44896;
assign w44898 = ~pi4870 & pi9040;
assign w44899 = ~pi4848 & ~pi9040;
assign w44900 = ~w44898 & ~w44899;
assign w44901 = pi2395 & ~w44900;
assign w44902 = ~pi2395 & w44900;
assign w44903 = ~w44901 & ~w44902;
assign w44904 = ~w44865 & ~w44894;
assign w44905 = w44865 & w44878;
assign w44906 = ~w44904 & ~w44905;
assign w44907 = w44885 & w44906;
assign w44908 = ~w44884 & w44894;
assign w44909 = w44884 & ~w44894;
assign w44910 = ~w44904 & ~w44909;
assign w44911 = w44878 & ~w44910;
assign w44912 = (~w44908 & w44910) | (~w44908 & w66558) | (w44910 & w66558);
assign w44913 = ~w44865 & ~w44871;
assign w44914 = ~w44912 & w44913;
assign w44915 = w44865 & ~w44894;
assign w44916 = (~w44878 & ~w44915) | (~w44878 & w64015) | (~w44915 & w64015);
assign w44917 = ~w44910 & w44916;
assign w44918 = w44878 & ~w44887;
assign w44919 = ~w44887 & w66559;
assign w44920 = ~w44886 & w44919;
assign w44921 = w44871 & ~w44884;
assign w44922 = ~w44894 & w44921;
assign w44923 = w44865 & w44894;
assign w44924 = w44887 & w44923;
assign w44925 = ~w44922 & ~w44924;
assign w44926 = ~w44917 & w44925;
assign w44927 = ~w44920 & w44926;
assign w44928 = w44887 & ~w44906;
assign w44929 = w44872 & ~w44928;
assign w44930 = w44927 & w44929;
assign w44931 = ~w44907 & ~w44914;
assign w44932 = (w44903 & w44930) | (w44903 & w66560) | (w44930 & w66560);
assign w44933 = ~w44903 & ~w44927;
assign w44934 = w44887 & w44894;
assign w44935 = ~w44922 & ~w44934;
assign w44936 = ~w44905 & ~w44917;
assign w44937 = ~w44935 & ~w44936;
assign w44938 = ~w44897 & ~w44937;
assign w44939 = ~w44933 & w44938;
assign w44940 = ~w44932 & w44939;
assign w44941 = pi2401 & w44940;
assign w44942 = ~pi2401 & ~w44940;
assign w44943 = ~w44941 & ~w44942;
assign w44944 = ~w44564 & w44574;
assign w44945 = ~w44755 & w44944;
assign w44946 = (~w44574 & ~w44583) | (~w44574 & w64016) | (~w44583 & w64016);
assign w44947 = w44561 & w44573;
assign w44948 = ~w44945 & ~w44947;
assign w44949 = ~w44946 & w44948;
assign w44950 = ~w44576 & ~w44947;
assign w44951 = ~w44565 & w44950;
assign w44952 = (w44547 & ~w44950) | (w44547 & w64017) | (~w44950 & w64017);
assign w44953 = (w44950 & w66561) | (w44950 & w66562) | (w66561 & w66562);
assign w44954 = ~w44750 & ~w44756;
assign w44955 = (w44954 & ~w44949) | (w44954 & w66563) | (~w44949 & w66563);
assign w44956 = w44528 & ~w44955;
assign w44957 = ~w44595 & w44748;
assign w44958 = w44562 & ~w44747;
assign w44959 = ~w44952 & ~w44958;
assign w44960 = ~w44528 & ~w44959;
assign w44961 = ~w44547 & w44592;
assign w44962 = ~w44735 & ~w44961;
assign w44963 = w44951 & ~w44962;
assign w44964 = ~w44957 & ~w44963;
assign w44965 = ~w44960 & w44964;
assign w44966 = ~w44956 & w44965;
assign w44967 = pi2460 & ~w44966;
assign w44968 = ~pi2460 & w44966;
assign w44969 = ~w44967 & ~w44968;
assign w44970 = ~pi4942 & pi9040;
assign w44971 = ~pi4827 & ~pi9040;
assign w44972 = ~w44970 & ~w44971;
assign w44973 = pi2370 & ~w44972;
assign w44974 = ~pi2370 & w44972;
assign w44975 = ~w44973 & ~w44974;
assign w44976 = ~pi4953 & pi9040;
assign w44977 = ~pi4938 & ~pi9040;
assign w44978 = ~w44976 & ~w44977;
assign w44979 = pi2393 & ~w44978;
assign w44980 = ~pi2393 & w44978;
assign w44981 = ~w44979 & ~w44980;
assign w44982 = ~pi4938 & pi9040;
assign w44983 = ~pi5211 & ~pi9040;
assign w44984 = ~w44982 & ~w44983;
assign w44985 = pi2360 & ~w44984;
assign w44986 = ~pi2360 & w44984;
assign w44987 = ~w44985 & ~w44986;
assign w44988 = w44981 & ~w44987;
assign w44989 = ~pi4956 & pi9040;
assign w44990 = ~pi5092 & ~pi9040;
assign w44991 = ~w44989 & ~w44990;
assign w44992 = pi2394 & ~w44991;
assign w44993 = ~pi2394 & w44991;
assign w44994 = ~w44992 & ~w44993;
assign w44995 = ~pi5277 & pi9040;
assign w44996 = ~pi4942 & ~pi9040;
assign w44997 = ~w44995 & ~w44996;
assign w44998 = pi2364 & ~w44997;
assign w44999 = ~pi2364 & w44997;
assign w45000 = ~w44998 & ~w44999;
assign w45001 = w44994 & ~w45000;
assign w45002 = w44988 & w45001;
assign w45003 = ~w44981 & ~w44987;
assign w45004 = ~w44994 & w45003;
assign w45005 = w44988 & w45000;
assign w45006 = ~w45004 & ~w45005;
assign w45007 = ~pi4848 & pi9040;
assign w45008 = ~pi4869 & ~pi9040;
assign w45009 = ~w45007 & ~w45008;
assign w45010 = pi2371 & ~w45009;
assign w45011 = ~pi2371 & w45009;
assign w45012 = ~w45010 & ~w45011;
assign w45013 = w45006 & ~w45012;
assign w45014 = w44987 & w45000;
assign w45015 = ~w44994 & w45000;
assign w45016 = ~w45014 & ~w45015;
assign w45017 = ~w44987 & ~w45000;
assign w45018 = ~w44981 & ~w45017;
assign w45019 = w45016 & w45018;
assign w45020 = w45012 & ~w45019;
assign w45021 = ~w45013 & ~w45020;
assign w45022 = w44981 & w44987;
assign w45023 = w45000 & w45012;
assign w45024 = w45022 & w45023;
assign w45025 = w44987 & ~w44994;
assign w45026 = ~w44981 & w44994;
assign w45027 = ~w45022 & ~w45026;
assign w45028 = ~w45014 & ~w45027;
assign w45029 = ~w44981 & ~w45000;
assign w45030 = w44981 & ~w44994;
assign w45031 = ~w45029 & ~w45030;
assign w45032 = w44987 & ~w45031;
assign w45033 = ~w45028 & w45032;
assign w45034 = w44987 & ~w45026;
assign w45035 = ~w45029 & ~w45034;
assign w45036 = ~w45033 & ~w45035;
assign w45037 = (~w45012 & w45033) | (~w45012 & w64018) | (w45033 & w64018);
assign w45038 = ~w45012 & w45027;
assign w45039 = w45025 & ~w45038;
assign w45040 = ~w45037 & w45039;
assign w45041 = w44975 & ~w45002;
assign w45042 = ~w45024 & w45041;
assign w45043 = ~w45021 & w45042;
assign w45044 = ~w45040 & w45043;
assign w45045 = w45014 & w45026;
assign w45046 = w45001 & w45022;
assign w45047 = ~w45045 & ~w45046;
assign w45048 = w45001 & w45003;
assign w45049 = ~w45006 & w45012;
assign w45050 = ~w44975 & ~w45048;
assign w45051 = w45047 & w45050;
assign w45052 = ~w45049 & w45051;
assign w45053 = ~w45044 & ~w45052;
assign w45054 = ~w44975 & w45006;
assign w45055 = ~w45028 & w45054;
assign w45056 = ~w44987 & w45001;
assign w45057 = ~w45045 & ~w45056;
assign w45058 = ~w45055 & w45057;
assign w45059 = ~w45012 & ~w45058;
assign w45060 = ~w45053 & w66564;
assign w45061 = (pi2407 & w45053) | (pi2407 & w66565) | (w45053 & w66565);
assign w45062 = ~w45060 & ~w45061;
assign w45063 = ~w44735 & ~w44949;
assign w45064 = ~w44528 & ~w45063;
assign w45065 = w44583 & ~w44589;
assign w45066 = w44596 & ~w45065;
assign w45067 = w44547 & ~w44561;
assign w45068 = w44555 & w45067;
assign w45069 = ~w44534 & w44737;
assign w45070 = w44534 & w44597;
assign w45071 = (~w44547 & w45069) | (~w44547 & w66566) | (w45069 & w66566);
assign w45072 = w44547 & ~w45070;
assign w45073 = ~w44950 & w45072;
assign w45074 = ~w44563 & ~w44582;
assign w45075 = ~w44594 & w45074;
assign w45076 = ~w45073 & w45075;
assign w45077 = (w44528 & ~w45076) | (w44528 & w66567) | (~w45076 & w66567);
assign w45078 = ~w45066 & ~w45068;
assign w45079 = ~w45077 & w45078;
assign w45080 = ~w45064 & w45079;
assign w45081 = pi2451 & ~w45080;
assign w45082 = ~pi2451 & w45080;
assign w45083 = ~w45081 & ~w45082;
assign w45084 = ~w44672 & ~w44709;
assign w45085 = ~w44614 & ~w44644;
assign w45086 = (w44627 & ~w45084) | (w44627 & w66568) | (~w45084 & w66568);
assign w45087 = (~w44662 & w44694) | (~w44662 & w66569) | (w44694 & w66569);
assign w45088 = w45084 & ~w45087;
assign w45089 = ~w45086 & ~w45088;
assign w45090 = w44627 & ~w44694;
assign w45091 = w44693 & ~w44717;
assign w45092 = ~w44620 & w44708;
assign w45093 = ~w44627 & ~w45092;
assign w45094 = ~w45091 & w45093;
assign w45095 = (w45084 & w45094) | (w45084 & w66570) | (w45094 & w66570);
assign w45096 = w44662 & ~w45095;
assign w45097 = ~w44641 & ~w44703;
assign w45098 = w44649 & w45097;
assign w45099 = ~w45089 & ~w45098;
assign w45100 = ~w45096 & w45099;
assign w45101 = pi2436 & ~w45100;
assign w45102 = ~pi2436 & w45100;
assign w45103 = ~w45101 & ~w45102;
assign w45104 = ~w44896 & ~w44911;
assign w45105 = w44885 & w44923;
assign w45106 = ~w44865 & w44871;
assign w45107 = ~w44872 & ~w45106;
assign w45108 = w44908 & ~w45107;
assign w45109 = w44885 & ~w44894;
assign w45110 = w44918 & ~w45109;
assign w45111 = ~w44884 & w45106;
assign w45112 = w44916 & ~w45111;
assign w45113 = ~w44905 & ~w45110;
assign w45114 = ~w45112 & w45113;
assign w45115 = ~w45105 & ~w45108;
assign w45116 = ~w45114 & w45115;
assign w45117 = ~w45104 & ~w45116;
assign w45118 = ~w44865 & w44885;
assign w45119 = (~w44878 & w45118) | (~w44878 & w66571) | (w45118 & w66571);
assign w45120 = ~w44878 & w44909;
assign w45121 = ~w44904 & ~w44922;
assign w45122 = (~w44919 & w45121) | (~w44919 & w66572) | (w45121 & w66572);
assign w45123 = ~w45106 & ~w45122;
assign w45124 = w44878 & ~w44904;
assign w45125 = ~w44923 & w45124;
assign w45126 = ~w45107 & w45125;
assign w45127 = w45125 & w45108;
assign w45128 = w44894 & w44913;
assign w45129 = w44913 & w66573;
assign w45130 = ~w44903 & ~w45129;
assign w45131 = ~w45119 & w45130;
assign w45132 = ~w45127 & w45131;
assign w45133 = ~w45123 & w45132;
assign w45134 = w44903 & ~w45105;
assign w45135 = w44913 & w45120;
assign w45136 = ~w44878 & ~w44935;
assign w45137 = ~w44924 & w45134;
assign w45138 = ~w45135 & w45137;
assign w45139 = ~w45126 & ~w45136;
assign w45140 = w45138 & w45139;
assign w45141 = ~w45133 & ~w45140;
assign w45142 = ~w45117 & ~w45141;
assign w45143 = ~pi2400 & w45142;
assign w45144 = pi2400 & ~w45142;
assign w45145 = ~w45143 & ~w45144;
assign w45146 = ~w44674 & w44703;
assign w45147 = ~w44645 & w44679;
assign w45148 = w44620 & ~w44691;
assign w45149 = w44683 & w45148;
assign w45150 = ~w44706 & ~w45147;
assign w45151 = ~w45149 & w45150;
assign w45152 = ~w44662 & ~w45151;
assign w45153 = w44634 & w44642;
assign w45154 = ~w44684 & ~w45153;
assign w45155 = w44662 & ~w45154;
assign w45156 = w44643 & w44681;
assign w45157 = w45093 & ~w45156;
assign w45158 = ~w44692 & ~w45157;
assign w45159 = ~w45146 & ~w45158;
assign w45160 = ~w45155 & w45159;
assign w45161 = ~w45152 & w45160;
assign w45162 = ~pi2443 & ~w45161;
assign w45163 = pi2443 & w45161;
assign w45164 = ~w45162 & ~w45163;
assign w45165 = ~pi4862 & pi9040;
assign w45166 = ~pi4866 & ~pi9040;
assign w45167 = ~w45165 & ~w45166;
assign w45168 = pi2370 & ~w45167;
assign w45169 = ~pi2370 & w45167;
assign w45170 = ~w45168 & ~w45169;
assign w45171 = ~pi4948 & pi9040;
assign w45172 = ~pi4758 & ~pi9040;
assign w45173 = ~w45171 & ~w45172;
assign w45174 = pi2385 & ~w45173;
assign w45175 = ~pi2385 & w45173;
assign w45176 = ~w45174 & ~w45175;
assign w45177 = w45170 & w45176;
assign w45178 = ~pi4954 & pi9040;
assign w45179 = ~pi4948 & ~pi9040;
assign w45180 = ~w45178 & ~w45179;
assign w45181 = pi2393 & ~w45180;
assign w45182 = ~pi2393 & w45180;
assign w45183 = ~w45181 & ~w45182;
assign w45184 = w45177 & ~w45183;
assign w45185 = ~pi5095 & pi9040;
assign w45186 = ~pi4761 & ~pi9040;
assign w45187 = ~w45185 & ~w45186;
assign w45188 = pi2352 & ~w45187;
assign w45189 = ~pi2352 & w45187;
assign w45190 = ~w45188 & ~w45189;
assign w45191 = ~w45184 & ~w45190;
assign w45192 = ~w45170 & ~w45183;
assign w45193 = w45170 & w45183;
assign w45194 = ~w45192 & ~w45193;
assign w45195 = ~pi5092 & pi9040;
assign w45196 = ~pi4865 & ~pi9040;
assign w45197 = ~w45195 & ~w45196;
assign w45198 = pi2398 & ~w45197;
assign w45199 = ~pi2398 & w45197;
assign w45200 = ~w45198 & ~w45199;
assign w45201 = w45176 & ~w45200;
assign w45202 = ~w45194 & w45201;
assign w45203 = w45190 & ~w45202;
assign w45204 = ~w45191 & ~w45203;
assign w45205 = ~w45194 & w45200;
assign w45206 = ~w45170 & ~w45200;
assign w45207 = ~w45176 & w45206;
assign w45208 = (~w45190 & w45205) | (~w45190 & w66574) | (w45205 & w66574);
assign w45209 = ~pi5295 & pi9040;
assign w45210 = ~pi4954 & ~pi9040;
assign w45211 = ~w45209 & ~w45210;
assign w45212 = pi2367 & ~w45211;
assign w45213 = ~pi2367 & w45211;
assign w45214 = ~w45212 & ~w45213;
assign w45215 = ~w45176 & ~w45183;
assign w45216 = w45206 & w45215;
assign w45217 = w45170 & w45200;
assign w45218 = ~w45206 & ~w45217;
assign w45219 = ~w45190 & ~w45200;
assign w45220 = w45183 & ~w45219;
assign w45221 = ~w45218 & ~w45220;
assign w45222 = w45183 & w45218;
assign w45223 = ~w45221 & ~w45222;
assign w45224 = w45190 & ~w45192;
assign w45225 = ~w45223 & w45224;
assign w45226 = ~w45214 & ~w45216;
assign w45227 = ~w45208 & w45226;
assign w45228 = ~w45225 & w45227;
assign w45229 = ~w45170 & ~w45176;
assign w45230 = ~w45177 & w45219;
assign w45231 = ~w45229 & w45230;
assign w45232 = ~w45176 & w45223;
assign w45233 = ~w45170 & w45200;
assign w45234 = w45176 & w45183;
assign w45235 = w45233 & w45234;
assign w45236 = w45214 & ~w45235;
assign w45237 = ~w45231 & w45236;
assign w45238 = ~w45232 & w45237;
assign w45239 = ~w45228 & ~w45238;
assign w45240 = ~w45204 & ~w45239;
assign w45241 = ~pi2449 & w45240;
assign w45242 = pi2449 & ~w45240;
assign w45243 = ~w45241 & ~w45242;
assign w45244 = ~w45190 & w45214;
assign w45245 = w45218 & w64019;
assign w45246 = ~w45183 & w45200;
assign w45247 = ~w45206 & ~w45246;
assign w45248 = ~w45245 & w45247;
assign w45249 = w45244 & w45248;
assign w45250 = w45214 & w45245;
assign w45251 = ~w45176 & ~w45214;
assign w45252 = w45246 & ~w45251;
assign w45253 = ~w45216 & ~w45252;
assign w45254 = ~w45250 & w45253;
assign w45255 = w45190 & ~w45254;
assign w45256 = w45206 & w45214;
assign w45257 = w45234 & w45256;
assign w45258 = ~w45215 & ~w45234;
assign w45259 = w45190 & w45200;
assign w45260 = w45218 & ~w45259;
assign w45261 = ~w45258 & ~w45260;
assign w45262 = ~w45206 & ~w45229;
assign w45263 = ~w45207 & ~w45262;
assign w45264 = (w45190 & ~w45258) | (w45190 & w64020) | (~w45258 & w64020);
assign w45265 = ~w45263 & w45264;
assign w45266 = ~w45260 & ~w45265;
assign w45267 = w45258 & ~w45266;
assign w45268 = ~w45214 & ~w45261;
assign w45269 = ~w45267 & w45268;
assign w45270 = ~w45249 & ~w45257;
assign w45271 = ~w45255 & w45270;
assign w45272 = ~w45269 & w45271;
assign w45273 = pi2441 & w45272;
assign w45274 = ~pi2441 & ~w45272;
assign w45275 = ~w45273 & ~w45274;
assign w45276 = w45183 & ~w45200;
assign w45277 = ~w45177 & ~w45276;
assign w45278 = ~w45190 & ~w45277;
assign w45279 = w45205 & w45278;
assign w45280 = (~w45190 & w45245) | (~w45190 & w66575) | (w45245 & w66575);
assign w45281 = ~w45193 & ~w45277;
assign w45282 = ~w45263 & ~w45281;
assign w45283 = ~w45191 & ~w45282;
assign w45284 = w45280 & ~w45282;
assign w45285 = (~w45214 & w45283) | (~w45214 & w66576) | (w45283 & w66576);
assign w45286 = ~w45284 & w45285;
assign w45287 = w45218 & w66577;
assign w45288 = (w45214 & w45265) | (w45214 & w66578) | (w45265 & w66578);
assign w45289 = ~w45263 & ~w45287;
assign w45290 = w45190 & ~w45289;
assign w45291 = w45247 & w45290;
assign w45292 = ~w45215 & w45244;
assign w45293 = ~w45218 & w45292;
assign w45294 = ~w45279 & ~w45293;
assign w45295 = ~w45288 & w45294;
assign w45296 = ~w45291 & w45295;
assign w45297 = ~w45286 & w45296;
assign w45298 = ~pi2445 & w45297;
assign w45299 = pi2445 & ~w45297;
assign w45300 = ~w45298 & ~w45299;
assign w45301 = ~pi4952 & pi9040;
assign w45302 = ~pi5090 & ~pi9040;
assign w45303 = ~w45301 & ~w45302;
assign w45304 = pi2376 & ~w45303;
assign w45305 = ~pi2376 & w45303;
assign w45306 = ~w45304 & ~w45305;
assign w45307 = ~pi5090 & pi9040;
assign w45308 = ~pi5210 & ~pi9040;
assign w45309 = ~w45307 & ~w45308;
assign w45310 = pi2365 & ~w45309;
assign w45311 = ~pi2365 & w45309;
assign w45312 = ~w45310 & ~w45311;
assign w45313 = w45306 & ~w45312;
assign w45314 = ~pi4824 & pi9040;
assign w45315 = ~pi4859 & ~pi9040;
assign w45316 = ~w45314 & ~w45315;
assign w45317 = pi2380 & ~w45316;
assign w45318 = ~pi2380 & w45316;
assign w45319 = ~w45317 & ~w45318;
assign w45320 = ~pi4939 & pi9040;
assign w45321 = ~pi5081 & ~pi9040;
assign w45322 = ~w45320 & ~w45321;
assign w45323 = pi2377 & ~w45322;
assign w45324 = ~pi2377 & w45322;
assign w45325 = ~w45323 & ~w45324;
assign w45326 = ~w45319 & ~w45325;
assign w45327 = w45313 & w45326;
assign w45328 = ~pi4859 & pi9040;
assign w45329 = ~pi4970 & ~pi9040;
assign w45330 = ~w45328 & ~w45329;
assign w45331 = pi2383 & ~w45330;
assign w45332 = ~pi2383 & w45330;
assign w45333 = ~w45331 & ~w45332;
assign w45334 = ~w45306 & ~w45319;
assign w45335 = ~w45312 & w45325;
assign w45336 = w45334 & w45335;
assign w45337 = ~pi5186 & pi9040;
assign w45338 = ~pi4820 & ~pi9040;
assign w45339 = ~w45337 & ~w45338;
assign w45340 = pi2397 & ~w45339;
assign w45341 = ~pi2397 & w45339;
assign w45342 = ~w45340 & ~w45341;
assign w45343 = ~w45325 & ~w45342;
assign w45344 = w45313 & w45343;
assign w45345 = w45312 & w45325;
assign w45346 = w45306 & w45345;
assign w45347 = w45345 & w45747;
assign w45348 = ~w45344 & ~w45347;
assign w45349 = ~w45336 & w45348;
assign w45350 = ~w45306 & w45312;
assign w45351 = w45326 & w45350;
assign w45352 = w45342 & ~w45351;
assign w45353 = ~w45312 & w45319;
assign w45354 = ~w45325 & ~w45353;
assign w45355 = ~w45353 & w64021;
assign w45356 = ~w45346 & ~w45355;
assign w45357 = ~w45352 & ~w45356;
assign w45358 = ~w45313 & w45342;
assign w45359 = w45306 & w45319;
assign w45360 = ~w45354 & ~w45359;
assign w45361 = w45306 & ~w45325;
assign w45362 = w45319 & w45361;
assign w45363 = ~w45360 & ~w45362;
assign w45364 = w45319 & w45358;
assign w45365 = ~w45363 & w45364;
assign w45366 = w45349 & ~w45357;
assign w45367 = ~w45365 & w45366;
assign w45368 = w45325 & w45342;
assign w45369 = w45353 & w45368;
assign w45370 = w45334 & w45345;
assign w45371 = w45312 & ~w45362;
assign w45372 = ~w45334 & ~w45361;
assign w45373 = ~w45312 & ~w45372;
assign w45374 = ~w45342 & ~w45373;
assign w45375 = ~w45371 & w45374;
assign w45376 = (~w45370 & ~w45363) | (~w45370 & w66579) | (~w45363 & w66579);
assign w45377 = ~w45375 & w45376;
assign w45378 = ~w45333 & ~w45377;
assign w45379 = ~w45327 & ~w45369;
assign w45380 = (w45379 & w45367) | (w45379 & w66580) | (w45367 & w66580);
assign w45381 = ~w45378 & w45380;
assign w45382 = pi2414 & ~w45381;
assign w45383 = ~pi2414 & w45381;
assign w45384 = ~w45382 & ~w45383;
assign w45385 = ~w45306 & ~w45312;
assign w45386 = w45342 & ~w45385;
assign w45387 = (w45325 & w45385) | (w45325 & w63429) | (w45385 & w63429);
assign w45388 = w45353 & ~w45387;
assign w45389 = (w45358 & w45388) | (w45358 & w66581) | (w45388 & w66581);
assign w45390 = w45319 & w45325;
assign w45391 = ~w45326 & ~w45390;
assign w45392 = ~w45306 & ~w45342;
assign w45393 = ~w45346 & ~w45392;
assign w45394 = ~w45391 & ~w45393;
assign w45395 = ~w45389 & ~w45394;
assign w45396 = ~w45374 & ~w45395;
assign w45397 = w45334 & w45368;
assign w45398 = ~w45388 & ~w45397;
assign w45399 = (~w45372 & w45388) | (~w45372 & w64022) | (w45388 & w64022);
assign w45400 = ~w45350 & ~w45359;
assign w45401 = w45358 & w45400;
assign w45402 = ~w45399 & ~w45401;
assign w45403 = w45312 & ~w45372;
assign w45404 = ~w45334 & w45335;
assign w45405 = ~w45359 & w45404;
assign w45406 = ~w45403 & ~w45405;
assign w45407 = w45342 & w45406;
assign w45408 = w45402 & w45407;
assign w45409 = ~w45349 & w45399;
assign w45410 = (w45333 & w45406) | (w45333 & w64023) | (w45406 & w64023);
assign w45411 = ~w45409 & w45410;
assign w45412 = ~w45408 & w45411;
assign w45413 = ~w45313 & ~w45350;
assign w45414 = w45319 & ~w45342;
assign w45415 = ~w45413 & w45414;
assign w45416 = ~w45333 & ~w45415;
assign w45417 = w45348 & w45416;
assign w45418 = w45402 & w45417;
assign w45419 = (~w45396 & w45412) | (~w45396 & w66582) | (w45412 & w66582);
assign w45420 = ~pi2419 & w45419;
assign w45421 = pi2419 & ~w45419;
assign w45422 = ~w45420 & ~w45421;
assign w45423 = ~w45000 & ~w45012;
assign w45424 = w45030 & ~w45423;
assign w45425 = ~w45005 & ~w45030;
assign w45426 = ~w45424 & ~w45425;
assign w45427 = w45038 & w45426;
assign w45428 = ~w44988 & w45016;
assign w45429 = ~w45032 & w45428;
assign w45430 = w45006 & w66583;
assign w45431 = ~w45429 & w45430;
assign w45432 = w44981 & ~w45017;
assign w45433 = ~w45029 & ~w45432;
assign w45434 = ~w44994 & w45433;
assign w45435 = ~w45426 & ~w45434;
assign w45436 = ~w45431 & w45435;
assign w45437 = ~w44975 & ~w45436;
assign w45438 = ~w45012 & w45429;
assign w45439 = (w44975 & w45438) | (w44975 & w66584) | (w45438 & w66584);
assign w45440 = ~w44975 & ~w45025;
assign w45441 = ~w45016 & ~w45440;
assign w45442 = ~w44975 & w45046;
assign w45443 = ~w45048 & ~w45441;
assign w45444 = (w45012 & ~w45443) | (w45012 & w66585) | (~w45443 & w66585);
assign w45445 = ~w45427 & ~w45444;
assign w45446 = ~w45439 & w45445;
assign w45447 = ~w45437 & w45446;
assign w45448 = pi2406 & ~w45447;
assign w45449 = ~pi2406 & w45447;
assign w45450 = ~w45448 & ~w45449;
assign w45451 = ~w44975 & w45012;
assign w45452 = ~w45033 & w66586;
assign w45453 = w45424 & w45440;
assign w45454 = w45014 & ~w45451;
assign w45455 = ~w45036 & w45454;
assign w45456 = ~w44994 & ~w45029;
assign w45457 = w45027 & ~w45456;
assign w45458 = ~w45423 & ~w45457;
assign w45459 = ~w45038 & ~w45458;
assign w45460 = w45000 & w45004;
assign w45461 = ~w45426 & ~w45460;
assign w45462 = ~w45459 & w45461;
assign w45463 = w44975 & ~w45462;
assign w45464 = ~w44975 & w45425;
assign w45465 = w45037 & w45464;
assign w45466 = ~w45452 & ~w45453;
assign w45467 = ~w45455 & w45466;
assign w45468 = ~w45463 & ~w45465;
assign w45469 = w45468 & w66587;
assign w45470 = (~pi2416 & ~w45468) | (~pi2416 & w66588) | (~w45468 & w66588);
assign w45471 = ~w45469 & ~w45470;
assign w45472 = w45184 & w45259;
assign w45473 = ~w45217 & w45234;
assign w45474 = ~w45290 & ~w45473;
assign w45475 = w45214 & ~w45474;
assign w45476 = w45219 & w45234;
assign w45477 = ~w45247 & w45282;
assign w45478 = ~w45190 & ~w45192;
assign w45479 = w45277 & ~w45478;
assign w45480 = w45176 & w45276;
assign w45481 = ~w45278 & ~w45480;
assign w45482 = ~w45479 & w45481;
assign w45483 = ~w45477 & ~w45482;
assign w45484 = ~w45214 & ~w45483;
assign w45485 = ~w45177 & ~w45281;
assign w45486 = w45244 & ~w45485;
assign w45487 = ~w45472 & ~w45476;
assign w45488 = ~w45486 & w45487;
assign w45489 = ~w45484 & w45488;
assign w45490 = (pi2446 & ~w45489) | (pi2446 & w66589) | (~w45489 & w66589);
assign w45491 = w45489 & w66590;
assign w45492 = ~w45490 & ~w45491;
assign w45493 = w44831 & w44843;
assign w45494 = w44779 & w44826;
assign w45495 = w44802 & w44808;
assign w45496 = ~w45494 & ~w45495;
assign w45497 = ~w44793 & ~w44839;
assign w45498 = w44816 & ~w45497;
assign w45499 = ~w45496 & ~w45498;
assign w45500 = w44780 & ~w44800;
assign w45501 = ~w44786 & w44844;
assign w45502 = ~w44840 & ~w45501;
assign w45503 = w44800 & ~w45502;
assign w45504 = ~w44816 & ~w44836;
assign w45505 = ~w45500 & w45504;
assign w45506 = ~w45503 & w45505;
assign w45507 = ~w44792 & w44827;
assign w45508 = ~w44845 & ~w45507;
assign w45509 = ~w44786 & ~w45508;
assign w45510 = w44780 & w44801;
assign w45511 = w44816 & ~w45510;
assign w45512 = ~w44841 & w45511;
assign w45513 = ~w44809 & w45512;
assign w45514 = ~w45509 & w45513;
assign w45515 = ~w45506 & ~w45514;
assign w45516 = ~w44794 & ~w45493;
assign w45517 = ~w45499 & w45516;
assign w45518 = ~w45515 & w45517;
assign w45519 = pi2412 & ~w45518;
assign w45520 = ~pi2412 & w45518;
assign w45521 = ~w45519 & ~w45520;
assign w45522 = w45343 & w45385;
assign w45523 = w45342 & w45362;
assign w45524 = w45306 & w45342;
assign w45525 = ~w45392 & ~w45524;
assign w45526 = ~w45391 & w45525;
assign w45527 = ~w45523 & ~w45526;
assign w45528 = w45335 & w45525;
assign w45529 = ~w45327 & ~w45528;
assign w45530 = ~w45312 & w45333;
assign w45531 = w45527 & w45530;
assign w45532 = w45529 & w45531;
assign w45533 = w45333 & w45390;
assign w45534 = w45527 & ~w45533;
assign w45535 = w45312 & ~w45534;
assign w45536 = ~w45333 & ~w45529;
assign w45537 = ~w45333 & ~w45335;
assign w45538 = w45391 & ~w45525;
assign w45539 = w45537 & w45538;
assign w45540 = ~w45522 & ~w45539;
assign w45541 = ~w45536 & w45540;
assign w45542 = ~w45532 & w45541;
assign w45543 = ~w45535 & w45542;
assign w45544 = pi2415 & ~w45543;
assign w45545 = ~pi2415 & w45543;
assign w45546 = ~w45544 & ~w45545;
assign w45547 = ~w44871 & w44919;
assign w45548 = ~w44888 & ~w44910;
assign w45549 = ~w45105 & ~w45548;
assign w45550 = ~w44878 & ~w45549;
assign w45551 = w44905 & w44922;
assign w45552 = w44925 & ~w45118;
assign w45553 = w44916 & ~w45552;
assign w45554 = w44878 & w45128;
assign w45555 = ~w44871 & w44909;
assign w45556 = w44865 & w45555;
assign w45557 = ~w45554 & ~w45556;
assign w45558 = w45134 & ~w45551;
assign w45559 = w45557 & w45558;
assign w45560 = ~w45553 & w45559;
assign w45561 = w44871 & ~w44912;
assign w45562 = w44906 & w44921;
assign w45563 = ~w44928 & ~w45135;
assign w45564 = w45563 & w66591;
assign w45565 = ~w45561 & w45564;
assign w45566 = ~w45560 & ~w45565;
assign w45567 = ~w45127 & ~w45547;
assign w45568 = ~w45550 & w45567;
assign w45569 = ~w45566 & w45568;
assign w45570 = pi2403 & ~w45569;
assign w45571 = ~pi2403 & w45569;
assign w45572 = ~w45570 & ~w45571;
assign w45573 = w44773 & ~w44835;
assign w45574 = ~w44820 & ~w44847;
assign w45575 = ~w44786 & ~w45574;
assign w45576 = w44779 & w44843;
assign w45577 = w44793 & ~w44827;
assign w45578 = ~w44816 & ~w45577;
assign w45579 = ~w45576 & w45578;
assign w45580 = ~w45575 & w45579;
assign w45581 = ~w44806 & w44816;
assign w45582 = ~w44780 & ~w44792;
assign w45583 = ~w45510 & ~w45582;
assign w45584 = w44786 & ~w45583;
assign w45585 = ~w44832 & ~w45494;
assign w45586 = ~w45501 & w45585;
assign w45587 = w45581 & w45586;
assign w45588 = ~w45584 & w45587;
assign w45589 = ~w45580 & ~w45588;
assign w45590 = ~w45573 & ~w45589;
assign w45591 = ~pi2405 & w45590;
assign w45592 = pi2405 & ~w45590;
assign w45593 = ~w45591 & ~w45592;
assign w45594 = ~w45114 & w66592;
assign w45595 = w44894 & w45118;
assign w45596 = ~w44915 & ~w44922;
assign w45597 = w44878 & ~w45596;
assign w45598 = w44903 & ~w45555;
assign w45599 = ~w45595 & w45598;
assign w45600 = ~w44896 & w45599;
assign w45601 = ~w45597 & w45600;
assign w45602 = ~w45594 & ~w45601;
assign w45603 = w44918 & ~w45557;
assign w45604 = ~w44920 & ~w45595;
assign w45605 = ~w45125 & ~w45604;
assign w45606 = ~w45135 & ~w45603;
assign w45607 = ~w45605 & w45606;
assign w45608 = ~w45602 & w45607;
assign w45609 = pi2411 & ~w45608;
assign w45610 = ~pi2411 & w45608;
assign w45611 = ~w45609 & ~w45610;
assign w45612 = ~pi4855 & pi9040;
assign w45613 = ~pi5186 & ~pi9040;
assign w45614 = ~w45612 & ~w45613;
assign w45615 = pi2386 & ~w45614;
assign w45616 = ~pi2386 & w45614;
assign w45617 = ~w45615 & ~w45616;
assign w45618 = ~pi4868 & pi9040;
assign w45619 = ~pi4855 & ~pi9040;
assign w45620 = ~w45618 & ~w45619;
assign w45621 = pi2399 & ~w45620;
assign w45622 = ~pi2399 & w45620;
assign w45623 = ~w45621 & ~w45622;
assign w45624 = w45617 & ~w45623;
assign w45625 = ~pi4826 & pi9040;
assign w45626 = ~pi4939 & ~pi9040;
assign w45627 = ~w45625 & ~w45626;
assign w45628 = pi2380 & ~w45627;
assign w45629 = ~pi2380 & w45627;
assign w45630 = ~w45628 & ~w45629;
assign w45631 = w45624 & w45630;
assign w45632 = ~pi5081 & pi9040;
assign w45633 = ~pi4759 & ~pi9040;
assign w45634 = ~w45632 & ~w45633;
assign w45635 = pi2395 & ~w45634;
assign w45636 = ~pi2395 & w45634;
assign w45637 = ~w45635 & ~w45636;
assign w45638 = w45631 & w45637;
assign w45639 = ~pi4893 & pi9040;
assign w45640 = ~pi4824 & ~pi9040;
assign w45641 = ~w45639 & ~w45640;
assign w45642 = pi2376 & ~w45641;
assign w45643 = ~pi2376 & w45641;
assign w45644 = ~w45642 & ~w45643;
assign w45645 = ~pi4819 & pi9040;
assign w45646 = ~pi4952 & ~pi9040;
assign w45647 = ~w45645 & ~w45646;
assign w45648 = pi2355 & ~w45647;
assign w45649 = ~pi2355 & w45647;
assign w45650 = ~w45648 & ~w45649;
assign w45651 = w45617 & ~w45650;
assign w45652 = w45617 & ~w45630;
assign w45653 = w45650 & ~w45652;
assign w45654 = w45637 & ~w45650;
assign w45655 = ~w45623 & ~w45654;
assign w45656 = ~w45651 & ~w45653;
assign w45657 = w45655 & w45656;
assign w45658 = w45623 & ~w45637;
assign w45659 = ~w45617 & ~w45630;
assign w45660 = ~w45658 & ~w45659;
assign w45661 = ~w45617 & ~w45637;
assign w45662 = w45630 & ~w45637;
assign w45663 = w45650 & ~w45662;
assign w45664 = ~w45660 & ~w45661;
assign w45665 = ~w45663 & w45664;
assign w45666 = ~w45657 & ~w45665;
assign w45667 = w45624 & ~w45637;
assign w45668 = w45650 & ~w45667;
assign w45669 = ~w45623 & w45662;
assign w45670 = w45623 & ~w45630;
assign w45671 = ~w45669 & ~w45670;
assign w45672 = w45668 & ~w45671;
assign w45673 = ~w45644 & ~w45672;
assign w45674 = w45623 & w45637;
assign w45675 = w45652 & w45674;
assign w45676 = w45650 & w45661;
assign w45677 = ~w45631 & ~w45675;
assign w45678 = ~w45676 & w45677;
assign w45679 = ~w45673 & ~w45678;
assign w45680 = ~w45630 & ~w45637;
assign w45681 = ~w45617 & w45630;
assign w45682 = ~w45652 & ~w45681;
assign w45683 = w45637 & w45682;
assign w45684 = w45682 & w66593;
assign w45685 = ~w45680 & ~w45684;
assign w45686 = w45668 & ~w45685;
assign w45687 = w45637 & w45681;
assign w45688 = ~w45667 & ~w45687;
assign w45689 = ~w45650 & ~w45688;
assign w45690 = ~w45686 & ~w45689;
assign w45691 = w45644 & ~w45690;
assign w45692 = ~w45617 & w45623;
assign w45693 = w45654 & w45692;
assign w45694 = ~w45638 & ~w45693;
assign w45695 = (w45694 & w45666) | (w45694 & w66594) | (w45666 & w66594);
assign w45696 = ~w45679 & w45695;
assign w45697 = ~w45691 & w45696;
assign w45698 = pi2409 & ~w45697;
assign w45699 = ~pi2409 & w45697;
assign w45700 = ~w45698 & ~w45699;
assign w45701 = w44826 & ~w44844;
assign w45702 = ~w44842 & w45701;
assign w45703 = ~w44805 & ~w44816;
assign w45704 = ~w44827 & w45703;
assign w45705 = ~w45702 & ~w45704;
assign w45706 = ~w44786 & ~w45705;
assign w45707 = w44792 & w45701;
assign w45708 = ~w44829 & ~w45707;
assign w45709 = ~w44800 & w44809;
assign w45710 = w44779 & w44847;
assign w45711 = ~w44816 & w45708;
assign w45712 = ~w45710 & w45711;
assign w45713 = ~w45709 & w45712;
assign w45714 = w44817 & w45708;
assign w45715 = ~w44849 & w45581;
assign w45716 = ~w45714 & w45715;
assign w45717 = (~w45706 & w45713) | (~w45706 & w66595) | (w45713 & w66595);
assign w45718 = ~pi2404 & w45717;
assign w45719 = pi2404 & ~w45717;
assign w45720 = ~w45718 & ~w45719;
assign w45721 = w45012 & w45433;
assign w45722 = w44975 & ~w45048;
assign w45723 = ~w45721 & w45722;
assign w45724 = ~w45001 & ~w45022;
assign w45725 = ~w45023 & w45724;
assign w45726 = w45016 & w45725;
assign w45727 = ~w44975 & ~w45024;
assign w45728 = w45047 & w45727;
assign w45729 = ~w45726 & w45728;
assign w45730 = ~w45723 & ~w45729;
assign w45731 = w44994 & w45022;
assign w45732 = w45012 & ~w45731;
assign w45733 = ~w45460 & w45732;
assign w45734 = w44975 & w45032;
assign w45735 = ~w45005 & ~w45012;
assign w45736 = ~w45734 & w45735;
assign w45737 = ~w45733 & ~w45736;
assign w45738 = ~w45730 & ~w45737;
assign w45739 = pi2422 & w45738;
assign w45740 = ~pi2422 & ~w45738;
assign w45741 = ~w45739 & ~w45740;
assign w45742 = w45350 & ~w45391;
assign w45743 = ~w45336 & ~w45742;
assign w45744 = w45398 & w45743;
assign w45745 = w45386 & w45744;
assign w45746 = (~w45333 & w45745) | (~w45333 & w66596) | (w45745 & w66596);
assign w45747 = w45306 & ~w45319;
assign w45748 = ~w45342 & w45747;
assign w45749 = ~w45537 & w45748;
assign w45750 = w45333 & ~w45744;
assign w45751 = ~w45409 & ~w45749;
assign w45752 = ~w45750 & w45751;
assign w45753 = ~w45746 & w45752;
assign w45754 = pi2427 & ~w45753;
assign w45755 = ~pi2427 & w45753;
assign w45756 = ~w45754 & ~w45755;
assign w45757 = w45658 & ~w45682;
assign w45758 = ~w45650 & w45757;
assign w45759 = ~w45630 & w45637;
assign w45760 = ~w45659 & ~w45674;
assign w45761 = ~w45759 & ~w45760;
assign w45762 = ~w45760 & w66597;
assign w45763 = w45659 & w45674;
assign w45764 = ~w45650 & w45682;
assign w45765 = (~w45637 & ~w45682) | (~w45637 & w66598) | (~w45682 & w66598);
assign w45766 = (~w45623 & ~w45682) | (~w45623 & w66599) | (~w45682 & w66599);
assign w45767 = ~w45765 & w45766;
assign w45768 = w45668 & ~w45761;
assign w45769 = ~w45659 & ~w45680;
assign w45770 = w45768 & w45769;
assign w45771 = ~w45762 & ~w45763;
assign w45772 = ~w45767 & w45771;
assign w45773 = ~w45770 & w45772;
assign w45774 = w45644 & ~w45773;
assign w45775 = ~w45623 & w45654;
assign w45776 = ~w45764 & ~w45775;
assign w45777 = ~w45623 & w45683;
assign w45778 = ~w45776 & ~w45777;
assign w45779 = ~w45644 & ~w45768;
assign w45780 = ~w45778 & w45779;
assign w45781 = w45624 & w45759;
assign w45782 = w45661 & w45670;
assign w45783 = ~w45781 & ~w45782;
assign w45784 = w45650 & ~w45783;
assign w45785 = ~w45758 & ~w45784;
assign w45786 = ~w45780 & w45785;
assign w45787 = ~w45774 & w45786;
assign w45788 = pi2410 & ~w45787;
assign w45789 = ~pi2410 & w45787;
assign w45790 = ~w45788 & ~w45789;
assign w45791 = w45623 & w45630;
assign w45792 = w45676 & w45791;
assign w45793 = w45617 & ~w45671;
assign w45794 = ~w45644 & w45684;
assign w45795 = ~w45793 & ~w45794;
assign w45796 = w45650 & ~w45795;
assign w45797 = ~w45630 & w45693;
assign w45798 = w45651 & w45662;
assign w45799 = ~w45669 & w45688;
assign w45800 = ~w45668 & ~w45799;
assign w45801 = ~w45644 & ~w45675;
assign w45802 = ~w45782 & ~w45798;
assign w45803 = w45801 & w45802;
assign w45804 = ~w45800 & w45803;
assign w45805 = ~w45617 & ~w45759;
assign w45806 = ~w45658 & w45805;
assign w45807 = w45663 & w45806;
assign w45808 = w45644 & ~w45775;
assign w45809 = ~w45757 & w45808;
assign w45810 = ~w45807 & w45809;
assign w45811 = ~w45804 & ~w45810;
assign w45812 = ~w45792 & ~w45797;
assign w45813 = ~w45796 & w45812;
assign w45814 = ~w45811 & w45813;
assign w45815 = pi2413 & ~w45814;
assign w45816 = ~pi2413 & w45814;
assign w45817 = ~w45815 & ~w45816;
assign w45818 = ~w45655 & w45805;
assign w45819 = w45653 & ~w45669;
assign w45820 = w45663 & ~w45759;
assign w45821 = ~w45650 & ~w45680;
assign w45822 = ~w45791 & w45821;
assign w45823 = ~w45820 & ~w45822;
assign w45824 = ~w45819 & w45823;
assign w45825 = ~w45644 & ~w45818;
assign w45826 = ~w45824 & w45825;
assign w45827 = w45760 & w45820;
assign w45828 = w45644 & ~w45763;
assign w45829 = ~w45798 & w45828;
assign w45830 = ~w45638 & w45829;
assign w45831 = ~w45827 & w45830;
assign w45832 = ~w45826 & ~w45831;
assign w45833 = w45777 & w45823;
assign w45834 = ~w45760 & w45806;
assign w45835 = ~w45781 & ~w45834;
assign w45836 = ~w45650 & ~w45835;
assign w45837 = ~w45792 & ~w45833;
assign w45838 = ~w45836 & w45837;
assign w45839 = ~w45832 & w45838;
assign w45840 = pi2418 & ~w45839;
assign w45841 = ~pi2418 & w45839;
assign w45842 = ~w45840 & ~w45841;
assign w45843 = ~pi5107 & pi9040;
assign w45844 = ~pi5101 & ~pi9040;
assign w45845 = ~w45843 & ~w45844;
assign w45846 = pi2456 & ~w45845;
assign w45847 = ~pi2456 & w45845;
assign w45848 = ~w45846 & ~w45847;
assign w45849 = ~pi4979 & pi9040;
assign w45850 = ~pi5290 & ~pi9040;
assign w45851 = ~w45849 & ~w45850;
assign w45852 = pi2424 & ~w45851;
assign w45853 = ~pi2424 & w45851;
assign w45854 = ~w45852 & ~w45853;
assign w45855 = ~w45848 & w45854;
assign w45856 = ~pi5418 & pi9040;
assign w45857 = ~pi5107 & ~pi9040;
assign w45858 = ~w45856 & ~w45857;
assign w45859 = pi2452 & ~w45858;
assign w45860 = ~pi2452 & w45858;
assign w45861 = ~w45859 & ~w45860;
assign w45862 = ~pi5046 & pi9040;
assign w45863 = ~pi5094 & ~pi9040;
assign w45864 = ~w45862 & ~w45863;
assign w45865 = pi2439 & ~w45864;
assign w45866 = ~pi2439 & w45864;
assign w45867 = ~w45865 & ~w45866;
assign w45868 = ~w45861 & ~w45867;
assign w45869 = w45855 & w45868;
assign w45870 = w45848 & ~w45861;
assign w45871 = ~pi5104 & pi9040;
assign w45872 = ~pi4989 & ~pi9040;
assign w45873 = ~w45871 & ~w45872;
assign w45874 = pi2440 & ~w45873;
assign w45875 = ~pi2440 & w45873;
assign w45876 = ~w45874 & ~w45875;
assign w45877 = w45867 & w45876;
assign w45878 = w45870 & w45877;
assign w45879 = w45854 & w45867;
assign w45880 = ~w45854 & ~w45867;
assign w45881 = ~w45870 & w45880;
assign w45882 = w45848 & ~w45854;
assign w45883 = w45861 & w45867;
assign w45884 = ~w45855 & ~w45879;
assign w45885 = ~w45880 & ~w45883;
assign w45886 = w45884 & w45885;
assign w45887 = w45861 & w45886;
assign w45888 = ~w45887 & w64024;
assign w45889 = ~pi5102 & pi9040;
assign w45890 = ~pi5053 & ~pi9040;
assign w45891 = ~w45889 & ~w45890;
assign w45892 = pi2461 & ~w45891;
assign w45893 = ~pi2461 & w45891;
assign w45894 = ~w45892 & ~w45893;
assign w45895 = ~w45876 & ~w45894;
assign w45896 = ~w45883 & w45895;
assign w45897 = ~w45888 & w45896;
assign w45898 = ~w45848 & w45867;
assign w45899 = ~w45884 & ~w45898;
assign w45900 = ~w45848 & ~w45854;
assign w45901 = ~w45868 & ~w45883;
assign w45902 = w45900 & w45901;
assign w45903 = w45881 & ~w45902;
assign w45904 = w45876 & ~w45894;
assign w45905 = (w45904 & w45903) | (w45904 & w66600) | (w45903 & w66600);
assign w45906 = (w45876 & w45887) | (w45876 & w64025) | (w45887 & w64025);
assign w45907 = w45854 & ~w45876;
assign w45908 = w45868 & w45907;
assign w45909 = w45855 & w45883;
assign w45910 = ~w45908 & ~w45909;
assign w45911 = ~w45902 & w45910;
assign w45912 = ~w45906 & w45911;
assign w45913 = w45854 & w45883;
assign w45914 = w45848 & w45880;
assign w45915 = ~w45913 & ~w45914;
assign w45916 = ~w45876 & ~w45915;
assign w45917 = ~w45861 & ~w45876;
assign w45918 = ~w45848 & w45917;
assign w45919 = ~w45879 & w45918;
assign w45920 = ~w45916 & ~w45919;
assign w45921 = (~w45870 & w45916) | (~w45870 & w66601) | (w45916 & w66601);
assign w45922 = (w45894 & ~w45912) | (w45894 & w66602) | (~w45912 & w66602);
assign w45923 = w45883 & ~w45894;
assign w45924 = w45900 & w45923;
assign w45925 = ~w45869 & ~w45878;
assign w45926 = ~w45924 & w45925;
assign w45927 = ~w45905 & w45926;
assign w45928 = ~w45897 & w45927;
assign w45929 = ~w45922 & w45928;
assign w45930 = ~pi2475 & ~w45929;
assign w45931 = pi2475 & w45929;
assign w45932 = ~w45930 & ~w45931;
assign w45933 = w45848 & w45854;
assign w45934 = ~w45877 & ~w45933;
assign w45935 = ~w45887 & w66603;
assign w45936 = w45854 & ~w45870;
assign w45937 = ~w45854 & ~w45861;
assign w45938 = ~w45900 & ~w45937;
assign w45939 = (~w45876 & w45870) | (~w45876 & w64026) | (w45870 & w64026);
assign w45940 = w45938 & w45939;
assign w45941 = w45910 & ~w45940;
assign w45942 = ~w45935 & w45941;
assign w45943 = w45861 & w45882;
assign w45944 = w45876 & ~w45943;
assign w45945 = w45855 & w45861;
assign w45946 = w45899 & ~w45945;
assign w45947 = w45944 & ~w45946;
assign w45948 = w45894 & ~w45940;
assign w45949 = w45920 & w45948;
assign w45950 = ~w45947 & w45949;
assign w45951 = ~w45911 & w45935;
assign w45952 = ~w45915 & w45944;
assign w45953 = ~w45937 & ~w45945;
assign w45954 = w45904 & ~w45953;
assign w45955 = w45880 & w45918;
assign w45956 = ~w45952 & ~w45955;
assign w45957 = ~w45954 & w45956;
assign w45958 = ~w45950 & w66604;
assign w45959 = (pi2474 & ~w45958) | (pi2474 & w64027) | (~w45958 & w64027);
assign w45960 = w45958 & w64028;
assign w45961 = ~w45959 & ~w45960;
assign w45962 = w45870 & w45880;
assign w45963 = ~w45914 & ~w45936;
assign w45964 = ~w45917 & w45938;
assign w45965 = ~w45945 & w45964;
assign w45966 = w45963 & w45965;
assign w45967 = ~w45848 & w45907;
assign w45968 = ~w45962 & ~w45967;
assign w45969 = ~w45902 & w45968;
assign w45970 = ~w45966 & w45969;
assign w45971 = (w45894 & ~w45970) | (w45894 & w66605) | (~w45970 & w66605);
assign w45972 = w45879 & w45918;
assign w45973 = w45904 & ~w45963;
assign w45974 = w45923 & w45933;
assign w45975 = ~w45854 & w45895;
assign w45976 = ~w45898 & w45975;
assign w45977 = ~w45914 & w45976;
assign w45978 = ~w45972 & ~w45974;
assign w45979 = ~w45973 & w45978;
assign w45980 = ~w45977 & w45979;
assign w45981 = ~w45951 & w45980;
assign w45982 = ~w45971 & w45981;
assign w45983 = ~pi2477 & w45982;
assign w45984 = pi2477 & ~w45982;
assign w45985 = ~w45983 & ~w45984;
assign w45986 = ~w45886 & ~w45909;
assign w45987 = ~w45913 & w45953;
assign w45988 = w45986 & ~w45987;
assign w45989 = ~w45894 & w45914;
assign w45990 = ~w45924 & ~w45989;
assign w45991 = (~w45876 & w45988) | (~w45876 & w66606) | (w45988 & w66606);
assign w45992 = w45876 & ~w45986;
assign w45993 = w45879 & w45917;
assign w45994 = ~w45869 & ~w45894;
assign w45995 = ~w45993 & w45994;
assign w45996 = ~w45992 & w45995;
assign w45997 = w45964 & w66607;
assign w45998 = w45884 & w45917;
assign w45999 = w45894 & ~w45962;
assign w46000 = ~w45998 & w45999;
assign w46001 = ~w45997 & w46000;
assign w46002 = ~w45996 & ~w46001;
assign w46003 = w45876 & w45953;
assign w46004 = ~w45912 & w46003;
assign w46005 = ~w45991 & ~w46002;
assign w46006 = w46005 & w66608;
assign w46007 = (pi2495 & ~w46005) | (pi2495 & w66609) | (~w46005 & w66609);
assign w46008 = ~w46006 & ~w46007;
assign w46009 = ~pi5458 & pi9040;
assign w46010 = ~pi5106 & ~pi9040;
assign w46011 = ~w46009 & ~w46010;
assign w46012 = pi2438 & ~w46011;
assign w46013 = ~pi2438 & w46011;
assign w46014 = ~w46012 & ~w46013;
assign w46015 = ~pi5097 & pi9040;
assign w46016 = ~pi5080 & ~pi9040;
assign w46017 = ~w46015 & ~w46016;
assign w46018 = pi2429 & ~w46017;
assign w46019 = ~pi2429 & w46017;
assign w46020 = ~w46018 & ~w46019;
assign w46021 = w46014 & w46020;
assign w46022 = ~pi5053 & pi9040;
assign w46023 = ~pi5281 & ~pi9040;
assign w46024 = ~w46022 & ~w46023;
assign w46025 = pi2459 & ~w46024;
assign w46026 = ~pi2459 & w46024;
assign w46027 = ~w46025 & ~w46026;
assign w46028 = ~pi4974 & pi9040;
assign w46029 = ~pi5332 & ~pi9040;
assign w46030 = ~w46028 & ~w46029;
assign w46031 = pi2433 & ~w46030;
assign w46032 = ~pi2433 & w46030;
assign w46033 = ~w46031 & ~w46032;
assign w46034 = w46027 & w46033;
assign w46035 = ~w46027 & ~w46033;
assign w46036 = ~w46034 & ~w46035;
assign w46037 = w46021 & ~w46036;
assign w46038 = w46014 & w46033;
assign w46039 = ~pi5057 & pi9040;
assign w46040 = ~pi5049 & ~pi9040;
assign w46041 = ~w46039 & ~w46040;
assign w46042 = pi2423 & ~w46041;
assign w46043 = ~pi2423 & w46041;
assign w46044 = ~w46042 & ~w46043;
assign w46045 = ~w46038 & ~w46044;
assign w46046 = w46020 & ~w46027;
assign w46047 = ~w46020 & w46027;
assign w46048 = ~w46046 & ~w46047;
assign w46049 = ~w46034 & ~w46048;
assign w46050 = w46045 & ~w46049;
assign w46051 = ~w46014 & ~w46033;
assign w46052 = w46027 & w46051;
assign w46053 = w46051 & w66610;
assign w46054 = ~w46014 & ~w46020;
assign w46055 = w46033 & w46054;
assign w46056 = (w46044 & ~w46054) | (w46044 & w66611) | (~w46054 & w66611);
assign w46057 = ~w46053 & w46056;
assign w46058 = (~w46037 & w46050) | (~w46037 & w66612) | (w46050 & w66612);
assign w46059 = ~pi5101 & pi9040;
assign w46060 = ~pi5097 & ~pi9040;
assign w46061 = ~w46059 & ~w46060;
assign w46062 = pi2458 & ~w46061;
assign w46063 = ~pi2458 & w46061;
assign w46064 = ~w46062 & ~w46063;
assign w46065 = ~w46058 & ~w46064;
assign w46066 = w46014 & ~w46033;
assign w46067 = w46014 & ~w46020;
assign w46068 = ~w46066 & ~w46067;
assign w46069 = w46027 & ~w46068;
assign w46070 = ~w46046 & ~w46066;
assign w46071 = w46020 & w46066;
assign w46072 = ~w46070 & ~w46071;
assign w46073 = w46044 & ~w46072;
assign w46074 = ~w46069 & w46073;
assign w46075 = ~w46014 & w46048;
assign w46076 = w46034 & w46067;
assign w46077 = ~w46044 & ~w46076;
assign w46078 = ~w46075 & w46077;
assign w46079 = ~w46074 & ~w46078;
assign w46080 = w46064 & w46079;
assign w46081 = w46014 & ~w46027;
assign w46082 = ~w46033 & ~w46067;
assign w46083 = ~w46081 & ~w46082;
assign w46084 = ~w46070 & w46083;
assign w46085 = ~w46036 & w46054;
assign w46086 = w46044 & ~w46085;
assign w46087 = ~w46084 & w46086;
assign w46088 = w46046 & w46066;
assign w46089 = ~w46044 & ~w46088;
assign w46090 = ~w46087 & ~w46089;
assign w46091 = ~w46065 & ~w46090;
assign w46092 = ~w46080 & w46091;
assign w46093 = ~pi2464 & w46092;
assign w46094 = pi2464 & ~w46092;
assign w46095 = ~w46093 & ~w46094;
assign w46096 = ~pi5332 & pi9040;
assign w46097 = ~pi5051 & ~pi9040;
assign w46098 = ~w46096 & ~w46097;
assign w46099 = pi2439 & ~w46098;
assign w46100 = ~pi2439 & w46098;
assign w46101 = ~w46099 & ~w46100;
assign w46102 = ~pi5281 & pi9040;
assign w46103 = ~pi5181 & ~pi9040;
assign w46104 = ~w46102 & ~w46103;
assign w46105 = pi2417 & ~w46104;
assign w46106 = ~pi2417 & w46104;
assign w46107 = ~w46105 & ~w46106;
assign w46108 = ~pi5342 & pi9040;
assign w46109 = ~pi5102 & ~pi9040;
assign w46110 = ~w46108 & ~w46109;
assign w46111 = pi2461 & ~w46110;
assign w46112 = ~pi2461 & w46110;
assign w46113 = ~w46111 & ~w46112;
assign w46114 = w46107 & ~w46113;
assign w46115 = ~w46107 & w46113;
assign w46116 = ~w46114 & ~w46115;
assign w46117 = ~pi5181 & pi9040;
assign w46118 = ~pi5104 & ~pi9040;
assign w46119 = ~w46117 & ~w46118;
assign w46120 = pi2455 & ~w46119;
assign w46121 = ~pi2455 & w46119;
assign w46122 = ~w46120 & ~w46121;
assign w46123 = w46101 & ~w46122;
assign w46124 = w46116 & w46123;
assign w46125 = ~pi5049 & pi9040;
assign w46126 = ~pi5458 & ~pi9040;
assign w46127 = ~w46125 & ~w46126;
assign w46128 = pi2438 & ~w46127;
assign w46129 = ~pi2438 & w46127;
assign w46130 = ~w46128 & ~w46129;
assign w46131 = ~w46101 & ~w46130;
assign w46132 = w46101 & w46130;
assign w46133 = ~w46131 & ~w46132;
assign w46134 = w46114 & w46133;
assign w46135 = ~w46131 & ~w46134;
assign w46136 = w46114 & w46131;
assign w46137 = w46122 & ~w46136;
assign w46138 = ~w46135 & w46137;
assign w46139 = ~pi4989 & pi9040;
assign w46140 = ~pi5418 & ~pi9040;
assign w46141 = ~w46139 & ~w46140;
assign w46142 = pi2429 & ~w46141;
assign w46143 = ~pi2429 & w46141;
assign w46144 = ~w46142 & ~w46143;
assign w46145 = ~w46122 & w46130;
assign w46146 = ~w46132 & ~w46145;
assign w46147 = w46116 & ~w46146;
assign w46148 = w46101 & ~w46130;
assign w46149 = ~w46136 & ~w46148;
assign w46150 = w46101 & ~w46113;
assign w46151 = ~w46130 & w46150;
assign w46152 = ~w46101 & w46107;
assign w46153 = w46113 & w46130;
assign w46154 = w46152 & w46153;
assign w46155 = ~w46122 & ~w46151;
assign w46156 = ~w46154 & w46155;
assign w46157 = ~w46149 & w46156;
assign w46158 = ~w46101 & w46115;
assign w46159 = ~w46145 & w46158;
assign w46160 = ~w46144 & ~w46147;
assign w46161 = ~w46159 & w46160;
assign w46162 = ~w46157 & w46161;
assign w46163 = ~w46107 & w46132;
assign w46164 = ~w46152 & ~w46163;
assign w46165 = w46113 & w46122;
assign w46166 = ~w46164 & w46165;
assign w46167 = ~w46113 & w46130;
assign w46168 = w46152 & w46167;
assign w46169 = ~w46113 & ~w46130;
assign w46170 = ~w46101 & ~w46107;
assign w46171 = w46169 & w46170;
assign w46172 = w46153 & w46170;
assign w46173 = ~w46150 & ~w46172;
assign w46174 = w46156 & ~w46173;
assign w46175 = w46144 & ~w46168;
assign w46176 = ~w46171 & w46175;
assign w46177 = ~w46166 & w46176;
assign w46178 = ~w46174 & w46177;
assign w46179 = ~w46162 & ~w46178;
assign w46180 = ~w46124 & ~w46138;
assign w46181 = ~w46179 & w46180;
assign w46182 = pi2465 & ~w46181;
assign w46183 = ~pi2465 & w46181;
assign w46184 = ~w46182 & ~w46183;
assign w46185 = ~pi5110 & pi9040;
assign w46186 = ~pi5327 & ~pi9040;
assign w46187 = ~w46185 & ~w46186;
assign w46188 = pi2462 & ~w46187;
assign w46189 = ~pi2462 & w46187;
assign w46190 = ~w46188 & ~w46189;
assign w46191 = ~pi5208 & pi9040;
assign w46192 = ~pi5542 & ~pi9040;
assign w46193 = ~w46191 & ~w46192;
assign w46194 = pi2448 & ~w46193;
assign w46195 = ~pi2448 & w46193;
assign w46196 = ~w46194 & ~w46195;
assign w46197 = ~pi5108 & pi9040;
assign w46198 = ~pi5291 & ~pi9040;
assign w46199 = ~w46197 & ~w46198;
assign w46200 = pi2432 & ~w46199;
assign w46201 = ~pi2432 & w46199;
assign w46202 = ~w46200 & ~w46201;
assign w46203 = w46196 & ~w46202;
assign w46204 = ~pi5206 & pi9040;
assign w46205 = ~pi5055 & ~pi9040;
assign w46206 = ~w46204 & ~w46205;
assign w46207 = pi2463 & ~w46206;
assign w46208 = ~pi2463 & w46206;
assign w46209 = ~w46207 & ~w46208;
assign w46210 = ~w46203 & ~w46209;
assign w46211 = ~pi5327 & pi9040;
assign w46212 = ~pi5103 & ~pi9040;
assign w46213 = ~w46211 & ~w46212;
assign w46214 = pi2426 & ~w46213;
assign w46215 = ~pi2426 & w46213;
assign w46216 = ~w46214 & ~w46215;
assign w46217 = ~pi5291 & pi9040;
assign w46218 = ~pi4971 & ~pi9040;
assign w46219 = ~w46217 & ~w46218;
assign w46220 = pi2453 & ~w46219;
assign w46221 = ~pi2453 & w46219;
assign w46222 = ~w46220 & ~w46221;
assign w46223 = w46216 & ~w46222;
assign w46224 = ~w46202 & ~w46223;
assign w46225 = w46216 & w46222;
assign w46226 = w46202 & ~w46225;
assign w46227 = ~w46224 & ~w46226;
assign w46228 = w46210 & w46227;
assign w46229 = ~w46196 & ~w46209;
assign w46230 = ~w46202 & w46216;
assign w46231 = ~w46196 & w46209;
assign w46232 = ~w46230 & w46231;
assign w46233 = ~w46203 & ~w46232;
assign w46234 = w46222 & ~w46233;
assign w46235 = ~w46225 & ~w46230;
assign w46236 = w46196 & ~w46222;
assign w46237 = w46202 & ~w46216;
assign w46238 = w46236 & w46237;
assign w46239 = ~w46229 & w46235;
assign w46240 = ~w46238 & w46239;
assign w46241 = ~w46234 & w46240;
assign w46242 = ~w46228 & ~w46241;
assign w46243 = w46190 & ~w46242;
assign w46244 = w46196 & w46209;
assign w46245 = ~w46216 & w46222;
assign w46246 = w46244 & w46245;
assign w46247 = w46203 & w46223;
assign w46248 = ~w46246 & ~w46247;
assign w46249 = ~w46196 & w46222;
assign w46250 = ~w46202 & w46249;
assign w46251 = w46248 & ~w46250;
assign w46252 = w46229 & w46235;
assign w46253 = w46202 & ~w46223;
assign w46254 = w46244 & w46253;
assign w46255 = ~w46252 & ~w46254;
assign w46256 = w46251 & w46255;
assign w46257 = ~w46190 & ~w46256;
assign w46258 = w46196 & ~w46245;
assign w46259 = ~w46245 & w66613;
assign w46260 = w46210 & w46245;
assign w46261 = ~w46259 & ~w46260;
assign w46262 = w46224 & ~w46261;
assign w46263 = w46209 & w46216;
assign w46264 = ~w46251 & w46263;
assign w46265 = ~w46262 & ~w46264;
assign w46266 = ~w46257 & w46265;
assign w46267 = ~w46243 & w46266;
assign w46268 = pi2476 & ~w46267;
assign w46269 = ~pi2476 & w46267;
assign w46270 = ~w46268 & ~w46269;
assign w46271 = w46107 & w46113;
assign w46272 = w46101 & w46107;
assign w46273 = ~w46271 & ~w46272;
assign w46274 = ~w46135 & ~w46273;
assign w46275 = ~w46113 & ~w46146;
assign w46276 = ~w46164 & w46275;
assign w46277 = w46101 & w46113;
assign w46278 = ~w46171 & ~w46277;
assign w46279 = w46122 & ~w46278;
assign w46280 = w46144 & ~w46172;
assign w46281 = ~w46276 & w46280;
assign w46282 = ~w46279 & w46281;
assign w46283 = ~w46274 & w46282;
assign w46284 = ~w46153 & ~w46169;
assign w46285 = ~w46107 & ~w46284;
assign w46286 = ~w46284 & w66614;
assign w46287 = ~w46136 & ~w46286;
assign w46288 = ~w46130 & ~w46287;
assign w46289 = w46133 & ~w46271;
assign w46290 = ~w46113 & w46272;
assign w46291 = w46122 & ~w46290;
assign w46292 = ~w46289 & ~w46291;
assign w46293 = w46170 & w46284;
assign w46294 = ~w46167 & ~w46293;
assign w46295 = w46146 & ~w46294;
assign w46296 = ~w46144 & ~w46154;
assign w46297 = ~w46292 & w46296;
assign w46298 = ~w46295 & w46297;
assign w46299 = ~w46288 & w46298;
assign w46300 = ~w46283 & ~w46299;
assign w46301 = pi2466 & w46300;
assign w46302 = ~pi2466 & ~w46300;
assign w46303 = ~w46301 & ~w46302;
assign w46304 = ~pi5100 & pi9040;
assign w46305 = ~pi5099 & ~pi9040;
assign w46306 = ~w46304 & ~w46305;
assign w46307 = pi2426 & ~w46306;
assign w46308 = ~pi2426 & w46306;
assign w46309 = ~w46307 & ~w46308;
assign w46310 = ~pi5106 & pi9040;
assign w46311 = ~pi5046 & ~pi9040;
assign w46312 = ~w46310 & ~w46311;
assign w46313 = pi2450 & ~w46312;
assign w46314 = ~pi2450 & w46312;
assign w46315 = ~w46313 & ~w46314;
assign w46316 = w46309 & ~w46315;
assign w46317 = ~pi5094 & pi9040;
assign w46318 = ~pi5036 & ~pi9040;
assign w46319 = ~w46317 & ~w46318;
assign w46320 = pi2442 & ~w46319;
assign w46321 = ~pi2442 & w46319;
assign w46322 = ~w46320 & ~w46321;
assign w46323 = ~pi5093 & pi9040;
assign w46324 = ~pi5342 & ~pi9040;
assign w46325 = ~w46323 & ~w46324;
assign w46326 = pi2456 & ~w46325;
assign w46327 = ~pi2456 & w46325;
assign w46328 = ~w46326 & ~w46327;
assign w46329 = w46322 & ~w46328;
assign w46330 = ~w46316 & w46329;
assign w46331 = w46309 & w46330;
assign w46332 = ~pi5290 & pi9040;
assign w46333 = ~pi5057 & ~pi9040;
assign w46334 = ~w46332 & ~w46333;
assign w46335 = pi2424 & ~w46334;
assign w46336 = ~pi2424 & w46334;
assign w46337 = ~w46335 & ~w46336;
assign w46338 = ~pi5099 & pi9040;
assign w46339 = ~pi4979 & ~pi9040;
assign w46340 = ~w46338 & ~w46339;
assign w46341 = pi2462 & ~w46340;
assign w46342 = ~pi2462 & w46340;
assign w46343 = ~w46341 & ~w46342;
assign w46344 = ~w46315 & w46343;
assign w46345 = ~w46309 & ~w46328;
assign w46346 = w46309 & w46328;
assign w46347 = ~w46345 & ~w46346;
assign w46348 = ~w46344 & ~w46347;
assign w46349 = w46315 & ~w46343;
assign w46350 = w46337 & ~w46349;
assign w46351 = ~w46348 & ~w46350;
assign w46352 = w46328 & w46343;
assign w46353 = ~w46309 & w46352;
assign w46354 = ~w46315 & ~w46343;
assign w46355 = w46345 & w46354;
assign w46356 = ~w46353 & ~w46355;
assign w46357 = w46322 & ~w46356;
assign w46358 = ~w46322 & w46344;
assign w46359 = (~w46358 & w46348) | (~w46358 & w66615) | (w46348 & w66615);
assign w46360 = ~w46357 & w46359;
assign w46361 = w46337 & ~w46360;
assign w46362 = ~w46309 & w46315;
assign w46363 = ~w46328 & ~w46343;
assign w46364 = w46309 & w46354;
assign w46365 = w46315 & w46352;
assign w46366 = ~w46364 & ~w46365;
assign w46367 = w46322 & ~w46345;
assign w46368 = ~w46363 & w46367;
assign w46369 = w46366 & w46368;
assign w46370 = w46362 & w46369;
assign w46371 = w46328 & w46354;
assign w46372 = w46322 & ~w46371;
assign w46373 = w46309 & w46322;
assign w46374 = w46315 & w46343;
assign w46375 = ~w46309 & w46374;
assign w46376 = ~w46328 & w46375;
assign w46377 = ~w46373 & ~w46376;
assign w46378 = ~w46372 & ~w46377;
assign w46379 = ~w46328 & w46343;
assign w46380 = w46309 & w46379;
assign w46381 = ~w46309 & w46363;
assign w46382 = ~w46380 & ~w46381;
assign w46383 = w46315 & ~w46382;
assign w46384 = ~w46328 & ~w46374;
assign w46385 = ~w46316 & w46384;
assign w46386 = ~w46309 & ~w46379;
assign w46387 = ~w46352 & ~w46386;
assign w46388 = ~w46353 & ~w46387;
assign w46389 = (w46322 & w46388) | (w46322 & w64029) | (w46388 & w64029);
assign w46390 = w46343 & w46389;
assign w46391 = ~w46353 & ~w46371;
assign w46392 = ~w46322 & ~w46391;
assign w46393 = ~w46322 & ~w46343;
assign w46394 = w46346 & w46393;
assign w46395 = ~w46364 & ~w46394;
assign w46396 = ~w46383 & w46395;
assign w46397 = ~w46392 & w46396;
assign w46398 = ~w46390 & w46397;
assign w46399 = ~w46337 & ~w46398;
assign w46400 = (~w46331 & ~w46369) | (~w46331 & w66616) | (~w46369 & w66616);
assign w46401 = ~w46378 & w46400;
assign w46402 = ~w46361 & w46401;
assign w46403 = (pi2489 & w46399) | (pi2489 & w66617) | (w46399 & w66617);
assign w46404 = ~w46399 & w66618;
assign w46405 = ~w46403 & ~w46404;
assign w46406 = w46122 & ~w46286;
assign w46407 = ~w46122 & ~w46290;
assign w46408 = ~w46101 & ~w46116;
assign w46409 = ~w46151 & ~w46153;
assign w46410 = ~w46408 & w46409;
assign w46411 = w46407 & ~w46410;
assign w46412 = w46272 & w46284;
assign w46413 = ~w46154 & ~w46412;
assign w46414 = (w46413 & w46411) | (w46413 & w66619) | (w46411 & w66619);
assign w46415 = w46144 & ~w46414;
assign w46416 = ~w46144 & ~w46285;
assign w46417 = w46413 & w46416;
assign w46418 = w46137 & ~w46417;
assign w46419 = ~w46144 & ~w46287;
assign w46420 = ~w46122 & w46413;
assign w46421 = ~w46419 & w46420;
assign w46422 = ~w46418 & ~w46421;
assign w46423 = ~w46415 & ~w46422;
assign w46424 = ~pi2468 & w46423;
assign w46425 = pi2468 & ~w46423;
assign w46426 = ~w46424 & ~w46425;
assign w46427 = ~w46196 & w46216;
assign w46428 = (w46209 & w46250) | (w46209 & w64030) | (w46250 & w64030);
assign w46429 = ~w46236 & ~w46249;
assign w46430 = w46226 & w46429;
assign w46431 = ~w46428 & ~w46430;
assign w46432 = w46231 & w46431;
assign w46433 = ~w46202 & w46246;
assign w46434 = ~w46209 & w46247;
assign w46435 = ~w46202 & ~w46209;
assign w46436 = ~w46429 & w46435;
assign w46437 = w46237 & w46429;
assign w46438 = w46229 & w46437;
assign w46439 = w46196 & w46202;
assign w46440 = w46225 & w46439;
assign w46441 = w46223 & w46231;
assign w46442 = w46190 & ~w46440;
assign w46443 = ~w46441 & w46442;
assign w46444 = w46248 & ~w46436;
assign w46445 = w46443 & w46444;
assign w46446 = ~w46438 & w46445;
assign w46447 = ~w46216 & ~w46222;
assign w46448 = ~w46196 & ~w46202;
assign w46449 = w46447 & w46448;
assign w46450 = ~w46190 & ~w46238;
assign w46451 = ~w46449 & w46450;
assign w46452 = w46209 & ~w46222;
assign w46453 = w46439 & w46452;
assign w46454 = ~w46244 & ~w46448;
assign w46455 = w46225 & ~w46454;
assign w46456 = w46202 & w46245;
assign w46457 = ~w46427 & ~w46456;
assign w46458 = ~w46209 & ~w46457;
assign w46459 = w46231 & w46447;
assign w46460 = ~w46453 & ~w46459;
assign w46461 = ~w46455 & w46460;
assign w46462 = w46451 & w46461;
assign w46463 = ~w46458 & w46462;
assign w46464 = ~w46446 & ~w46463;
assign w46465 = ~w46433 & ~w46434;
assign w46466 = ~w46432 & w46465;
assign w46467 = ~w46464 & w46466;
assign w46468 = ~pi2473 & w46467;
assign w46469 = pi2473 & ~w46467;
assign w46470 = ~w46468 & ~w46469;
assign w46471 = w46316 & w46352;
assign w46472 = w46315 & w46328;
assign w46473 = w46309 & ~w46472;
assign w46474 = ~w46384 & w46473;
assign w46475 = ~w46389 & ~w46474;
assign w46476 = w46337 & ~w46475;
assign w46477 = w46329 & w46383;
assign w46478 = ~w46353 & ~w46364;
assign w46479 = (~w46375 & w46478) | (~w46375 & w66620) | (w46478 & w66620);
assign w46480 = ~w46322 & ~w46479;
assign w46481 = w46309 & ~w46349;
assign w46482 = ~w46322 & w46354;
assign w46483 = w46386 & ~w46482;
assign w46484 = (~w46329 & w46483) | (~w46329 & w66621) | (w46483 & w66621);
assign w46485 = ~w46330 & ~w46337;
assign w46486 = ~w46484 & w46485;
assign w46487 = (~w46471 & ~w46369) | (~w46471 & w66622) | (~w46369 & w66622);
assign w46488 = ~w46477 & w46487;
assign w46489 = ~w46480 & ~w46486;
assign w46490 = w46488 & w46489;
assign w46491 = ~w46476 & w46490;
assign w46492 = pi2496 & ~w46491;
assign w46493 = ~pi2496 & w46491;
assign w46494 = ~w46492 & ~w46493;
assign w46495 = ~w46316 & ~w46362;
assign w46496 = ~w46382 & ~w46495;
assign w46497 = (~w46337 & ~w46366) | (~w46337 & w66623) | (~w46366 & w66623);
assign w46498 = ~w46496 & ~w46497;
assign w46499 = w46322 & ~w46498;
assign w46500 = w46344 & w46347;
assign w46501 = ~w46374 & ~w46482;
assign w46502 = ~w46347 & ~w46373;
assign w46503 = ~w46501 & w46502;
assign w46504 = ~w46369 & ~w46500;
assign w46505 = ~w46503 & w46504;
assign w46506 = w46337 & ~w46505;
assign w46507 = ~w46322 & ~w46500;
assign w46508 = w46351 & w46507;
assign w46509 = ~w46499 & ~w46508;
assign w46510 = ~w46506 & w46509;
assign w46511 = ~pi2502 & w46510;
assign w46512 = pi2502 & ~w46510;
assign w46513 = ~w46511 & ~w46512;
assign w46514 = w46020 & ~w46038;
assign w46515 = ~w46027 & ~w46067;
assign w46516 = ~w46514 & w46515;
assign w46517 = ~w46079 & w46516;
assign w46518 = ~w46014 & w46033;
assign w46519 = ~w46027 & w46518;
assign w46520 = w46044 & w46519;
assign w46521 = ~w46054 & ~w46071;
assign w46522 = w46036 & ~w46521;
assign w46523 = ~w46036 & ~w46044;
assign w46524 = w46514 & w46523;
assign w46525 = ~w46035 & w46044;
assign w46526 = w46014 & w46525;
assign w46527 = ~w46072 & w46526;
assign w46528 = w46064 & ~w46520;
assign w46529 = ~w46522 & w46528;
assign w46530 = ~w46524 & ~w46527;
assign w46531 = w46529 & w46530;
assign w46532 = w46044 & ~w46067;
assign w46533 = ~w46048 & ~w46082;
assign w46534 = ~w46532 & w46533;
assign w46535 = ~w46072 & w66624;
assign w46536 = ~w46075 & ~w46516;
assign w46537 = ~w46518 & ~w46536;
assign w46538 = (~w46064 & ~w46045) | (~w46064 & w66625) | (~w46045 & w66625);
assign w46539 = ~w46534 & w46538;
assign w46540 = ~w46535 & w46539;
assign w46541 = ~w46537 & w46540;
assign w46542 = ~w46531 & ~w46541;
assign w46543 = ~w46542 & w66626;
assign w46544 = (pi2471 & w46542) | (pi2471 & w66627) | (w46542 & w66627);
assign w46545 = ~w46543 & ~w46544;
assign w46546 = ~pi5343 & pi9040;
assign w46547 = ~pi5042 & ~pi9040;
assign w46548 = ~w46546 & ~w46547;
assign w46549 = pi2454 & ~w46548;
assign w46550 = ~pi2454 & w46548;
assign w46551 = ~w46549 & ~w46550;
assign w46552 = ~pi4976 & pi9040;
assign w46553 = ~pi5206 & ~pi9040;
assign w46554 = ~w46552 & ~w46553;
assign w46555 = pi2447 & ~w46554;
assign w46556 = ~pi2447 & w46554;
assign w46557 = ~w46555 & ~w46556;
assign w46558 = ~pi5082 & pi9040;
assign w46559 = ~pi5056 & ~pi9040;
assign w46560 = ~w46558 & ~w46559;
assign w46561 = pi2457 & ~w46560;
assign w46562 = ~pi2457 & w46560;
assign w46563 = ~w46561 & ~w46562;
assign w46564 = w46557 & w46563;
assign w46565 = ~pi5180 & pi9040;
assign w46566 = ~pi5178 & ~pi9040;
assign w46567 = ~w46565 & ~w46566;
assign w46568 = pi2437 & ~w46567;
assign w46569 = ~pi2437 & w46567;
assign w46570 = ~w46568 & ~w46569;
assign w46571 = ~pi5088 & pi9040;
assign w46572 = ~pi5108 & ~pi9040;
assign w46573 = ~w46571 & ~w46572;
assign w46574 = pi2435 & ~w46573;
assign w46575 = ~pi2435 & w46573;
assign w46576 = ~w46574 & ~w46575;
assign w46577 = w46570 & ~w46576;
assign w46578 = w46564 & w46577;
assign w46579 = w46563 & ~w46570;
assign w46580 = ~w46557 & ~w46576;
assign w46581 = w46579 & w46580;
assign w46582 = ~w46578 & ~w46581;
assign w46583 = ~w46557 & w46576;
assign w46584 = ~w46570 & w46583;
assign w46585 = ~w46570 & ~w46576;
assign w46586 = ~w46563 & w46585;
assign w46587 = (~w46570 & ~w46585) | (~w46570 & w46579) | (~w46585 & w46579);
assign w46588 = w46557 & ~w46587;
assign w46589 = ~w46584 & ~w46588;
assign w46590 = ~pi5096 & pi9040;
assign w46591 = ~pi5088 & ~pi9040;
assign w46592 = ~w46590 & ~w46591;
assign w46593 = pi2434 & ~w46592;
assign w46594 = ~pi2434 & w46592;
assign w46595 = ~w46593 & ~w46594;
assign w46596 = ~w46589 & ~w46595;
assign w46597 = w46583 & w46579;
assign w46598 = w46582 & ~w46597;
assign w46599 = ~w46596 & w46598;
assign w46600 = ~w46551 & ~w46599;
assign w46601 = w46557 & w46576;
assign w46602 = ~w46570 & w46601;
assign w46603 = w46601 & w46579;
assign w46604 = w46570 & w46583;
assign w46605 = ~w46563 & w46580;
assign w46606 = ~w46604 & ~w46605;
assign w46607 = w46551 & ~w46606;
assign w46608 = w46582 & ~w46607;
assign w46609 = ~w46595 & ~w46603;
assign w46610 = w46608 & w46609;
assign w46611 = w46551 & ~w46583;
assign w46612 = (w46608 & w64031) | (w46608 & w64032) | (w64031 & w64032);
assign w46613 = w46595 & ~w46597;
assign w46614 = ~w46612 & w46613;
assign w46615 = ~w46610 & ~w46614;
assign w46616 = ~w46615 & w66628;
assign w46617 = (~pi2470 & w46615) | (~pi2470 & w66629) | (w46615 & w66629);
assign w46618 = ~w46616 & ~w46617;
assign w46619 = ~pi5179 & pi9040;
assign w46620 = ~pi5091 & ~pi9040;
assign w46621 = ~w46619 & ~w46620;
assign w46622 = pi2448 & ~w46621;
assign w46623 = ~pi2448 & w46621;
assign w46624 = ~w46622 & ~w46623;
assign w46625 = ~pi5042 & pi9040;
assign w46626 = ~pi5047 & ~pi9040;
assign w46627 = ~w46625 & ~w46626;
assign w46628 = pi2434 & ~w46627;
assign w46629 = ~pi2434 & w46627;
assign w46630 = ~w46628 & ~w46629;
assign w46631 = w46624 & ~w46630;
assign w46632 = ~pi5047 & pi9040;
assign w46633 = ~pi5048 & ~pi9040;
assign w46634 = ~w46632 & ~w46633;
assign w46635 = pi2421 & ~w46634;
assign w46636 = ~pi2421 & w46634;
assign w46637 = ~w46635 & ~w46636;
assign w46638 = w46631 & ~w46637;
assign w46639 = ~w46624 & ~w46630;
assign w46640 = w46637 & w46639;
assign w46641 = ~w46638 & ~w46640;
assign w46642 = ~pi5103 & pi9040;
assign w46643 = ~pi5179 & ~pi9040;
assign w46644 = ~w46642 & ~w46643;
assign w46645 = pi2435 & ~w46644;
assign w46646 = ~pi2435 & w46644;
assign w46647 = ~w46645 & ~w46646;
assign w46648 = ~w46637 & ~w46647;
assign w46649 = ~w46624 & w46630;
assign w46650 = w46648 & w46649;
assign w46651 = w46641 & ~w46650;
assign w46652 = ~w46630 & ~w46647;
assign w46653 = ~pi5056 & pi9040;
assign w46654 = ~pi5096 & ~pi9040;
assign w46655 = ~w46653 & ~w46654;
assign w46656 = pi2430 & ~w46655;
assign w46657 = ~pi2430 & w46655;
assign w46658 = ~w46656 & ~w46657;
assign w46659 = ~w46652 & w46658;
assign w46660 = ~w46639 & w46659;
assign w46661 = ~w46651 & w46660;
assign w46662 = ~w46631 & ~w46649;
assign w46663 = w46648 & w46662;
assign w46664 = w46631 & w46637;
assign w46665 = ~w46624 & w46647;
assign w46666 = w46630 & w46665;
assign w46667 = ~w46664 & ~w46666;
assign w46668 = ~w46663 & w46667;
assign w46669 = ~pi5339 & pi9040;
assign w46670 = ~pi5082 & ~pi9040;
assign w46671 = ~w46669 & ~w46670;
assign w46672 = pi2453 & ~w46671;
assign w46673 = ~pi2453 & w46671;
assign w46674 = ~w46672 & ~w46673;
assign w46675 = ~w46668 & ~w46674;
assign w46676 = w46637 & w46647;
assign w46677 = ~w46648 & ~w46676;
assign w46678 = ~w46631 & w46677;
assign w46679 = w46641 & ~w46678;
assign w46680 = ~w46674 & ~w46679;
assign w46681 = ~w46662 & w46677;
assign w46682 = ~w46649 & ~w46681;
assign w46683 = w46668 & w46682;
assign w46684 = ~w46680 & w46683;
assign w46685 = (~w46658 & w46684) | (~w46658 & w66630) | (w46684 & w66630);
assign w46686 = w46639 & w46659;
assign w46687 = w46624 & ~w46658;
assign w46688 = w46630 & w46637;
assign w46689 = ~w46647 & w46688;
assign w46690 = ~w46687 & w46689;
assign w46691 = ~w46641 & w46658;
assign w46692 = (~w46674 & ~w46659) | (~w46674 & w66631) | (~w46659 & w66631);
assign w46693 = ~w46690 & w46692;
assign w46694 = ~w46691 & w46693;
assign w46695 = w46658 & w46679;
assign w46696 = ~w46650 & w46674;
assign w46697 = (w46696 & ~w46679) | (w46696 & w66632) | (~w46679 & w66632);
assign w46698 = ~w46694 & ~w46697;
assign w46699 = ~w46661 & ~w46698;
assign w46700 = ~w46685 & w46699;
assign w46701 = pi2490 & ~w46700;
assign w46702 = ~pi2490 & w46700;
assign w46703 = ~w46701 & ~w46702;
assign w46704 = w46148 & w46271;
assign w46705 = w46156 & ~w46293;
assign w46706 = ~w46115 & ~w46130;
assign w46707 = ~w46150 & w46706;
assign w46708 = ~w46163 & ~w46707;
assign w46709 = w46122 & w46708;
assign w46710 = ~w46705 & ~w46709;
assign w46711 = w46122 & ~w46168;
assign w46712 = w46113 & w46163;
assign w46713 = w46407 & ~w46712;
assign w46714 = ~w46711 & ~w46713;
assign w46715 = w46144 & ~w46704;
assign w46716 = ~w46714 & w46715;
assign w46717 = ~w46710 & w46716;
assign w46718 = ~w46133 & w46705;
assign w46719 = ~w46165 & ~w46277;
assign w46720 = w46708 & ~w46719;
assign w46721 = ~w46134 & ~w46144;
assign w46722 = ~w46720 & w46721;
assign w46723 = ~w46718 & w46722;
assign w46724 = ~w46717 & ~w46723;
assign w46725 = ~pi2467 & w46724;
assign w46726 = pi2467 & ~w46724;
assign w46727 = ~w46725 & ~w46726;
assign w46728 = w46231 & w46455;
assign w46729 = w46244 & w46447;
assign w46730 = w46202 & w46216;
assign w46731 = w46429 & w46730;
assign w46732 = w46190 & ~w46729;
assign w46733 = ~w46260 & w46732;
assign w46734 = ~w46434 & ~w46731;
assign w46735 = w46733 & w46734;
assign w46736 = ~w46728 & w46735;
assign w46737 = ~w46209 & w46222;
assign w46738 = ~w46452 & ~w46737;
assign w46739 = w46230 & ~w46738;
assign w46740 = ~w46234 & ~w46739;
assign w46741 = ~w46438 & w46451;
assign w46742 = w46740 & w46741;
assign w46743 = ~w46736 & ~w46742;
assign w46744 = ~w46449 & ~w46731;
assign w46745 = ~w46209 & ~w46744;
assign w46746 = ~w46433 & ~w46453;
assign w46747 = ~w46745 & w46746;
assign w46748 = ~w46743 & w46747;
assign w46749 = ~pi2480 & w46748;
assign w46750 = pi2480 & ~w46748;
assign w46751 = ~w46749 & ~w46750;
assign w46752 = ~pi5109 & pi9040;
assign w46753 = ~pi4976 & ~pi9040;
assign w46754 = ~w46752 & ~w46753;
assign w46755 = pi2458 & ~w46754;
assign w46756 = ~pi2458 & w46754;
assign w46757 = ~w46755 & ~w46756;
assign w46758 = ~pi5178 & pi9040;
assign w46759 = ~pi5343 & ~pi9040;
assign w46760 = ~w46758 & ~w46759;
assign w46761 = pi2433 & ~w46760;
assign w46762 = ~pi2433 & w46760;
assign w46763 = ~w46761 & ~w46762;
assign w46764 = ~w46757 & w46763;
assign w46765 = ~pi4971 & pi9040;
assign w46766 = ~pi5447 & ~pi9040;
assign w46767 = ~w46765 & ~w46766;
assign w46768 = pi2437 & ~w46767;
assign w46769 = ~pi2437 & w46767;
assign w46770 = ~w46768 & ~w46769;
assign w46771 = w46757 & w46770;
assign w46772 = ~pi5105 & pi9040;
assign w46773 = ~pi5180 & ~pi9040;
assign w46774 = ~w46772 & ~w46773;
assign w46775 = pi2428 & ~w46774;
assign w46776 = ~pi2428 & w46774;
assign w46777 = ~w46775 & ~w46776;
assign w46778 = ~w46771 & ~w46777;
assign w46779 = ~pi5542 & pi9040;
assign w46780 = ~pi5110 & ~pi9040;
assign w46781 = ~w46779 & ~w46780;
assign w46782 = pi2444 & ~w46781;
assign w46783 = ~pi2444 & w46781;
assign w46784 = ~w46782 & ~w46783;
assign w46785 = w46770 & w46784;
assign w46786 = w46763 & ~w46770;
assign w46787 = ~w46763 & w46770;
assign w46788 = ~w46786 & ~w46787;
assign w46789 = w46757 & w46788;
assign w46790 = (~w46785 & ~w46788) | (~w46785 & w66633) | (~w46788 & w66633);
assign w46791 = w46778 & ~w46790;
assign w46792 = ~w46770 & ~w46777;
assign w46793 = ~w46757 & ~w46792;
assign w46794 = (~w46763 & w46793) | (~w46763 & w66634) | (w46793 & w66634);
assign w46795 = w46763 & ~w46784;
assign w46796 = w46757 & w46795;
assign w46797 = ~w46757 & w46777;
assign w46798 = ~w46770 & w46784;
assign w46799 = w46797 & w46798;
assign w46800 = ~w46796 & ~w46799;
assign w46801 = ~w46794 & w46800;
assign w46802 = ~w46791 & w46801;
assign w46803 = w46764 & ~w46802;
assign w46804 = ~pi5048 & pi9040;
assign w46805 = ~pi5209 & ~pi9040;
assign w46806 = ~w46804 & ~w46805;
assign w46807 = pi2447 & ~w46806;
assign w46808 = ~pi2447 & w46806;
assign w46809 = ~w46807 & ~w46808;
assign w46810 = w46763 & w46770;
assign w46811 = w46777 & w46810;
assign w46812 = w46809 & ~w46811;
assign w46813 = w46757 & ~w46777;
assign w46814 = w46786 & w46813;
assign w46815 = ~w46764 & ~w46797;
assign w46816 = w46770 & w46813;
assign w46817 = w46813 & w46787;
assign w46818 = w46815 & ~w46817;
assign w46819 = w46784 & ~w46818;
assign w46820 = ~w46784 & ~w46813;
assign w46821 = w46815 & w46820;
assign w46822 = w46812 & ~w46814;
assign w46823 = ~w46821 & w46822;
assign w46824 = ~w46819 & w46823;
assign w46825 = w46763 & ~w46792;
assign w46826 = ~w46757 & ~w46770;
assign w46827 = ~w46771 & ~w46826;
assign w46828 = ~w46784 & ~w46825;
assign w46829 = ~w46827 & w46828;
assign w46830 = ~w46788 & w46827;
assign w46831 = w46777 & w46830;
assign w46832 = w46784 & w46789;
assign w46833 = ~w46809 & ~w46829;
assign w46834 = ~w46831 & ~w46832;
assign w46835 = w46833 & w46834;
assign w46836 = ~w46824 & ~w46835;
assign w46837 = ~w46803 & ~w46836;
assign w46838 = ~pi2501 & w46837;
assign w46839 = pi2501 & ~w46837;
assign w46840 = ~w46838 & ~w46839;
assign w46841 = w46372 & ~w46380;
assign w46842 = ~w46473 & ~w46500;
assign w46843 = w46841 & ~w46842;
assign w46844 = w46337 & ~w46394;
assign w46845 = ~w46471 & w46844;
assign w46846 = ~w46376 & w46845;
assign w46847 = ~w46843 & w46846;
assign w46848 = w46362 & ~w46379;
assign w46849 = ~w46322 & ~w46363;
assign w46850 = ~w46472 & w46849;
assign w46851 = ~w46353 & w46850;
assign w46852 = ~w46841 & ~w46851;
assign w46853 = ~w46337 & ~w46848;
assign w46854 = ~w46852 & w46853;
assign w46855 = ~w46847 & ~w46854;
assign w46856 = w46330 & w46344;
assign w46857 = ~w46344 & ~w46356;
assign w46858 = w46316 & w46379;
assign w46859 = ~w46857 & ~w46858;
assign w46860 = ~w46322 & ~w46859;
assign w46861 = ~w46370 & ~w46856;
assign w46862 = ~w46860 & w46861;
assign w46863 = ~w46855 & w46862;
assign w46864 = pi2509 & ~w46863;
assign w46865 = ~pi2509 & w46863;
assign w46866 = ~w46864 & ~w46865;
assign w46867 = ~w46665 & ~w46688;
assign w46868 = ~w46658 & ~w46867;
assign w46869 = (w46674 & ~w46649) | (w46674 & w66635) | (~w46649 & w66635);
assign w46870 = w46868 & w46869;
assign w46871 = ~w46647 & w46675;
assign w46872 = w46637 & w46665;
assign w46873 = ~w46658 & w46872;
assign w46874 = w46630 & ~w46665;
assign w46875 = w46674 & w46676;
assign w46876 = ~w46874 & w46875;
assign w46877 = ~w46652 & ~w46658;
assign w46878 = w46867 & ~w46877;
assign w46879 = ~w46674 & ~w46872;
assign w46880 = ~w46868 & w46879;
assign w46881 = ~w46878 & w46880;
assign w46882 = w46624 & w46690;
assign w46883 = w46658 & w46674;
assign w46884 = ~w46651 & w46883;
assign w46885 = ~w46873 & ~w46876;
assign w46886 = ~w46870 & w46885;
assign w46887 = ~w46882 & w46886;
assign w46888 = ~w46881 & ~w46884;
assign w46889 = w46887 & w46888;
assign w46890 = ~w46871 & w46889;
assign w46891 = pi2492 & ~w46890;
assign w46892 = ~pi2492 & w46890;
assign w46893 = ~w46891 & ~w46892;
assign w46894 = ~w46563 & w46570;
assign w46895 = w46580 & ~w46894;
assign w46896 = ~w46603 & ~w46895;
assign w46897 = ~w46551 & ~w46896;
assign w46898 = ~w46557 & ~w46894;
assign w46899 = w46557 & w46894;
assign w46900 = w46894 & w46601;
assign w46901 = w46551 & w46570;
assign w46902 = ~w46586 & ~w46901;
assign w46903 = (~w46898 & ~w46902) | (~w46898 & w66636) | (~w46902 & w66636);
assign w46904 = ~w46897 & ~w46903;
assign w46905 = w46595 & ~w46904;
assign w46906 = ~w46563 & w46576;
assign w46907 = ~w46604 & ~w46906;
assign w46908 = w46551 & ~w46563;
assign w46909 = ~w46894 & ~w46908;
assign w46910 = ~w46907 & w46909;
assign w46911 = ~w46579 & ~w46901;
assign w46912 = w46898 & w46911;
assign w46913 = w46595 & ~w46912;
assign w46914 = w46910 & ~w46913;
assign w46915 = ~w46581 & ~w46899;
assign w46916 = w46551 & ~w46915;
assign w46917 = ~w46577 & ~w46584;
assign w46918 = ~w46563 & ~w46917;
assign w46919 = ~w46551 & ~w46602;
assign w46920 = ~w46564 & ~w46584;
assign w46921 = w46919 & ~w46920;
assign w46922 = w46551 & w46603;
assign w46923 = ~w46918 & ~w46921;
assign w46924 = ~w46922 & w46923;
assign w46925 = ~w46595 & ~w46924;
assign w46926 = ~w46914 & ~w46916;
assign w46927 = ~w46905 & w46926;
assign w46928 = ~w46925 & w46927;
assign w46929 = pi2479 & w46928;
assign w46930 = ~pi2479 & ~w46928;
assign w46931 = ~w46929 & ~w46930;
assign w46932 = ~w46209 & w46437;
assign w46933 = ~w46237 & w46737;
assign w46934 = ~w46258 & w46933;
assign w46935 = w46196 & w46227;
assign w46936 = ~w46253 & w46259;
assign w46937 = w46431 & ~w46936;
assign w46938 = w46203 & ~w46216;
assign w46939 = w46431 & w66637;
assign w46940 = ~w46934 & ~w46935;
assign w46941 = ~w46432 & w46940;
assign w46942 = (~w46190 & ~w46941) | (~w46190 & w66638) | (~w46941 & w66638);
assign w46943 = w46190 & ~w46937;
assign w46944 = ~w46238 & ~w46731;
assign w46945 = w46209 & ~w46944;
assign w46946 = ~w46932 & ~w46945;
assign w46947 = ~w46943 & w46946;
assign w46948 = ~w46942 & w46947;
assign w46949 = pi2497 & w46948;
assign w46950 = ~pi2497 & ~w46948;
assign w46951 = ~w46949 & ~w46950;
assign w46952 = w46044 & ~w46052;
assign w46953 = ~w46084 & w46089;
assign w46954 = ~w46952 & ~w46953;
assign w46955 = ~w46027 & w46066;
assign w46956 = w46044 & ~w46955;
assign w46957 = ~w46083 & w46956;
assign w46958 = w46034 & ~w46067;
assign w46959 = ~w46086 & w46958;
assign w46960 = w46538 & ~w46957;
assign w46961 = ~w46959 & w46960;
assign w46962 = ~w46076 & ~w46519;
assign w46963 = ~w46021 & ~w46955;
assign w46964 = w46044 & ~w46071;
assign w46965 = ~w46963 & w46964;
assign w46966 = w46027 & w46068;
assign w46967 = ~w46044 & ~w46072;
assign w46968 = ~w46966 & w46967;
assign w46969 = ~w46053 & w46064;
assign w46970 = w46962 & w46969;
assign w46971 = ~w46965 & w46970;
assign w46972 = ~w46968 & w46971;
assign w46973 = ~w46961 & ~w46972;
assign w46974 = ~w46954 & ~w46973;
assign w46975 = ~pi2478 & w46974;
assign w46976 = pi2478 & ~w46974;
assign w46977 = ~w46975 & ~w46976;
assign w46978 = w46785 & w46797;
assign w46979 = ~w46792 & ~w46978;
assign w46980 = w46764 & ~w46979;
assign w46981 = (~w46816 & ~w46830) | (~w46816 & w66639) | (~w46830 & w66639);
assign w46982 = ~w46795 & ~w46981;
assign w46983 = ~w46796 & w46820;
assign w46984 = ~w46787 & ~w46797;
assign w46985 = w46983 & w46984;
assign w46986 = ~w46980 & ~w46985;
assign w46987 = ~w46982 & w46986;
assign w46988 = ~w46809 & ~w46987;
assign w46989 = ~w46795 & ~w46799;
assign w46990 = ~w46825 & ~w46989;
assign w46991 = ~w46802 & w46809;
assign w46992 = ~w46757 & ~w46788;
assign w46993 = ~w46789 & ~w46992;
assign w46994 = w46777 & ~w46993;
assign w46995 = ~w46784 & w46830;
assign w46996 = w46994 & w46995;
assign w46997 = w46771 & w46820;
assign w46998 = ~w46763 & w46784;
assign w46999 = (~w46998 & ~w46820) | (~w46998 & w66640) | (~w46820 & w66640);
assign w47000 = ~w46763 & ~w46813;
assign w47001 = ~w46999 & ~w47000;
assign w47002 = ~w46990 & ~w47001;
assign w47003 = ~w46996 & w47002;
assign w47004 = ~w46991 & w47003;
assign w47005 = (pi2483 & ~w47004) | (pi2483 & w66641) | (~w47004 & w66641);
assign w47006 = w47004 & w66642;
assign w47007 = ~w47005 & ~w47006;
assign w47008 = w46770 & w46998;
assign w47009 = ~w46771 & ~w46784;
assign w47010 = ~w46816 & ~w47009;
assign w47011 = w46788 & ~w47010;
assign w47012 = w46764 & w46798;
assign w47013 = ~w47008 & ~w47012;
assign w47014 = ~w47011 & w47013;
assign w47015 = w46778 & ~w46992;
assign w47016 = w47014 & w47015;
assign w47017 = (w46809 & w47016) | (w46809 & w66643) | (w47016 & w66643);
assign w47018 = ~w46796 & ~w46811;
assign w47019 = w46777 & w47018;
assign w47020 = w46993 & w47019;
assign w47021 = w47014 & ~w47020;
assign w47022 = ~w46796 & w46812;
assign w47023 = ~w47021 & ~w47022;
assign w47024 = ~w47017 & ~w47023;
assign w47025 = ~pi2494 & w47024;
assign w47026 = pi2494 & ~w47024;
assign w47027 = ~w47025 & ~w47026;
assign w47028 = w46624 & ~w46647;
assign w47029 = w46667 & ~w47028;
assign w47030 = w46639 & ~w46676;
assign w47031 = w46674 & ~w47030;
assign w47032 = ~w46660 & w47031;
assign w47033 = w47029 & w47032;
assign w47034 = w46883 & ~w47029;
assign w47035 = w46652 & w46695;
assign w47036 = ~w46630 & w46687;
assign w47037 = ~w46666 & ~w46677;
assign w47038 = ~w47036 & w47037;
assign w47039 = ~w46681 & ~w47038;
assign w47040 = (~w46650 & w46651) | (~w46650 & w66644) | (w46651 & w66644);
assign w47041 = ~w47039 & w47040;
assign w47042 = ~w46674 & ~w47041;
assign w47043 = ~w46882 & ~w47033;
assign w47044 = ~w47034 & w47043;
assign w47045 = ~w47035 & w47044;
assign w47046 = (pi2485 & ~w47045) | (pi2485 & w66645) | (~w47045 & w66645);
assign w47047 = w47045 & w66646;
assign w47048 = ~w47046 & ~w47047;
assign w47049 = ~w46691 & ~w46695;
assign w47050 = w47039 & ~w47049;
assign w47051 = ~w46640 & ~w46689;
assign w47052 = (~w46883 & ~w47051) | (~w46883 & w66647) | (~w47051 & w66647);
assign w47053 = w46631 & ~w46677;
assign w47054 = w46874 & ~w47028;
assign w47055 = ~w46686 & ~w47054;
assign w47056 = ~w46637 & ~w47055;
assign w47057 = ~w47052 & ~w47053;
assign w47058 = ~w47056 & w47057;
assign w47059 = w46660 & ~w47054;
assign w47060 = ~w46637 & w46639;
assign w47061 = ~w47036 & ~w47060;
assign w47062 = ~w46868 & w47061;
assign w47063 = ~w46647 & ~w47062;
assign w47064 = ~w46658 & ~w47028;
assign w47065 = ~w46640 & w47064;
assign w47066 = w46662 & w47065;
assign w47067 = ~w46674 & ~w47059;
assign w47068 = ~w47066 & w47067;
assign w47069 = ~w47063 & w47068;
assign w47070 = ~w47058 & ~w47069;
assign w47071 = ~w47070 & w66648;
assign w47072 = (pi2503 & w47070) | (pi2503 & w66649) | (w47070 & w66649);
assign w47073 = ~w47071 & ~w47072;
assign w47074 = ~w46055 & w46963;
assign w47075 = ~w46064 & ~w47074;
assign w47076 = w46051 & w46064;
assign w47077 = w46962 & ~w47076;
assign w47078 = ~w46020 & ~w47077;
assign w47079 = ~w47075 & ~w47078;
assign w47080 = w46044 & ~w47079;
assign w47081 = ~w46014 & w46020;
assign w47082 = ~w46045 & ~w47081;
assign w47083 = w46034 & ~w47082;
assign w47084 = w46014 & w46049;
assign w47085 = ~w47083 & ~w47084;
assign w47086 = w46064 & ~w47085;
assign w47087 = ~w46064 & w47081;
assign w47088 = ~w46525 & w47087;
assign w47089 = ~w46048 & ~w46066;
assign w47090 = ~w46044 & ~w47089;
assign w47091 = w47074 & w47090;
assign w47092 = ~w47088 & ~w47091;
assign w47093 = ~w47086 & w47092;
assign w47094 = ~w47080 & w47093;
assign w47095 = pi2484 & ~w47094;
assign w47096 = ~pi2484 & w47094;
assign w47097 = ~w47095 & ~w47096;
assign w47098 = (~w47012 & ~w46830) | (~w47012 & w66650) | (~w46830 & w66650);
assign w47099 = ~w46777 & ~w47098;
assign w47100 = ~w46786 & ~w46979;
assign w47101 = ~w46997 & ~w47012;
assign w47102 = w47018 & w47101;
assign w47103 = (~w46809 & ~w47102) | (~w46809 & w66651) | (~w47102 & w66651);
assign w47104 = ~w46819 & w46993;
assign w47105 = ~w46982 & w47104;
assign w47106 = ~w46983 & ~w46993;
assign w47107 = w46809 & ~w47106;
assign w47108 = ~w47105 & w47107;
assign w47109 = ~w47001 & ~w47099;
assign w47110 = ~w47103 & w47109;
assign w47111 = ~w47108 & w47110;
assign w47112 = pi2488 & ~w47111;
assign w47113 = ~pi2488 & w47111;
assign w47114 = ~w47112 & ~w47113;
assign w47115 = w46583 & ~w46909;
assign w47116 = ~w46578 & ~w46900;
assign w47117 = w46611 & w47116;
assign w47118 = w46557 & w46586;
assign w47119 = ~w46557 & w46577;
assign w47120 = ~w46597 & ~w47119;
assign w47121 = ~w47118 & w47120;
assign w47122 = w47117 & w47121;
assign w47123 = ~w46595 & ~w47115;
assign w47124 = ~w47122 & w47123;
assign w47125 = w46595 & w47116;
assign w47126 = w46570 & w46605;
assign w47127 = ~w46611 & ~w46908;
assign w47128 = ~w46586 & ~w47127;
assign w47129 = ~w46576 & w46579;
assign w47130 = w46919 & ~w47129;
assign w47131 = ~w47128 & ~w47130;
assign w47132 = ~w46910 & ~w47126;
assign w47133 = w47125 & w47132;
assign w47134 = ~w47131 & w47133;
assign w47135 = w47116 & w47121;
assign w47136 = ~w46551 & ~w47125;
assign w47137 = ~w47135 & w47136;
assign w47138 = (~w47137 & w47134) | (~w47137 & w66652) | (w47134 & w66652);
assign w47139 = ~pi2486 & w47138;
assign w47140 = pi2486 & ~w47138;
assign w47141 = ~w47139 & ~w47140;
assign w47142 = ~w46551 & w46604;
assign w47143 = w46601 & ~w46911;
assign w47144 = ~w46578 & ~w46586;
assign w47145 = ~w46912 & w47144;
assign w47146 = ~w47143 & w47145;
assign w47147 = ~w46595 & ~w47146;
assign w47148 = ~w47126 & ~w47143;
assign w47149 = w47117 & ~w47148;
assign w47150 = w46551 & ~w46917;
assign w47151 = ~w46585 & ~w46906;
assign w47152 = ~w46551 & w46557;
assign w47153 = ~w47151 & w47152;
assign w47154 = ~w46581 & ~w47153;
assign w47155 = ~w47150 & w47154;
assign w47156 = w46595 & ~w47155;
assign w47157 = ~w47142 & ~w47147;
assign w47158 = ~w47149 & ~w47156;
assign w47159 = w47157 & w47158;
assign w47160 = pi2500 & ~w47159;
assign w47161 = ~pi2500 & w47159;
assign w47162 = ~w47160 & ~w47161;
assign w47163 = ~pi5506 & pi9040;
assign w47164 = ~pi5215 & ~pi9040;
assign w47165 = ~w47163 & ~w47164;
assign w47166 = pi2482 & ~w47165;
assign w47167 = ~pi2482 & w47165;
assign w47168 = ~w47166 & ~w47167;
assign w47169 = ~pi5284 & pi9040;
assign w47170 = ~pi5430 & ~pi9040;
assign w47171 = ~w47169 & ~w47170;
assign w47172 = pi2524 & ~w47171;
assign w47173 = ~pi2524 & w47171;
assign w47174 = ~w47172 & ~w47173;
assign w47175 = w47168 & w47174;
assign w47176 = ~pi5289 & pi9040;
assign w47177 = ~pi5340 & ~pi9040;
assign w47178 = ~w47176 & ~w47177;
assign w47179 = pi2521 & ~w47178;
assign w47180 = ~pi2521 & w47178;
assign w47181 = ~w47179 & ~w47180;
assign w47182 = ~pi5738 & pi9040;
assign w47183 = ~pi5456 & ~pi9040;
assign w47184 = ~w47182 & ~w47183;
assign w47185 = pi2507 & ~w47184;
assign w47186 = ~pi2507 & w47184;
assign w47187 = ~w47185 & ~w47186;
assign w47188 = w47181 & ~w47187;
assign w47189 = w47175 & w47188;
assign w47190 = ~pi5205 & pi9040;
assign w47191 = ~pi5294 & ~pi9040;
assign w47192 = ~w47190 & ~w47191;
assign w47193 = pi2525 & ~w47192;
assign w47194 = ~pi2525 & w47192;
assign w47195 = ~w47193 & ~w47194;
assign w47196 = ~pi5286 & pi9040;
assign w47197 = ~pi5738 & ~pi9040;
assign w47198 = ~w47196 & ~w47197;
assign w47199 = pi2514 & ~w47198;
assign w47200 = ~pi2514 & w47198;
assign w47201 = ~w47199 & ~w47200;
assign w47202 = ~w47181 & w47201;
assign w47203 = ~w47168 & w47174;
assign w47204 = ~w47181 & ~w47187;
assign w47205 = w47181 & w47187;
assign w47206 = ~w47204 & ~w47205;
assign w47207 = w47203 & ~w47206;
assign w47208 = ~w47168 & ~w47174;
assign w47209 = ~w47175 & w47201;
assign w47210 = ~w47208 & w47209;
assign w47211 = ~w47207 & ~w47210;
assign w47212 = ~w47202 & ~w47211;
assign w47213 = w47187 & ~w47201;
assign w47214 = ~w47202 & ~w47213;
assign w47215 = w47208 & ~w47214;
assign w47216 = ~w47189 & w47195;
assign w47217 = ~w47215 & w47216;
assign w47218 = ~w47212 & w47217;
assign w47219 = w47174 & ~w47181;
assign w47220 = ~w47174 & w47187;
assign w47221 = ~w47219 & ~w47220;
assign w47222 = w47210 & ~w47221;
assign w47223 = w47201 & ~w47203;
assign w47224 = w47205 & w47223;
assign w47225 = ~w47201 & ~w47219;
assign w47226 = w47168 & ~w47201;
assign w47227 = (~w47187 & ~w47226) | (~w47187 & w66653) | (~w47226 & w66653);
assign w47228 = w47225 & w47227;
assign w47229 = ~w47181 & w47226;
assign w47230 = ~w47195 & ~w47229;
assign w47231 = ~w47224 & w47230;
assign w47232 = ~w47222 & w47231;
assign w47233 = ~w47228 & w47232;
assign w47234 = ~w47218 & ~w47233;
assign w47235 = w47174 & ~w47201;
assign w47236 = ~w47187 & ~w47235;
assign w47237 = w47209 & w66654;
assign w47238 = ~w47201 & w47208;
assign w47239 = ~w47181 & w47238;
assign w47240 = ~w47174 & w47181;
assign w47241 = w47226 & w47240;
assign w47242 = ~w47239 & ~w47241;
assign w47243 = ~w47237 & w47242;
assign w47244 = ~w47181 & w47236;
assign w47245 = w47243 & w47244;
assign w47246 = ~w47168 & w47201;
assign w47247 = ~w47226 & ~w47246;
assign w47248 = w47187 & w47219;
assign w47249 = ~w47247 & w47248;
assign w47250 = ~w47245 & ~w47249;
assign w47251 = ~w47234 & w47250;
assign w47252 = pi2536 & ~w47251;
assign w47253 = ~pi2536 & w47251;
assign w47254 = ~w47252 & ~w47253;
assign w47255 = w47220 & w47237;
assign w47256 = ~w47219 & ~w47226;
assign w47257 = w47175 & ~w47225;
assign w47258 = w47187 & ~w47257;
assign w47259 = ~w47256 & w47258;
assign w47260 = w47168 & ~w47181;
assign w47261 = w47174 & ~w47187;
assign w47262 = ~w47201 & ~w47261;
assign w47263 = w47260 & ~w47262;
assign w47264 = ~w47205 & w47238;
assign w47265 = w47240 & w47246;
assign w47266 = ~w47195 & ~w47265;
assign w47267 = ~w47263 & ~w47264;
assign w47268 = w47266 & w47267;
assign w47269 = ~w47259 & w47268;
assign w47270 = ~w47220 & ~w47261;
assign w47271 = ~w47188 & w47246;
assign w47272 = ~w47270 & ~w47271;
assign w47273 = w47168 & w47240;
assign w47274 = ~w47229 & w47270;
assign w47275 = ~w47273 & w47274;
assign w47276 = ~w47272 & ~w47275;
assign w47277 = w47174 & w47181;
assign w47278 = w47247 & w47277;
assign w47279 = w47195 & ~w47278;
assign w47280 = ~w47276 & w47279;
assign w47281 = ~w47269 & ~w47280;
assign w47282 = ~w47239 & ~w47278;
assign w47283 = ~w47187 & ~w47282;
assign w47284 = w47205 & w47246;
assign w47285 = ~w47255 & ~w47284;
assign w47286 = ~w47283 & w47285;
assign w47287 = ~w47281 & w47286;
assign w47288 = pi2538 & ~w47287;
assign w47289 = ~pi2538 & w47287;
assign w47290 = ~w47288 & ~w47289;
assign w47291 = ~pi5341 & pi9040;
assign w47292 = ~pi5284 & ~pi9040;
assign w47293 = ~w47291 & ~w47292;
assign w47294 = pi2522 & ~w47293;
assign w47295 = ~pi2522 & w47293;
assign w47296 = ~w47294 & ~w47295;
assign w47297 = ~pi5630 & pi9040;
assign w47298 = ~pi5422 & ~pi9040;
assign w47299 = ~w47297 & ~w47298;
assign w47300 = pi2527 & ~w47299;
assign w47301 = ~pi2527 & w47299;
assign w47302 = ~w47300 & ~w47301;
assign w47303 = w47296 & w47302;
assign w47304 = ~pi5545 & pi9040;
assign w47305 = ~pi5289 & ~pi9040;
assign w47306 = ~w47304 & ~w47305;
assign w47307 = pi2493 & ~w47306;
assign w47308 = ~pi2493 & w47306;
assign w47309 = ~w47307 & ~w47308;
assign w47310 = ~pi5456 & pi9040;
assign w47311 = ~pi5461 & ~pi9040;
assign w47312 = ~w47310 & ~w47311;
assign w47313 = pi2469 & ~w47312;
assign w47314 = ~pi2469 & w47312;
assign w47315 = ~w47313 & ~w47314;
assign w47316 = w47309 & w47315;
assign w47317 = ~w47309 & ~w47315;
assign w47318 = ~w47316 & ~w47317;
assign w47319 = ~pi5292 & pi9040;
assign w47320 = ~pi5630 & ~pi9040;
assign w47321 = ~w47319 & ~w47320;
assign w47322 = pi2506 & ~w47321;
assign w47323 = ~pi2506 & w47321;
assign w47324 = ~w47322 & ~w47323;
assign w47325 = w47318 & w47324;
assign w47326 = w47318 & w66655;
assign w47327 = w47302 & ~w47324;
assign w47328 = ~w47296 & ~w47324;
assign w47329 = ~w47327 & ~w47328;
assign w47330 = w47316 & ~w47329;
assign w47331 = ~w47326 & ~w47330;
assign w47332 = ~pi5215 & pi9040;
assign w47333 = ~pi5545 & ~pi9040;
assign w47334 = ~w47332 & ~w47333;
assign w47335 = pi2517 & ~w47334;
assign w47336 = ~pi2517 & w47334;
assign w47337 = ~w47335 & ~w47336;
assign w47338 = ~w47296 & ~w47315;
assign w47339 = w47324 & ~w47338;
assign w47340 = ~w47302 & w47309;
assign w47341 = ~w47296 & ~w47340;
assign w47342 = ~w47296 & ~w47318;
assign w47343 = ~w47318 & w64034;
assign w47344 = (~w47315 & w47318) | (~w47315 & w66656) | (w47318 & w66656);
assign w47345 = w47341 & ~w47344;
assign w47346 = w47309 & ~w47324;
assign w47347 = ~w47302 & ~w47346;
assign w47348 = ~w47339 & w47347;
assign w47349 = ~w47345 & w47348;
assign w47350 = w47296 & ~w47324;
assign w47351 = ~w47315 & w47350;
assign w47352 = w47350 & w47317;
assign w47353 = ~w47337 & ~w47352;
assign w47354 = w47331 & w47353;
assign w47355 = ~w47349 & w47354;
assign w47356 = w47296 & w47340;
assign w47357 = w47337 & ~w47356;
assign w47358 = w47302 & ~w47309;
assign w47359 = ~w47315 & w47324;
assign w47360 = w47358 & w47359;
assign w47361 = ~w47338 & ~w47358;
assign w47362 = ~w47317 & ~w47324;
assign w47363 = ~w47361 & w47362;
assign w47364 = ~w47360 & ~w47363;
assign w47365 = w47357 & w47364;
assign w47366 = ~w47345 & w47365;
assign w47367 = ~w47355 & ~w47366;
assign w47368 = ~w47296 & w47360;
assign w47369 = w47296 & w47318;
assign w47370 = ~w47342 & ~w47369;
assign w47371 = (~w47351 & ~w47370) | (~w47351 & w66657) | (~w47370 & w66657);
assign w47372 = ~w47302 & ~w47371;
assign w47373 = w47302 & w47309;
assign w47374 = w47328 & w47373;
assign w47375 = ~w47368 & ~w47374;
assign w47376 = ~w47372 & w47375;
assign w47377 = ~w47367 & w47376;
assign w47378 = pi2540 & w47377;
assign w47379 = ~pi2540 & ~w47377;
assign w47380 = ~w47378 & ~w47379;
assign w47381 = ~w47243 & ~w47270;
assign w47382 = w47204 & ~w47247;
assign w47383 = w47247 & w66658;
assign w47384 = w47203 & w47213;
assign w47385 = w47188 & w47238;
assign w47386 = w47195 & ~w47384;
assign w47387 = ~w47382 & w47386;
assign w47388 = ~w47385 & w47387;
assign w47389 = ~w47222 & ~w47383;
assign w47390 = w47388 & w47389;
assign w47391 = ~w47188 & w47238;
assign w47392 = w47236 & ~w47273;
assign w47393 = ~w47258 & ~w47392;
assign w47394 = w47266 & ~w47284;
assign w47395 = ~w47391 & w47394;
assign w47396 = ~w47393 & w47395;
assign w47397 = ~w47390 & ~w47396;
assign w47398 = ~w47381 & ~w47397;
assign w47399 = ~pi2532 & w47398;
assign w47400 = pi2532 & ~w47398;
assign w47401 = ~w47399 & ~w47400;
assign w47402 = w47303 & ~w47364;
assign w47403 = (~w47302 & w47342) | (~w47302 & w66659) | (w47342 & w66659);
assign w47404 = w47296 & w47315;
assign w47405 = ~w47338 & ~w47404;
assign w47406 = w47373 & ~w47405;
assign w47407 = w47325 & w47405;
assign w47408 = ~w47406 & ~w47407;
assign w47409 = (~w47337 & ~w47408) | (~w47337 & w66660) | (~w47408 & w66660);
assign w47410 = ~w47309 & ~w47328;
assign w47411 = w47347 & ~w47410;
assign w47412 = w47316 & w47328;
assign w47413 = ~w47410 & ~w47412;
assign w47414 = w47302 & ~w47413;
assign w47415 = w47309 & w47351;
assign w47416 = w47324 & w47404;
assign w47417 = ~w47411 & ~w47416;
assign w47418 = ~w47415 & w47417;
assign w47419 = ~w47414 & w47418;
assign w47420 = w47337 & ~w47419;
assign w47421 = ~w47402 & ~w47409;
assign w47422 = ~w47420 & w47421;
assign w47423 = ~pi2553 & w47422;
assign w47424 = pi2553 & ~w47422;
assign w47425 = ~w47423 & ~w47424;
assign w47426 = ~pi5214 & pi9040;
assign w47427 = ~pi5506 & ~pi9040;
assign w47428 = ~w47426 & ~w47427;
assign w47429 = pi2517 & ~w47428;
assign w47430 = ~pi2517 & w47428;
assign w47431 = ~w47429 & ~w47430;
assign w47432 = ~pi5347 & pi9040;
assign w47433 = ~pi5338 & ~pi9040;
assign w47434 = ~w47432 & ~w47433;
assign w47435 = pi2481 & ~w47434;
assign w47436 = ~pi2481 & w47434;
assign w47437 = ~w47435 & ~w47436;
assign w47438 = ~w47431 & ~w47437;
assign w47439 = ~pi5544 & pi9040;
assign w47440 = ~pi5205 & ~pi9040;
assign w47441 = ~w47439 & ~w47440;
assign w47442 = pi2469 & ~w47441;
assign w47443 = ~pi2469 & w47441;
assign w47444 = ~w47442 & ~w47443;
assign w47445 = ~pi5287 & pi9040;
assign w47446 = ~pi5346 & ~pi9040;
assign w47447 = ~w47445 & ~w47446;
assign w47448 = pi2526 & ~w47447;
assign w47449 = ~pi2526 & w47447;
assign w47450 = ~w47448 & ~w47449;
assign w47451 = ~w47444 & w47450;
assign w47452 = ~w47437 & ~w47451;
assign w47453 = ~pi5430 & pi9040;
assign w47454 = ~pi5544 & ~pi9040;
assign w47455 = ~w47453 & ~w47454;
assign w47456 = pi2515 & ~w47455;
assign w47457 = ~pi2515 & w47455;
assign w47458 = ~w47456 & ~w47457;
assign w47459 = (~w47458 & w47451) | (~w47458 & w64036) | (w47451 & w64036);
assign w47460 = ~w47437 & w47459;
assign w47461 = ~w47431 & w47450;
assign w47462 = w47458 & w47461;
assign w47463 = w47461 & w47528;
assign w47464 = ~w47460 & ~w47463;
assign w47465 = w47438 & ~w47464;
assign w47466 = w47444 & ~w47458;
assign w47467 = w47431 & w47466;
assign w47468 = ~w47431 & ~w47451;
assign w47469 = ~w47444 & w47458;
assign w47470 = w47468 & w47469;
assign w47471 = ~w47467 & ~w47470;
assign w47472 = w47437 & ~w47471;
assign w47473 = ~pi5212 & pi9040;
assign w47474 = ~pi5347 & ~pi9040;
assign w47475 = ~w47473 & ~w47474;
assign w47476 = pi2513 & ~w47475;
assign w47477 = ~pi2513 & w47475;
assign w47478 = ~w47476 & ~w47477;
assign w47479 = w47452 & w47458;
assign w47480 = ~w47438 & ~w47479;
assign w47481 = ~w47468 & ~w47480;
assign w47482 = w47431 & w47450;
assign w47483 = w47469 & w47482;
assign w47484 = ~w47444 & ~w47461;
assign w47485 = w47444 & w47450;
assign w47486 = ~w47484 & ~w47485;
assign w47487 = ~w47484 & w66661;
assign w47488 = (~w47478 & ~w47483) | (~w47478 & w66662) | (~w47483 & w66662);
assign w47489 = ~w47487 & w47488;
assign w47490 = w47464 & w47489;
assign w47491 = ~w47481 & w47490;
assign w47492 = w47431 & ~w47450;
assign w47493 = w47450 & ~w47458;
assign w47494 = ~w47492 & ~w47493;
assign w47495 = ~w47450 & w47458;
assign w47496 = ~w47484 & ~w47495;
assign w47497 = ~w47437 & w47494;
assign w47498 = ~w47496 & w47497;
assign w47499 = ~w47431 & ~w47466;
assign w47500 = w47437 & w47444;
assign w47501 = ~w47444 & w47492;
assign w47502 = ~w47458 & w47501;
assign w47503 = ~w47500 & ~w47502;
assign w47504 = ~w47499 & ~w47503;
assign w47505 = w47466 & w47482;
assign w47506 = w47478 & ~w47505;
assign w47507 = ~w47498 & w47506;
assign w47508 = ~w47504 & w47507;
assign w47509 = ~w47491 & ~w47508;
assign w47510 = ~w47465 & ~w47472;
assign w47511 = ~w47509 & w47510;
assign w47512 = pi2552 & ~w47511;
assign w47513 = ~pi2552 & w47511;
assign w47514 = ~w47512 & ~w47513;
assign w47515 = w47468 & ~w47495;
assign w47516 = w47437 & ~w47478;
assign w47517 = w47515 & w47516;
assign w47518 = w47468 & w66663;
assign w47519 = w47431 & w47459;
assign w47520 = w47444 & ~w47492;
assign w47521 = (~w47501 & w47515) | (~w47501 & w66664) | (w47515 & w66664);
assign w47522 = w47437 & ~w47521;
assign w47523 = ~w47444 & w47462;
assign w47524 = ~w47518 & ~w47523;
assign w47525 = ~w47519 & w47524;
assign w47526 = ~w47522 & w47525;
assign w47527 = w47478 & ~w47526;
assign w47528 = w47444 & w47458;
assign w47529 = w47492 & w47528;
assign w47530 = ~w47483 & ~w47529;
assign w47531 = ~w47470 & w47530;
assign w47532 = ~w47450 & ~w47458;
assign w47533 = (~w47437 & ~w47484) | (~w47437 & w66665) | (~w47484 & w66665);
assign w47534 = ~w47468 & w47533;
assign w47535 = w47531 & ~w47534;
assign w47536 = ~w47478 & ~w47535;
assign w47537 = ~w47523 & w47531;
assign w47538 = (~w47517 & w47537) | (~w47517 & w66666) | (w47537 & w66666);
assign w47539 = ~w47536 & w47538;
assign w47540 = ~w47527 & w47539;
assign w47541 = pi2546 & ~w47540;
assign w47542 = ~pi2546 & w47540;
assign w47543 = ~w47541 & ~w47542;
assign w47544 = ~pi5298 & pi9040;
assign w47545 = ~pi5288 & ~pi9040;
assign w47546 = ~w47544 & ~w47545;
assign w47547 = pi2516 & ~w47546;
assign w47548 = ~pi2516 & w47546;
assign w47549 = ~w47547 & ~w47548;
assign w47550 = ~pi5213 & pi9040;
assign w47551 = ~pi5330 & ~pi9040;
assign w47552 = ~w47550 & ~w47551;
assign w47553 = pi2504 & ~w47552;
assign w47554 = ~pi2504 & w47552;
assign w47555 = ~w47553 & ~w47554;
assign w47556 = ~pi5736 & pi9040;
assign w47557 = ~pi5378 & ~pi9040;
assign w47558 = ~w47556 & ~w47557;
assign w47559 = pi2487 & ~w47558;
assign w47560 = ~pi2487 & w47558;
assign w47561 = ~w47559 & ~w47560;
assign w47562 = ~w47555 & w47561;
assign w47563 = ~pi5297 & pi9040;
assign w47564 = ~pi5296 & ~pi9040;
assign w47565 = ~w47563 & ~w47564;
assign w47566 = pi2472 & ~w47565;
assign w47567 = ~pi2472 & w47565;
assign w47568 = ~w47566 & ~w47567;
assign w47569 = w47562 & w47568;
assign w47570 = ~w47555 & ~w47561;
assign w47571 = ~pi5283 & pi9040;
assign w47572 = ~pi5298 & ~pi9040;
assign w47573 = ~w47571 & ~w47572;
assign w47574 = pi2520 & ~w47573;
assign w47575 = ~pi2520 & w47573;
assign w47576 = ~w47574 & ~w47575;
assign w47577 = w47568 & w47576;
assign w47578 = ~w47568 & ~w47576;
assign w47579 = ~w47577 & ~w47578;
assign w47580 = w47570 & w47579;
assign w47581 = ~pi5583 & pi9040;
assign w47582 = ~pi5213 & ~pi9040;
assign w47583 = ~w47581 & ~w47582;
assign w47584 = pi2518 & ~w47583;
assign w47585 = ~pi2518 & w47583;
assign w47586 = ~w47584 & ~w47585;
assign w47587 = w47555 & ~w47576;
assign w47588 = ~w47561 & w47587;
assign w47589 = w47561 & ~w47568;
assign w47590 = ~w47555 & ~w47576;
assign w47591 = ~w47589 & w47590;
assign w47592 = w47555 & w47576;
assign w47593 = w47561 & w47592;
assign w47594 = ~w47588 & ~w47591;
assign w47595 = ~w47593 & w47594;
assign w47596 = (w47586 & ~w47579) | (w47586 & w64037) | (~w47579 & w64037);
assign w47597 = (~w47569 & w47595) | (~w47569 & w64038) | (w47595 & w64038);
assign w47598 = w47555 & w47589;
assign w47599 = ~w47569 & ~w47598;
assign w47600 = ~w47586 & ~w47599;
assign w47601 = ~w47568 & ~w47586;
assign w47602 = w47587 & w47601;
assign w47603 = w47555 & ~w47561;
assign w47604 = w47577 & w47603;
assign w47605 = ~w47602 & ~w47604;
assign w47606 = w47555 & ~w47568;
assign w47607 = w47586 & ~w47606;
assign w47608 = w47568 & ~w47603;
assign w47609 = w47607 & ~w47608;
assign w47610 = w47576 & w47586;
assign w47611 = ~w47555 & w47610;
assign w47612 = w47561 & w47578;
assign w47613 = ~w47611 & ~w47612;
assign w47614 = ~w47562 & ~w47613;
assign w47615 = w47605 & ~w47609;
assign w47616 = ~w47600 & w47615;
assign w47617 = ~w47614 & w47616;
assign w47618 = ~w47562 & ~w47568;
assign w47619 = (~w47586 & ~w47618) | (~w47586 & w66667) | (~w47618 & w66667);
assign w47620 = w47568 & w47592;
assign w47621 = ~w47612 & ~w47620;
assign w47622 = w47599 & w47621;
assign w47623 = w47619 & w47622;
assign w47624 = (~w47623 & ~w47617) | (~w47623 & w64039) | (~w47617 & w64039);
assign w47625 = w47549 & ~w47624;
assign w47626 = w47561 & ~w47602;
assign w47627 = w47590 & w47601;
assign w47628 = w47610 & w66668;
assign w47629 = ~w47561 & ~w47628;
assign w47630 = ~w47627 & w47629;
assign w47631 = ~w47626 & ~w47630;
assign w47632 = (~w47549 & ~w47616) | (~w47549 & w66669) | (~w47616 & w66669);
assign w47633 = w47607 & ~w47621;
assign w47634 = ~w47631 & ~w47633;
assign w47635 = ~w47632 & w47634;
assign w47636 = (pi2544 & w47625) | (pi2544 & w66670) | (w47625 & w66670);
assign w47637 = ~w47625 & w66671;
assign w47638 = ~w47636 & ~w47637;
assign w47639 = ~pi5546 & pi9040;
assign w47640 = pi5204 & ~pi9040;
assign w47641 = ~w47639 & ~w47640;
assign w47642 = pi2504 & ~w47641;
assign w47643 = ~pi2504 & w47641;
assign w47644 = ~w47642 & ~w47643;
assign w47645 = ~pi5344 & pi9040;
assign w47646 = ~pi5736 & ~pi9040;
assign w47647 = ~w47645 & ~w47646;
assign w47648 = pi2487 & ~w47647;
assign w47649 = ~pi2487 & w47647;
assign w47650 = ~w47648 & ~w47649;
assign w47651 = ~pi5543 & pi9040;
assign w47652 = ~pi5429 & ~pi9040;
assign w47653 = ~w47651 & ~w47652;
assign w47654 = pi2525 & ~w47653;
assign w47655 = ~pi2525 & w47653;
assign w47656 = ~w47654 & ~w47655;
assign w47657 = ~w47650 & w47656;
assign w47658 = ~pi5203 & pi9040;
assign w47659 = ~pi5584 & ~pi9040;
assign w47660 = ~w47658 & ~w47659;
assign w47661 = pi2524 & ~w47660;
assign w47662 = ~pi2524 & w47660;
assign w47663 = ~w47661 & ~w47662;
assign w47664 = ~pi5335 & pi9040;
assign w47665 = ~pi5337 & ~pi9040;
assign w47666 = ~w47664 & ~w47665;
assign w47667 = pi2523 & ~w47666;
assign w47668 = ~pi2523 & w47666;
assign w47669 = ~w47667 & ~w47668;
assign w47670 = w47663 & ~w47669;
assign w47671 = ~w47663 & w47669;
assign w47672 = ~w47670 & ~w47671;
assign w47673 = w47657 & ~w47672;
assign w47674 = w47650 & w47656;
assign w47675 = ~pi5584 & pi9040;
assign w47676 = ~pi5345 & ~pi9040;
assign w47677 = ~w47675 & ~w47676;
assign w47678 = pi2510 & ~w47677;
assign w47679 = ~pi2510 & w47677;
assign w47680 = ~w47678 & ~w47679;
assign w47681 = w47663 & w47680;
assign w47682 = w47674 & ~w47681;
assign w47683 = w47672 & w47682;
assign w47684 = ~w47673 & ~w47683;
assign w47685 = w47656 & ~w47669;
assign w47686 = ~w47670 & ~w47674;
assign w47687 = (w47680 & w47686) | (w47680 & w66672) | (w47686 & w66672);
assign w47688 = w47656 & w47663;
assign w47689 = ~w47650 & ~w47688;
assign w47690 = w47687 & ~w47689;
assign w47691 = ~w47656 & ~w47663;
assign w47692 = ~w47650 & w47691;
assign w47693 = w47650 & w47663;
assign w47694 = ~w47656 & w47693;
assign w47695 = ~w47692 & ~w47694;
assign w47696 = ~w47669 & ~w47680;
assign w47697 = ~w47695 & w47696;
assign w47698 = w47684 & ~w47697;
assign w47699 = (~w47644 & ~w47698) | (~w47644 & w66673) | (~w47698 & w66673);
assign w47700 = ~w47688 & ~w47691;
assign w47701 = ~w47650 & w47669;
assign w47702 = ~w47700 & w47701;
assign w47703 = ~w47650 & w47663;
assign w47704 = w47656 & w47703;
assign w47705 = w47680 & ~w47704;
assign w47706 = ~w47702 & w47705;
assign w47707 = ~w47656 & w47669;
assign w47708 = w47695 & w47707;
assign w47709 = ~w47680 & ~w47708;
assign w47710 = w47681 & ~w47685;
assign w47711 = ~w47706 & ~w47710;
assign w47712 = ~w47709 & w47711;
assign w47713 = w47684 & w47695;
assign w47714 = w47709 & ~w47713;
assign w47715 = w47687 & ~w47692;
assign w47716 = w47644 & ~w47715;
assign w47717 = ~w47714 & w47716;
assign w47718 = ~w47699 & ~w47712;
assign w47719 = ~w47717 & w47718;
assign w47720 = ~pi2547 & ~w47719;
assign w47721 = pi2547 & w47719;
assign w47722 = ~w47720 & ~w47721;
assign w47723 = ~w47175 & w47195;
assign w47724 = ~w47270 & ~w47723;
assign w47725 = w47247 & ~w47724;
assign w47726 = w47220 & w47246;
assign w47727 = ~w47725 & ~w47726;
assign w47728 = w47181 & ~w47727;
assign w47729 = ~w47174 & w47260;
assign w47730 = w47227 & ~w47729;
assign w47731 = ~w47181 & w47208;
assign w47732 = w47187 & ~w47241;
assign w47733 = ~w47731 & w47732;
assign w47734 = ~w47730 & ~w47733;
assign w47735 = ~w47237 & ~w47383;
assign w47736 = (~w47195 & w47734) | (~w47195 & w66674) | (w47734 & w66674);
assign w47737 = ~w47208 & w47213;
assign w47738 = ~w47202 & ~w47246;
assign w47739 = w47730 & ~w47738;
assign w47740 = ~w47737 & ~w47739;
assign w47741 = w47195 & ~w47240;
assign w47742 = ~w47740 & w47741;
assign w47743 = ~w47728 & ~w47736;
assign w47744 = ~w47742 & w47743;
assign w47745 = pi2542 & w47744;
assign w47746 = ~pi2542 & ~w47744;
assign w47747 = ~w47745 & ~w47746;
assign w47748 = ~w47682 & ~w47686;
assign w47749 = ~w47673 & w47748;
assign w47750 = ~w47650 & w47672;
assign w47751 = w47700 & ~w47750;
assign w47752 = w47705 & ~w47751;
assign w47753 = ~w47751 & w66675;
assign w47754 = ~w47680 & ~w47688;
assign w47755 = w47650 & w47754;
assign w47756 = ~w47708 & w47755;
assign w47757 = ~w47702 & ~w47749;
assign w47758 = ~w47756 & w47757;
assign w47759 = (w47644 & ~w47758) | (w47644 & w66676) | (~w47758 & w66676);
assign w47760 = w47650 & ~w47669;
assign w47761 = ~w47701 & ~w47760;
assign w47762 = ~w47691 & w47754;
assign w47763 = w47754 & w66677;
assign w47764 = ~w47710 & ~w47763;
assign w47765 = ~w47761 & ~w47764;
assign w47766 = ~w47657 & w47671;
assign w47767 = w47715 & w47766;
assign w47768 = ~w47663 & w47674;
assign w47769 = ~w47650 & ~w47669;
assign w47770 = ~w47700 & w47769;
assign w47771 = ~w47768 & ~w47770;
assign w47772 = w47705 & ~w47771;
assign w47773 = w47656 & w47696;
assign w47774 = (~w47773 & ~w47695) | (~w47773 & w66678) | (~w47695 & w66678);
assign w47775 = (~w47644 & w47772) | (~w47644 & w66679) | (w47772 & w66679);
assign w47776 = ~w47765 & ~w47767;
assign w47777 = ~w47775 & w47776;
assign w47778 = ~w47759 & w47777;
assign w47779 = pi2541 & w47778;
assign w47780 = ~pi2541 & ~w47778;
assign w47781 = ~w47779 & ~w47780;
assign w47782 = w47346 & w47404;
assign w47783 = w47302 & ~w47350;
assign w47784 = w47405 & w47783;
assign w47785 = w47303 & w47317;
assign w47786 = ~w47782 & ~w47785;
assign w47787 = ~w47784 & w47786;
assign w47788 = w47327 & w47787;
assign w47789 = (~w47415 & ~w47370) | (~w47415 & w66680) | (~w47370 & w66680);
assign w47790 = ~w47788 & w47789;
assign w47791 = w47337 & ~w47790;
assign w47792 = w47357 & ~w47416;
assign w47793 = ~w47302 & ~w47316;
assign w47794 = ~w47405 & w47793;
assign w47795 = ~w47343 & ~w47794;
assign w47796 = w47787 & w47795;
assign w47797 = ~w47792 & ~w47796;
assign w47798 = ~w47791 & ~w47797;
assign w47799 = ~pi2549 & w47798;
assign w47800 = pi2549 & ~w47798;
assign w47801 = ~w47799 & ~w47800;
assign w47802 = ~pi5288 & pi9040;
assign w47803 = ~pi5335 & ~pi9040;
assign w47804 = ~w47802 & ~w47803;
assign w47805 = pi2499 & ~w47804;
assign w47806 = ~pi2499 & w47804;
assign w47807 = ~w47805 & ~w47806;
assign w47808 = ~pi5641 & pi9040;
assign w47809 = ~pi5344 & ~pi9040;
assign w47810 = ~w47808 & ~w47809;
assign w47811 = pi2508 & ~w47810;
assign w47812 = ~pi2508 & w47810;
assign w47813 = ~w47811 & ~w47812;
assign w47814 = ~w47807 & ~w47813;
assign w47815 = ~pi5345 & pi9040;
assign w47816 = ~pi5336 & ~pi9040;
assign w47817 = ~w47815 & ~w47816;
assign w47818 = pi2519 & ~w47817;
assign w47819 = ~pi2519 & w47817;
assign w47820 = ~w47818 & ~w47819;
assign w47821 = ~pi5204 & pi9040;
assign w47822 = ~pi5583 & ~pi9040;
assign w47823 = ~w47821 & ~w47822;
assign w47824 = pi2522 & ~w47823;
assign w47825 = ~pi2522 & w47823;
assign w47826 = ~w47824 & ~w47825;
assign w47827 = w47820 & ~w47826;
assign w47828 = ~w47820 & w47826;
assign w47829 = ~w47813 & w47828;
assign w47830 = ~w47827 & ~w47829;
assign w47831 = w47814 & w47830;
assign w47832 = ~w47807 & w47813;
assign w47833 = w47827 & w47832;
assign w47834 = w47807 & ~w47813;
assign w47835 = w47828 & w47834;
assign w47836 = ~w47833 & ~w47835;
assign w47837 = ~w47831 & w47836;
assign w47838 = ~pi5296 & pi9040;
assign w47839 = ~pi5628 & ~pi9040;
assign w47840 = ~w47838 & ~w47839;
assign w47841 = pi2512 & ~w47840;
assign w47842 = ~pi2512 & w47840;
assign w47843 = ~w47841 & ~w47842;
assign w47844 = ~w47837 & w47843;
assign w47845 = w47807 & ~w47820;
assign w47846 = ~w47826 & w47845;
assign w47847 = w47820 & w47834;
assign w47848 = w47834 & w47884;
assign w47849 = ~w47846 & ~w47848;
assign w47850 = ~w47843 & ~w47849;
assign w47851 = w47813 & w47850;
assign w47852 = w47814 & w47826;
assign w47853 = (w47843 & ~w47814) | (w47843 & w66681) | (~w47814 & w66681);
assign w47854 = w47834 & w47827;
assign w47855 = w47853 & ~w47854;
assign w47856 = ~w47807 & w47827;
assign w47857 = ~w47826 & ~w47843;
assign w47858 = ~w47813 & ~w47843;
assign w47859 = ~w47857 & ~w47858;
assign w47860 = ~w47856 & ~w47859;
assign w47861 = ~w47855 & ~w47860;
assign w47862 = ~pi5334 & pi9040;
assign w47863 = ~pi5641 & ~pi9040;
assign w47864 = ~w47862 & ~w47863;
assign w47865 = pi2493 & ~w47864;
assign w47866 = ~pi2493 & w47864;
assign w47867 = ~w47865 & ~w47866;
assign w47868 = w47813 & ~w47826;
assign w47869 = w47845 & ~w47868;
assign w47870 = ~w47845 & w47868;
assign w47871 = w47843 & ~w47870;
assign w47872 = ~w47869 & w47871;
assign w47873 = w47814 & ~w47820;
assign w47874 = ~w47847 & ~w47873;
assign w47875 = ~w47843 & w47874;
assign w47876 = ~w47872 & ~w47875;
assign w47877 = w47807 & w47813;
assign w47878 = w47807 & ~w47843;
assign w47879 = ~w47877 & ~w47878;
assign w47880 = ~w47827 & ~w47879;
assign w47881 = ~w47876 & w47880;
assign w47882 = ~w47861 & ~w47867;
assign w47883 = ~w47881 & w47882;
assign w47884 = w47820 & w47826;
assign w47885 = w47832 & w47884;
assign w47886 = w47867 & ~w47885;
assign w47887 = ~w47876 & w47886;
assign w47888 = ~w47883 & ~w47887;
assign w47889 = ~w47844 & ~w47851;
assign w47890 = ~w47888 & w66682;
assign w47891 = (~pi2535 & w47888) | (~pi2535 & w66683) | (w47888 & w66683);
assign w47892 = ~w47890 & ~w47891;
assign w47893 = w47578 & w47603;
assign w47894 = w47589 & w47610;
assign w47895 = ~w47591 & ~w47620;
assign w47896 = ~w47586 & ~w47895;
assign w47897 = (w47568 & ~w47587) | (w47568 & w66684) | (~w47587 & w66684);
assign w47898 = ~w47618 & ~w47897;
assign w47899 = w47562 & w47576;
assign w47900 = ~w47898 & ~w47899;
assign w47901 = w47586 & ~w47900;
assign w47902 = w47549 & ~w47580;
assign w47903 = w47605 & ~w47896;
assign w47904 = w47902 & w47903;
assign w47905 = ~w47901 & w47904;
assign w47906 = w47570 & w47577;
assign w47907 = w47619 & ~w47897;
assign w47908 = ~w47549 & ~w47906;
assign w47909 = (w47908 & w47595) | (w47908 & w66685) | (w47595 & w66685);
assign w47910 = ~w47907 & w47909;
assign w47911 = ~w47893 & ~w47894;
assign w47912 = (w47911 & w47905) | (w47911 & w66686) | (w47905 & w66686);
assign w47913 = pi2528 & w47912;
assign w47914 = ~pi2528 & ~w47912;
assign w47915 = ~w47913 & ~w47914;
assign w47916 = w47685 & w47693;
assign w47917 = ~w47686 & w47754;
assign w47918 = ~w47670 & ~w47688;
assign w47919 = ~w47761 & ~w47918;
assign w47920 = ~w47917 & ~w47919;
assign w47921 = (~w47644 & w47752) | (~w47644 & w66687) | (w47752 & w66687);
assign w47922 = ~w47656 & w47760;
assign w47923 = ~w47702 & ~w47922;
assign w47924 = w47687 & ~w47923;
assign w47925 = ~w47681 & ~w47694;
assign w47926 = ~w47752 & w64040;
assign w47927 = ~w47696 & ~w47762;
assign w47928 = w47686 & ~w47927;
assign w47929 = (w47644 & w47926) | (w47644 & w66688) | (w47926 & w66688);
assign w47930 = ~w47763 & ~w47916;
assign w47931 = ~w47924 & w47930;
assign w47932 = ~w47921 & w47931;
assign w47933 = ~w47929 & w47932;
assign w47934 = pi2533 & w47933;
assign w47935 = ~pi2533 & ~w47933;
assign w47936 = ~w47934 & ~w47935;
assign w47937 = ~w47324 & ~w47338;
assign w47938 = w47341 & w47361;
assign w47939 = ~w47359 & ~w47937;
assign w47940 = ~w47938 & w47939;
assign w47941 = ~w47356 & ~w47785;
assign w47942 = ~w47940 & w47941;
assign w47943 = ~w47337 & ~w47942;
assign w47944 = w47362 & w47405;
assign w47945 = w47793 & w47944;
assign w47946 = ~w47337 & w47793;
assign w47947 = ~w47346 & ~w47783;
assign w47948 = ~w47946 & w47947;
assign w47949 = w47370 & w47948;
assign w47950 = w47331 & ~w47414;
assign w47951 = w47337 & ~w47370;
assign w47952 = ~w47950 & w47951;
assign w47953 = ~w47374 & ~w47945;
assign w47954 = ~w47949 & w47953;
assign w47955 = ~w47943 & w47954;
assign w47956 = ~w47952 & w47955;
assign w47957 = pi2545 & ~w47956;
assign w47958 = ~pi2545 & w47956;
assign w47959 = ~w47957 & ~w47958;
assign w47960 = w47586 & w47598;
assign w47961 = w47562 & ~w47579;
assign w47962 = ~w47586 & w47603;
assign w47963 = ~w47960 & ~w47962;
assign w47964 = ~w47961 & w47963;
assign w47965 = ~w47614 & w47902;
assign w47966 = w47964 & w47965;
assign w47967 = w47555 & ~w47589;
assign w47968 = w47561 & w47590;
assign w47969 = ~w47967 & ~w47968;
assign w47970 = (~w47586 & ~w47592) | (~w47586 & w66689) | (~w47592 & w66689);
assign w47971 = ~w47969 & ~w47970;
assign w47972 = ~w47561 & w47590;
assign w47973 = ~w47899 & ~w47972;
assign w47974 = ~w47586 & ~w47973;
assign w47975 = ~w47549 & ~w47971;
assign w47976 = ~w47974 & w47975;
assign w47977 = ~w47966 & ~w47976;
assign w47978 = w47592 & w47601;
assign w47979 = w47629 & ~w47978;
assign w47980 = ~w47626 & ~w47979;
assign w47981 = ~w47977 & ~w47980;
assign w47982 = ~pi2530 & w47981;
assign w47983 = pi2530 & ~w47981;
assign w47984 = ~w47982 & ~w47983;
assign w47985 = ~w47680 & ~w47760;
assign w47986 = ~w47771 & w47985;
assign w47987 = ~w47703 & ~w47760;
assign w47988 = w47705 & ~w47922;
assign w47989 = ~w47987 & w47988;
assign w47990 = w47657 & w47671;
assign w47991 = ~w47680 & w47694;
assign w47992 = ~w47644 & ~w47916;
assign w47993 = ~w47990 & w47992;
assign w47994 = ~w47991 & w47993;
assign w47995 = ~w47989 & w47994;
assign w47996 = ~w47657 & ~w47760;
assign w47997 = ~w47680 & ~w47768;
assign w47998 = ~w47996 & w47997;
assign w47999 = ~w47988 & ~w47998;
assign w48000 = w47644 & ~w47766;
assign w48001 = ~w47999 & w48000;
assign w48002 = ~w47995 & ~w48001;
assign w48003 = ~w47753 & ~w47986;
assign w48004 = ~w47767 & w48003;
assign w48005 = ~w48002 & w48004;
assign w48006 = pi2568 & w48005;
assign w48007 = ~pi2568 & ~w48005;
assign w48008 = ~w48006 & ~w48007;
assign w48009 = w47606 & w47610;
assign w48010 = ~w47592 & w47601;
assign w48011 = (~w48010 & w47621) | (~w48010 & w66690) | (w47621 & w66690);
assign w48012 = ~w47967 & ~w48011;
assign w48013 = w47561 & w47577;
assign w48014 = ~w48009 & ~w48013;
assign w48015 = ~w48012 & w48014;
assign w48016 = w47549 & ~w48015;
assign w48017 = ~w47588 & w47970;
assign w48018 = (w47586 & ~w47587) | (w47586 & w66691) | (~w47587 & w66691);
assign w48019 = w47973 & w48018;
assign w48020 = w47568 & ~w48017;
assign w48021 = ~w48019 & w48020;
assign w48022 = ~w47604 & w48018;
assign w48023 = ~w47586 & ~w47906;
assign w48024 = ~w47968 & w48023;
assign w48025 = ~w48022 & ~w48024;
assign w48026 = ~w47893 & ~w47978;
assign w48027 = ~w47628 & w48026;
assign w48028 = (~w47549 & w48025) | (~w47549 & w66692) | (w48025 & w66692);
assign w48029 = ~w47627 & ~w48021;
assign w48030 = ~w48028 & w48029;
assign w48031 = ~w48016 & w48030;
assign w48032 = pi2531 & ~w48031;
assign w48033 = ~pi2531 & w48031;
assign w48034 = ~w48032 & ~w48033;
assign w48035 = ~w47505 & ~w47529;
assign w48036 = ~w47516 & ~w48035;
assign w48037 = w47520 & w47532;
assign w48038 = ~w47444 & w47532;
assign w48039 = (w47437 & ~w47461) | (w47437 & w64036) | (~w47461 & w64036);
assign w48040 = ~w48038 & w48039;
assign w48041 = ~w47533 & ~w48040;
assign w48042 = w47464 & ~w48037;
assign w48043 = (w47478 & ~w48042) | (w47478 & w66693) | (~w48042 & w66693);
assign w48044 = w47486 & w47494;
assign w48045 = ~w47502 & ~w48044;
assign w48046 = (~w47437 & w48044) | (~w47437 & w66694) | (w48044 & w66694);
assign w48047 = ~w47458 & w47461;
assign w48048 = ~w47460 & w48047;
assign w48049 = ~w48046 & ~w48048;
assign w48050 = ~w47478 & ~w48049;
assign w48051 = ~w47461 & w47516;
assign w48052 = w48035 & w48051;
assign w48053 = (~w48036 & ~w48045) | (~w48036 & w66695) | (~w48045 & w66695);
assign w48054 = ~w48043 & w48053;
assign w48055 = ~w48050 & w48054;
assign w48056 = pi2562 & ~w48055;
assign w48057 = ~pi2562 & w48055;
assign w48058 = ~w48056 & ~w48057;
assign w48059 = w47438 & w47485;
assign w48060 = ~w47499 & ~w47500;
assign w48061 = ~w47482 & w47500;
assign w48062 = ~w47469 & ~w48061;
assign w48063 = ~w48060 & w48062;
assign w48064 = w47530 & ~w48038;
assign w48065 = ~w48063 & w48064;
assign w48066 = ~w47478 & ~w48065;
assign w48067 = w47494 & ~w47499;
assign w48068 = w47478 & w47486;
assign w48069 = ~w48067 & ~w48068;
assign w48070 = w47437 & ~w48069;
assign w48071 = w47431 & w47493;
assign w48072 = ~w47501 & ~w48071;
assign w48073 = ~w47437 & ~w48072;
assign w48074 = ~w47470 & ~w48073;
assign w48075 = w47478 & ~w48074;
assign w48076 = ~w48059 & ~w48066;
assign w48077 = ~w48070 & ~w48075;
assign w48078 = w48076 & w48077;
assign w48079 = pi2574 & ~w48078;
assign w48080 = ~pi2574 & w48078;
assign w48081 = ~w48079 & ~w48080;
assign w48082 = ~pi5207 & pi9040;
assign w48083 = ~pi5543 & ~pi9040;
assign w48084 = ~w48082 & ~w48083;
assign w48085 = pi2491 & ~w48084;
assign w48086 = ~pi2491 & w48084;
assign w48087 = ~w48085 & ~w48086;
assign w48088 = ~pi5378 & pi9040;
assign w48089 = ~pi5358 & ~pi9040;
assign w48090 = ~w48088 & ~w48089;
assign w48091 = pi2508 & ~w48090;
assign w48092 = ~pi2508 & w48090;
assign w48093 = ~w48091 & ~w48092;
assign w48094 = ~pi5421 & pi9040;
assign w48095 = ~pi5203 & ~pi9040;
assign w48096 = ~w48094 & ~w48095;
assign w48097 = pi2505 & ~w48096;
assign w48098 = ~pi2505 & w48096;
assign w48099 = ~w48097 & ~w48098;
assign w48100 = w48093 & ~w48099;
assign w48101 = ~pi5628 & pi9040;
assign w48102 = ~pi5285 & ~pi9040;
assign w48103 = ~w48101 & ~w48102;
assign w48104 = pi2520 & ~w48103;
assign w48105 = ~pi2520 & w48103;
assign w48106 = ~w48104 & ~w48105;
assign w48107 = ~w48093 & ~w48106;
assign w48108 = ~w48100 & ~w48107;
assign w48109 = ~pi5337 & pi9040;
assign w48110 = ~pi5334 & ~pi9040;
assign w48111 = ~w48109 & ~w48110;
assign w48112 = pi2516 & ~w48111;
assign w48113 = ~pi2516 & w48111;
assign w48114 = ~w48112 & ~w48113;
assign w48115 = w48108 & w48114;
assign w48116 = w48099 & ~w48114;
assign w48117 = w48107 & w48116;
assign w48118 = ~w48115 & ~w48117;
assign w48119 = ~pi5285 & pi9040;
assign w48120 = pi5546 & ~pi9040;
assign w48121 = ~w48119 & ~w48120;
assign w48122 = pi2499 & ~w48121;
assign w48123 = ~pi2499 & w48121;
assign w48124 = ~w48122 & ~w48123;
assign w48125 = (~w48124 & w48115) | (~w48124 & w66696) | (w48115 & w66696);
assign w48126 = ~w48099 & w48114;
assign w48127 = w48106 & ~w48116;
assign w48128 = ~w48126 & w48127;
assign w48129 = ~w48125 & ~w48128;
assign w48130 = ~w48087 & ~w48129;
assign w48131 = w48093 & w48106;
assign w48132 = w48099 & w48114;
assign w48133 = w48131 & w48132;
assign w48134 = ~w48087 & w48093;
assign w48135 = ~w48099 & ~w48106;
assign w48136 = w48114 & w48135;
assign w48137 = ~w48134 & w48136;
assign w48138 = w48087 & ~w48106;
assign w48139 = w48100 & ~w48114;
assign w48140 = ~w48138 & w48139;
assign w48141 = ~w48133 & ~w48137;
assign w48142 = (~w48124 & ~w48141) | (~w48124 & w66697) | (~w48141 & w66697);
assign w48143 = w48087 & ~w48117;
assign w48144 = ~w48107 & ~w48116;
assign w48145 = ~w48131 & ~w48144;
assign w48146 = w48143 & w48145;
assign w48147 = w48099 & ~w48106;
assign w48148 = w48093 & ~w48114;
assign w48149 = w48147 & w48148;
assign w48150 = w48106 & ~w48114;
assign w48151 = ~w48136 & ~w48150;
assign w48152 = w48134 & ~w48151;
assign w48153 = w48087 & w48114;
assign w48154 = w48100 & w48106;
assign w48155 = ~w48147 & ~w48154;
assign w48156 = w48153 & ~w48155;
assign w48157 = ~w48093 & ~w48114;
assign w48158 = w48135 & w48157;
assign w48159 = ~w48149 & ~w48158;
assign w48160 = ~w48152 & w48159;
assign w48161 = ~w48156 & w48160;
assign w48162 = w48124 & ~w48161;
assign w48163 = ~w48142 & ~w48146;
assign w48164 = ~w48130 & w48163;
assign w48165 = ~w48162 & w48164;
assign w48166 = pi2534 & ~w48165;
assign w48167 = ~pi2534 & w48165;
assign w48168 = ~w48166 & ~w48167;
assign w48169 = w48100 & ~w48151;
assign w48170 = w48106 & w48114;
assign w48171 = ~w48158 & ~w48170;
assign w48172 = w48087 & ~w48171;
assign w48173 = ~w48087 & w48149;
assign w48174 = ~w48093 & w48099;
assign w48175 = w48118 & w48174;
assign w48176 = w48124 & ~w48173;
assign w48177 = ~w48169 & w48176;
assign w48178 = ~w48172 & w48177;
assign w48179 = ~w48175 & w48178;
assign w48180 = ~w48087 & w48132;
assign w48181 = w48099 & w48106;
assign w48182 = w48093 & w48114;
assign w48183 = w48147 & w48182;
assign w48184 = ~w48093 & w48150;
assign w48185 = ~w48183 & ~w48184;
assign w48186 = ~w48181 & ~w48185;
assign w48187 = w48138 & w48148;
assign w48188 = ~w48107 & ~w48131;
assign w48189 = ~w48116 & ~w48136;
assign w48190 = ~w48188 & ~w48189;
assign w48191 = ~w48087 & ~w48188;
assign w48192 = ~w48124 & ~w48180;
assign w48193 = ~w48187 & w48192;
assign w48194 = ~w48191 & w48193;
assign w48195 = ~w48186 & ~w48190;
assign w48196 = w48194 & w48195;
assign w48197 = ~w48179 & ~w48196;
assign w48198 = pi2529 & w48197;
assign w48199 = ~pi2529 & ~w48197;
assign w48200 = ~w48198 & ~w48199;
assign w48201 = ~w48157 & ~w48182;
assign w48202 = ~w48099 & ~w48201;
assign w48203 = ~w48201 & w66698;
assign w48204 = w48087 & ~w48203;
assign w48205 = w48106 & w48116;
assign w48206 = ~w48087 & ~w48205;
assign w48207 = ~w48182 & ~w48184;
assign w48208 = w48189 & w48207;
assign w48209 = w48206 & ~w48208;
assign w48210 = w48181 & w48201;
assign w48211 = ~w48183 & ~w48210;
assign w48212 = (w48211 & w48209) | (w48211 & w66699) | (w48209 & w66699);
assign w48213 = w48124 & ~w48212;
assign w48214 = ~w48124 & ~w48202;
assign w48215 = w48211 & w48214;
assign w48216 = w48143 & ~w48215;
assign w48217 = ~w48117 & ~w48203;
assign w48218 = ~w48124 & ~w48217;
assign w48219 = ~w48087 & w48211;
assign w48220 = ~w48218 & w48219;
assign w48221 = ~w48216 & ~w48220;
assign w48222 = ~w48213 & ~w48221;
assign w48223 = ~pi2539 & w48222;
assign w48224 = pi2539 & ~w48222;
assign w48225 = ~w48223 & ~w48224;
assign w48226 = ~w47836 & ~w47843;
assign w48227 = w47827 & w47871;
assign w48228 = ~w47814 & ~w47878;
assign w48229 = w47884 & ~w48228;
assign w48230 = w47813 & ~w47820;
assign w48231 = ~w47826 & ~w47832;
assign w48232 = ~w48230 & ~w48231;
assign w48233 = (w47843 & ~w48230) | (w47843 & w66700) | (~w48230 & w66700);
assign w48234 = ~w48232 & w48233;
assign w48235 = w47832 & w47857;
assign w48236 = ~w47867 & ~w48235;
assign w48237 = ~w48229 & w48236;
assign w48238 = ~w48234 & w48237;
assign w48239 = ~w47829 & ~w47885;
assign w48240 = w47826 & w47832;
assign w48241 = ~w47873 & ~w48240;
assign w48242 = w47807 & w47868;
assign w48243 = (~w47843 & ~w47868) | (~w47843 & w66701) | (~w47868 & w66701);
assign w48244 = w48241 & w48243;
assign w48245 = ~w47877 & w48233;
assign w48246 = ~w47847 & ~w48242;
assign w48247 = w47843 & ~w48246;
assign w48248 = ~w48244 & ~w48245;
assign w48249 = ~w47854 & w47867;
assign w48250 = w48239 & w48249;
assign w48251 = (w48250 & ~w48248) | (w48250 & w66702) | (~w48248 & w66702);
assign w48252 = ~w48238 & ~w48251;
assign w48253 = ~w48226 & ~w48227;
assign w48254 = ~w47851 & w48253;
assign w48255 = ~w48252 & w48254;
assign w48256 = pi2573 & w48255;
assign w48257 = ~pi2573 & ~w48255;
assign w48258 = ~w48256 & ~w48257;
assign w48259 = w47828 & ~w47879;
assign w48260 = w47813 & w47820;
assign w48261 = w47858 & w47884;
assign w48262 = ~w48260 & ~w48261;
assign w48263 = ~w47807 & ~w48262;
assign w48264 = ~w47826 & ~w47874;
assign w48265 = w48236 & ~w48259;
assign w48266 = ~w48247 & w48265;
assign w48267 = ~w48263 & ~w48264;
assign w48268 = w48266 & w48267;
assign w48269 = ~w47832 & ~w47834;
assign w48270 = ~w47828 & ~w48260;
assign w48271 = w47813 & w47845;
assign w48272 = ~w47833 & ~w48271;
assign w48273 = w47843 & ~w48270;
assign w48274 = w48272 & w48273;
assign w48275 = (w47867 & w47830) | (w47867 & w66703) | (w47830 & w66703);
assign w48276 = ~w48274 & w48275;
assign w48277 = ~w47850 & w48276;
assign w48278 = ~w48268 & ~w48277;
assign w48279 = ~w47820 & w47859;
assign w48280 = ~w48228 & w48279;
assign w48281 = ~w48278 & ~w48280;
assign w48282 = pi2567 & w48281;
assign w48283 = ~pi2567 & ~w48281;
assign w48284 = ~w48282 & ~w48283;
assign w48285 = ~pi5346 & pi9040;
assign w48286 = ~pi5333 & ~pi9040;
assign w48287 = ~w48285 & ~w48286;
assign w48288 = pi2513 & ~w48287;
assign w48289 = ~pi2513 & w48287;
assign w48290 = ~w48288 & ~w48289;
assign w48291 = ~pi5338 & pi9040;
assign w48292 = ~pi5662 & ~pi9040;
assign w48293 = ~w48291 & ~w48292;
assign w48294 = pi2526 & ~w48293;
assign w48295 = ~pi2526 & w48293;
assign w48296 = ~w48294 & ~w48295;
assign w48297 = ~w48290 & ~w48296;
assign w48298 = w48290 & ~w48296;
assign w48299 = ~pi5333 & pi9040;
assign w48300 = ~pi5212 & ~pi9040;
assign w48301 = ~w48299 & ~w48300;
assign w48302 = pi2514 & ~w48301;
assign w48303 = ~pi2514 & w48301;
assign w48304 = ~w48302 & ~w48303;
assign w48305 = ~w48290 & ~w48304;
assign w48306 = ~pi5340 & pi9040;
assign w48307 = ~pi5348 & ~pi9040;
assign w48308 = ~w48306 & ~w48307;
assign w48309 = pi2511 & ~w48308;
assign w48310 = ~pi2511 & w48308;
assign w48311 = ~w48309 & ~w48310;
assign w48312 = ~w48305 & w48311;
assign w48313 = ~w48298 & w48312;
assign w48314 = ~w48296 & ~w48311;
assign w48315 = w48297 & w48304;
assign w48316 = w48314 & ~w48315;
assign w48317 = ~w48313 & ~w48316;
assign w48318 = ~pi5662 & pi9040;
assign w48319 = ~pi5341 & ~pi9040;
assign w48320 = ~w48318 & ~w48319;
assign w48321 = pi2498 & ~w48320;
assign w48322 = ~pi2498 & w48320;
assign w48323 = ~w48321 & ~w48322;
assign w48324 = ~w48317 & ~w48323;
assign w48325 = ~w48317 & w66704;
assign w48326 = w48305 & ~w48311;
assign w48327 = w48290 & w48304;
assign w48328 = w48296 & w48327;
assign w48329 = ~w48326 & ~w48328;
assign w48330 = ~w48296 & w48304;
assign w48331 = w48296 & ~w48304;
assign w48332 = ~w48330 & ~w48331;
assign w48333 = ~w48305 & ~w48327;
assign w48334 = ~w48311 & ~w48323;
assign w48335 = w48332 & w48334;
assign w48336 = w48333 & w48335;
assign w48337 = w48329 & ~w48336;
assign w48338 = w48317 & ~w48337;
assign w48339 = ~w48296 & w48311;
assign w48340 = ~w48333 & w48339;
assign w48341 = ~w48290 & w48311;
assign w48342 = ~w48331 & ~w48341;
assign w48343 = ~w48297 & w48323;
assign w48344 = w48332 & w48343;
assign w48345 = w48290 & w48311;
assign w48346 = (~w48342 & w48344) | (~w48342 & w66705) | (w48344 & w66705);
assign w48347 = w48290 & ~w48311;
assign w48348 = ~w48323 & ~w48347;
assign w48349 = w48314 & w48333;
assign w48350 = ~w48348 & w48349;
assign w48351 = ~w48340 & ~w48350;
assign w48352 = ~w48346 & w48351;
assign w48353 = ~w48338 & w48352;
assign w48354 = ~pi5294 & pi9040;
assign w48355 = ~pi5292 & ~pi9040;
assign w48356 = ~w48354 & ~w48355;
assign w48357 = pi2482 & ~w48356;
assign w48358 = ~pi2482 & w48356;
assign w48359 = ~w48357 & ~w48358;
assign w48360 = ~w48353 & ~w48359;
assign w48361 = w48296 & w48311;
assign w48362 = w48359 & w48361;
assign w48363 = w48305 & w48362;
assign w48364 = ~w48305 & ~w48342;
assign w48365 = (~w48330 & w48342) | (~w48330 & w66706) | (w48342 & w66706);
assign w48366 = ~w48323 & w48359;
assign w48367 = ~w48365 & w48366;
assign w48368 = ~w48331 & ~w48345;
assign w48369 = w48361 & w48368;
assign w48370 = w48359 & ~w48369;
assign w48371 = w48344 & w48370;
assign w48372 = ~w48296 & ~w48304;
assign w48373 = ~w48323 & ~w48372;
assign w48374 = w48290 & w48332;
assign w48375 = ~w48304 & w48323;
assign w48376 = ~w48290 & ~w48375;
assign w48377 = ~w48332 & w48376;
assign w48378 = ~w48374 & ~w48377;
assign w48379 = w48378 & w66707;
assign w48380 = ~w48363 & ~w48367;
assign w48381 = ~w48371 & w48380;
assign w48382 = ~w48325 & ~w48379;
assign w48383 = w48381 & w48382;
assign w48384 = ~w48360 & w66708;
assign w48385 = (pi2555 & w48360) | (pi2555 & w66709) | (w48360 & w66709);
assign w48386 = ~w48384 & ~w48385;
assign w48387 = ~w48137 & w48191;
assign w48388 = ~w48093 & ~w48126;
assign w48389 = ~w48150 & w48388;
assign w48390 = ~w48131 & w48153;
assign w48391 = ~w48389 & w48390;
assign w48392 = ~w48387 & ~w48391;
assign w48393 = ~w48124 & ~w48392;
assign w48394 = ~w48154 & ~w48389;
assign w48395 = w48392 & ~w48394;
assign w48396 = w48135 & w48201;
assign w48397 = w48185 & ~w48396;
assign w48398 = ~w48087 & ~w48397;
assign w48399 = (w48124 & w48395) | (w48124 & w66710) | (w48395 & w66710);
assign w48400 = w48108 & w48215;
assign w48401 = w48087 & ~w48149;
assign w48402 = w48100 & w48170;
assign w48403 = w48206 & ~w48402;
assign w48404 = ~w48401 & ~w48403;
assign w48405 = ~w48393 & ~w48404;
assign w48406 = ~w48400 & w48405;
assign w48407 = (pi2543 & ~w48406) | (pi2543 & w66711) | (~w48406 & w66711);
assign w48408 = w48406 & w66712;
assign w48409 = ~w48407 & ~w48408;
assign w48410 = w48314 & ~w48333;
assign w48411 = ~w48364 & ~w48410;
assign w48412 = ~w48296 & ~w48411;
assign w48413 = w48323 & ~w48368;
assign w48414 = w48311 & w48331;
assign w48415 = ~w48368 & ~w48414;
assign w48416 = ~w48343 & ~w48415;
assign w48417 = ~w48413 & ~w48416;
assign w48418 = ~w48412 & ~w48417;
assign w48419 = ~w48359 & ~w48418;
assign w48420 = ~w48312 & ~w48326;
assign w48421 = w48375 & w48420;
assign w48422 = w48370 & ~w48421;
assign w48423 = ~w48414 & ~w48422;
assign w48424 = w48413 & ~w48423;
assign w48425 = w48290 & ~w48372;
assign w48426 = w48366 & ~w48425;
assign w48427 = w48420 & w48426;
assign w48428 = ~w48327 & w48362;
assign w48429 = ~w48427 & ~w48428;
assign w48430 = ~w48379 & w48429;
assign w48431 = ~w48419 & w48430;
assign w48432 = w48431 & w66713;
assign w48433 = (~pi2550 & ~w48431) | (~pi2550 & w66714) | (~w48431 & w66714);
assign w48434 = ~w48432 & ~w48433;
assign w48435 = w48328 & w48413;
assign w48436 = w48323 & ~w48411;
assign w48437 = ~w48314 & w48323;
assign w48438 = w48298 & w48437;
assign w48439 = ~w48348 & ~w48438;
assign w48440 = ~w48333 & w48437;
assign w48441 = ~w48350 & ~w48440;
assign w48442 = ~w48324 & w48441;
assign w48443 = (~w48436 & ~w48442) | (~w48436 & w64041) | (~w48442 & w64041);
assign w48444 = ~w48359 & ~w48443;
assign w48445 = ~w48336 & ~w48435;
assign w48446 = (w48445 & w48442) | (w48445 & w66715) | (w48442 & w66715);
assign w48447 = (pi2551 & w48444) | (pi2551 & w66716) | (w48444 & w66716);
assign w48448 = ~w48444 & w66717;
assign w48449 = ~w48447 & ~w48448;
assign w48450 = ~w48323 & ~w48342;
assign w48451 = (w48450 & ~w48351) | (w48450 & w66718) | (~w48351 & w66718);
assign w48452 = ~w48311 & ~w48378;
assign w48453 = w48422 & ~w48452;
assign w48454 = ~w48315 & w48329;
assign w48455 = ~w48373 & ~w48454;
assign w48456 = (~w48359 & ~w48378) | (~w48359 & w66719) | (~w48378 & w66719);
assign w48457 = ~w48455 & w48456;
assign w48458 = ~w48453 & ~w48457;
assign w48459 = ~w48438 & ~w48451;
assign w48460 = ~w48458 & w48459;
assign w48461 = pi2556 & w48460;
assign w48462 = ~pi2556 & ~w48460;
assign w48463 = ~w48461 & ~w48462;
assign w48464 = w47872 & ~w48239;
assign w48465 = ~w47846 & ~w47878;
assign w48466 = ~w47813 & ~w48465;
assign w48467 = ~w47852 & w48245;
assign w48468 = w47843 & ~w48467;
assign w48469 = ~w48466 & ~w48468;
assign w48470 = ~w47867 & ~w48469;
assign w48471 = w47814 & w47853;
assign w48472 = ~w47848 & ~w48261;
assign w48473 = w48272 & w48472;
assign w48474 = ~w48471 & w48473;
assign w48475 = w47867 & ~w48474;
assign w48476 = ~w48232 & ~w48241;
assign w48477 = ~w47833 & ~w47847;
assign w48478 = (~w47843 & w48476) | (~w47843 & w66720) | (w48476 & w66720);
assign w48479 = ~w48464 & ~w48478;
assign w48480 = ~w48475 & w48479;
assign w48481 = ~w48470 & w48480;
assign w48482 = pi2588 & w48481;
assign w48483 = ~pi2588 & ~w48481;
assign w48484 = ~w48482 & ~w48483;
assign w48485 = ~pi5608 & pi9040;
assign w48486 = ~pi5882 & ~pi9040;
assign w48487 = ~w48485 & ~w48486;
assign w48488 = pi2575 & ~w48487;
assign w48489 = ~pi2575 & w48487;
assign w48490 = ~w48488 & ~w48489;
assign w48491 = ~pi5532 & pi9040;
assign w48492 = ~pi5618 & ~pi9040;
assign w48493 = ~w48491 & ~w48492;
assign w48494 = pi2537 & ~w48493;
assign w48495 = ~pi2537 & w48493;
assign w48496 = ~w48494 & ~w48495;
assign w48497 = ~pi5562 & pi9040;
assign w48498 = ~pi5626 & ~pi9040;
assign w48499 = ~w48497 & ~w48498;
assign w48500 = pi2578 & ~w48499;
assign w48501 = ~pi2578 & w48499;
assign w48502 = ~w48500 & ~w48501;
assign w48503 = ~w48496 & w48502;
assign w48504 = ~pi5459 & pi9040;
assign w48505 = ~pi5530 & ~pi9040;
assign w48506 = ~w48504 & ~w48505;
assign w48507 = pi2577 & ~w48506;
assign w48508 = ~pi2577 & w48506;
assign w48509 = ~w48507 & ~w48508;
assign w48510 = w48503 & w48509;
assign w48511 = ~pi5634 & pi9040;
assign w48512 = ~pi5793 & ~pi9040;
assign w48513 = ~w48511 & ~w48512;
assign w48514 = pi2569 & ~w48513;
assign w48515 = ~pi2569 & w48513;
assign w48516 = ~w48514 & ~w48515;
assign w48517 = (~w48516 & ~w48503) | (~w48516 & w66721) | (~w48503 & w66721);
assign w48518 = ~w48496 & w48509;
assign w48519 = w48496 & ~w48509;
assign w48520 = ~w48518 & ~w48519;
assign w48521 = ~pi5537 & pi9040;
assign w48522 = ~pi5619 & ~pi9040;
assign w48523 = ~w48521 & ~w48522;
assign w48524 = pi2570 & ~w48523;
assign w48525 = ~pi2570 & w48523;
assign w48526 = ~w48524 & ~w48525;
assign w48527 = ~w48502 & w48526;
assign w48528 = ~w48496 & ~w48502;
assign w48529 = ~w48527 & ~w48528;
assign w48530 = w48520 & ~w48529;
assign w48531 = w48517 & ~w48530;
assign w48532 = w48496 & w48502;
assign w48533 = w48526 & w48532;
assign w48534 = ~w48528 & ~w48533;
assign w48535 = w48520 & w48534;
assign w48536 = w48502 & ~w48509;
assign w48537 = w48526 & w48536;
assign w48538 = ~w48502 & ~w48526;
assign w48539 = w48496 & w48538;
assign w48540 = ~w48537 & ~w48539;
assign w48541 = w48516 & w48540;
assign w48542 = ~w48535 & w48541;
assign w48543 = ~w48542 & w66722;
assign w48544 = w48510 & ~w48526;
assign w48545 = w48526 & w48528;
assign w48546 = (w48516 & ~w48528) | (w48516 & w66723) | (~w48528 & w66723);
assign w48547 = ~w48544 & w48546;
assign w48548 = w48496 & w48526;
assign w48549 = ~w48516 & ~w48548;
assign w48550 = w48509 & w48538;
assign w48551 = w48549 & ~w48550;
assign w48552 = ~w48547 & ~w48551;
assign w48553 = ~w48533 & ~w48536;
assign w48554 = (~w48553 & w48542) | (~w48553 & w64042) | (w48542 & w64042);
assign w48555 = (~w48490 & w48554) | (~w48490 & w66724) | (w48554 & w66724);
assign w48556 = ~w48509 & ~w48526;
assign w48557 = w48509 & w48526;
assign w48558 = ~w48556 & ~w48557;
assign w48559 = w48528 & ~w48558;
assign w48560 = ~w48519 & ~w48540;
assign w48561 = (w48516 & w48560) | (w48516 & w66725) | (w48560 & w66725);
assign w48562 = w48502 & ~w48516;
assign w48563 = w48496 & w48556;
assign w48564 = w48562 & w48563;
assign w48565 = ~w48561 & ~w48564;
assign w48566 = ~w48543 & w48565;
assign w48567 = ~w48555 & w48566;
assign w48568 = pi2598 & ~w48567;
assign w48569 = ~pi2598 & w48567;
assign w48570 = ~w48568 & ~w48569;
assign w48571 = ~pi5449 & pi9040;
assign w48572 = ~pi5685 & ~pi9040;
assign w48573 = ~w48571 & ~w48572;
assign w48574 = pi2578 & ~w48573;
assign w48575 = ~pi2578 & w48573;
assign w48576 = ~w48574 & ~w48575;
assign w48577 = ~pi5547 & pi9040;
assign w48578 = ~pi5625 & ~pi9040;
assign w48579 = ~w48577 & ~w48578;
assign w48580 = pi2576 & ~w48579;
assign w48581 = ~pi2576 & w48579;
assign w48582 = ~w48580 & ~w48581;
assign w48583 = ~pi5802 & pi9040;
assign w48584 = ~pi5636 & ~pi9040;
assign w48585 = ~w48583 & ~w48584;
assign w48586 = pi2563 & ~w48585;
assign w48587 = ~pi2563 & w48585;
assign w48588 = ~w48586 & ~w48587;
assign w48589 = ~w48582 & w48588;
assign w48590 = ~pi5552 & pi9040;
assign w48591 = ~pi5450 & ~pi9040;
assign w48592 = ~w48590 & ~w48591;
assign w48593 = pi2554 & ~w48592;
assign w48594 = ~pi2554 & w48592;
assign w48595 = ~w48593 & ~w48594;
assign w48596 = ~pi5464 & pi9040;
assign w48597 = ~pi5633 & ~pi9040;
assign w48598 = ~w48596 & ~w48597;
assign w48599 = pi2589 & ~w48598;
assign w48600 = ~pi2589 & w48598;
assign w48601 = ~w48599 & ~w48600;
assign w48602 = (~w48601 & ~w48589) | (~w48601 & w66726) | (~w48589 & w66726);
assign w48603 = w48582 & w48595;
assign w48604 = ~pi5625 & pi9040;
assign w48605 = ~pi5449 & ~pi9040;
assign w48606 = ~w48604 & ~w48605;
assign w48607 = pi2537 & ~w48606;
assign w48608 = ~pi2537 & w48606;
assign w48609 = ~w48607 & ~w48608;
assign w48610 = ~w48588 & w48609;
assign w48611 = w48603 & w48610;
assign w48612 = w48602 & ~w48611;
assign w48613 = w48588 & ~w48595;
assign w48614 = ~w48582 & ~w48609;
assign w48615 = w48582 & w48609;
assign w48616 = ~w48614 & ~w48615;
assign w48617 = w48613 & ~w48616;
assign w48618 = ~w48603 & ~w48617;
assign w48619 = w48612 & ~w48618;
assign w48620 = w48582 & ~w48588;
assign w48621 = ~w48601 & w48609;
assign w48622 = ~w48595 & w48620;
assign w48623 = ~w48621 & w48622;
assign w48624 = ~w48619 & ~w48623;
assign w48625 = ~w48576 & ~w48624;
assign w48626 = w48595 & ~w48601;
assign w48627 = w48595 & w48609;
assign w48628 = w48582 & w48588;
assign w48629 = w48621 & ~w48628;
assign w48630 = (~w48576 & w48629) | (~w48576 & w66727) | (w48629 & w66727);
assign w48631 = ~w48626 & ~w48630;
assign w48632 = ~w48589 & ~w48620;
assign w48633 = ~w48631 & w48632;
assign w48634 = ~w48582 & ~w48595;
assign w48635 = w48588 & ~w48609;
assign w48636 = w48634 & w48635;
assign w48637 = w48601 & ~w48636;
assign w48638 = ~w48595 & ~w48609;
assign w48639 = ~w48627 & ~w48638;
assign w48640 = w48589 & w48639;
assign w48641 = ~w48638 & ~w48640;
assign w48642 = w48637 & ~w48641;
assign w48643 = ~w48603 & ~w48634;
assign w48644 = w48629 & w48643;
assign w48645 = w48582 & w48601;
assign w48646 = ~w48611 & ~w48613;
assign w48647 = w48645 & ~w48646;
assign w48648 = ~w48610 & ~w48635;
assign w48649 = w48634 & w48648;
assign w48650 = ~w48644 & ~w48649;
assign w48651 = ~w48647 & w48650;
assign w48652 = w48576 & ~w48651;
assign w48653 = ~w48633 & ~w48642;
assign w48654 = ~w48652 & w48653;
assign w48655 = ~w48625 & w48654;
assign w48656 = ~pi2605 & w48655;
assign w48657 = pi2605 & ~w48655;
assign w48658 = ~w48656 & ~w48657;
assign w48659 = w48613 & w48615;
assign w48660 = w48595 & w48616;
assign w48661 = w48616 & w66728;
assign w48662 = ~w48659 & ~w48661;
assign w48663 = ~w48588 & ~w48616;
assign w48664 = ~w48616 & w66729;
assign w48665 = w48601 & ~w48664;
assign w48666 = ~w48634 & w48648;
assign w48667 = w48632 & ~w48666;
assign w48668 = w48602 & ~w48660;
assign w48669 = ~w48667 & w48668;
assign w48670 = (w48662 & w48669) | (w48662 & w66730) | (w48669 & w66730);
assign w48671 = w48576 & ~w48670;
assign w48672 = ~w48576 & ~w48663;
assign w48673 = w48662 & w48672;
assign w48674 = w48637 & ~w48673;
assign w48675 = ~w48636 & ~w48664;
assign w48676 = ~w48576 & ~w48675;
assign w48677 = ~w48601 & w48662;
assign w48678 = ~w48676 & w48677;
assign w48679 = ~w48674 & ~w48678;
assign w48680 = ~w48671 & ~w48679;
assign w48681 = ~pi2614 & w48680;
assign w48682 = pi2614 & ~w48680;
assign w48683 = ~w48681 & ~w48682;
assign w48684 = w48609 & w48634;
assign w48685 = w48588 & w48684;
assign w48686 = ~w48601 & w48685;
assign w48687 = w48643 & ~w48648;
assign w48688 = w48601 & ~w48685;
assign w48689 = ~w48603 & ~w48649;
assign w48690 = w48688 & ~w48689;
assign w48691 = w48576 & ~w48687;
assign w48692 = ~w48686 & w48691;
assign w48693 = ~w48690 & w48692;
assign w48694 = ~w48610 & w48643;
assign w48695 = ~w48588 & w48694;
assign w48696 = ~w48601 & ~w48639;
assign w48697 = ~w48628 & ~w48661;
assign w48698 = ~w48645 & ~w48697;
assign w48699 = w48601 & w48684;
assign w48700 = ~w48576 & ~w48617;
assign w48701 = ~w48696 & ~w48699;
assign w48702 = w48700 & w48701;
assign w48703 = ~w48695 & w48702;
assign w48704 = ~w48698 & w48703;
assign w48705 = ~w48693 & ~w48704;
assign w48706 = pi2603 & w48705;
assign w48707 = ~pi2603 & ~w48705;
assign w48708 = ~w48706 & ~w48707;
assign w48709 = w48503 & w48558;
assign w48710 = w48496 & ~w48502;
assign w48711 = ~w48558 & ~w48562;
assign w48712 = ~w48548 & ~w48710;
assign w48713 = ~w48709 & w48712;
assign w48714 = w48516 & ~w48556;
assign w48715 = ~w48516 & ~w48538;
assign w48716 = w48520 & ~w48715;
assign w48717 = w48519 & w48527;
assign w48718 = ~w48716 & ~w48717;
assign w48719 = ~w48538 & w48714;
assign w48720 = ~w48718 & w48719;
assign w48721 = (w48490 & ~w48713) | (w48490 & w66731) | (~w48713 & w66731);
assign w48722 = ~w48720 & w48721;
assign w48723 = w48509 & w48710;
assign w48724 = ~w48526 & w48532;
assign w48725 = ~w48510 & ~w48724;
assign w48726 = w48516 & ~w48725;
assign w48727 = ~w48516 & w48539;
assign w48728 = w48537 & ~w48716;
assign w48729 = w48559 & ~w48714;
assign w48730 = ~w48490 & ~w48723;
assign w48731 = ~w48544 & w48730;
assign w48732 = ~w48727 & w48731;
assign w48733 = ~w48726 & ~w48728;
assign w48734 = ~w48729 & w48733;
assign w48735 = w48732 & w48734;
assign w48736 = ~w48533 & ~w48539;
assign w48737 = w48516 & ~w48723;
assign w48738 = ~w48736 & w48737;
assign w48739 = ~w48503 & ~w48516;
assign w48740 = ~w48518 & w48739;
assign w48741 = w48736 & w48740;
assign w48742 = ~w48738 & ~w48741;
assign w48743 = ~w48509 & ~w48534;
assign w48744 = w48742 & w48743;
assign w48745 = (~w48744 & w48735) | (~w48744 & w66732) | (w48735 & w66732);
assign w48746 = ~pi2623 & w48745;
assign w48747 = pi2623 & ~w48745;
assign w48748 = ~w48746 & ~w48747;
assign w48749 = w48549 & w48560;
assign w48750 = w48520 & w48527;
assign w48751 = ~w48709 & ~w48750;
assign w48752 = w48742 & w48751;
assign w48753 = w48490 & ~w48752;
assign w48754 = w48490 & ~w48518;
assign w48755 = ~w48519 & w48526;
assign w48756 = ~w48563 & ~w48754;
assign w48757 = ~w48755 & w48756;
assign w48758 = w48737 & w48757;
assign w48759 = ~w48528 & ~w48562;
assign w48760 = w48557 & ~w48759;
assign w48761 = ~w48727 & ~w48760;
assign w48762 = ~w48490 & ~w48761;
assign w48763 = ~w48564 & ~w48749;
assign w48764 = ~w48758 & ~w48762;
assign w48765 = w48763 & w48764;
assign w48766 = ~w48753 & w48765;
assign w48767 = pi2641 & ~w48766;
assign w48768 = ~pi2641 & w48766;
assign w48769 = ~w48767 & ~w48768;
assign w48770 = ~w48612 & ~w48688;
assign w48771 = ~w48603 & w48639;
assign w48772 = ~w48666 & ~w48771;
assign w48773 = w48603 & w48635;
assign w48774 = w48639 & w48694;
assign w48775 = ~w48588 & ~w48595;
assign w48776 = w48616 & w48775;
assign w48777 = (~w48601 & w48774) | (~w48601 & w66733) | (w48774 & w66733);
assign w48778 = w48576 & ~w48773;
assign w48779 = (w48778 & ~w48772) | (w48778 & w66734) | (~w48772 & w66734);
assign w48780 = ~w48777 & w48779;
assign w48781 = ~w48603 & ~w48645;
assign w48782 = ~w48772 & ~w48781;
assign w48783 = w48696 & ~w48776;
assign w48784 = ~w48576 & ~w48640;
assign w48785 = ~w48783 & w48784;
assign w48786 = ~w48782 & w48785;
assign w48787 = ~w48780 & ~w48786;
assign w48788 = ~w48770 & ~w48787;
assign w48789 = ~pi2619 & w48788;
assign w48790 = pi2619 & ~w48788;
assign w48791 = ~w48789 & ~w48790;
assign w48792 = ~pi5793 & pi9040;
assign w48793 = ~pi5460 & ~pi9040;
assign w48794 = ~w48792 & ~w48793;
assign w48795 = pi2572 & ~w48794;
assign w48796 = ~pi2572 & w48794;
assign w48797 = ~w48795 & ~w48796;
assign w48798 = ~pi5618 & pi9040;
assign w48799 = ~pi5537 & ~pi9040;
assign w48800 = ~w48798 & ~w48799;
assign w48801 = pi2559 & ~w48800;
assign w48802 = ~pi2559 & w48800;
assign w48803 = ~w48801 & ~w48802;
assign w48804 = ~w48797 & ~w48803;
assign w48805 = ~pi5450 & pi9040;
assign w48806 = ~pi5802 & ~pi9040;
assign w48807 = ~w48805 & ~w48806;
assign w48808 = pi2560 & ~w48807;
assign w48809 = ~pi2560 & w48807;
assign w48810 = ~w48808 & ~w48809;
assign w48811 = ~pi5878 & pi9040;
assign w48812 = ~pi5552 & ~pi9040;
assign w48813 = ~w48811 & ~w48812;
assign w48814 = pi2585 & ~w48813;
assign w48815 = ~pi2585 & w48813;
assign w48816 = ~w48814 & ~w48815;
assign w48817 = ~w48810 & ~w48816;
assign w48818 = ~pi5636 & pi9040;
assign w48819 = ~pi5608 & ~pi9040;
assign w48820 = ~w48818 & ~w48819;
assign w48821 = pi2554 & ~w48820;
assign w48822 = ~pi2554 & w48820;
assign w48823 = ~w48821 & ~w48822;
assign w48824 = w48817 & ~w48823;
assign w48825 = w48804 & w48824;
assign w48826 = w48810 & w48823;
assign w48827 = w48803 & ~w48810;
assign w48828 = ~w48826 & ~w48827;
assign w48829 = (w48797 & w48828) | (w48797 & w64043) | (w48828 & w64043);
assign w48830 = ~w48803 & w48810;
assign w48831 = ~w48816 & ~w48823;
assign w48832 = w48830 & w48831;
assign w48833 = w48829 & ~w48832;
assign w48834 = w48804 & w48826;
assign w48835 = ~w48797 & ~w48834;
assign w48836 = ~w48827 & ~w48830;
assign w48837 = w48816 & ~w48826;
assign w48838 = w48836 & w48837;
assign w48839 = w48835 & ~w48838;
assign w48840 = ~w48797 & w48816;
assign w48841 = ~w48810 & w48816;
assign w48842 = w48823 & w48841;
assign w48843 = w48840 & ~w48842;
assign w48844 = w48803 & ~w48826;
assign w48845 = ~w48841 & w48844;
assign w48846 = (~w48845 & w48839) | (~w48845 & w66735) | (w48839 & w66735);
assign w48847 = ~pi5541 & pi9040;
assign w48848 = ~pi5532 & ~pi9040;
assign w48849 = ~w48847 & ~w48848;
assign w48850 = pi2576 & ~w48849;
assign w48851 = ~pi2576 & w48849;
assign w48852 = ~w48850 & ~w48851;
assign w48853 = ~w48833 & w48852;
assign w48854 = ~w48846 & w48853;
assign w48855 = w48797 & ~w48810;
assign w48856 = w48810 & ~w48823;
assign w48857 = w48816 & w48856;
assign w48858 = ~w48855 & ~w48857;
assign w48859 = ~w48803 & ~w48858;
assign w48860 = ~w48836 & w48840;
assign w48861 = w48797 & w48823;
assign w48862 = w48817 & w48861;
assign w48863 = w48804 & w48856;
assign w48864 = w48810 & ~w48816;
assign w48865 = w48803 & w48823;
assign w48866 = w48864 & w48865;
assign w48867 = ~w48863 & ~w48866;
assign w48868 = w48797 & w48803;
assign w48869 = w48864 & w48868;
assign w48870 = ~w48862 & ~w48869;
assign w48871 = ~w48860 & w48870;
assign w48872 = w48867 & w48871;
assign w48873 = ~w48859 & w48872;
assign w48874 = ~w48852 & ~w48873;
assign w48875 = ~w48803 & ~w48823;
assign w48876 = w48817 & ~w48865;
assign w48877 = ~w48875 & w48876;
assign w48878 = w48867 & ~w48877;
assign w48879 = w48816 & w48875;
assign w48880 = ~w48862 & ~w48879;
assign w48881 = ~w48878 & ~w48880;
assign w48882 = w48803 & w48826;
assign w48883 = w48841 & w48875;
assign w48884 = ~w48882 & ~w48883;
assign w48885 = w48797 & ~w48884;
assign w48886 = ~w48825 & ~w48885;
assign w48887 = ~w48881 & w48886;
assign w48888 = ~w48854 & w48887;
assign w48889 = ~w48874 & w48888;
assign w48890 = pi2596 & ~w48889;
assign w48891 = ~pi2596 & w48889;
assign w48892 = ~w48890 & ~w48891;
assign w48893 = ~pi5538 & pi9040;
assign w48894 = ~pi5533 & ~pi9040;
assign w48895 = ~w48893 & ~w48894;
assign w48896 = pi2561 & ~w48895;
assign w48897 = ~pi2561 & w48895;
assign w48898 = ~w48896 & ~w48897;
assign w48899 = ~pi5740 & pi9040;
assign w48900 = ~pi5794 & ~pi9040;
assign w48901 = ~w48899 & ~w48900;
assign w48902 = pi2557 & ~w48901;
assign w48903 = ~pi2557 & w48901;
assign w48904 = ~w48902 & ~w48903;
assign w48905 = w48898 & ~w48904;
assign w48906 = ~pi5606 & pi9040;
assign w48907 = ~pi5616 & ~pi9040;
assign w48908 = ~w48906 & ~w48907;
assign w48909 = pi2566 & ~w48908;
assign w48910 = ~pi2566 & w48908;
assign w48911 = ~w48909 & ~w48910;
assign w48912 = ~w48905 & ~w48911;
assign w48913 = ~pi5631 & pi9040;
assign w48914 = ~pi5454 & ~pi9040;
assign w48915 = ~w48913 & ~w48914;
assign w48916 = pi2587 & ~w48915;
assign w48917 = ~pi2587 & w48915;
assign w48918 = ~w48916 & ~w48917;
assign w48919 = w48904 & w48918;
assign w48920 = ~w48898 & w48904;
assign w48921 = ~w48919 & ~w48920;
assign w48922 = ~pi5616 & pi9040;
assign w48923 = ~pi5536 & ~pi9040;
assign w48924 = ~w48922 & ~w48923;
assign w48925 = pi2583 & ~w48924;
assign w48926 = ~pi2583 & w48924;
assign w48927 = ~w48925 & ~w48926;
assign w48928 = w48921 & w48927;
assign w48929 = ~w48904 & ~w48918;
assign w48930 = ~w48898 & w48919;
assign w48931 = ~w48929 & ~w48930;
assign w48932 = ~pi5549 & pi9040;
assign w48933 = ~pi5809 & ~pi9040;
assign w48934 = ~w48932 & ~w48933;
assign w48935 = pi2571 & ~w48934;
assign w48936 = ~pi2571 & w48934;
assign w48937 = ~w48935 & ~w48936;
assign w48938 = ~w48898 & ~w48918;
assign w48939 = w48927 & w48938;
assign w48940 = ~w48937 & ~w48939;
assign w48941 = w48931 & w48940;
assign w48942 = ~w48928 & ~w48941;
assign w48943 = w48912 & ~w48942;
assign w48944 = w48918 & w48927;
assign w48945 = ~w48904 & w48944;
assign w48946 = w48944 & w66736;
assign w48947 = ~w48918 & w48927;
assign w48948 = ~w48905 & ~w48929;
assign w48949 = ~w48947 & ~w48948;
assign w48950 = ~w48948 & w66737;
assign w48951 = w48898 & w48918;
assign w48952 = ~w48938 & ~w48951;
assign w48953 = w48904 & ~w48952;
assign w48954 = w48898 & w48929;
assign w48955 = ~w48953 & ~w48954;
assign w48956 = ~w48927 & w48954;
assign w48957 = w48911 & ~w48956;
assign w48958 = ~w48955 & w48957;
assign w48959 = (~w48911 & ~w48919) | (~w48911 & w64044) | (~w48919 & w64044);
assign w48960 = w48904 & ~w48927;
assign w48961 = ~w48959 & w48960;
assign w48962 = w48937 & ~w48946;
assign w48963 = ~w48950 & w48962;
assign w48964 = ~w48961 & w48963;
assign w48965 = ~w48958 & w48964;
assign w48966 = w48921 & w66738;
assign w48967 = ~w48937 & ~w48966;
assign w48968 = w48904 & w48944;
assign w48969 = ~w48898 & w48968;
assign w48970 = w48967 & ~w48969;
assign w48971 = ~w48904 & w48939;
assign w48972 = w48911 & w48949;
assign w48973 = ~w48971 & ~w48972;
assign w48974 = w48970 & w48973;
assign w48975 = ~w48965 & ~w48974;
assign w48976 = ~w48943 & ~w48975;
assign w48977 = ~pi2601 & w48976;
assign w48978 = pi2601 & ~w48976;
assign w48979 = ~w48977 & ~w48978;
assign w48980 = ~pi5936 & pi9040;
assign w48981 = ~pi5453 & ~pi9040;
assign w48982 = ~w48980 & ~w48981;
assign w48983 = pi2590 & ~w48982;
assign w48984 = ~pi2590 & w48982;
assign w48985 = ~w48983 & ~w48984;
assign w48986 = ~pi5540 & pi9040;
assign w48987 = ~pi5734 & ~pi9040;
assign w48988 = ~w48986 & ~w48987;
assign w48989 = pi2584 & ~w48988;
assign w48990 = ~pi2584 & w48988;
assign w48991 = ~w48989 & ~w48990;
assign w48992 = ~pi5734 & pi9040;
assign w48993 = ~pi5548 & ~pi9040;
assign w48994 = ~w48992 & ~w48993;
assign w48995 = pi2564 & ~w48994;
assign w48996 = ~pi2564 & w48994;
assign w48997 = ~w48995 & ~w48996;
assign w48998 = w48991 & ~w48997;
assign w48999 = ~pi5452 & pi9040;
assign w49000 = ~pi5535 & ~pi9040;
assign w49001 = ~w48999 & ~w49000;
assign w49002 = pi2579 & ~w49001;
assign w49003 = ~pi2579 & w49001;
assign w49004 = ~w49002 & ~w49003;
assign w49005 = ~pi5809 & pi9040;
assign w49006 = ~pi5455 & ~pi9040;
assign w49007 = ~w49005 & ~w49006;
assign w49008 = pi2580 & ~w49007;
assign w49009 = ~pi2580 & w49007;
assign w49010 = ~w49008 & ~w49009;
assign w49011 = ~w49004 & w49010;
assign w49012 = w48998 & w49011;
assign w49013 = ~w48985 & ~w49012;
assign w49014 = ~w48997 & ~w49010;
assign w49015 = ~w49004 & w49014;
assign w49016 = w48997 & ~w49010;
assign w49017 = w49004 & w49016;
assign w49018 = ~w49015 & ~w49017;
assign w49019 = ~w48991 & ~w49018;
assign w49020 = w48991 & ~w49004;
assign w49021 = w49016 & w49020;
assign w49022 = w48985 & ~w49021;
assign w49023 = ~w49019 & w49022;
assign w49024 = ~w49013 & ~w49023;
assign w49025 = w48991 & ~w49010;
assign w49026 = w48985 & w48997;
assign w49027 = w49025 & w49026;
assign w49028 = ~w48985 & ~w48991;
assign w49029 = w49014 & w49028;
assign w49030 = w49004 & w49029;
assign w49031 = ~w48991 & w49010;
assign w49032 = ~w48997 & ~w49028;
assign w49033 = w49031 & w49032;
assign w49034 = ~w48991 & w48997;
assign w49035 = ~w48998 & ~w49034;
assign w49036 = ~w48985 & ~w49035;
assign w49037 = ~w49004 & w49036;
assign w49038 = w48997 & w49010;
assign w49039 = w49004 & ~w49038;
assign w49040 = ~w48997 & w49010;
assign w49041 = ~w49004 & ~w49040;
assign w49042 = ~w49039 & ~w49041;
assign w49043 = w48991 & w49042;
assign w49044 = ~pi5670 & pi9040;
assign w49045 = ~pi5733 & ~pi9040;
assign w49046 = ~w49044 & ~w49045;
assign w49047 = pi2581 & ~w49046;
assign w49048 = ~pi2581 & w49046;
assign w49049 = ~w49047 & ~w49048;
assign w49050 = ~w49027 & w49049;
assign w49051 = ~w49030 & w49050;
assign w49052 = ~w49033 & w49051;
assign w49053 = ~w49037 & ~w49043;
assign w49054 = w49052 & w49053;
assign w49055 = w49035 & w49039;
assign w49056 = w49014 & ~w49020;
assign w49057 = ~w49055 & w49056;
assign w49058 = ~w49049 & ~w49057;
assign w49059 = w48985 & w49004;
assign w49060 = w48998 & w49059;
assign w49061 = w49011 & w49034;
assign w49062 = ~w49017 & ~w49031;
assign w49063 = ~w48985 & ~w49062;
assign w49064 = w48985 & ~w49040;
assign w49065 = ~w49025 & ~w49034;
assign w49066 = w49064 & w49065;
assign w49067 = ~w49060 & ~w49061;
assign w49068 = ~w49066 & w49067;
assign w49069 = ~w49063 & w49068;
assign w49070 = w49058 & w49069;
assign w49071 = ~w49054 & ~w49070;
assign w49072 = ~w49024 & ~w49071;
assign w49073 = ~pi2592 & w49072;
assign w49074 = pi2592 & ~w49072;
assign w49075 = ~w49073 & ~w49074;
assign w49076 = w48985 & w49011;
assign w49077 = ~w49035 & w49076;
assign w49078 = ~w49011 & ~w49025;
assign w49079 = w49032 & w49078;
assign w49080 = ~w49020 & ~w49079;
assign w49081 = ~w48985 & ~w49021;
assign w49082 = ~w49080 & w49081;
assign w49083 = w49016 & w49081;
assign w49084 = (w49041 & w49082) | (w49041 & w66739) | (w49082 & w66739);
assign w49085 = w49028 & ~w49061;
assign w49086 = ~w49042 & w49085;
assign w49087 = w48991 & ~w49040;
assign w49088 = w49059 & w49087;
assign w49089 = ~w49004 & w49034;
assign w49090 = ~w49012 & ~w49049;
assign w49091 = ~w49027 & ~w49089;
assign w49092 = w49090 & w49091;
assign w49093 = ~w49088 & w49092;
assign w49094 = ~w49086 & w49093;
assign w49095 = ~w49018 & w49025;
assign w49096 = w49013 & w49042;
assign w49097 = w49049 & ~w49079;
assign w49098 = ~w49095 & w49097;
assign w49099 = ~w49096 & w49098;
assign w49100 = ~w49094 & ~w49099;
assign w49101 = ~w49077 & ~w49084;
assign w49102 = ~w49100 & w49101;
assign w49103 = pi2593 & w49102;
assign w49104 = ~pi2593 & ~w49102;
assign w49105 = ~w49103 & ~w49104;
assign w49106 = w48905 & w48927;
assign w49107 = ~w48898 & ~w48927;
assign w49108 = ~w48911 & w49107;
assign w49109 = ~w49106 & ~w49108;
assign w49110 = w48918 & ~w49109;
assign w49111 = (w48937 & w49109) | (w48937 & w66740) | (w49109 & w66740);
assign w49112 = ~w48911 & w48927;
assign w49113 = ~w48930 & w66741;
assign w49114 = ~w48920 & ~w48927;
assign w49115 = w48952 & w49114;
assign w49116 = ~w49113 & ~w49115;
assign w49117 = ~w49111 & ~w49116;
assign w49118 = w48911 & w48969;
assign w49119 = ~w49110 & ~w49118;
assign w49120 = ~w48937 & ~w49119;
assign w49121 = ~w48939 & ~w48960;
assign w49122 = w48911 & ~w48920;
assign w49123 = ~w49121 & w49122;
assign w49124 = ~w48931 & w49112;
assign w49125 = w48898 & w48911;
assign w49126 = ~w49106 & w49125;
assign w49127 = w48912 & w48929;
assign w49128 = ~w48952 & w48960;
assign w49129 = ~w49126 & ~w49127;
assign w49130 = ~w49128 & w49129;
assign w49131 = ~w49124 & w49130;
assign w49132 = w48937 & ~w49131;
assign w49133 = ~w49117 & ~w49123;
assign w49134 = ~w49120 & w49133;
assign w49135 = ~w49132 & w49134;
assign w49136 = pi2607 & ~w49135;
assign w49137 = ~pi2607 & w49135;
assign w49138 = ~w49136 & ~w49137;
assign w49139 = w48528 & w48546;
assign w49140 = (w48557 & w48549) | (w48557 & w66742) | (w48549 & w66742);
assign w49141 = ~w48536 & ~w48550;
assign w49142 = w48496 & ~w49141;
assign w49143 = ~w49139 & ~w49140;
assign w49144 = ~w49142 & w49143;
assign w49145 = w48490 & ~w49144;
assign w49146 = w48503 & ~w48714;
assign w49147 = ~w48532 & ~w48545;
assign w49148 = ~w48563 & w49147;
assign w49149 = w48516 & ~w49148;
assign w49150 = ~w49146 & ~w49149;
assign w49151 = ~w48490 & ~w49150;
assign w49152 = w48516 & ~w48750;
assign w49153 = w48517 & w48718;
assign w49154 = ~w49152 & ~w49153;
assign w49155 = ~w49145 & ~w49154;
assign w49156 = ~w49151 & w49155;
assign w49157 = ~pi2652 & w49156;
assign w49158 = pi2652 & ~w49156;
assign w49159 = ~w49157 & ~w49158;
assign w49160 = w48817 & w48865;
assign w49161 = (w48828 & w66743) | (w48828 & w66744) | (w66743 & w66744);
assign w49162 = ~w48824 & ~w48842;
assign w49163 = ~w48857 & w49162;
assign w49164 = (w48868 & ~w49162) | (w48868 & w66745) | (~w49162 & w66745);
assign w49165 = ~w48839 & ~w49161;
assign w49166 = (~w49160 & ~w49165) | (~w49160 & w66746) | (~w49165 & w66746);
assign w49167 = ~w48852 & ~w49166;
assign w49168 = ~w48803 & w48816;
assign w49169 = w48861 & w49168;
assign w49170 = (w48797 & w48838) | (w48797 & w64045) | (w48838 & w64045);
assign w49171 = ~w48810 & ~w48823;
assign w49172 = ~w48882 & ~w49171;
assign w49173 = w48839 & ~w49172;
assign w49174 = w48878 & ~w49170;
assign w49175 = ~w49173 & w49174;
assign w49176 = ~w48832 & ~w49169;
assign w49177 = (w49176 & w49175) | (w49176 & w66747) | (w49175 & w66747);
assign w49178 = ~w49167 & w49177;
assign w49179 = pi2600 & ~w49178;
assign w49180 = ~pi2600 & w49178;
assign w49181 = ~w49179 & ~w49180;
assign w49182 = ~w48816 & w48834;
assign w49183 = w48816 & w48865;
assign w49184 = w48797 & ~w49168;
assign w49185 = ~w49183 & ~w49184;
assign w49186 = w49162 & w49185;
assign w49187 = ~w48855 & ~w49186;
assign w49188 = w48816 & w49171;
assign w49189 = w48797 & w49188;
assign w49190 = ~w48852 & ~w49189;
assign w49191 = ~w48881 & w49190;
assign w49192 = w48841 & w48865;
assign w49193 = w48810 & ~w48840;
assign w49194 = ~w49184 & w49193;
assign w49195 = w48852 & ~w49192;
assign w49196 = ~w48877 & w49195;
assign w49197 = w48880 & ~w49194;
assign w49198 = w49196 & w49197;
assign w49199 = (~w49198 & ~w49191) | (~w49198 & w66748) | (~w49191 & w66748);
assign w49200 = ~w49182 & ~w49199;
assign w49201 = ~pi2609 & w49200;
assign w49202 = pi2609 & ~w49200;
assign w49203 = ~w49201 & ~w49202;
assign w49204 = w49004 & w49010;
assign w49205 = w49035 & w49204;
assign w49206 = w49014 & w66749;
assign w49207 = (~w48985 & ~w49035) | (~w48985 & w64046) | (~w49035 & w64046);
assign w49208 = ~w49206 & w49207;
assign w49209 = ~w49022 & ~w49208;
assign w49210 = w49011 & w66750;
assign w49211 = ~w48991 & ~w49011;
assign w49212 = w49026 & w49211;
assign w49213 = ~w49035 & w49064;
assign w49214 = ~w49011 & ~w49020;
assign w49215 = w48997 & ~w49214;
assign w49216 = ~w49213 & w49215;
assign w49217 = ~w49029 & ~w49210;
assign w49218 = ~w49212 & w49217;
assign w49219 = ~w49216 & w49218;
assign w49220 = w49058 & w49219;
assign w49221 = ~w49211 & w49213;
assign w49222 = ~w49205 & ~w49221;
assign w49223 = ~w48985 & w49012;
assign w49224 = w49049 & ~w49223;
assign w49225 = ~w49083 & w49224;
assign w49226 = w49222 & w49225;
assign w49227 = ~w49220 & ~w49226;
assign w49228 = ~w49060 & ~w49209;
assign w49229 = ~w49227 & w49228;
assign w49230 = pi2594 & ~w49229;
assign w49231 = ~pi2594 & w49229;
assign w49232 = ~w49230 & ~w49231;
assign w49233 = ~pi5539 & pi9040;
assign w49234 = ~pi5722 & ~pi9040;
assign w49235 = ~w49233 & ~w49234;
assign w49236 = pi2561 & ~w49235;
assign w49237 = ~pi2561 & w49235;
assign w49238 = ~w49236 & ~w49237;
assign w49239 = ~pi5624 & pi9040;
assign w49240 = ~pi5808 & ~pi9040;
assign w49241 = ~w49239 & ~w49240;
assign w49242 = pi2570 & ~w49241;
assign w49243 = ~pi2570 & w49241;
assign w49244 = ~w49242 & ~w49243;
assign w49245 = w49238 & ~w49244;
assign w49246 = ~pi5536 & pi9040;
assign w49247 = ~pi5539 & ~pi9040;
assign w49248 = ~w49246 & ~w49247;
assign w49249 = pi2586 & ~w49248;
assign w49250 = ~pi2586 & w49248;
assign w49251 = ~w49249 & ~w49250;
assign w49252 = w49245 & w49251;
assign w49253 = ~pi5455 & pi9040;
assign w49254 = ~pi5936 & ~pi9040;
assign w49255 = ~w49253 & ~w49254;
assign w49256 = pi2582 & ~w49255;
assign w49257 = ~pi2582 & w49255;
assign w49258 = ~w49256 & ~w49257;
assign w49259 = ~w49238 & ~w49258;
assign w49260 = ~pi5722 & pi9040;
assign w49261 = ~pi5609 & ~pi9040;
assign w49262 = ~w49260 & ~w49261;
assign w49263 = pi2575 & ~w49262;
assign w49264 = ~pi2575 & w49262;
assign w49265 = ~w49263 & ~w49264;
assign w49266 = ~w49244 & ~w49265;
assign w49267 = ~w49259 & w49266;
assign w49268 = w49244 & ~w49251;
assign w49269 = w49265 & w49268;
assign w49270 = ~w49267 & ~w49269;
assign w49271 = ~w49238 & ~w49265;
assign w49272 = w49251 & w49258;
assign w49273 = w49271 & w49272;
assign w49274 = w49244 & w49265;
assign w49275 = w49259 & w49274;
assign w49276 = ~w49251 & ~w49258;
assign w49277 = w49266 & w49276;
assign w49278 = ~w49275 & ~w49277;
assign w49279 = ~w49258 & ~w49268;
assign w49280 = w49238 & w49265;
assign w49281 = ~w49271 & ~w49280;
assign w49282 = w49279 & w49281;
assign w49283 = w49278 & w49282;
assign w49284 = w49270 & ~w49273;
assign w49285 = ~w49283 & w49284;
assign w49286 = ~pi5453 & pi9040;
assign w49287 = ~pi5631 & ~pi9040;
assign w49288 = ~w49286 & ~w49287;
assign w49289 = pi2557 & ~w49288;
assign w49290 = ~pi2557 & w49288;
assign w49291 = ~w49289 & ~w49290;
assign w49292 = (w49291 & ~w49285) | (w49291 & w66751) | (~w49285 & w66751);
assign w49293 = w49279 & w49280;
assign w49294 = w49258 & w49281;
assign w49295 = w49244 & w49251;
assign w49296 = w49281 & w64047;
assign w49297 = ~w49293 & ~w49296;
assign w49298 = ~w49244 & ~w49258;
assign w49299 = ~w49265 & ~w49298;
assign w49300 = w49259 & w49299;
assign w49301 = ~w49251 & ~w49280;
assign w49302 = w49244 & w49258;
assign w49303 = w49301 & ~w49302;
assign w49304 = w49285 & w49303;
assign w49305 = w49297 & ~w49300;
assign w49306 = (~w49291 & w49304) | (~w49291 & w66752) | (w49304 & w66752);
assign w49307 = ~w49238 & w49244;
assign w49308 = w49276 & w49307;
assign w49309 = w49238 & w49258;
assign w49310 = ~w49251 & w49309;
assign w49311 = w49244 & w49281;
assign w49312 = ~w49244 & ~w49281;
assign w49313 = ~w49311 & ~w49312;
assign w49314 = w49310 & w49313;
assign w49315 = ~w49244 & w49273;
assign w49316 = w49251 & w49265;
assign w49317 = w49298 & w49316;
assign w49318 = ~w49308 & ~w49317;
assign w49319 = ~w49315 & w49318;
assign w49320 = ~w49314 & w49319;
assign w49321 = ~w49292 & w49320;
assign w49322 = ~w49306 & w49321;
assign w49323 = ~pi2597 & w49322;
assign w49324 = pi2597 & ~w49322;
assign w49325 = ~w49323 & ~w49324;
assign w49326 = ~pi5742 & pi9040;
assign w49327 = ~pi5464 & ~pi9040;
assign w49328 = ~w49326 & ~w49327;
assign w49329 = pi2560 & ~w49328;
assign w49330 = ~pi2560 & w49328;
assign w49331 = ~w49329 & ~w49330;
assign w49332 = ~pi5626 & pi9040;
assign w49333 = ~pi5634 & ~pi9040;
assign w49334 = ~w49332 & ~w49333;
assign w49335 = pi2585 & ~w49334;
assign w49336 = ~pi2585 & w49334;
assign w49337 = ~w49335 & ~w49336;
assign w49338 = ~pi5687 & pi9040;
assign w49339 = ~pi5541 & ~pi9040;
assign w49340 = ~w49338 & ~w49339;
assign w49341 = pi2580 & ~w49340;
assign w49342 = ~pi2580 & w49340;
assign w49343 = ~w49341 & ~w49342;
assign w49344 = ~w49337 & ~w49343;
assign w49345 = ~pi5619 & pi9040;
assign w49346 = ~pi5459 & ~pi9040;
assign w49347 = ~w49345 & ~w49346;
assign w49348 = pi2581 & ~w49347;
assign w49349 = ~pi2581 & w49347;
assign w49350 = ~w49348 & ~w49349;
assign w49351 = w49344 & ~w49350;
assign w49352 = ~w49337 & w49350;
assign w49353 = w49343 & w49352;
assign w49354 = ~w49351 & ~w49353;
assign w49355 = ~pi5530 & pi9040;
assign w49356 = ~pi5878 & ~pi9040;
assign w49357 = ~w49355 & ~w49356;
assign w49358 = pi2591 & ~w49357;
assign w49359 = ~pi2591 & w49357;
assign w49360 = ~w49358 & ~w49359;
assign w49361 = ~w49354 & w49360;
assign w49362 = w49337 & ~w49360;
assign w49363 = ~w49350 & w49362;
assign w49364 = ~w49343 & ~w49352;
assign w49365 = w49337 & w49343;
assign w49366 = w49350 & ~w49365;
assign w49367 = w49364 & w49366;
assign w49368 = ~pi5633 & pi9040;
assign w49369 = ~pi5562 & ~pi9040;
assign w49370 = ~w49368 & ~w49369;
assign w49371 = pi2548 & ~w49370;
assign w49372 = ~pi2548 & w49370;
assign w49373 = ~w49371 & ~w49372;
assign w49374 = (~w49373 & w49367) | (~w49373 & w66753) | (w49367 & w66753);
assign w49375 = w49350 & w49373;
assign w49376 = w49337 & w49373;
assign w49377 = ~w49350 & ~w49376;
assign w49378 = (w49365 & w49377) | (w49365 & w66754) | (w49377 & w66754);
assign w49379 = w49343 & ~w49360;
assign w49380 = w49350 & w49360;
assign w49381 = ~w49337 & ~w49379;
assign w49382 = ~w49380 & w49381;
assign w49383 = w49375 & w49382;
assign w49384 = ~w49361 & ~w49378;
assign w49385 = w49384 & w66755;
assign w49386 = ~w49331 & ~w49385;
assign w49387 = ~w49350 & w49360;
assign w49388 = ~w49344 & ~w49365;
assign w49389 = w49387 & w49388;
assign w49390 = (w49373 & ~w49362) | (w49373 & w49375) | (~w49362 & w49375);
assign w49391 = w49364 & ~w49387;
assign w49392 = w49390 & w49391;
assign w49393 = (w49331 & w49392) | (w49331 & w66756) | (w49392 & w66756);
assign w49394 = w49331 & ~w49376;
assign w49395 = ~w49350 & w49379;
assign w49396 = ~w49394 & w49395;
assign w49397 = w49344 & w49380;
assign w49398 = w49350 & ~w49360;
assign w49399 = w49331 & w49398;
assign w49400 = ~w49397 & ~w49399;
assign w49401 = ~w49373 & ~w49400;
assign w49402 = w49337 & w49380;
assign w49403 = (w49373 & ~w49379) | (w49373 & w49375) | (~w49379 & w49375);
assign w49404 = ~w49402 & w49403;
assign w49405 = ~w49351 & w49404;
assign w49406 = w49360 & w49388;
assign w49407 = w49405 & w49406;
assign w49408 = ~w49396 & ~w49401;
assign w49409 = ~w49393 & w49408;
assign w49410 = ~w49407 & w49409;
assign w49411 = ~w49386 & w49410;
assign w49412 = pi2604 & ~w49411;
assign w49413 = ~pi2604 & w49411;
assign w49414 = ~w49412 & ~w49413;
assign w49415 = ~w48939 & w48959;
assign w49416 = ~w48918 & w49107;
assign w49417 = ~w48945 & ~w49416;
assign w49418 = w48911 & w49417;
assign w49419 = ~w49415 & ~w49418;
assign w49420 = w48951 & w48960;
assign w49421 = ~w48966 & ~w49420;
assign w49422 = ~w48956 & ~w49110;
assign w49423 = ~w49419 & w49422;
assign w49424 = (w48937 & ~w49423) | (w48937 & w64048) | (~w49423 & w64048);
assign w49425 = (~w48954 & w49417) | (~w48954 & w66757) | (w49417 & w66757);
assign w49426 = ~w48937 & ~w49425;
assign w49427 = w49421 & ~w49426;
assign w49428 = ~w48911 & ~w49427;
assign w49429 = ~w48912 & ~w48954;
assign w49430 = ~w48945 & ~w49128;
assign w49431 = w49429 & w49430;
assign w49432 = w48967 & w49431;
assign w49433 = ~w49424 & ~w49432;
assign w49434 = w49433 & w66758;
assign w49435 = (~pi2615 & ~w49433) | (~pi2615 & w66759) | (~w49433 & w66759);
assign w49436 = ~w49434 & ~w49435;
assign w49437 = ~pi5808 & pi9040;
assign w49438 = ~pi5540 & ~pi9040;
assign w49439 = ~w49437 & ~w49438;
assign w49440 = pi2564 & ~w49439;
assign w49441 = ~pi2564 & w49439;
assign w49442 = ~w49440 & ~w49441;
assign w49443 = ~pi5454 & pi9040;
assign w49444 = ~pi5538 & ~pi9040;
assign w49445 = ~w49443 & ~w49444;
assign w49446 = pi2587 & ~w49445;
assign w49447 = ~pi2587 & w49445;
assign w49448 = ~w49446 & ~w49447;
assign w49449 = ~pi5609 & pi9040;
assign w49450 = ~pi5668 & ~pi9040;
assign w49451 = ~w49449 & ~w49450;
assign w49452 = pi2571 & ~w49451;
assign w49453 = ~pi2571 & w49451;
assign w49454 = ~w49452 & ~w49453;
assign w49455 = ~pi5535 & pi9040;
assign w49456 = ~pi5624 & ~pi9040;
assign w49457 = ~w49455 & ~w49456;
assign w49458 = pi2584 & ~w49457;
assign w49459 = ~pi2584 & w49457;
assign w49460 = ~w49458 & ~w49459;
assign w49461 = w49454 & ~w49460;
assign w49462 = ~w49448 & w49461;
assign w49463 = w49454 & w49460;
assign w49464 = w49448 & w49463;
assign w49465 = ~w49462 & ~w49464;
assign w49466 = ~w49454 & ~w49460;
assign w49467 = ~pi5794 & pi9040;
assign w49468 = ~pi5549 & ~pi9040;
assign w49469 = ~w49467 & ~w49468;
assign w49470 = pi2565 & ~w49469;
assign w49471 = ~pi2565 & w49469;
assign w49472 = ~w49470 & ~w49471;
assign w49473 = w49466 & w49472;
assign w49474 = ~w49454 & ~w49472;
assign w49475 = w49460 & w49474;
assign w49476 = ~w49473 & ~w49475;
assign w49477 = w49454 & w49472;
assign w49478 = ~w49448 & w49477;
assign w49479 = w49448 & ~w49460;
assign w49480 = ~w49454 & w49479;
assign w49481 = ~w49478 & ~w49480;
assign w49482 = w49476 & w49481;
assign w49483 = w49482 & w63431;
assign w49484 = ~w49477 & ~w49479;
assign w49485 = ~w49448 & ~w49454;
assign w49486 = ~pi5668 & pi9040;
assign w49487 = ~pi5670 & ~pi9040;
assign w49488 = ~w49486 & ~w49487;
assign w49489 = pi2558 & ~w49488;
assign w49490 = ~pi2558 & w49488;
assign w49491 = ~w49489 & ~w49490;
assign w49492 = ~w49485 & ~w49491;
assign w49493 = w49484 & w49492;
assign w49494 = (~w49442 & w49483) | (~w49442 & w64049) | (w49483 & w64049);
assign w49495 = w49460 & ~w49491;
assign w49496 = w49485 & w49495;
assign w49497 = ~w49462 & ~w49496;
assign w49498 = ~w49472 & ~w49497;
assign w49499 = (w49442 & w49498) | (w49442 & w66760) | (w49498 & w66760);
assign w49500 = w49448 & w49472;
assign w49501 = ~w49454 & w49500;
assign w49502 = (w49501 & w49494) | (w49501 & w66761) | (w49494 & w66761);
assign w49503 = (~w49485 & ~w49465) | (~w49485 & w64050) | (~w49465 & w64050);
assign w49504 = w49442 & ~w49491;
assign w49505 = w49503 & w49504;
assign w49506 = w49448 & w49491;
assign w49507 = w49474 & w49506;
assign w49508 = w49461 & w49500;
assign w49509 = ~w49454 & w49460;
assign w49510 = ~w49500 & ~w49509;
assign w49511 = ~w49448 & ~w49472;
assign w49512 = ~w49461 & ~w49511;
assign w49513 = w49510 & w49512;
assign w49514 = ~w49507 & ~w49508;
assign w49515 = ~w49513 & w49514;
assign w49516 = ~w49498 & w49515;
assign w49517 = ~w49442 & ~w49516;
assign w49518 = w49466 & w49511;
assign w49519 = ~w49448 & w49460;
assign w49520 = w49472 & w49519;
assign w49521 = w49442 & ~w49466;
assign w49522 = ~w49518 & ~w49520;
assign w49523 = (w49522 & w49503) | (w49522 & w66762) | (w49503 & w66762);
assign w49524 = w49491 & ~w49523;
assign w49525 = ~w49505 & ~w49517;
assign w49526 = ~w49524 & w49525;
assign w49527 = (pi2618 & ~w49526) | (pi2618 & w66763) | (~w49526 & w66763);
assign w49528 = w49526 & w66764;
assign w49529 = ~w49527 & ~w49528;
assign w49530 = ~w49491 & ~w49509;
assign w49531 = ~w49464 & ~w49474;
assign w49532 = w49530 & ~w49531;
assign w49533 = w49500 & w49532;
assign w49534 = ~w49511 & ~w49530;
assign w49535 = w49482 & w63432;
assign w49536 = (~w49491 & ~w49477) | (~w49491 & w64051) | (~w49477 & w64051);
assign w49537 = ~w49495 & ~w49536;
assign w49538 = ~w49482 & w49537;
assign w49539 = ~w49535 & ~w49538;
assign w49540 = w49491 & ~w49510;
assign w49541 = w49476 & w49540;
assign w49542 = (w49539 & w66765) | (w49539 & w66766) | (w66765 & w66766);
assign w49543 = ~w49442 & ~w49539;
assign w49544 = w49491 & ~w49509;
assign w49545 = w49511 & w49544;
assign w49546 = ~w49507 & ~w49545;
assign w49547 = w49503 & ~w49546;
assign w49548 = ~w49533 & ~w49547;
assign w49549 = ~w49543 & w49548;
assign w49550 = (pi2620 & ~w49549) | (pi2620 & w66767) | (~w49549 & w66767);
assign w49551 = w49549 & w66768;
assign w49552 = ~w49550 & ~w49551;
assign w49553 = ~w48832 & ~w48834;
assign w49554 = (~w49171 & ~w49553) | (~w49171 & w66769) | (~w49553 & w66769);
assign w49555 = w48804 & ~w49554;
assign w49556 = w48878 & w49163;
assign w49557 = w48810 & w48835;
assign w49558 = w49556 & w49557;
assign w49559 = w48830 & w48861;
assign w49560 = ~w48883 & ~w49183;
assign w49561 = (w48852 & ~w49560) | (w48852 & w66770) | (~w49560 & w66770);
assign w49562 = ~w49160 & ~w49188;
assign w49563 = ~w48797 & ~w49562;
assign w49564 = w49161 & ~w49556;
assign w49565 = w49553 & ~w49563;
assign w49566 = (~w48852 & w49564) | (~w48852 & w66771) | (w49564 & w66771);
assign w49567 = ~w49164 & ~w49561;
assign w49568 = ~w49555 & w49567;
assign w49569 = ~w49558 & w49568;
assign w49570 = ~w49566 & w49569;
assign w49571 = pi2608 & ~w49570;
assign w49572 = ~pi2608 & w49570;
assign w49573 = ~w49571 & ~w49572;
assign w49574 = ~w49270 & ~w49278;
assign w49575 = w49280 & w49298;
assign w49576 = ~w49299 & ~w49575;
assign w49577 = w49251 & ~w49576;
assign w49578 = w49297 & ~w49577;
assign w49579 = ~w49313 & ~w49578;
assign w49580 = ~w49251 & ~w49274;
assign w49581 = ~w49251 & w49258;
assign w49582 = w49265 & w49581;
assign w49583 = w49245 & ~w49582;
assign w49584 = ~w49298 & ~w49309;
assign w49585 = ~w49583 & ~w49584;
assign w49586 = w49313 & w49580;
assign w49587 = ~w49585 & w49586;
assign w49588 = ~w49579 & ~w49587;
assign w49589 = w49291 & ~w49588;
assign w49590 = w49291 & ~w49310;
assign w49591 = ~w49300 & w49590;
assign w49592 = ~w49576 & w66772;
assign w49593 = w49271 & w49295;
assign w49594 = ~w49269 & ~w49593;
assign w49595 = ~w49592 & w49594;
assign w49596 = ~w49591 & ~w49595;
assign w49597 = ~w49291 & w49585;
assign w49598 = ~w49317 & ~w49574;
assign w49599 = ~w49597 & w49598;
assign w49600 = ~w49596 & w49599;
assign w49601 = (pi2611 & w49589) | (pi2611 & w66773) | (w49589 & w66773);
assign w49602 = ~w49589 & w66774;
assign w49603 = ~w49601 & ~w49602;
assign w49604 = ~w49463 & w49500;
assign w49605 = w49442 & ~w49519;
assign w49606 = ~w49484 & ~w49604;
assign w49607 = ~w49605 & w49606;
assign w49608 = ~w49499 & ~w49607;
assign w49609 = w49491 & ~w49608;
assign w49610 = ~w49477 & ~w49480;
assign w49611 = w49504 & ~w49610;
assign w49612 = ~w49460 & ~w49491;
assign w49613 = ~w49442 & ~w49612;
assign w49614 = w49604 & ~w49613;
assign w49615 = ~w49611 & ~w49614;
assign w49616 = ~w49494 & w49615;
assign w49617 = ~w49609 & w49616;
assign w49618 = pi2621 & ~w49617;
assign w49619 = ~pi2621 & w49617;
assign w49620 = ~w49618 & ~w49619;
assign w49621 = ~w49343 & ~w49373;
assign w49622 = w49380 & w49621;
assign w49623 = w49388 & w49398;
assign w49624 = ~w49352 & w64053;
assign w49625 = ~w49623 & w66775;
assign w49626 = (~w49354 & w64054) | (~w49354 & w64055) | (w64054 & w64055);
assign w49627 = ~w49367 & w63434;
assign w49628 = w49343 & ~w49350;
assign w49629 = ~w49366 & ~w49628;
assign w49630 = (w49373 & w49366) | (w49373 & w63435) | (w49366 & w63435);
assign w49631 = ~w49382 & w49630;
assign w49632 = ~w49627 & ~w49631;
assign w49633 = ~w49626 & ~w49632;
assign w49634 = ~w49337 & w49373;
assign w49635 = (w49634 & w49623) | (w49634 & w64056) | (w49623 & w64056);
assign w49636 = ~w49628 & ~w49635;
assign w49637 = (~w49625 & ~w49633) | (~w49625 & w64057) | (~w49633 & w64057);
assign w49638 = ~w49331 & ~w49637;
assign w49639 = (w49331 & w49632) | (w49331 & w66776) | (w49632 & w66776);
assign w49640 = w49361 & w49373;
assign w49641 = w49362 & ~w49621;
assign w49642 = w49629 & w49641;
assign w49643 = ~w49622 & ~w49642;
assign w49644 = ~w49640 & w49643;
assign w49645 = ~w49639 & w49644;
assign w49646 = (pi2606 & w49638) | (pi2606 & w66777) | (w49638 & w66777);
assign w49647 = ~w49638 & w66778;
assign w49648 = ~w49646 & ~w49647;
assign w49649 = ~w49373 & w49389;
assign w49650 = ~w49388 & ~w49398;
assign w49651 = ~w49623 & ~w49650;
assign w49652 = ~w49373 & ~w49651;
assign w49653 = (~w49331 & w49652) | (~w49331 & w66779) | (w49652 & w66779);
assign w49654 = ~w49344 & ~w49404;
assign w49655 = ~w49382 & ~w49654;
assign w49656 = ~w49360 & ~w49373;
assign w49657 = ~w49388 & w66780;
assign w49658 = ~w49367 & w66781;
assign w49659 = w49331 & ~w49623;
assign w49660 = ~w49657 & w49659;
assign w49661 = ~w49658 & w49660;
assign w49662 = ~w49655 & w49661;
assign w49663 = ~w49635 & ~w49649;
assign w49664 = (w49663 & w49662) | (w49663 & w66782) | (w49662 & w66782);
assign w49665 = ~pi2612 & w49664;
assign w49666 = pi2612 & ~w49664;
assign w49667 = ~w49665 & ~w49666;
assign w49668 = (w49059 & w49221) | (w49059 & w66783) | (w49221 & w66783);
assign w49669 = (~w49015 & w49018) | (~w49015 & w66784) | (w49018 & w66784);
assign w49670 = w48985 & ~w49669;
assign w49671 = ~w49031 & ~w49089;
assign w49672 = w49036 & ~w49671;
assign w49673 = (~w49021 & ~w49042) | (~w49021 & w66785) | (~w49042 & w66785);
assign w49674 = ~w49672 & w49673;
assign w49675 = ~w49670 & w49674;
assign w49676 = ~w49049 & ~w49675;
assign w49677 = (~w49049 & ~w49207) | (~w49049 & w66786) | (~w49207 & w66786);
assign w49678 = w49055 & ~w49677;
assign w49679 = w48985 & ~w49671;
assign w49680 = (w49049 & w49082) | (w49049 & w66787) | (w49082 & w66787);
assign w49681 = ~w49668 & ~w49678;
assign w49682 = ~w49680 & w49681;
assign w49683 = ~w49676 & w49682;
assign w49684 = ~pi2599 & ~w49683;
assign w49685 = pi2599 & w49683;
assign w49686 = ~w49684 & ~w49685;
assign w49687 = ~w48911 & ~w49429;
assign w49688 = w48957 & ~w48968;
assign w49689 = ~w49687 & ~w49688;
assign w49690 = w48952 & w49122;
assign w49691 = ~w48911 & ~w48944;
assign w49692 = ~w48921 & w49691;
assign w49693 = w48937 & ~w48971;
assign w49694 = ~w49690 & ~w49692;
assign w49695 = w49693 & w49694;
assign w49696 = w48898 & w49112;
assign w49697 = ~w49107 & ~w49696;
assign w49698 = ~w48904 & ~w49697;
assign w49699 = w48919 & w49125;
assign w49700 = ~w49416 & ~w49699;
assign w49701 = ~w49698 & w49700;
assign w49702 = w48970 & w49701;
assign w49703 = ~w49695 & ~w49702;
assign w49704 = ~w49689 & ~w49703;
assign w49705 = ~pi2635 & w49704;
assign w49706 = pi2635 & ~w49704;
assign w49707 = ~w49705 & ~w49706;
assign w49708 = ~w49285 & w49295;
assign w49709 = ~w49281 & ~w49302;
assign w49710 = w49580 & w49709;
assign w49711 = ~w49245 & ~w49307;
assign w49712 = w49316 & w49711;
assign w49713 = w49294 & ~w49711;
assign w49714 = ~w49291 & ~w49712;
assign w49715 = ~w49710 & w49714;
assign w49716 = ~w49713 & w49715;
assign w49717 = w49238 & w49302;
assign w49718 = w49291 & ~w49717;
assign w49719 = w49278 & ~w49582;
assign w49720 = w49718 & w49719;
assign w49721 = ~w49577 & w49720;
assign w49722 = ~w49716 & ~w49721;
assign w49723 = ~w49708 & ~w49722;
assign w49724 = ~pi2602 & w49723;
assign w49725 = pi2602 & ~w49723;
assign w49726 = ~w49724 & ~w49725;
assign w49727 = w49500 & w49509;
assign w49728 = w49466 & ~w49506;
assign w49729 = ~w49466 & ~w49485;
assign w49730 = w49465 & w49729;
assign w49731 = ~w49472 & ~w49728;
assign w49732 = ~w49730 & w49731;
assign w49733 = ~w49474 & ~w49477;
assign w49734 = w49612 & w49733;
assign w49735 = w49442 & ~w49727;
assign w49736 = ~w49734 & w49735;
assign w49737 = ~w49732 & w49736;
assign w49738 = w49491 & w49730;
assign w49739 = ~w49442 & ~w49496;
assign w49740 = ~w49518 & w49739;
assign w49741 = ~w49532 & w49740;
assign w49742 = ~w49738 & w49741;
assign w49743 = ~w49737 & ~w49742;
assign w49744 = ~w49448 & w49473;
assign w49745 = w49491 & ~w49508;
assign w49746 = ~w49744 & w49745;
assign w49747 = ~w49536 & ~w49746;
assign w49748 = ~w49743 & ~w49747;
assign w49749 = ~pi2627 & w49748;
assign w49750 = pi2627 & ~w49748;
assign w49751 = ~w49749 & ~w49750;
assign w49752 = w49265 & w49296;
assign w49753 = w49301 & w49711;
assign w49754 = ~w49259 & ~w49298;
assign w49755 = w49709 & w49754;
assign w49756 = ~w49252 & ~w49593;
assign w49757 = ~w49753 & w49756;
assign w49758 = ~w49755 & w49757;
assign w49759 = ~w49752 & w49758;
assign w49760 = ~w49269 & w49718;
assign w49761 = ~w49759 & ~w49760;
assign w49762 = w49258 & ~w49313;
assign w49763 = (~w49258 & ~w49758) | (~w49258 & w66788) | (~w49758 & w66788);
assign w49764 = w49291 & ~w49762;
assign w49765 = ~w49763 & w49764;
assign w49766 = ~w49761 & ~w49765;
assign w49767 = ~pi2595 & w49766;
assign w49768 = pi2595 & ~w49766;
assign w49769 = ~w49767 & ~w49768;
assign w49770 = w49405 & w66789;
assign w49771 = ~w49365 & ~w49630;
assign w49772 = w49350 & w49362;
assign w49773 = ~w49377 & ~w49772;
assign w49774 = (~w49397 & w49771) | (~w49397 & w66790) | (w49771 & w66790);
assign w49775 = w49331 & ~w49774;
assign w49776 = ~w49353 & w49390;
assign w49777 = ~w49352 & ~w49362;
assign w49778 = ~w49367 & w64058;
assign w49779 = (~w49624 & w49778) | (~w49624 & w66791) | (w49778 & w66791);
assign w49780 = ~w49331 & ~w49779;
assign w49781 = w49354 & ~w49360;
assign w49782 = ~w49374 & ~w49656;
assign w49783 = ~w49781 & ~w49782;
assign w49784 = ~w49383 & ~w49770;
assign w49785 = ~w49783 & w49784;
assign w49786 = ~w49775 & ~w49780;
assign w49787 = w49785 & w49786;
assign w49788 = pi2622 & ~w49787;
assign w49789 = ~pi2622 & w49787;
assign w49790 = ~w49788 & ~w49789;
assign w49791 = ~pi5737 & pi9040;
assign w49792 = ~pi5873 & ~pi9040;
assign w49793 = ~w49791 & ~w49792;
assign w49794 = pi2639 & ~w49793;
assign w49795 = ~pi2639 & w49793;
assign w49796 = ~w49794 & ~w49795;
assign w49797 = ~pi5810 & pi9040;
assign w49798 = ~pi6011 & ~pi9040;
assign w49799 = ~w49797 & ~w49798;
assign w49800 = pi2645 & ~w49799;
assign w49801 = ~pi2645 & w49799;
assign w49802 = ~w49800 & ~w49801;
assign w49803 = w49796 & w49802;
assign w49804 = ~w49796 & ~w49802;
assign w49805 = ~w49803 & ~w49804;
assign w49806 = ~pi5849 & pi9040;
assign w49807 = ~pi5781 & ~pi9040;
assign w49808 = ~w49806 & ~w49807;
assign w49809 = pi2631 & ~w49808;
assign w49810 = ~pi2631 & w49808;
assign w49811 = ~w49809 & ~w49810;
assign w49812 = ~pi6011 & pi9040;
assign w49813 = ~pi5932 & ~pi9040;
assign w49814 = ~w49812 & ~w49813;
assign w49815 = pi2640 & ~w49814;
assign w49816 = ~pi2640 & w49814;
assign w49817 = ~w49815 & ~w49816;
assign w49818 = ~w49811 & ~w49817;
assign w49819 = ~pi5811 & pi9040;
assign w49820 = ~pi5910 & ~pi9040;
assign w49821 = ~w49819 & ~w49820;
assign w49822 = pi2613 & ~w49821;
assign w49823 = ~pi2613 & w49821;
assign w49824 = ~w49822 & ~w49823;
assign w49825 = ~w49796 & w49824;
assign w49826 = ~w49802 & ~w49824;
assign w49827 = ~w49825 & ~w49826;
assign w49828 = w49818 & w49827;
assign w49829 = ~w49796 & ~w49824;
assign w49830 = ~w49811 & ~w49829;
assign w49831 = ~w49828 & w49830;
assign w49832 = ~w49805 & w49831;
assign w49833 = w49811 & ~w49824;
assign w49834 = ~w49805 & w49833;
assign w49835 = w49802 & w49811;
assign w49836 = w49825 & w49835;
assign w49837 = w49817 & ~w49836;
assign w49838 = ~w49834 & w49837;
assign w49839 = ~w49802 & ~w49811;
assign w49840 = w49825 & w49839;
assign w49841 = w49796 & w49824;
assign w49842 = ~w49833 & ~w49841;
assign w49843 = w49802 & ~w49842;
assign w49844 = w49817 & ~w49840;
assign w49845 = ~w49843 & w49844;
assign w49846 = ~w49804 & w49845;
assign w49847 = w49838 & ~w49846;
assign w49848 = ~pi5934 & pi9040;
assign w49849 = ~pi6018 & ~pi9040;
assign w49850 = ~w49848 & ~w49849;
assign w49851 = pi2649 & ~w49850;
assign w49852 = ~pi2649 & w49850;
assign w49853 = ~w49851 & ~w49852;
assign w49854 = w49811 & w49841;
assign w49855 = (~w49817 & ~w49841) | (~w49817 & w49818) | (~w49841 & w49818);
assign w49856 = w49836 & w49855;
assign w49857 = ~w49802 & ~w49829;
assign w49858 = w49833 & w49857;
assign w49859 = (~w49853 & ~w49827) | (~w49853 & w66792) | (~w49827 & w66792);
assign w49860 = ~w49858 & w49859;
assign w49861 = ~w49856 & w49860;
assign w49862 = ~w49847 & w49861;
assign w49863 = w49818 & w49825;
assign w49864 = w49841 & w66793;
assign w49865 = ~w49863 & ~w49864;
assign w49866 = w49802 & ~w49811;
assign w49867 = w49829 & ~w49866;
assign w49868 = w49855 & ~w49867;
assign w49869 = w49803 & ~w49824;
assign w49870 = w49829 & w49866;
assign w49871 = ~w49869 & ~w49870;
assign w49872 = w49837 & w49871;
assign w49873 = ~w49868 & ~w49872;
assign w49874 = w49796 & ~w49811;
assign w49875 = w49826 & w49874;
assign w49876 = ~w49834 & ~w49875;
assign w49877 = ~w49802 & ~w49876;
assign w49878 = w49853 & w49865;
assign w49879 = ~w49873 & w49878;
assign w49880 = ~w49877 & w49879;
assign w49881 = ~w49862 & ~w49880;
assign w49882 = ~w49881 & w66794;
assign w49883 = (pi2669 & w49881) | (pi2669 & w66795) | (w49881 & w66795);
assign w49884 = ~w49882 & ~w49883;
assign w49885 = ~w49817 & ~w49824;
assign w49886 = ~w49854 & ~w49885;
assign w49887 = ~w49805 & ~w49886;
assign w49888 = w49824 & w49866;
assign w49889 = w49817 & ~w49826;
assign w49890 = ~w49869 & w49889;
assign w49891 = ~w49888 & w49890;
assign w49892 = ~w49887 & ~w49891;
assign w49893 = ~w49853 & ~w49892;
assign w49894 = w49817 & w49824;
assign w49895 = ~w49885 & ~w49894;
assign w49896 = w49805 & w49895;
assign w49897 = w49831 & w49896;
assign w49898 = w49818 & w49841;
assign w49899 = ~w49802 & w49898;
assign w49900 = w49796 & ~w49894;
assign w49901 = w49866 & ~w49900;
assign w49902 = w49857 & w49895;
assign w49903 = ~w49901 & ~w49902;
assign w49904 = w49876 & w49903;
assign w49905 = w49853 & ~w49904;
assign w49906 = ~w49897 & ~w49899;
assign w49907 = ~w49893 & w49906;
assign w49908 = ~w49905 & w49907;
assign w49909 = pi2670 & ~w49908;
assign w49910 = ~pi2670 & w49908;
assign w49911 = ~w49909 & ~w49910;
assign w49912 = ~pi5745 & pi9040;
assign w49913 = ~pi5727 & ~pi9040;
assign w49914 = ~w49912 & ~w49913;
assign w49915 = pi2613 & ~w49914;
assign w49916 = ~pi2613 & w49914;
assign w49917 = ~w49915 & ~w49916;
assign w49918 = ~pi5727 & pi9040;
assign w49919 = ~pi5814 & ~pi9040;
assign w49920 = ~w49918 & ~w49919;
assign w49921 = pi2625 & ~w49920;
assign w49922 = ~pi2625 & w49920;
assign w49923 = ~w49921 & ~w49922;
assign w49924 = ~pi5812 & pi9040;
assign w49925 = ~pi6158 & ~pi9040;
assign w49926 = ~w49924 & ~w49925;
assign w49927 = pi2654 & ~w49926;
assign w49928 = ~pi2654 & w49926;
assign w49929 = ~w49927 & ~w49928;
assign w49930 = w49923 & ~w49929;
assign w49931 = ~pi6037 & pi9040;
assign w49932 = ~pi5791 & ~pi9040;
assign w49933 = ~w49931 & ~w49932;
assign w49934 = pi2634 & ~w49933;
assign w49935 = ~pi2634 & w49933;
assign w49936 = ~w49934 & ~w49935;
assign w49937 = ~pi5879 & pi9040;
assign w49938 = ~pi5747 & ~pi9040;
assign w49939 = ~w49937 & ~w49938;
assign w49940 = pi2645 & ~w49939;
assign w49941 = ~pi2645 & w49939;
assign w49942 = ~w49940 & ~w49941;
assign w49943 = ~pi5944 & pi9040;
assign w49944 = ~pi5891 & ~pi9040;
assign w49945 = ~w49943 & ~w49944;
assign w49946 = pi2651 & ~w49945;
assign w49947 = ~pi2651 & w49945;
assign w49948 = ~w49946 & ~w49947;
assign w49949 = w49942 & w49948;
assign w49950 = ~w49923 & w49949;
assign w49951 = ~w49936 & ~w49950;
assign w49952 = ~w49923 & w49948;
assign w49953 = w49923 & ~w49948;
assign w49954 = ~w49952 & ~w49953;
assign w49955 = w49951 & ~w49954;
assign w49956 = w49942 & ~w49948;
assign w49957 = w49923 & w49956;
assign w49958 = ~w49955 & ~w49957;
assign w49959 = ~w49936 & ~w49948;
assign w49960 = ~w49929 & ~w49959;
assign w49961 = ~w49923 & ~w49948;
assign w49962 = ~w49942 & w49961;
assign w49963 = (w49936 & ~w49961) | (w49936 & w64059) | (~w49961 & w64059);
assign w49964 = w49960 & ~w49963;
assign w49965 = w49936 & w49950;
assign w49966 = ~w49964 & ~w49965;
assign w49967 = w49923 & w49949;
assign w49968 = ~w49929 & ~w49942;
assign w49969 = w49952 & w49968;
assign w49970 = w49936 & ~w49969;
assign w49971 = ~w49967 & w49970;
assign w49972 = w49929 & ~w49942;
assign w49973 = ~w49961 & ~w49972;
assign w49974 = ~w49948 & ~w49973;
assign w49975 = w49971 & ~w49974;
assign w49976 = ~w49929 & w49953;
assign w49977 = ~w49950 & ~w49976;
assign w49978 = ~w49936 & w49977;
assign w49979 = ~w49942 & w49948;
assign w49980 = ~w49929 & w49942;
assign w49981 = ~w49979 & ~w49980;
assign w49982 = w49923 & ~w49968;
assign w49983 = ~w49981 & w49982;
assign w49984 = (~w49983 & w49975) | (~w49983 & w63436) | (w49975 & w63436);
assign w49985 = ~w49929 & w49966;
assign w49986 = w49984 & w49985;
assign w49987 = (~w49917 & w49986) | (~w49917 & w64060) | (w49986 & w64060);
assign w49988 = w49949 & w49930;
assign w49989 = w49917 & ~w49984;
assign w49990 = w49929 & w49948;
assign w49991 = ~w49936 & w49990;
assign w49992 = w49956 & w49960;
assign w49993 = ~w49991 & ~w49992;
assign w49994 = ~w49923 & ~w49993;
assign w49995 = w49954 & w49972;
assign w49996 = w49936 & w49995;
assign w49997 = ~w49988 & ~w49996;
assign w49998 = ~w49994 & w49997;
assign w49999 = ~w49989 & w49998;
assign w50000 = ~w49987 & w49999;
assign w50001 = pi2671 & ~w50000;
assign w50002 = ~pi2671 & w50000;
assign w50003 = ~w50001 & ~w50002;
assign w50004 = ~w49811 & ~w49894;
assign w50005 = ~w49803 & ~w49874;
assign w50006 = ~w50004 & ~w50005;
assign w50007 = ~w49840 & ~w49898;
assign w50008 = ~w49818 & ~w49870;
assign w50009 = w50007 & ~w50008;
assign w50010 = ~w50006 & ~w50009;
assign w50011 = w49853 & ~w50010;
assign w50012 = w49824 & ~w49839;
assign w50013 = w49805 & w50012;
assign w50014 = ~w49830 & ~w50013;
assign w50015 = ~w50013 & w66796;
assign w50016 = ~w49817 & ~w50015;
assign w50017 = ~w49838 & ~w50016;
assign w50018 = w49845 & ~w50006;
assign w50019 = ~w49839 & w49885;
assign w50020 = w49805 & w50019;
assign w50021 = w50007 & ~w50020;
assign w50022 = (w50021 & ~w50018) | (w50021 & w66797) | (~w50018 & w66797);
assign w50023 = ~w49853 & ~w50022;
assign w50024 = ~w50011 & ~w50017;
assign w50025 = ~w50023 & w50024;
assign w50026 = ~pi2679 & w50025;
assign w50027 = pi2679 & ~w50025;
assign w50028 = ~w50026 & ~w50027;
assign w50029 = w49818 & w49867;
assign w50030 = ~w49900 & ~w50004;
assign w50031 = w49845 & ~w50030;
assign w50032 = w49802 & w49833;
assign w50033 = ~w49888 & ~w50032;
assign w50034 = ~w49817 & ~w50033;
assign w50035 = w49811 & ~w49817;
assign w50036 = ~w49835 & ~w49874;
assign w50037 = ~w50035 & w50036;
assign w50038 = w50012 & w50037;
assign w50039 = w49865 & ~w50034;
assign w50040 = ~w50038 & w50039;
assign w50041 = (~w49853 & ~w50040) | (~w49853 & w66798) | (~w50040 & w66798);
assign w50042 = w49827 & w50035;
assign w50043 = w49818 & ~w49869;
assign w50044 = ~w49899 & w50043;
assign w50045 = w49853 & ~w50042;
assign w50046 = ~w49845 & w50045;
assign w50047 = ~w50044 & w50046;
assign w50048 = ~w49854 & ~w49870;
assign w50049 = w49817 & ~w50048;
assign w50050 = ~w50029 & ~w50049;
assign w50051 = ~w49897 & w50050;
assign w50052 = ~w50047 & w50051;
assign w50053 = ~w50041 & w50052;
assign w50054 = pi2677 & ~w50053;
assign w50055 = ~pi2677 & w50053;
assign w50056 = ~w50054 & ~w50055;
assign w50057 = ~pi5862 & pi9040;
assign w50058 = ~pi5732 & ~pi9040;
assign w50059 = ~w50057 & ~w50058;
assign w50060 = pi2639 & ~w50059;
assign w50061 = ~pi2639 & w50059;
assign w50062 = ~w50060 & ~w50061;
assign w50063 = ~pi5873 & pi9040;
assign w50064 = ~pi5811 & ~pi9040;
assign w50065 = ~w50063 & ~w50064;
assign w50066 = pi2629 & ~w50065;
assign w50067 = ~pi2629 & w50065;
assign w50068 = ~w50066 & ~w50067;
assign w50069 = ~w50062 & ~w50068;
assign w50070 = ~pi5871 & pi9040;
assign w50071 = ~pi5804 & ~pi9040;
assign w50072 = ~w50070 & ~w50071;
assign w50073 = pi2610 & ~w50072;
assign w50074 = ~pi2610 & w50072;
assign w50075 = ~w50073 & ~w50074;
assign w50076 = ~pi5804 & pi9040;
assign w50077 = ~pi5862 & ~pi9040;
assign w50078 = ~w50076 & ~w50077;
assign w50079 = pi2649 & ~w50078;
assign w50080 = ~pi2649 & w50078;
assign w50081 = ~w50079 & ~w50080;
assign w50082 = w50075 & w50081;
assign w50083 = w50062 & w50068;
assign w50084 = ~w50069 & ~w50083;
assign w50085 = ~w50082 & w50084;
assign w50086 = w50075 & w50085;
assign w50087 = ~w50069 & ~w50086;
assign w50088 = ~pi5781 & pi9040;
assign w50089 = ~pi5934 & ~pi9040;
assign w50090 = ~w50088 & ~w50089;
assign w50091 = pi2653 & ~w50090;
assign w50092 = ~pi2653 & w50090;
assign w50093 = ~w50091 & ~w50092;
assign w50094 = w50069 & ~w50081;
assign w50095 = w50069 & w66799;
assign w50096 = w50093 & ~w50095;
assign w50097 = ~w50087 & w50096;
assign w50098 = ~w50075 & ~w50081;
assign w50099 = ~w50082 & ~w50098;
assign w50100 = w50062 & ~w50093;
assign w50101 = ~w50099 & w50100;
assign w50102 = ~w50068 & ~w50081;
assign w50103 = w50062 & w50102;
assign w50104 = (~w50093 & ~w50102) | (~w50093 & w66800) | (~w50102 & w66800);
assign w50105 = ~w50083 & w50104;
assign w50106 = ~w50095 & ~w50100;
assign w50107 = w50105 & ~w50106;
assign w50108 = ~pi5725 & pi9040;
assign w50109 = ~pi5871 & ~pi9040;
assign w50110 = ~w50108 & ~w50109;
assign w50111 = pi2638 & ~w50110;
assign w50112 = ~pi2638 & w50110;
assign w50113 = ~w50111 & ~w50112;
assign w50114 = ~w50062 & ~w50075;
assign w50115 = w50081 & w50093;
assign w50116 = w50069 & w50099;
assign w50117 = ~w50115 & ~w50116;
assign w50118 = w50114 & ~w50117;
assign w50119 = ~w50062 & w50093;
assign w50120 = w50068 & ~w50119;
assign w50121 = ~w50099 & w50120;
assign w50122 = ~w50113 & ~w50121;
assign w50123 = ~w50107 & w50122;
assign w50124 = ~w50118 & w50123;
assign w50125 = w50069 & w50098;
assign w50126 = ~w50062 & w50075;
assign w50127 = ~w50075 & w50083;
assign w50128 = ~w50126 & ~w50127;
assign w50129 = w50115 & ~w50128;
assign w50130 = w50068 & ~w50081;
assign w50131 = w50126 & w50130;
assign w50132 = w50068 & w50081;
assign w50133 = w50084 & w66801;
assign w50134 = (~w50130 & ~w50084) | (~w50130 & w66802) | (~w50084 & w66802);
assign w50135 = ~w50133 & ~w50134;
assign w50136 = ~w50093 & w50135;
assign w50137 = w50113 & ~w50125;
assign w50138 = ~w50131 & w50137;
assign w50139 = ~w50129 & w50138;
assign w50140 = ~w50136 & w50139;
assign w50141 = ~w50124 & ~w50140;
assign w50142 = ~w50097 & ~w50101;
assign w50143 = ~w50141 & w50142;
assign w50144 = pi2656 & ~w50143;
assign w50145 = ~pi2656 & w50143;
assign w50146 = ~w50144 & ~w50145;
assign w50147 = ~pi5800 & pi9040;
assign w50148 = ~pi5951 & ~pi9040;
assign w50149 = ~w50147 & ~w50148;
assign w50150 = pi2643 & ~w50149;
assign w50151 = ~pi2643 & w50149;
assign w50152 = ~w50150 & ~w50151;
assign w50153 = ~pi6002 & pi9040;
assign w50154 = ~pi5746 & ~pi9040;
assign w50155 = ~w50153 & ~w50154;
assign w50156 = pi2655 & ~w50155;
assign w50157 = ~pi2655 & w50155;
assign w50158 = ~w50156 & ~w50157;
assign w50159 = w50152 & w50158;
assign w50160 = ~pi5741 & pi9040;
assign w50161 = ~pi5884 & ~pi9040;
assign w50162 = ~w50160 & ~w50161;
assign w50163 = pi2644 & ~w50162;
assign w50164 = ~pi2644 & w50162;
assign w50165 = ~w50163 & ~w50164;
assign w50166 = ~pi6146 & pi9040;
assign w50167 = ~pi5799 & ~pi9040;
assign w50168 = ~w50166 & ~w50167;
assign w50169 = pi2637 & ~w50168;
assign w50170 = ~pi2637 & w50168;
assign w50171 = ~w50169 & ~w50170;
assign w50172 = ~pi5881 & pi9040;
assign w50173 = ~pi5800 & ~pi9040;
assign w50174 = ~w50172 & ~w50173;
assign w50175 = pi2625 & ~w50174;
assign w50176 = ~pi2625 & w50174;
assign w50177 = ~w50175 & ~w50176;
assign w50178 = ~w50171 & w50177;
assign w50179 = w50152 & w50178;
assign w50180 = w50178 & w50191;
assign w50181 = ~w50171 & ~w50177;
assign w50182 = w50158 & w50178;
assign w50183 = (~w50152 & ~w50178) | (~w50152 & w66803) | (~w50178 & w66803);
assign w50184 = ~w50181 & ~w50183;
assign w50185 = w50152 & ~w50171;
assign w50186 = ~w50152 & w50171;
assign w50187 = ~w50185 & ~w50186;
assign w50188 = w50171 & w50177;
assign w50189 = w50165 & ~w50188;
assign w50190 = w50187 & w50189;
assign w50191 = w50152 & ~w50165;
assign w50192 = w50171 & ~w50177;
assign w50193 = w50191 & ~w50192;
assign w50194 = ~w50179 & ~w50193;
assign w50195 = ~w50158 & w50194;
assign w50196 = ~w50165 & w50186;
assign w50197 = ~w50152 & w50177;
assign w50198 = w50158 & ~w50197;
assign w50199 = ~w50196 & w50198;
assign w50200 = (~w50190 & w50195) | (~w50190 & w64061) | (w50195 & w64061);
assign w50201 = ~w50152 & w50158;
assign w50202 = ~w50191 & ~w50201;
assign w50203 = ~w50184 & ~w50202;
assign w50204 = w50200 & w50203;
assign w50205 = (~w50180 & ~w50200) | (~w50180 & w66804) | (~w50200 & w66804);
assign w50206 = ~w50159 & ~w50205;
assign w50207 = w50159 & w50194;
assign w50208 = w50194 & w66805;
assign w50209 = ~w50165 & ~w50178;
assign w50210 = ~w50189 & ~w50209;
assign w50211 = w50152 & w50210;
assign w50212 = ~w50158 & ~w50197;
assign w50213 = w50190 & w50212;
assign w50214 = w50190 & w64062;
assign w50215 = ~w50152 & w50181;
assign w50216 = (w50158 & ~w50188) | (w50158 & w50201) | (~w50188 & w50201);
assign w50217 = ~w50215 & w50216;
assign w50218 = w50187 & w50217;
assign w50219 = ~pi5874 & pi9040;
assign w50220 = ~pi6028 & ~pi9040;
assign w50221 = ~w50219 & ~w50220;
assign w50222 = pi2651 & ~w50221;
assign w50223 = ~pi2651 & w50221;
assign w50224 = ~w50222 & ~w50223;
assign w50225 = ~w50158 & ~w50165;
assign w50226 = (w50224 & w50187) | (w50224 & w64063) | (w50187 & w64063);
assign w50227 = ~w50211 & w50226;
assign w50228 = w50227 & w66806;
assign w50229 = w50165 & w50192;
assign w50230 = w50212 & ~w50229;
assign w50231 = ~w50217 & ~w50230;
assign w50232 = w50186 & w64064;
assign w50233 = w50152 & w50181;
assign w50234 = w50181 & w66807;
assign w50235 = w50158 & w50165;
assign w50236 = w50185 & w50235;
assign w50237 = w50181 & w66808;
assign w50238 = ~w50224 & ~w50236;
assign w50239 = ~w50232 & w50238;
assign w50240 = ~w50234 & ~w50237;
assign w50241 = w50239 & w50240;
assign w50242 = ~w50231 & w50241;
assign w50243 = (~w50208 & w50228) | (~w50208 & w64065) | (w50228 & w64065);
assign w50244 = w50243 & w66809;
assign w50245 = (pi2663 & ~w50243) | (pi2663 & w66810) | (~w50243 & w66810);
assign w50246 = ~w50244 & ~w50245;
assign w50247 = ~pi5814 & pi9040;
assign w50248 = ~pi5725 & ~pi9040;
assign w50249 = ~w50247 & ~w50248;
assign w50250 = pi2647 & ~w50249;
assign w50251 = ~pi2647 & w50249;
assign w50252 = ~w50250 & ~w50251;
assign w50253 = ~pi5891 & pi9040;
assign w50254 = ~pi5849 & ~pi9040;
assign w50255 = ~w50253 & ~w50254;
assign w50256 = pi2638 & ~w50255;
assign w50257 = ~pi2638 & w50255;
assign w50258 = ~w50256 & ~w50257;
assign w50259 = ~pi5791 & pi9040;
assign w50260 = ~pi5745 & ~pi9040;
assign w50261 = ~w50259 & ~w50260;
assign w50262 = pi2629 & ~w50261;
assign w50263 = ~pi2629 & w50261;
assign w50264 = ~w50262 & ~w50263;
assign w50265 = ~w50258 & w50264;
assign w50266 = ~pi5932 & pi9040;
assign w50267 = ~pi5879 & ~pi9040;
assign w50268 = ~w50266 & ~w50267;
assign w50269 = pi2650 & ~w50268;
assign w50270 = ~pi2650 & w50268;
assign w50271 = ~w50269 & ~w50270;
assign w50272 = ~pi5747 & pi9040;
assign w50273 = ~pi6037 & ~pi9040;
assign w50274 = ~w50272 & ~w50273;
assign w50275 = pi2626 & ~w50274;
assign w50276 = ~pi2626 & w50274;
assign w50277 = ~w50275 & ~w50276;
assign w50278 = w50271 & w50277;
assign w50279 = w50265 & w50278;
assign w50280 = w50258 & ~w50271;
assign w50281 = w50264 & ~w50277;
assign w50282 = ~w50280 & ~w50281;
assign w50283 = w50258 & w50281;
assign w50284 = ~w50258 & ~w50264;
assign w50285 = ~w50283 & ~w50284;
assign w50286 = ~w50264 & ~w50277;
assign w50287 = ~w50271 & ~w50277;
assign w50288 = w50265 & ~w50287;
assign w50289 = ~pi6158 & pi9040;
assign w50290 = ~pi5944 & ~pi9040;
assign w50291 = ~w50289 & ~w50290;
assign w50292 = pi2630 & ~w50291;
assign w50293 = ~pi2630 & w50291;
assign w50294 = ~w50292 & ~w50293;
assign w50295 = ~w50288 & w50294;
assign w50296 = w50258 & ~w50264;
assign w50297 = ~w50286 & ~w50296;
assign w50298 = w50295 & w50297;
assign w50299 = w50285 & w50298;
assign w50300 = (w50294 & ~w50287) | (w50294 & w50988) | (~w50287 & w50988);
assign w50301 = (~w50300 & ~w50298) | (~w50300 & w64066) | (~w50298 & w64066);
assign w50302 = w50258 & w50271;
assign w50303 = ~w50258 & ~w50271;
assign w50304 = ~w50302 & ~w50303;
assign w50305 = ~w50264 & ~w50294;
assign w50306 = ~w50304 & w50305;
assign w50307 = ~w50279 & ~w50306;
assign w50308 = (w50307 & w50301) | (w50307 & w66811) | (w50301 & w66811);
assign w50309 = w50252 & ~w50308;
assign w50310 = ~w50264 & w50271;
assign w50311 = ~w50281 & ~w50310;
assign w50312 = ~w50258 & w50311;
assign w50313 = ~w50283 & ~w50312;
assign w50314 = (~w50294 & w50312) | (~w50294 & w66812) | (w50312 & w66812);
assign w50315 = w50280 & w50314;
assign w50316 = ~w50278 & ~w50287;
assign w50317 = w50284 & ~w50316;
assign w50318 = w50264 & ~w50271;
assign w50319 = ~w50265 & ~w50277;
assign w50320 = ~w50318 & ~w50319;
assign w50321 = ~w50282 & w50320;
assign w50322 = (w50294 & w50321) | (w50294 & w66813) | (w50321 & w66813);
assign w50323 = w50280 & ~w50300;
assign w50324 = ~w50258 & ~w50277;
assign w50325 = w50271 & w50324;
assign w50326 = ~w50277 & ~w50294;
assign w50327 = ~w50305 & ~w50326;
assign w50328 = ~w50325 & ~w50327;
assign w50329 = w50286 & w50302;
assign w50330 = (w50294 & ~w50284) | (w50294 & w66814) | (~w50284 & w66814);
assign w50331 = ~w50329 & w50330;
assign w50332 = ~w50328 & ~w50331;
assign w50333 = w50264 & w50302;
assign w50334 = w50277 & w50333;
assign w50335 = ~w50323 & ~w50334;
assign w50336 = ~w50332 & w50335;
assign w50337 = ~w50252 & ~w50336;
assign w50338 = ~w50315 & ~w50322;
assign w50339 = ~w50337 & w50338;
assign w50340 = ~w50309 & w50339;
assign w50341 = pi2658 & ~w50340;
assign w50342 = ~pi2658 & w50340;
assign w50343 = ~w50341 & ~w50342;
assign w50344 = w50158 & ~w50232;
assign w50345 = ~w50180 & w50344;
assign w50346 = ~w50191 & w50192;
assign w50347 = ~w50193 & ~w50346;
assign w50348 = w50209 & ~w50347;
assign w50349 = ~w50158 & ~w50348;
assign w50350 = ~w50345 & ~w50349;
assign w50351 = w50195 & w50210;
assign w50352 = w50181 & ~w50202;
assign w50353 = w50184 & w50189;
assign w50354 = w50224 & ~w50352;
assign w50355 = ~w50351 & w66815;
assign w50356 = w50177 & w50187;
assign w50357 = w50187 & w66816;
assign w50358 = ~w50212 & ~w50357;
assign w50359 = w50183 & ~w50358;
assign w50360 = ~w50196 & ~w50224;
assign w50361 = ~w50180 & w50360;
assign w50362 = ~w50207 & w50361;
assign w50363 = ~w50359 & w50362;
assign w50364 = ~w50355 & ~w50363;
assign w50365 = ~w50350 & ~w50364;
assign w50366 = pi2660 & ~w50365;
assign w50367 = ~pi2660 & w50365;
assign w50368 = ~w50366 & ~w50367;
assign w50369 = ~w50075 & w50103;
assign w50370 = w50126 & w50132;
assign w50371 = ~w50085 & ~w50093;
assign w50372 = (w50093 & ~w50083) | (w50093 & w66817) | (~w50083 & w66817);
assign w50373 = w50130 & w50372;
assign w50374 = ~w50113 & ~w50370;
assign w50375 = ~w50116 & w50374;
assign w50376 = ~w50369 & w50375;
assign w50377 = ~w50371 & ~w50373;
assign w50378 = w50376 & w50377;
assign w50379 = ~w50075 & w50135;
assign w50380 = ~w50102 & ~w50132;
assign w50381 = ~w50068 & w50082;
assign w50382 = ~w50094 & ~w50381;
assign w50383 = w50372 & w50382;
assign w50384 = w50126 & w50380;
assign w50385 = ~w50383 & w50384;
assign w50386 = w50125 & w50372;
assign w50387 = ~w50086 & ~w50115;
assign w50388 = w50062 & ~w50387;
assign w50389 = w50113 & ~w50386;
assign w50390 = ~w50385 & w50389;
assign w50391 = ~w50379 & w50390;
assign w50392 = (~w50378 & ~w50391) | (~w50378 & w66818) | (~w50391 & w66818);
assign w50393 = ~pi2657 & w50392;
assign w50394 = pi2657 & ~w50392;
assign w50395 = ~w50393 & ~w50394;
assign w50396 = w50171 & ~w50201;
assign w50397 = ~w50189 & w50396;
assign w50398 = ~w50165 & ~w50346;
assign w50399 = w50397 & w50398;
assign w50400 = w50186 & w50344;
assign w50401 = ~w50182 & ~w50215;
assign w50402 = ~w50235 & ~w50401;
assign w50403 = ~w50234 & ~w50399;
assign w50404 = w50403 & w66819;
assign w50405 = ~w50224 & ~w50404;
assign w50406 = ~w50232 & ~w50233;
assign w50407 = w50158 & ~w50406;
assign w50408 = ~w50357 & ~w50407;
assign w50409 = (w50224 & w50407) | (w50224 & w66820) | (w50407 & w66820);
assign w50410 = ~w50180 & ~w50346;
assign w50411 = w50224 & ~w50410;
assign w50412 = ~w50237 & ~w50357;
assign w50413 = ~w50411 & w50412;
assign w50414 = ~w50158 & ~w50413;
assign w50415 = ~w50208 & ~w50236;
assign w50416 = ~w50409 & w50415;
assign w50417 = ~w50414 & w50416;
assign w50418 = ~w50405 & w50417;
assign w50419 = pi2664 & ~w50418;
assign w50420 = ~pi2664 & w50418;
assign w50421 = ~w50419 & ~w50420;
assign w50422 = w50062 & w50075;
assign w50423 = w50380 & w50422;
assign w50424 = ~w50370 & ~w50423;
assign w50425 = ~w50075 & ~w50380;
assign w50426 = ~w50113 & ~w50425;
assign w50427 = w50424 & w50426;
assign w50428 = w50096 & ~w50427;
assign w50429 = ~w50380 & w66821;
assign w50430 = ~w50095 & ~w50429;
assign w50431 = ~w50113 & ~w50430;
assign w50432 = ~w50093 & w50424;
assign w50433 = ~w50431 & w50432;
assign w50434 = ~w50428 & ~w50433;
assign w50435 = w50093 & w50429;
assign w50436 = ~w50062 & w50099;
assign w50437 = ~w50093 & ~w50132;
assign w50438 = ~w50369 & w50437;
assign w50439 = ~w50436 & w50438;
assign w50440 = w50424 & ~w50435;
assign w50441 = ~w50439 & w50440;
assign w50442 = w50113 & ~w50441;
assign w50443 = ~w50434 & ~w50442;
assign w50444 = ~pi2666 & w50443;
assign w50445 = pi2666 & ~w50443;
assign w50446 = ~w50444 & ~w50445;
assign w50447 = ~pi6045 & pi9040;
assign w50448 = ~pi5933 & ~pi9040;
assign w50449 = ~w50447 & ~w50448;
assign w50450 = pi2648 & ~w50449;
assign w50451 = ~pi2648 & w50449;
assign w50452 = ~w50450 & ~w50451;
assign w50453 = ~pi6016 & pi9040;
assign w50454 = ~pi5797 & ~pi9040;
assign w50455 = ~w50453 & ~w50454;
assign w50456 = pi2647 & ~w50455;
assign w50457 = ~pi2647 & w50455;
assign w50458 = ~w50456 & ~w50457;
assign w50459 = w50452 & w50458;
assign w50460 = ~pi5883 & pi9040;
assign w50461 = ~pi6146 & ~pi9040;
assign w50462 = ~w50460 & ~w50461;
assign w50463 = pi2633 & ~w50462;
assign w50464 = ~pi2633 & w50462;
assign w50465 = ~w50463 & ~w50464;
assign w50466 = ~pi5723 & pi9040;
assign w50467 = ~pi5807 & ~pi9040;
assign w50468 = ~w50466 & ~w50467;
assign w50469 = pi2626 & ~w50468;
assign w50470 = ~pi2626 & w50468;
assign w50471 = ~w50469 & ~w50470;
assign w50472 = ~w50465 & ~w50471;
assign w50473 = w50459 & w50472;
assign w50474 = ~pi5933 & pi9040;
assign w50475 = ~pi5743 & ~pi9040;
assign w50476 = ~w50474 & ~w50475;
assign w50477 = pi2632 & ~w50476;
assign w50478 = ~pi2632 & w50476;
assign w50479 = ~w50477 & ~w50478;
assign w50480 = w50458 & ~w50471;
assign w50481 = w50465 & ~w50480;
assign w50482 = ~w50458 & w50471;
assign w50483 = w50481 & ~w50482;
assign w50484 = ~pi5839 & pi9040;
assign w50485 = ~pi6036 & ~pi9040;
assign w50486 = ~w50484 & ~w50485;
assign w50487 = pi2624 & ~w50486;
assign w50488 = ~pi2624 & w50486;
assign w50489 = ~w50487 & ~w50488;
assign w50490 = w50458 & w50489;
assign w50491 = ~w50458 & ~w50489;
assign w50492 = ~w50490 & ~w50491;
assign w50493 = w50483 & w50492;
assign w50494 = w50483 & w66822;
assign w50495 = w50472 & w50490;
assign w50496 = ~w50494 & ~w50495;
assign w50497 = w50458 & ~w50465;
assign w50498 = ~w50481 & ~w50497;
assign w50499 = w50458 & w50471;
assign w50500 = ~w50452 & ~w50499;
assign w50501 = ~w50471 & w50489;
assign w50502 = w50471 & ~w50489;
assign w50503 = ~w50501 & ~w50502;
assign w50504 = w50500 & w50503;
assign w50505 = ~w50465 & w50502;
assign w50506 = ~w50504 & ~w50505;
assign w50507 = w50498 & ~w50506;
assign w50508 = w50452 & w50489;
assign w50509 = (w50508 & ~w50481) | (w50508 & w66823) | (~w50481 & w66823);
assign w50510 = ~w50498 & w50509;
assign w50511 = ~w50507 & ~w50510;
assign w50512 = (~w50479 & ~w50511) | (~w50479 & w66824) | (~w50511 & w66824);
assign w50513 = w50465 & ~w50489;
assign w50514 = w50452 & ~w50458;
assign w50515 = w50513 & w50514;
assign w50516 = ~w50480 & ~w50508;
assign w50517 = ~w50465 & ~w50490;
assign w50518 = ~w50516 & w50517;
assign w50519 = ~w50515 & ~w50518;
assign w50520 = ~w50452 & w50499;
assign w50521 = w50452 & w50501;
assign w50522 = w50472 & ~w50489;
assign w50523 = ~w50458 & ~w50471;
assign w50524 = ~w50522 & w50523;
assign w50525 = ~w50521 & ~w50524;
assign w50526 = ~w50518 & w66825;
assign w50527 = w50525 & w50526;
assign w50528 = w50479 & ~w50527;
assign w50529 = (~w50502 & ~w50481) | (~w50502 & w63331) | (~w50481 & w63331);
assign w50530 = ~w50513 & ~w50529;
assign w50531 = ~w50452 & w50530;
assign w50532 = ~w50471 & w50515;
assign w50533 = ~w50473 & ~w50532;
assign w50534 = ~w50531 & w50533;
assign w50535 = ~w50528 & w50534;
assign w50536 = ~w50512 & w50535;
assign w50537 = pi2661 & ~w50536;
assign w50538 = ~pi2661 & w50536;
assign w50539 = ~w50537 & ~w50538;
assign w50540 = ~w50356 & w50397;
assign w50541 = ~w50211 & ~w50540;
assign w50542 = (~w50224 & w50204) | (~w50224 & w66826) | (w50204 & w66826);
assign w50543 = w50235 & ~w50408;
assign w50544 = (~w50213 & w50200) | (~w50213 & w66827) | (w50200 & w66827);
assign w50545 = ~w50543 & w50544;
assign w50546 = ~w50542 & w50545;
assign w50547 = pi2678 & w50546;
assign w50548 = ~pi2678 & ~w50546;
assign w50549 = ~w50547 & ~w50548;
assign w50550 = w49952 & w49972;
assign w50551 = ~w49936 & w50550;
assign w50552 = ~w49923 & ~w49942;
assign w50553 = ~w49973 & ~w50552;
assign w50554 = w49981 & w50553;
assign w50555 = w49966 & ~w50554;
assign w50556 = w49917 & ~w50555;
assign w50557 = ~w49983 & ~w50554;
assign w50558 = ~w49923 & w49929;
assign w50559 = w49956 & ~w50558;
assign w50560 = w49951 & ~w50559;
assign w50561 = ~w49971 & ~w50560;
assign w50562 = ~w49976 & ~w49995;
assign w50563 = ~w50561 & w50562;
assign w50564 = ~w49917 & ~w50563;
assign w50565 = (~w50551 & w50557) | (~w50551 & w66828) | (w50557 & w66828);
assign w50566 = ~w50556 & w50565;
assign w50567 = ~w50564 & w50566;
assign w50568 = pi2673 & ~w50567;
assign w50569 = ~pi2673 & w50567;
assign w50570 = ~w50568 & ~w50569;
assign w50571 = w50465 & w50489;
assign w50572 = (~w50514 & w50524) | (~w50514 & w64067) | (w50524 & w64067);
assign w50573 = (~w50520 & w50572) | (~w50520 & w66829) | (w50572 & w66829);
assign w50574 = w50571 & ~w50573;
assign w50575 = w50502 & w50514;
assign w50576 = ~w50520 & ~w50575;
assign w50577 = (~w50479 & ~w50576) | (~w50479 & w66830) | (~w50576 & w66830);
assign w50578 = (w50517 & w50572) | (w50517 & w66831) | (w50572 & w66831);
assign w50579 = ~w50458 & ~w50503;
assign w50580 = w50480 & w50513;
assign w50581 = ~w50579 & ~w50580;
assign w50582 = (~w50452 & w50579) | (~w50452 & w66832) | (w50579 & w66832);
assign w50583 = ~w50458 & ~w50472;
assign w50584 = w50452 & w50503;
assign w50585 = w50583 & w50584;
assign w50586 = ~w50582 & ~w50585;
assign w50587 = w50496 & w50586;
assign w50588 = w50479 & ~w50587;
assign w50589 = ~w50473 & ~w50577;
assign w50590 = ~w50578 & w50589;
assign w50591 = ~w50574 & w50590;
assign w50592 = ~w50588 & w50591;
assign w50593 = pi2667 & ~w50592;
assign w50594 = ~pi2667 & w50592;
assign w50595 = ~w50593 & ~w50594;
assign w50596 = w50082 & w50083;
assign w50597 = w50114 & w50380;
assign w50598 = w50104 & ~w50597;
assign w50599 = ~w50597 & w66833;
assign w50600 = ~w50098 & w50133;
assign w50601 = ~w50083 & w50115;
assign w50602 = ~w50381 & w50601;
assign w50603 = ~w50596 & ~w50602;
assign w50604 = ~w50599 & w50603;
assign w50605 = ~w50600 & w50604;
assign w50606 = ~w50113 & ~w50605;
assign w50607 = w50093 & ~w50131;
assign w50608 = ~w50101 & ~w50607;
assign w50609 = ~w50105 & w50608;
assign w50610 = w50082 & w50084;
assign w50611 = w50598 & ~w50610;
assign w50612 = w50113 & ~w50383;
assign w50613 = ~w50611 & w50612;
assign w50614 = ~w50609 & ~w50613;
assign w50615 = ~w50606 & w50614;
assign w50616 = pi2665 & ~w50615;
assign w50617 = ~pi2665 & w50615;
assign w50618 = ~w50616 & ~w50617;
assign w50619 = ~pi5951 & pi9040;
assign w50620 = ~pi5723 & ~pi9040;
assign w50621 = ~w50619 & ~w50620;
assign w50622 = pi2616 & ~w50621;
assign w50623 = ~pi2616 & w50621;
assign w50624 = ~w50622 & ~w50623;
assign w50625 = ~pi5797 & pi9040;
assign w50626 = ~pi6045 & ~pi9040;
assign w50627 = ~w50625 & ~w50626;
assign w50628 = pi2636 & ~w50627;
assign w50629 = ~pi2636 & w50627;
assign w50630 = ~w50628 & ~w50629;
assign w50631 = ~w50624 & ~w50630;
assign w50632 = ~pi5803 & pi9040;
assign w50633 = ~pi6033 & ~pi9040;
assign w50634 = ~w50632 & ~w50633;
assign w50635 = pi2628 & ~w50634;
assign w50636 = ~pi2628 & w50634;
assign w50637 = ~w50635 & ~w50636;
assign w50638 = ~pi5844 & pi9040;
assign w50639 = ~pi5874 & ~pi9040;
assign w50640 = ~w50638 & ~w50639;
assign w50641 = pi2643 & ~w50640;
assign w50642 = ~pi2643 & w50640;
assign w50643 = ~w50641 & ~w50642;
assign w50644 = ~w50637 & ~w50643;
assign w50645 = w50637 & w50643;
assign w50646 = ~w50644 & ~w50645;
assign w50647 = w50631 & ~w50646;
assign w50648 = ~w50637 & w50643;
assign w50649 = w50624 & w50648;
assign w50650 = w50637 & ~w50643;
assign w50651 = w50630 & w50650;
assign w50652 = ~w50649 & ~w50651;
assign w50653 = ~w50647 & w50652;
assign w50654 = ~pi5801 & pi9040;
assign w50655 = ~pi5806 & ~pi9040;
assign w50656 = ~w50654 & ~w50655;
assign w50657 = pi2637 & ~w50656;
assign w50658 = ~pi2637 & w50656;
assign w50659 = ~w50657 & ~w50658;
assign w50660 = ~pi5884 & pi9040;
assign w50661 = ~pi5735 & ~pi9040;
assign w50662 = ~w50660 & ~w50661;
assign w50663 = pi2617 & ~w50662;
assign w50664 = ~pi2617 & w50662;
assign w50665 = ~w50663 & ~w50664;
assign w50666 = ~w50659 & ~w50665;
assign w50667 = ~w50653 & w50666;
assign w50668 = w50659 & w50665;
assign w50669 = w50649 & w50668;
assign w50670 = ~w50643 & ~w50665;
assign w50671 = ~w50650 & ~w50665;
assign w50672 = ~w50659 & ~w50671;
assign w50673 = w50624 & w50637;
assign w50674 = w50630 & w50673;
assign w50675 = ~w50670 & w50674;
assign w50676 = ~w50672 & w50675;
assign w50677 = ~w50648 & w50668;
assign w50678 = w50659 & ~w50665;
assign w50679 = ~w50647 & w50678;
assign w50680 = ~w50677 & ~w50679;
assign w50681 = ~w50646 & ~w50665;
assign w50682 = ~w50631 & ~w50681;
assign w50683 = ~w50680 & ~w50682;
assign w50684 = w50630 & w50644;
assign w50685 = ~w50673 & ~w50684;
assign w50686 = ~w50651 & w50685;
assign w50687 = w50685 & w66834;
assign w50688 = w50624 & w50630;
assign w50689 = ~w50631 & ~w50688;
assign w50690 = w50650 & ~w50689;
assign w50691 = ~w50624 & ~w50637;
assign w50692 = w50630 & w50665;
assign w50693 = w50691 & w50692;
assign w50694 = ~w50690 & ~w50693;
assign w50695 = w50687 & ~w50694;
assign w50696 = w50624 & ~w50643;
assign w50697 = ~w50624 & w50643;
assign w50698 = ~w50696 & ~w50697;
assign w50699 = ~w50637 & ~w50698;
assign w50700 = w50685 & ~w50699;
assign w50701 = w50670 & ~w50673;
assign w50702 = ~w50674 & ~w50701;
assign w50703 = w50672 & w50702;
assign w50704 = ~w50700 & w50703;
assign w50705 = ~w50669 & ~w50676;
assign w50706 = ~w50667 & w50705;
assign w50707 = ~w50704 & w50706;
assign w50708 = ~w50683 & ~w50695;
assign w50709 = w50707 & w50708;
assign w50710 = pi2688 & ~w50709;
assign w50711 = ~pi2688 & w50709;
assign w50712 = ~w50710 & ~w50711;
assign w50713 = ~w50630 & w50665;
assign w50714 = ~w50650 & w50713;
assign w50715 = w50698 & w50714;
assign w50716 = w50637 & w50715;
assign w50717 = ~w50695 & ~w50699;
assign w50718 = w50668 & ~w50717;
assign w50719 = ~w50630 & ~w50653;
assign w50720 = ~w50645 & w50688;
assign w50721 = w50665 & ~w50720;
assign w50722 = ~w50686 & w50721;
assign w50723 = ~w50719 & ~w50722;
assign w50724 = ~w50659 & ~w50723;
assign w50725 = ~w50630 & ~w50637;
assign w50726 = w50666 & ~w50725;
assign w50727 = w50686 & w50726;
assign w50728 = w50678 & ~w50685;
assign w50729 = ~w50659 & ~w50670;
assign w50730 = w50720 & ~w50729;
assign w50731 = ~w50716 & ~w50730;
assign w50732 = ~w50728 & w50731;
assign w50733 = ~w50727 & w50732;
assign w50734 = ~w50724 & w50733;
assign w50735 = w50734 & w66835;
assign w50736 = (pi2685 & ~w50734) | (pi2685 & w66836) | (~w50734 & w66836);
assign w50737 = ~w50735 & ~w50736;
assign w50738 = ~pi5743 & pi9040;
assign w50739 = ~pi5883 & ~pi9040;
assign w50740 = ~w50738 & ~w50739;
assign w50741 = pi2642 & ~w50740;
assign w50742 = ~pi2642 & w50740;
assign w50743 = ~w50741 & ~w50742;
assign w50744 = ~pi5806 & pi9040;
assign w50745 = ~pi5844 & ~pi9040;
assign w50746 = ~w50744 & ~w50745;
assign w50747 = pi2632 & ~w50746;
assign w50748 = ~pi2632 & w50746;
assign w50749 = ~w50747 & ~w50748;
assign w50750 = ~pi6036 & pi9040;
assign w50751 = ~pi5877 & ~pi9040;
assign w50752 = ~w50750 & ~w50751;
assign w50753 = pi2636 & ~w50752;
assign w50754 = ~pi2636 & w50752;
assign w50755 = ~w50753 & ~w50754;
assign w50756 = ~pi5877 & pi9040;
assign w50757 = ~pi6002 & ~pi9040;
assign w50758 = ~w50756 & ~w50757;
assign w50759 = pi2646 & ~w50758;
assign w50760 = ~pi2646 & w50758;
assign w50761 = ~w50759 & ~w50760;
assign w50762 = ~w50755 & w50761;
assign w50763 = ~pi6033 & pi9040;
assign w50764 = ~pi5839 & ~pi9040;
assign w50765 = ~w50763 & ~w50764;
assign w50766 = pi2624 & ~w50765;
assign w50767 = ~pi2624 & w50765;
assign w50768 = ~w50766 & ~w50767;
assign w50769 = w50755 & ~w50768;
assign w50770 = ~w50749 & ~w50762;
assign w50771 = ~w50769 & w50770;
assign w50772 = w50770 & w66837;
assign w50773 = ~w50749 & w50761;
assign w50774 = ~w50755 & ~w50768;
assign w50775 = w50773 & w50774;
assign w50776 = ~w50772 & ~w50775;
assign w50777 = ~pi5799 & pi9040;
assign w50778 = ~pi5801 & ~pi9040;
assign w50779 = ~w50777 & ~w50778;
assign w50780 = pi2628 & ~w50779;
assign w50781 = ~pi2628 & w50779;
assign w50782 = ~w50780 & ~w50781;
assign w50783 = w50749 & w50761;
assign w50784 = w50769 & w50783;
assign w50785 = ~w50755 & w50768;
assign w50786 = w50783 & w50785;
assign w50787 = ~w50782 & ~w50784;
assign w50788 = ~w50786 & w50787;
assign w50789 = w50776 & w50788;
assign w50790 = ~w50749 & w50769;
assign w50791 = w50769 & w50773;
assign w50792 = w50761 & ~w50774;
assign w50793 = w50749 & ~w50792;
assign w50794 = ~w50749 & w50768;
assign w50795 = w50762 & w50794;
assign w50796 = ~w50793 & ~w50795;
assign w50797 = w50743 & ~w50796;
assign w50798 = ~w50743 & w50771;
assign w50799 = w50749 & w50755;
assign w50800 = ~w50761 & ~w50768;
assign w50801 = w50743 & w50768;
assign w50802 = ~w50800 & ~w50801;
assign w50803 = w50799 & ~w50802;
assign w50804 = w50782 & ~w50791;
assign w50805 = ~w50803 & w50804;
assign w50806 = ~w50798 & w50805;
assign w50807 = ~w50797 & w50806;
assign w50808 = ~w50789 & ~w50807;
assign w50809 = w50774 & ~w50783;
assign w50810 = w50749 & w50809;
assign w50811 = w50749 & w50768;
assign w50812 = ~w50790 & ~w50811;
assign w50813 = ~w50810 & w50812;
assign w50814 = ~w50782 & ~w50813;
assign w50815 = ~w50768 & w50773;
assign w50816 = ~w50786 & ~w50815;
assign w50817 = ~w50814 & w50816;
assign w50818 = ~w50743 & ~w50817;
assign w50819 = ~w50808 & ~w50818;
assign w50820 = ~pi2659 & w50819;
assign w50821 = pi2659 & ~w50819;
assign w50822 = ~w50820 & ~w50821;
assign w50823 = ~w49936 & w50554;
assign w50824 = ~w49977 & w49981;
assign w50825 = w49942 & w49990;
assign w50826 = ~w49976 & ~w50825;
assign w50827 = w49963 & w50826;
assign w50828 = ~w49936 & ~w49969;
assign w50829 = ~w49988 & w50828;
assign w50830 = ~w50553 & w50829;
assign w50831 = (~w50824 & w50830) | (~w50824 & w64068) | (w50830 & w64068);
assign w50832 = ~w49917 & ~w50831;
assign w50833 = w49936 & ~w49956;
assign w50834 = ~w49990 & w50833;
assign w50835 = w49923 & w49936;
assign w50836 = w49979 & ~w50835;
assign w50837 = ~w49979 & ~w50558;
assign w50838 = ~w50836 & ~w50837;
assign w50839 = w50834 & w50838;
assign w50840 = ~w49930 & ~w50558;
assign w50841 = (w49979 & ~w50840) | (w49979 & w66838) | (~w50840 & w66838);
assign w50842 = w50840 & w66839;
assign w50843 = ~w49929 & ~w49936;
assign w50844 = ~w49957 & ~w49962;
assign w50845 = w50843 & ~w50844;
assign w50846 = w49942 & w50827;
assign w50847 = ~w50841 & ~w50842;
assign w50848 = ~w50845 & w50847;
assign w50849 = ~w50846 & w50848;
assign w50850 = w49917 & ~w50849;
assign w50851 = ~w50823 & ~w50839;
assign w50852 = ~w50832 & w50851;
assign w50853 = w50852 & w66840;
assign w50854 = (~pi2681 & ~w50852) | (~pi2681 & w66841) | (~w50852 & w66841);
assign w50855 = ~w50853 & ~w50854;
assign w50856 = ~w50530 & w50581;
assign w50857 = (w50856 & w64069) | (w50856 & w64070) | (w64069 & w64070);
assign w50858 = w50459 & w50503;
assign w50859 = ~w50479 & ~w50858;
assign w50860 = ~w50493 & w50859;
assign w50861 = ~w50857 & w50860;
assign w50862 = w50497 & w50502;
assign w50863 = ~w50495 & ~w50583;
assign w50864 = w50452 & ~w50863;
assign w50865 = w50471 & w50571;
assign w50866 = w50479 & ~w50865;
assign w50867 = ~w50452 & ~w50497;
assign w50868 = ~w50583 & w50867;
assign w50869 = ~w50862 & w50866;
assign w50870 = ~w50868 & w50869;
assign w50871 = ~w50864 & w50870;
assign w50872 = w50482 & ~w50519;
assign w50873 = (~w50872 & w50861) | (~w50872 & w66842) | (w50861 & w66842);
assign w50874 = ~pi2662 & w50873;
assign w50875 = pi2662 & ~w50873;
assign w50876 = ~w50874 & ~w50875;
assign w50877 = w50631 & w50644;
assign w50878 = w50630 & w50646;
assign w50879 = ~w50630 & w50643;
assign w50880 = w50637 & w50879;
assign w50881 = ~w50878 & ~w50880;
assign w50882 = (w50665 & w50878) | (w50665 & w66843) | (w50878 & w66843);
assign w50883 = w50671 & ~w50696;
assign w50884 = w50881 & w50883;
assign w50885 = ~w50659 & ~w50877;
assign w50886 = ~w50882 & w50885;
assign w50887 = ~w50884 & w50886;
assign w50888 = w50648 & w50688;
assign w50889 = ~w50690 & w66844;
assign w50890 = w50881 & ~w50889;
assign w50891 = ~w50691 & w50701;
assign w50892 = w50659 & ~w50888;
assign w50893 = ~w50891 & w50892;
assign w50894 = ~w50890 & w50893;
assign w50895 = ~w50887 & ~w50894;
assign w50896 = ~w50687 & ~w50882;
assign w50897 = w50696 & ~w50896;
assign w50898 = ~w50630 & ~w50665;
assign w50899 = w50673 & w50898;
assign w50900 = ~w50897 & ~w50899;
assign w50901 = ~w50895 & w50900;
assign w50902 = pi2696 & ~w50901;
assign w50903 = ~pi2696 & w50901;
assign w50904 = ~w50902 & ~w50903;
assign w50905 = ~w50749 & ~w50801;
assign w50906 = ~w50749 & w50755;
assign w50907 = w50761 & w50768;
assign w50908 = w50906 & w50907;
assign w50909 = ~w50743 & ~w50761;
assign w50910 = w50769 & w50909;
assign w50911 = ~w50908 & ~w50910;
assign w50912 = w50905 & ~w50911;
assign w50913 = w50749 & ~w50769;
assign w50914 = ~w50743 & w50761;
assign w50915 = ~w50906 & w50914;
assign w50916 = ~w50913 & w50915;
assign w50917 = ~w50773 & w50801;
assign w50918 = w50755 & ~w50761;
assign w50919 = w50811 & w50918;
assign w50920 = w50776 & w50809;
assign w50921 = w50782 & ~w50917;
assign w50922 = ~w50919 & w50921;
assign w50923 = ~w50916 & w50922;
assign w50924 = ~w50912 & w50923;
assign w50925 = ~w50920 & w50924;
assign w50926 = ~w50785 & ~w50790;
assign w50927 = ~w50761 & ~w50926;
assign w50928 = ~w50784 & ~w50915;
assign w50929 = ~w50916 & ~w50928;
assign w50930 = ~w50743 & w50790;
assign w50931 = ~w50782 & w50911;
assign w50932 = ~w50930 & w50931;
assign w50933 = ~w50927 & ~w50929;
assign w50934 = w50932 & w50933;
assign w50935 = ~w50773 & ~w50811;
assign w50936 = w50743 & ~w50792;
assign w50937 = ~w50935 & w50936;
assign w50938 = (~w50937 & w50925) | (~w50937 & w66845) | (w50925 & w66845);
assign w50939 = ~pi2676 & w50938;
assign w50940 = pi2676 & ~w50938;
assign w50941 = ~w50939 & ~w50940;
assign w50942 = ~w50646 & w50689;
assign w50943 = w50648 & ~w50665;
assign w50944 = ~w50689 & w50943;
assign w50945 = ~w50942 & ~w50944;
assign w50946 = w50694 & w50945;
assign w50947 = ~w50659 & ~w50946;
assign w50948 = w50644 & w50659;
assign w50949 = w50688 & w50948;
assign w50950 = w50652 & ~w50879;
assign w50951 = w50668 & ~w50950;
assign w50952 = ~w50644 & w50678;
assign w50953 = w50950 & w50952;
assign w50954 = ~w50715 & ~w50949;
assign w50955 = ~w50951 & w50954;
assign w50956 = ~w50953 & w50955;
assign w50957 = ~w50947 & w50956;
assign w50958 = pi2682 & ~w50957;
assign w50959 = ~pi2682 & w50957;
assign w50960 = ~w50958 & ~w50959;
assign w50961 = ~w50786 & ~w50919;
assign w50962 = ~w50755 & w50794;
assign w50963 = w50794 & w66846;
assign w50964 = w50743 & ~w50918;
assign w50965 = ~w50800 & ~w50906;
assign w50966 = w50964 & ~w50965;
assign w50967 = ~w50768 & w50915;
assign w50968 = w50782 & w50911;
assign w50969 = ~w50963 & ~w50966;
assign w50970 = ~w50967 & w50969;
assign w50971 = w50968 & w50970;
assign w50972 = ~w50906 & ~w50962;
assign w50973 = ~w50810 & w50972;
assign w50974 = ~w50743 & ~w50782;
assign w50975 = (w50974 & w50973) | (w50974 & w66847) | (w50973 & w66847);
assign w50976 = (w50961 & w50971) | (w50961 & w66848) | (w50971 & w66848);
assign w50977 = w50961 & w50973;
assign w50978 = ~w50749 & w50918;
assign w50979 = ~w50930 & w50978;
assign w50980 = w50743 & ~w50782;
assign w50981 = ~w50979 & w50980;
assign w50982 = ~w50977 & w50981;
assign w50983 = ~w50976 & ~w50982;
assign w50984 = pi2680 & w50983;
assign w50985 = ~pi2680 & ~w50983;
assign w50986 = ~w50984 & ~w50985;
assign w50987 = w50280 & w50332;
assign w50988 = ~w50264 & w50294;
assign w50989 = w50303 & w50988;
assign w50990 = ~w50252 & ~w50989;
assign w50991 = w50258 & ~w50316;
assign w50992 = ~w50327 & w50991;
assign w50993 = w50311 & w66849;
assign w50994 = ~w50285 & w50316;
assign w50995 = ~w50271 & w50277;
assign w50996 = ~w50264 & w50995;
assign w50997 = ~w50333 & ~w50996;
assign w50998 = w50294 & ~w50997;
assign w50999 = ~w50992 & ~w50993;
assign w51000 = ~w50994 & ~w50998;
assign w51001 = w50999 & w51000;
assign w51002 = w50286 & ~w50304;
assign w51003 = w50294 & ~w50311;
assign w51004 = ~w50988 & w50995;
assign w51005 = ~w51003 & ~w51004;
assign w51006 = w50258 & ~w51005;
assign w51007 = ~w50278 & ~w50281;
assign w51008 = ~w50258 & ~w51007;
assign w51009 = ~w50295 & w51008;
assign w51010 = ~w51002 & ~w51009;
assign w51011 = ~w51006 & w51010;
assign w51012 = ~w50252 & ~w51011;
assign w51013 = (~w50987 & w51001) | (~w50987 & w66850) | (w51001 & w66850);
assign w51014 = ~w51012 & w51013;
assign w51015 = pi2675 & w51014;
assign w51016 = ~pi2675 & ~w51014;
assign w51017 = ~w51015 & ~w51016;
assign w51018 = w49954 & w49968;
assign w51019 = ~w49951 & ~w50843;
assign w51020 = ~w51018 & ~w51019;
assign w51021 = w49956 & w50558;
assign w51022 = w49970 & ~w51021;
assign w51023 = ~w51020 & ~w51022;
assign w51024 = ~w49942 & ~w49953;
assign w51025 = w50834 & ~w51024;
assign w51026 = ~w49936 & w49957;
assign w51027 = w49917 & ~w50550;
assign w51028 = ~w49988 & w51027;
assign w51029 = ~w51026 & w51028;
assign w51030 = ~w51025 & w51029;
assign w51031 = ~w49950 & ~w49981;
assign w51032 = ~w49936 & ~w51031;
assign w51033 = ~w49917 & ~w49992;
assign w51034 = ~w50838 & w51033;
assign w51035 = ~w51032 & w51034;
assign w51036 = ~w51030 & ~w51035;
assign w51037 = ~w51023 & ~w51036;
assign w51038 = ~pi2689 & w51037;
assign w51039 = pi2689 & ~w51037;
assign w51040 = ~w51038 & ~w51039;
assign w51041 = ~w50458 & ~w50465;
assign w51042 = w50517 & w50584;
assign w51043 = (~w51042 & w50856) | (~w51042 & w66851) | (w50856 & w66851);
assign w51044 = w50479 & ~w51043;
assign w51045 = ~w50520 & w50866;
assign w51046 = w50856 & w64071;
assign w51047 = ~w50521 & ~w50575;
assign w51048 = ~w50504 & w51047;
assign w51049 = ~w50494 & w51048;
assign w51050 = (~w51045 & w51046) | (~w51045 & w66852) | (w51046 & w66852);
assign w51051 = ~w51044 & ~w51050;
assign w51052 = ~pi2672 & w51051;
assign w51053 = pi2672 & ~w51051;
assign w51054 = ~w51052 & ~w51053;
assign w51055 = w50321 & ~w50327;
assign w51056 = w50300 & ~w50320;
assign w51057 = ~w50330 & ~w51007;
assign w51058 = w50313 & w51057;
assign w51059 = ~w50252 & ~w51056;
assign w51060 = ~w51058 & w51059;
assign w51061 = ~w50279 & ~w50329;
assign w51062 = ~w50996 & w51061;
assign w51063 = w51061 & w66853;
assign w51064 = ~w50299 & w66854;
assign w51065 = ~w51060 & ~w51064;
assign w51066 = w50286 & w51003;
assign w51067 = ~w51055 & ~w51066;
assign w51068 = ~w50315 & w51067;
assign w51069 = ~w51065 & w51068;
assign w51070 = ~pi2693 & ~w51069;
assign w51071 = pi2693 & w51069;
assign w51072 = ~w51070 & ~w51071;
assign w51073 = w50993 & ~w51062;
assign w51074 = w50252 & w50280;
assign w51075 = ~w50296 & ~w51002;
assign w51076 = ~w51074 & ~w51075;
assign w51077 = w50265 & w50316;
assign w51078 = ~w51076 & ~w51077;
assign w51079 = ~w50294 & ~w51078;
assign w51080 = w50280 & w50286;
assign w51081 = (~w51080 & ~w50295) | (~w51080 & w66855) | (~w50295 & w66855);
assign w51082 = ~w50252 & ~w51081;
assign w51083 = w50258 & w50318;
assign w51084 = ~w50305 & ~w50318;
assign w51085 = ~w50296 & w51084;
assign w51086 = w50278 & ~w51085;
assign w51087 = w50324 & w51084;
assign w51088 = ~w51083 & ~w51087;
assign w51089 = ~w51086 & w51088;
assign w51090 = w50252 & ~w51089;
assign w51091 = ~w51073 & ~w51082;
assign w51092 = ~w51090 & w51091;
assign w51093 = ~w51079 & w51092;
assign w51094 = pi2698 & w51093;
assign w51095 = ~pi2698 & ~w51093;
assign w51096 = ~w51094 & ~w51095;
assign w51097 = ~w50799 & ~w50963;
assign w51098 = w50964 & ~w51097;
assign w51099 = w50799 & w50801;
assign w51100 = ~w50774 & ~w50905;
assign w51101 = ~w50800 & ~w50907;
assign w51102 = ~w51100 & ~w51101;
assign w51103 = w50788 & ~w51099;
assign w51104 = ~w51102 & w51103;
assign w51105 = w50743 & ~w50926;
assign w51106 = ~w50775 & w50782;
assign w51107 = ~w51105 & w51106;
assign w51108 = ~w51104 & ~w51107;
assign w51109 = w50782 & w50793;
assign w51110 = ~w50794 & ~w51109;
assign w51111 = ~w50743 & ~w50785;
assign w51112 = ~w51110 & w51111;
assign w51113 = ~w51098 & ~w51112;
assign w51114 = ~w51108 & w51113;
assign w51115 = pi2687 & ~w51114;
assign w51116 = ~pi2687 & w51114;
assign w51117 = ~w51115 & ~w51116;
assign w51118 = ~pi6079 & pi9040;
assign w51119 = ~pi6265 & ~pi9040;
assign w51120 = ~w51118 & ~w51119;
assign w51121 = pi2717 & ~w51120;
assign w51122 = ~pi2717 & w51120;
assign w51123 = ~w51121 & ~w51122;
assign w51124 = ~pi6086 & pi9040;
assign w51125 = ~pi6121 & ~pi9040;
assign w51126 = ~w51124 & ~w51125;
assign w51127 = pi2711 & ~w51126;
assign w51128 = ~pi2711 & w51126;
assign w51129 = ~w51127 & ~w51128;
assign w51130 = ~pi6266 & pi9040;
assign w51131 = ~pi6029 & ~pi9040;
assign w51132 = ~w51130 & ~w51131;
assign w51133 = pi2683 & ~w51132;
assign w51134 = ~pi2683 & w51132;
assign w51135 = ~w51133 & ~w51134;
assign w51136 = w51129 & ~w51135;
assign w51137 = ~pi6072 & pi9040;
assign w51138 = ~pi6046 & ~pi9040;
assign w51139 = ~w51137 & ~w51138;
assign w51140 = pi2695 & ~w51139;
assign w51141 = ~pi2695 & w51139;
assign w51142 = ~w51140 & ~w51141;
assign w51143 = ~pi5952 & pi9040;
assign w51144 = ~pi6275 & ~pi9040;
assign w51145 = ~w51143 & ~w51144;
assign w51146 = pi2710 & ~w51145;
assign w51147 = ~pi2710 & w51145;
assign w51148 = ~w51146 & ~w51147;
assign w51149 = w51142 & ~w51148;
assign w51150 = ~pi6074 & pi9040;
assign w51151 = ~pi6068 & ~pi9040;
assign w51152 = ~w51150 & ~w51151;
assign w51153 = pi2714 & ~w51152;
assign w51154 = ~pi2714 & w51152;
assign w51155 = ~w51153 & ~w51154;
assign w51156 = ~w51149 & ~w51155;
assign w51157 = ~w51136 & ~w51156;
assign w51158 = ~w51135 & ~w51155;
assign w51159 = w51157 & w51158;
assign w51160 = ~w51129 & w51142;
assign w51161 = w51135 & ~w51142;
assign w51162 = ~w51135 & w51142;
assign w51163 = ~w51161 & ~w51162;
assign w51164 = (~w51160 & w51163) | (~w51160 & w64072) | (w51163 & w64072);
assign w51165 = w51135 & w51142;
assign w51166 = w51155 & w51165;
assign w51167 = ~w51135 & w51148;
assign w51168 = ~w51142 & w51167;
assign w51169 = w51167 & w66856;
assign w51170 = ~w51148 & w51158;
assign w51171 = w51135 & ~w51148;
assign w51172 = ~w51142 & w51171;
assign w51173 = ~w51170 & ~w51172;
assign w51174 = ~w51166 & ~w51169;
assign w51175 = w51173 & w51174;
assign w51176 = w51164 & w51175;
assign w51177 = ~w51159 & ~w51176;
assign w51178 = w51123 & ~w51177;
assign w51179 = ~w51157 & ~w51173;
assign w51180 = ~w51167 & ~w51171;
assign w51181 = ~w51164 & ~w51180;
assign w51182 = w51148 & w51155;
assign w51183 = w51129 & ~w51162;
assign w51184 = ~w51161 & ~w51183;
assign w51185 = (w51182 & w51183) | (w51182 & w66857) | (w51183 & w66857);
assign w51186 = ~w51179 & ~w51185;
assign w51187 = (~w51123 & ~w51186) | (~w51123 & w66858) | (~w51186 & w66858);
assign w51188 = w51155 & w51180;
assign w51189 = w51142 & w51155;
assign w51190 = w51148 & w51163;
assign w51191 = (~w51155 & w51190) | (~w51155 & w66859) | (w51190 & w66859);
assign w51192 = ~w51189 & ~w51191;
assign w51193 = ~w51129 & ~w51188;
assign w51194 = ~w51192 & w51193;
assign w51195 = ~w51187 & ~w51194;
assign w51196 = ~w51178 & w51195;
assign w51197 = pi2729 & w51196;
assign w51198 = ~pi2729 & ~w51196;
assign w51199 = ~w51197 & ~w51198;
assign w51200 = ~w51129 & ~w51142;
assign w51201 = w51180 & w51200;
assign w51202 = w51129 & w51161;
assign w51203 = w51161 & w64073;
assign w51204 = w51155 & ~w51203;
assign w51205 = ~w51201 & w51204;
assign w51206 = w51160 & w51167;
assign w51207 = ~w51155 & ~w51206;
assign w51208 = ~w51205 & ~w51207;
assign w51209 = ~w51129 & ~w51155;
assign w51210 = ~w51180 & w51209;
assign w51211 = ~w51163 & w51188;
assign w51212 = w51129 & w51180;
assign w51213 = w51129 & ~w51158;
assign w51214 = ~w51162 & ~w51213;
assign w51215 = ~w51190 & ~w51214;
assign w51216 = w51212 & ~w51215;
assign w51217 = w51123 & ~w51206;
assign w51218 = ~w51210 & w51217;
assign w51219 = ~w51211 & w51218;
assign w51220 = ~w51216 & w51219;
assign w51221 = w51136 & w51182;
assign w51222 = ~w51135 & w51200;
assign w51223 = ~w51148 & w51222;
assign w51224 = w51163 & w51188;
assign w51225 = ~w51149 & ~w51202;
assign w51226 = w51160 & w51171;
assign w51227 = w51155 & ~w51226;
assign w51228 = ~w51225 & ~w51227;
assign w51229 = ~w51123 & ~w51169;
assign w51230 = ~w51221 & ~w51223;
assign w51231 = ~w51224 & w51230;
assign w51232 = ~w51228 & w51229;
assign w51233 = w51231 & w51232;
assign w51234 = ~w51220 & ~w51233;
assign w51235 = ~w51208 & ~w51234;
assign w51236 = ~pi2731 & w51235;
assign w51237 = pi2731 & ~w51235;
assign w51238 = ~w51236 & ~w51237;
assign w51239 = w51185 & w51200;
assign w51240 = (~w51202 & w51164) | (~w51202 & w66860) | (w51164 & w66860);
assign w51241 = w51156 & ~w51240;
assign w51242 = w51180 & w64074;
assign w51243 = ~w51168 & ~w51226;
assign w51244 = w51155 & ~w51243;
assign w51245 = w51123 & ~w51242;
assign w51246 = ~w51244 & w51245;
assign w51247 = ~w51241 & w51246;
assign w51248 = w51171 & w51227;
assign w51249 = w51180 & w51214;
assign w51250 = ~w51158 & w51160;
assign w51251 = ~w51166 & w51250;
assign w51252 = w51229 & ~w51251;
assign w51253 = ~w51248 & ~w51249;
assign w51254 = w51252 & w51253;
assign w51255 = ~w51247 & ~w51254;
assign w51256 = ~w51223 & ~w51242;
assign w51257 = ~w51155 & ~w51256;
assign w51258 = ~w51221 & ~w51239;
assign w51259 = ~w51257 & w51258;
assign w51260 = ~w51255 & w51259;
assign w51261 = pi2747 & ~w51260;
assign w51262 = ~pi2747 & w51260;
assign w51263 = ~w51261 & ~w51262;
assign w51264 = ~pi6094 & pi9040;
assign w51265 = ~pi5963 & ~pi9040;
assign w51266 = ~w51264 & ~w51265;
assign w51267 = pi2668 & ~w51266;
assign w51268 = ~pi2668 & w51266;
assign w51269 = ~w51267 & ~w51268;
assign w51270 = ~pi6043 & pi9040;
assign w51271 = ~pi6166 & ~pi9040;
assign w51272 = ~w51270 & ~w51271;
assign w51273 = pi2709 & ~w51272;
assign w51274 = ~pi2709 & w51272;
assign w51275 = ~w51273 & ~w51274;
assign w51276 = w51269 & w51275;
assign w51277 = ~pi6025 & pi9040;
assign w51278 = ~pi6167 & ~pi9040;
assign w51279 = ~w51277 & ~w51278;
assign w51280 = pi2692 & ~w51279;
assign w51281 = ~pi2692 & w51279;
assign w51282 = ~w51280 & ~w51281;
assign w51283 = w51276 & ~w51282;
assign w51284 = ~pi5964 & pi9040;
assign w51285 = ~pi6017 & ~pi9040;
assign w51286 = ~w51284 & ~w51285;
assign w51287 = pi2702 & ~w51286;
assign w51288 = ~pi2702 & w51286;
assign w51289 = ~w51287 & ~w51288;
assign w51290 = (w51289 & ~w51276) | (w51289 & w51806) | (~w51276 & w51806);
assign w51291 = w51269 & ~w51275;
assign w51292 = ~pi6165 & pi9040;
assign w51293 = ~pi6089 & ~pi9040;
assign w51294 = ~w51292 & ~w51293;
assign w51295 = pi2700 & ~w51294;
assign w51296 = ~pi2700 & w51294;
assign w51297 = ~w51295 & ~w51296;
assign w51298 = ~w51275 & w51297;
assign w51299 = w51275 & ~w51297;
assign w51300 = ~w51298 & ~w51299;
assign w51301 = w51282 & w51300;
assign w51302 = w51300 & w66861;
assign w51303 = w51290 & ~w51302;
assign w51304 = w51282 & ~w51297;
assign w51305 = ~w51275 & ~w51282;
assign w51306 = ~w51304 & ~w51305;
assign w51307 = ~w51269 & w51306;
assign w51308 = ~w51269 & ~w51275;
assign w51309 = ~w51282 & w51300;
assign w51310 = (~w51308 & ~w51300) | (~w51308 & w64075) | (~w51300 & w64075);
assign w51311 = w51307 & ~w51310;
assign w51312 = w51269 & ~w51306;
assign w51313 = ~w51311 & w66862;
assign w51314 = ~pi6039 & pi9040;
assign w51315 = ~pi6204 & ~pi9040;
assign w51316 = ~w51314 & ~w51315;
assign w51317 = pi2716 & ~w51316;
assign w51318 = ~pi2716 & w51316;
assign w51319 = ~w51317 & ~w51318;
assign w51320 = ~w51303 & w51319;
assign w51321 = ~w51313 & w51320;
assign w51322 = ~w51269 & w51275;
assign w51323 = w51282 & w51322;
assign w51324 = w51289 & ~w51305;
assign w51325 = ~w51323 & w51324;
assign w51326 = ~w51282 & w51297;
assign w51327 = ~w51304 & ~w51326;
assign w51328 = ~w51283 & ~w51308;
assign w51329 = w51327 & w51328;
assign w51330 = ~w51269 & ~w51282;
assign w51331 = ~w51326 & ~w51330;
assign w51332 = w51290 & ~w51331;
assign w51333 = w51322 & w51304;
assign w51334 = ~w51332 & ~w51333;
assign w51335 = w51269 & ~w51327;
assign w51336 = w51289 & ~w51298;
assign w51337 = ~w51291 & w51336;
assign w51338 = ~w51307 & ~w51335;
assign w51339 = ~w51337 & w51338;
assign w51340 = ~w51334 & w51339;
assign w51341 = ~w51289 & ~w51297;
assign w51342 = w51330 & w51341;
assign w51343 = ~w51275 & w51342;
assign w51344 = ~w51282 & ~w51289;
assign w51345 = ~w51269 & ~w51344;
assign w51346 = ~w51283 & ~w51345;
assign w51347 = ~w51311 & w66863;
assign w51348 = w51282 & w51291;
assign w51349 = ~w51341 & w51348;
assign w51350 = w51334 & ~w51349;
assign w51351 = ~w51347 & w51350;
assign w51352 = ~w51319 & ~w51351;
assign w51353 = (~w51343 & ~w51329) | (~w51343 & w66864) | (~w51329 & w66864);
assign w51354 = ~w51340 & w51353;
assign w51355 = ~w51321 & w51354;
assign w51356 = (pi2726 & ~w51355) | (pi2726 & w66865) | (~w51355 & w66865);
assign w51357 = w51355 & w66866;
assign w51358 = ~w51356 & ~w51357;
assign w51359 = ~pi6073 & pi9040;
assign w51360 = ~pi6179 & ~pi9040;
assign w51361 = ~w51359 & ~w51360;
assign w51362 = pi2701 & ~w51361;
assign w51363 = ~pi2701 & w51361;
assign w51364 = ~w51362 & ~w51363;
assign w51365 = ~pi6017 & pi9040;
assign w51366 = ~pi6040 & ~pi9040;
assign w51367 = ~w51365 & ~w51366;
assign w51368 = pi2694 & ~w51367;
assign w51369 = ~pi2694 & w51367;
assign w51370 = ~w51368 & ~w51369;
assign w51371 = w51364 & ~w51370;
assign w51372 = ~pi6010 & pi9040;
assign w51373 = ~pi6039 & ~pi9040;
assign w51374 = ~w51372 & ~w51373;
assign w51375 = pi2708 & ~w51374;
assign w51376 = ~pi2708 & w51374;
assign w51377 = ~w51375 & ~w51376;
assign w51378 = ~pi6007 & pi9040;
assign w51379 = ~pi6094 & ~pi9040;
assign w51380 = ~w51378 & ~w51379;
assign w51381 = pi2718 & ~w51380;
assign w51382 = ~pi2718 & w51380;
assign w51383 = ~w51381 & ~w51382;
assign w51384 = w51377 & w51383;
assign w51385 = w51371 & w51384;
assign w51386 = w51377 & ~w51383;
assign w51387 = ~w51364 & w51386;
assign w51388 = w51386 & w51398;
assign w51389 = ~w51385 & ~w51388;
assign w51390 = ~pi6145 & pi9040;
assign w51391 = ~pi6093 & ~pi9040;
assign w51392 = ~w51390 & ~w51391;
assign w51393 = pi2690 & ~w51392;
assign w51394 = ~pi2690 & w51392;
assign w51395 = ~w51393 & ~w51394;
assign w51396 = ~w51364 & w51370;
assign w51397 = w51383 & w51396;
assign w51398 = ~w51364 & ~w51370;
assign w51399 = ~w51377 & ~w51383;
assign w51400 = w51398 & w51399;
assign w51401 = (~w51395 & ~w51396) | (~w51395 & w66867) | (~w51396 & w66867);
assign w51402 = ~w51400 & w51401;
assign w51403 = w51389 & w51402;
assign w51404 = w51370 & ~w51383;
assign w51405 = w51364 & ~w51377;
assign w51406 = w51404 & ~w51405;
assign w51407 = w51364 & ~w51404;
assign w51408 = w51370 & w51377;
assign w51409 = ~w51386 & ~w51408;
assign w51410 = w51407 & w51409;
assign w51411 = w51395 & ~w51406;
assign w51412 = ~w51410 & w51411;
assign w51413 = ~w51403 & ~w51412;
assign w51414 = ~w51395 & w51404;
assign w51415 = w51405 & w51414;
assign w51416 = ~w51413 & ~w51415;
assign w51417 = ~pi6048 & pi9040;
assign w51418 = ~pi6025 & ~pi9040;
assign w51419 = ~w51417 & ~w51418;
assign w51420 = pi2699 & ~w51419;
assign w51421 = ~pi2699 & w51419;
assign w51422 = ~w51420 & ~w51421;
assign w51423 = ~w51416 & w51422;
assign w51424 = ~w51377 & w51383;
assign w51425 = w51371 & w51424;
assign w51426 = w51386 & w51396;
assign w51427 = ~w51425 & ~w51426;
assign w51428 = w51377 & w51398;
assign w51429 = (w51395 & ~w51398) | (w51395 & w66868) | (~w51398 & w66868);
assign w51430 = ~w51371 & ~w51384;
assign w51431 = ~w51429 & ~w51430;
assign w51432 = ~w51400 & w51427;
assign w51433 = ~w51431 & w51432;
assign w51434 = w51395 & ~w51433;
assign w51435 = w51396 & w51424;
assign w51436 = w51429 & ~w51435;
assign w51437 = w51364 & w51377;
assign w51438 = ~w51395 & ~w51437;
assign w51439 = ~w51370 & w51424;
assign w51440 = w51438 & ~w51439;
assign w51441 = ~w51436 & ~w51440;
assign w51442 = w51364 & w51370;
assign w51443 = ~w51383 & w51405;
assign w51444 = ~w51384 & ~w51443;
assign w51445 = (w51442 & w51443) | (w51442 & w66869) | (w51443 & w66869);
assign w51446 = ~w51414 & ~w51445;
assign w51447 = ~w51441 & w51446;
assign w51448 = ~w51422 & ~w51447;
assign w51449 = ~w51434 & ~w51448;
assign w51450 = ~w51423 & w51449;
assign w51451 = pi2721 & ~w51450;
assign w51452 = ~pi2721 & w51450;
assign w51453 = ~w51451 & ~w51452;
assign w51454 = ~pi6044 & pi9040;
assign w51455 = ~pi6139 & ~pi9040;
assign w51456 = ~w51454 & ~w51455;
assign w51457 = pi2674 & ~w51456;
assign w51458 = ~pi2674 & w51456;
assign w51459 = ~w51457 & ~w51458;
assign w51460 = ~pi6029 & pi9040;
assign w51461 = ~pi6183 & ~pi9040;
assign w51462 = ~w51460 & ~w51461;
assign w51463 = pi2708 & ~w51462;
assign w51464 = ~pi2708 & w51462;
assign w51465 = ~w51463 & ~w51464;
assign w51466 = ~w51459 & w51465;
assign w51467 = ~pi6265 & pi9040;
assign w51468 = ~pi5956 & ~pi9040;
assign w51469 = ~w51467 & ~w51468;
assign w51470 = pi2699 & ~w51469;
assign w51471 = ~pi2699 & w51469;
assign w51472 = ~w51470 & ~w51471;
assign w51473 = ~pi6142 & pi9040;
assign w51474 = ~pi6241 & ~pi9040;
assign w51475 = ~w51473 & ~w51474;
assign w51476 = pi2707 & ~w51475;
assign w51477 = ~pi2707 & w51475;
assign w51478 = ~w51476 & ~w51477;
assign w51479 = w51472 & ~w51478;
assign w51480 = w51466 & w51479;
assign w51481 = ~pi6047 & pi9040;
assign w51482 = ~pi6072 & ~pi9040;
assign w51483 = ~w51481 & ~w51482;
assign w51484 = pi2713 & ~w51483;
assign w51485 = ~pi2713 & w51483;
assign w51486 = ~w51484 & ~w51485;
assign w51487 = ~w51480 & w51486;
assign w51488 = w51459 & w51478;
assign w51489 = w51465 & w51488;
assign w51490 = ~w51465 & ~w51478;
assign w51491 = ~w51472 & ~w51490;
assign w51492 = ~pi6032 & pi9040;
assign w51493 = ~pi5965 & ~pi9040;
assign w51494 = ~w51492 & ~w51493;
assign w51495 = pi2719 & ~w51494;
assign w51496 = ~pi2719 & w51494;
assign w51497 = ~w51495 & ~w51496;
assign w51498 = ~w51479 & ~w51497;
assign w51499 = ~w51491 & w51498;
assign w51500 = w51459 & w51472;
assign w51501 = ~w51478 & w51500;
assign w51502 = w51500 & w51490;
assign w51503 = ~w51491 & ~w51502;
assign w51504 = w51497 & ~w51503;
assign w51505 = ~w51489 & ~w51499;
assign w51506 = ~w51504 & w51505;
assign w51507 = w51487 & w51506;
assign w51508 = w51459 & ~w51465;
assign w51509 = ~w51466 & ~w51508;
assign w51510 = w51497 & w51509;
assign w51511 = w51509 & w66870;
assign w51512 = ~w51459 & ~w51472;
assign w51513 = ~w51500 & ~w51512;
assign w51514 = ~w51465 & ~w51513;
assign w51515 = ~w51472 & ~w51478;
assign w51516 = w51466 & w51515;
assign w51517 = (~w51497 & w51514) | (~w51497 & w66871) | (w51514 & w66871);
assign w51518 = ~w51509 & ~w51512;
assign w51519 = ~w51465 & w51472;
assign w51520 = w51478 & ~w51519;
assign w51521 = w51518 & w51520;
assign w51522 = ~w51511 & ~w51521;
assign w51523 = ~w51517 & w51522;
assign w51524 = w51522 & w66872;
assign w51525 = ~w51507 & ~w51524;
assign w51526 = ~w51459 & w51490;
assign w51527 = w51497 & w51515;
assign w51528 = ~w51526 & ~w51527;
assign w51529 = w51513 & ~w51528;
assign w51530 = ~w51508 & ~w51520;
assign w51531 = ~w51465 & ~w51472;
assign w51532 = ~w51530 & w51531;
assign w51533 = w51478 & w51497;
assign w51534 = w51512 & w51533;
assign w51535 = w51465 & ~w51497;
assign w51536 = w51472 & w51535;
assign w51537 = ~w51534 & ~w51536;
assign w51538 = ~w51529 & w51537;
assign w51539 = ~w51532 & w51538;
assign w51540 = w51465 & w51497;
assign w51541 = ~w51539 & w51540;
assign w51542 = ~w51525 & ~w51541;
assign w51543 = ~pi2735 & w51542;
assign w51544 = pi2735 & ~w51542;
assign w51545 = ~w51543 & ~w51544;
assign w51546 = (~w51149 & w51164) | (~w51149 & w66873) | (w51164 & w66873);
assign w51547 = w51217 & ~w51546;
assign w51548 = ~w51169 & ~w51547;
assign w51549 = w51155 & ~w51548;
assign w51550 = (~w51123 & ~w51156) | (~w51123 & w66874) | (~w51156 & w66874);
assign w51551 = ~w51165 & ~w51550;
assign w51552 = ~w51189 & ~w51551;
assign w51553 = w51212 & ~w51552;
assign w51554 = (~w51123 & w51163) | (~w51123 & w64076) | (w51163 & w64076);
assign w51555 = ~w51242 & w51554;
assign w51556 = w51148 & ~w51555;
assign w51557 = w51204 & ~w51222;
assign w51558 = (~w51158 & ~w51156) | (~w51158 & w66875) | (~w51156 & w66875);
assign w51559 = ~w51557 & w51558;
assign w51560 = ~w51556 & ~w51559;
assign w51561 = w51148 & ~w51155;
assign w51562 = w51184 & w51561;
assign w51563 = w51123 & ~w51562;
assign w51564 = ~w51560 & ~w51563;
assign w51565 = ~w51553 & ~w51564;
assign w51566 = (pi2750 & ~w51565) | (pi2750 & w66876) | (~w51565 & w66876);
assign w51567 = w51565 & w66877;
assign w51568 = ~w51566 & ~w51567;
assign w51569 = ~pi6166 & pi9040;
assign w51570 = ~pi6073 & ~pi9040;
assign w51571 = ~w51569 & ~w51570;
assign w51572 = pi2717 & ~w51571;
assign w51573 = ~pi2717 & w51571;
assign w51574 = ~w51572 & ~w51573;
assign w51575 = ~pi5963 & pi9040;
assign w51576 = ~pi6124 & ~pi9040;
assign w51577 = ~w51575 & ~w51576;
assign w51578 = pi2695 & ~w51577;
assign w51579 = ~pi2695 & w51577;
assign w51580 = ~w51578 & ~w51579;
assign w51581 = ~w51574 & w51580;
assign w51582 = ~pi6167 & pi9040;
assign w51583 = ~pi6010 & ~pi9040;
assign w51584 = ~w51582 & ~w51583;
assign w51585 = pi2715 & ~w51584;
assign w51586 = ~pi2715 & w51584;
assign w51587 = ~w51585 & ~w51586;
assign w51588 = ~w51574 & ~w51587;
assign w51589 = ~pi6034 & pi9040;
assign w51590 = ~pi6075 & ~pi9040;
assign w51591 = ~w51589 & ~w51590;
assign w51592 = pi2709 & ~w51591;
assign w51593 = ~pi2709 & w51591;
assign w51594 = ~w51592 & ~w51593;
assign w51595 = w51588 & w51594;
assign w51596 = w51574 & ~w51594;
assign w51597 = w51580 & w51596;
assign w51598 = ~w51595 & ~w51597;
assign w51599 = ~pi6093 & pi9040;
assign w51600 = ~pi6030 & ~pi9040;
assign w51601 = ~w51599 & ~w51600;
assign w51602 = pi2697 & ~w51601;
assign w51603 = ~pi2697 & w51601;
assign w51604 = ~w51602 & ~w51603;
assign w51605 = ~w51598 & w51604;
assign w51606 = ~w51598 & w66878;
assign w51607 = ~w51574 & w51587;
assign w51608 = w51580 & w51594;
assign w51609 = ~w51580 & ~w51594;
assign w51610 = ~w51608 & ~w51609;
assign w51611 = w51607 & w51610;
assign w51612 = w51574 & ~w51587;
assign w51613 = ~w51604 & ~w51612;
assign w51614 = ~w51580 & ~w51596;
assign w51615 = ~w51587 & ~w51594;
assign w51616 = ~w51574 & ~w51615;
assign w51617 = w51614 & ~w51616;
assign w51618 = w51604 & ~w51617;
assign w51619 = (~w51613 & w51617) | (~w51613 & w66879) | (w51617 & w66879);
assign w51620 = ~w51611 & ~w51619;
assign w51621 = ~pi6040 & pi9040;
assign w51622 = ~pi6165 & ~pi9040;
assign w51623 = ~w51621 & ~w51622;
assign w51624 = pi2692 & ~w51623;
assign w51625 = ~pi2692 & w51623;
assign w51626 = ~w51624 & ~w51625;
assign w51627 = ~w51620 & w51626;
assign w51628 = w51574 & w51604;
assign w51629 = ~w51574 & ~w51594;
assign w51630 = ~w51615 & ~w51629;
assign w51631 = w51580 & ~w51607;
assign w51632 = ~w51630 & ~w51631;
assign w51633 = w51628 & w51632;
assign w51634 = w51574 & ~w51580;
assign w51635 = w51594 & w51634;
assign w51636 = ~w51595 & ~w51635;
assign w51637 = ~w51604 & ~w51636;
assign w51638 = w51580 & w51588;
assign w51639 = ~w51574 & ~w51604;
assign w51640 = ~w51628 & ~w51639;
assign w51641 = w51608 & ~w51640;
assign w51642 = w51587 & ~w51594;
assign w51643 = ~w51581 & ~w51634;
assign w51644 = w51642 & w51643;
assign w51645 = ~w51638 & ~w51641;
assign w51646 = ~w51644 & w51645;
assign w51647 = ~w51633 & ~w51637;
assign w51648 = w51646 & w51647;
assign w51649 = ~w51626 & ~w51648;
assign w51650 = w51604 & ~w51609;
assign w51651 = ~w51587 & ~w51604;
assign w51652 = ~w51634 & ~w51651;
assign w51653 = w51640 & ~w51652;
assign w51654 = (w51642 & w51653) | (w51642 & w66880) | (w51653 & w66880);
assign w51655 = w51587 & w51614;
assign w51656 = w51587 & w51594;
assign w51657 = ~w51581 & ~w51656;
assign w51658 = ~w51607 & ~w51657;
assign w51659 = w51650 & ~w51658;
assign w51660 = ~w51658 & w66881;
assign w51661 = w51655 & w51660;
assign w51662 = ~w51606 & ~w51654;
assign w51663 = ~w51661 & w51662;
assign w51664 = ~w51627 & w51663;
assign w51665 = ~w51649 & w51664;
assign w51666 = pi2725 & ~w51665;
assign w51667 = ~pi2725 & w51665;
assign w51668 = ~w51666 & ~w51667;
assign w51669 = w51276 & w51304;
assign w51670 = w51331 & ~w51669;
assign w51671 = w51324 & ~w51670;
assign w51672 = (w51319 & w51339) | (w51319 & w66882) | (w51339 & w66882);
assign w51673 = w51289 & w51297;
assign w51674 = w51322 & w51673;
assign w51675 = w51291 & w51326;
assign w51676 = (~w51289 & w51307) | (~w51289 & w66883) | (w51307 & w66883);
assign w51677 = ~w51333 & w51336;
assign w51678 = ~w51339 & w64077;
assign w51679 = ~w51675 & ~w51676;
assign w51680 = (~w51319 & w51678) | (~w51319 & w66884) | (w51678 & w66884);
assign w51681 = w51304 & w51308;
assign w51682 = ~w51674 & ~w51681;
assign w51683 = ~w51672 & w51682;
assign w51684 = ~w51680 & w51683;
assign w51685 = pi2720 & ~w51684;
assign w51686 = ~pi2720 & w51684;
assign w51687 = ~w51685 & ~w51686;
assign w51688 = ~w51497 & ~w51500;
assign w51689 = w51518 & w51688;
assign w51690 = ~w51516 & ~w51689;
assign w51691 = w51506 & ~w51690;
assign w51692 = ~w51465 & w51534;
assign w51693 = w51488 & w51536;
assign w51694 = ~w51478 & w51497;
assign w51695 = w51519 & w51694;
assign w51696 = ~w51693 & ~w51695;
assign w51697 = w51465 & w51513;
assign w51698 = w51513 & w64078;
assign w51699 = w51501 & ~w51535;
assign w51700 = ~w51698 & ~w51699;
assign w51701 = w51498 & w51530;
assign w51702 = ~w51486 & ~w51516;
assign w51703 = ~w51701 & w51702;
assign w51704 = w51700 & w51703;
assign w51705 = w51497 & w51508;
assign w51706 = w51486 & ~w51705;
assign w51707 = w51538 & w66885;
assign w51708 = ~w51704 & ~w51707;
assign w51709 = ~w51692 & w51696;
assign w51710 = ~w51691 & w51709;
assign w51711 = ~w51708 & w51710;
assign w51712 = pi2732 & ~w51711;
assign w51713 = ~pi2732 & w51711;
assign w51714 = ~w51712 & ~w51713;
assign w51715 = ~pi6089 & pi9040;
assign w51716 = ~pi6007 & ~pi9040;
assign w51717 = ~w51715 & ~w51716;
assign w51718 = pi2700 & ~w51717;
assign w51719 = ~pi2700 & w51717;
assign w51720 = ~w51718 & ~w51719;
assign w51721 = ~pi6075 & pi9040;
assign w51722 = ~pi6048 & ~pi9040;
assign w51723 = ~w51721 & ~w51722;
assign w51724 = pi2704 & ~w51723;
assign w51725 = ~pi2704 & w51723;
assign w51726 = ~w51724 & ~w51725;
assign w51727 = ~w51720 & w51726;
assign w51728 = ~pi6124 & pi9040;
assign w51729 = ~pi5950 & ~pi9040;
assign w51730 = ~w51728 & ~w51729;
assign w51731 = pi2701 & ~w51730;
assign w51732 = ~pi2701 & w51730;
assign w51733 = ~w51731 & ~w51732;
assign w51734 = ~pi6173 & pi9040;
assign w51735 = ~pi6043 & ~pi9040;
assign w51736 = ~w51734 & ~w51735;
assign w51737 = pi2684 & ~w51736;
assign w51738 = ~pi2684 & w51736;
assign w51739 = ~w51737 & ~w51738;
assign w51740 = ~w51733 & ~w51739;
assign w51741 = w51727 & w51740;
assign w51742 = ~pi6088 & pi9040;
assign w51743 = ~pi5964 & ~pi9040;
assign w51744 = ~w51742 & ~w51743;
assign w51745 = pi2716 & ~w51744;
assign w51746 = ~pi2716 & w51744;
assign w51747 = ~w51745 & ~w51746;
assign w51748 = w51733 & ~w51747;
assign w51749 = ~w51727 & ~w51739;
assign w51750 = w51748 & w51749;
assign w51751 = w51720 & w51733;
assign w51752 = w51739 & w51747;
assign w51753 = w51751 & w51752;
assign w51754 = ~pi6204 & pi9040;
assign w51755 = ~pi6170 & ~pi9040;
assign w51756 = ~w51754 & ~w51755;
assign w51757 = pi2694 & ~w51756;
assign w51758 = ~pi2694 & w51756;
assign w51759 = ~w51757 & ~w51758;
assign w51760 = ~w51753 & ~w51759;
assign w51761 = ~w51720 & ~w51739;
assign w51762 = ~w51733 & w51747;
assign w51763 = w51726 & w51747;
assign w51764 = ~w51762 & ~w51763;
assign w51765 = w51761 & ~w51764;
assign w51766 = ~w51750 & w51760;
assign w51767 = ~w51765 & w51766;
assign w51768 = w51720 & w51739;
assign w51769 = ~w51761 & ~w51768;
assign w51770 = (~w51740 & ~w51769) | (~w51740 & w66886) | (~w51769 & w66886);
assign w51771 = (w51740 & w51769) | (w51740 & w66887) | (w51769 & w66887);
assign w51772 = ~w51770 & ~w51771;
assign w51773 = w51739 & ~w51747;
assign w51774 = ~w51720 & w51733;
assign w51775 = w51773 & w51774;
assign w51776 = w51759 & ~w51775;
assign w51777 = ~w51772 & w51776;
assign w51778 = ~w51767 & ~w51777;
assign w51779 = ~w51720 & ~w51733;
assign w51780 = ~w51751 & ~w51779;
assign w51781 = w51773 & w51780;
assign w51782 = w51747 & w51779;
assign w51783 = ~w51781 & ~w51782;
assign w51784 = w51726 & ~w51783;
assign w51785 = ~w51739 & w51747;
assign w51786 = w51774 & w51785;
assign w51787 = ~w51747 & w51751;
assign w51788 = ~w51786 & ~w51787;
assign w51789 = w51759 & ~w51788;
assign w51790 = ~w51773 & ~w51785;
assign w51791 = w51720 & w51790;
assign w51792 = ~w51748 & ~w51762;
assign w51793 = ~w51739 & w51792;
assign w51794 = ~w51759 & ~w51793;
assign w51795 = ~w51781 & w66888;
assign w51796 = w51794 & w51795;
assign w51797 = ~w51789 & ~w51791;
assign w51798 = ~w51796 & w51797;
assign w51799 = ~w51726 & ~w51798;
assign w51800 = ~w51741 & ~w51784;
assign w51801 = ~w51778 & w51800;
assign w51802 = ~w51799 & w51801;
assign w51803 = pi2728 & ~w51802;
assign w51804 = ~pi2728 & w51802;
assign w51805 = ~w51803 & ~w51804;
assign w51806 = w51282 & w51289;
assign w51807 = ~w51300 & w51806;
assign w51808 = ~w51307 & w51807;
assign w51809 = w51310 & w51344;
assign w51810 = w51297 & ~w51806;
assign w51811 = w51345 & w51810;
assign w51812 = ~w51319 & ~w51681;
assign w51813 = ~w51811 & w51812;
assign w51814 = ~w51808 & w51813;
assign w51815 = ~w51809 & w51814;
assign w51816 = w51276 & w51297;
assign w51817 = w51307 & ~w51810;
assign w51818 = w51319 & ~w51816;
assign w51819 = ~w51817 & w51818;
assign w51820 = w51269 & w51301;
assign w51821 = ~w51330 & ~w51333;
assign w51822 = w51319 & ~w51821;
assign w51823 = ~w51289 & ~w51820;
assign w51824 = ~w51822 & w51823;
assign w51825 = w51269 & w51309;
assign w51826 = w51289 & ~w51669;
assign w51827 = ~w51825 & w51826;
assign w51828 = ~w51824 & ~w51827;
assign w51829 = (~w51342 & w51815) | (~w51342 & w66889) | (w51815 & w66889);
assign w51830 = ~w51828 & w51829;
assign w51831 = pi2722 & ~w51830;
assign w51832 = ~pi2722 & w51830;
assign w51833 = ~w51831 & ~w51832;
assign w51834 = ~pi6121 & pi9040;
assign w51835 = ~pi6047 & ~pi9040;
assign w51836 = ~w51834 & ~w51835;
assign w51837 = pi2674 & ~w51836;
assign w51838 = ~pi2674 & w51836;
assign w51839 = ~w51837 & ~w51838;
assign w51840 = ~pi5956 & pi9040;
assign w51841 = ~pi6266 & ~pi9040;
assign w51842 = ~w51840 & ~w51841;
assign w51843 = pi2712 & ~w51842;
assign w51844 = ~pi2712 & w51842;
assign w51845 = ~w51843 & ~w51844;
assign w51846 = w51839 & ~w51845;
assign w51847 = ~pi6046 & pi9040;
assign w51848 = ~pi5991 & ~pi9040;
assign w51849 = ~w51847 & ~w51848;
assign w51850 = pi2713 & ~w51849;
assign w51851 = ~pi2713 & w51849;
assign w51852 = ~w51850 & ~w51851;
assign w51853 = w51846 & w51852;
assign w51854 = ~pi6256 & pi9040;
assign w51855 = ~pi6142 & ~pi9040;
assign w51856 = ~w51854 & ~w51855;
assign w51857 = pi2703 & ~w51856;
assign w51858 = ~pi2703 & w51856;
assign w51859 = ~w51857 & ~w51858;
assign w51860 = w51845 & ~w51859;
assign w51861 = ~w51839 & w51860;
assign w51862 = w51860 & w66890;
assign w51863 = ~w51853 & ~w51862;
assign w51864 = ~pi6139 & pi9040;
assign w51865 = ~pi5952 & ~pi9040;
assign w51866 = ~w51864 & ~w51865;
assign w51867 = pi2686 & ~w51866;
assign w51868 = ~pi2686 & w51866;
assign w51869 = ~w51867 & ~w51868;
assign w51870 = ~w51863 & w51869;
assign w51871 = ~w51852 & w51859;
assign w51872 = w51839 & w51871;
assign w51873 = ~w51845 & w51859;
assign w51874 = ~w51872 & ~w51873;
assign w51875 = ~w51845 & w51869;
assign w51876 = ~w51846 & ~w51875;
assign w51877 = ~w51874 & w51876;
assign w51878 = w51839 & ~w51859;
assign w51879 = ~w51852 & w51878;
assign w51880 = w51878 & w66891;
assign w51881 = w51852 & w51859;
assign w51882 = w51845 & w51881;
assign w51883 = ~w51880 & ~w51882;
assign w51884 = w51869 & ~w51883;
assign w51885 = ~w51839 & w51884;
assign w51886 = ~w51839 & w51859;
assign w51887 = ~w51878 & ~w51886;
assign w51888 = ~w51881 & ~w51887;
assign w51889 = ~w51887 & w66892;
assign w51890 = w51852 & w51886;
assign w51891 = (~w51869 & ~w51886) | (~w51869 & w66893) | (~w51886 & w66893);
assign w51892 = w51845 & w51852;
assign w51893 = ~w51886 & ~w51892;
assign w51894 = w51891 & ~w51893;
assign w51895 = ~pi6068 & pi9040;
assign w51896 = ~pi6171 & ~pi9040;
assign w51897 = ~w51895 & ~w51896;
assign w51898 = pi2705 & ~w51897;
assign w51899 = ~pi2705 & w51897;
assign w51900 = ~w51898 & ~w51899;
assign w51901 = (~w51900 & w51874) | (~w51900 & w66894) | (w51874 & w66894);
assign w51902 = ~w51889 & ~w51894;
assign w51903 = w51901 & w51902;
assign w51904 = ~w51885 & w51903;
assign w51905 = w51846 & w51881;
assign w51906 = ~w51846 & ~w51852;
assign w51907 = ~w51839 & w51845;
assign w51908 = w51859 & w51907;
assign w51909 = ~w51906 & ~w51908;
assign w51910 = ~w51869 & ~w51871;
assign w51911 = ~w51909 & w51910;
assign w51912 = ~w51839 & ~w51859;
assign w51913 = ~w51845 & w51912;
assign w51914 = w51912 & w64079;
assign w51915 = w51877 & w51891;
assign w51916 = w51845 & ~w51852;
assign w51917 = w51839 & w51869;
assign w51918 = ~w51916 & w51917;
assign w51919 = w51900 & ~w51918;
assign w51920 = w51919 & w66895;
assign w51921 = ~w51911 & w51920;
assign w51922 = ~w51915 & w51921;
assign w51923 = ~w51904 & ~w51922;
assign w51924 = ~w51870 & ~w51923;
assign w51925 = ~pi2745 & w51924;
assign w51926 = pi2745 & ~w51924;
assign w51927 = ~w51925 & ~w51926;
assign w51928 = ~w51275 & ~w51806;
assign w51929 = w51307 & w51928;
assign w51930 = ~w51674 & w51821;
assign w51931 = ~w51309 & ~w51930;
assign w51932 = ~w51282 & ~w51673;
assign w51933 = w51928 & ~w51932;
assign w51934 = ~w51825 & ~w51933;
assign w51935 = ~w51931 & w51934;
assign w51936 = w51319 & ~w51935;
assign w51937 = (~w51326 & w51325) | (~w51326 & w66896) | (w51325 & w66896);
assign w51938 = ~w51289 & w51309;
assign w51939 = ~w51937 & ~w51938;
assign w51940 = ~w51319 & ~w51939;
assign w51941 = (~w51929 & ~w51339) | (~w51929 & w66897) | (~w51339 & w66897);
assign w51942 = ~w51940 & w51941;
assign w51943 = ~w51936 & w51942;
assign w51944 = pi2723 & ~w51943;
assign w51945 = ~pi2723 & w51943;
assign w51946 = ~w51944 & ~w51945;
assign w51947 = w51510 & ~w51528;
assign w51948 = ~w51514 & ~w51697;
assign w51949 = w51478 & w51948;
assign w51950 = w51487 & ~w51947;
assign w51951 = ~w51949 & w51950;
assign w51952 = ~w51504 & w51700;
assign w51953 = w51466 & ~w51952;
assign w51954 = w51478 & w51514;
assign w51955 = ~w51486 & ~w51705;
assign w51956 = ~w51954 & w51955;
assign w51957 = ~w51953 & w51956;
assign w51958 = ~w51501 & ~w51688;
assign w51959 = ~w51489 & ~w51536;
assign w51960 = w51486 & w51959;
assign w51961 = w51509 & ~w51958;
assign w51962 = ~w51960 & w51961;
assign w51963 = (~w51962 & w51957) | (~w51962 & w66898) | (w51957 & w66898);
assign w51964 = ~pi2734 & w51963;
assign w51965 = pi2734 & ~w51963;
assign w51966 = ~w51964 & ~w51965;
assign w51967 = w51726 & ~w51774;
assign w51968 = ~w51752 & w51780;
assign w51969 = ~w51967 & ~w51968;
assign w51970 = w51720 & ~w51792;
assign w51971 = w51771 & ~w51970;
assign w51972 = ~w51727 & ~w51768;
assign w51973 = w51748 & ~w51972;
assign w51974 = w51773 & w51779;
assign w51975 = ~w51759 & ~w51974;
assign w51976 = ~w51973 & w51975;
assign w51977 = ~w51969 & w51976;
assign w51978 = ~w51971 & w51977;
assign w51979 = ~w51740 & ~w51774;
assign w51980 = ~w51783 & w51979;
assign w51981 = (~w51726 & w51769) | (~w51726 & w66899) | (w51769 & w66899);
assign w51982 = ~w51751 & w51981;
assign w51983 = w51748 & w51982;
assign w51984 = w51720 & w51763;
assign w51985 = ~w51739 & w51751;
assign w51986 = ~w51741 & ~w51985;
assign w51987 = ~w51747 & ~w51986;
assign w51988 = w51759 & ~w51786;
assign w51989 = ~w51984 & w51988;
assign w51990 = ~w51987 & w51989;
assign w51991 = ~w51980 & w51990;
assign w51992 = ~w51983 & w51991;
assign w51993 = ~w51978 & ~w51992;
assign w51994 = ~pi2724 & w51993;
assign w51995 = pi2724 & ~w51993;
assign w51996 = ~w51994 & ~w51995;
assign w51997 = ~w51852 & ~w51886;
assign w51998 = ~w51860 & w51997;
assign w51999 = w51997 & w66900;
assign w52000 = ~w51887 & w51892;
assign w52001 = ~w51862 & ~w52000;
assign w52002 = ~w51999 & w52001;
assign w52003 = ~w51861 & w51891;
assign w52004 = ~w51997 & w52003;
assign w52005 = (~w51900 & ~w52002) | (~w51900 & w66901) | (~w52002 & w66901);
assign w52006 = ~w51852 & w51908;
assign w52007 = w52001 & ~w52006;
assign w52008 = w51891 & ~w52007;
assign w52009 = ~w51869 & w51998;
assign w52010 = w51869 & ~w51871;
assign w52011 = ~w51890 & ~w52010;
assign w52012 = w52001 & w66902;
assign w52013 = ~w52006 & ~w52009;
assign w52014 = ~w52012 & w52013;
assign w52015 = w51900 & ~w52014;
assign w52016 = ~w52005 & ~w52008;
assign w52017 = ~w52015 & w52016;
assign w52018 = ~pi2730 & w52017;
assign w52019 = pi2730 & ~w52017;
assign w52020 = ~w52018 & ~w52019;
assign w52021 = w51608 & w51612;
assign w52022 = ~w51596 & w51643;
assign w52023 = ~w51632 & ~w52022;
assign w52024 = ~w51595 & ~w51626;
assign w52025 = ~w52023 & ~w52024;
assign w52026 = ~w51644 & ~w52025;
assign w52027 = w51604 & ~w52026;
assign w52028 = ~w51615 & ~w51656;
assign w52029 = w51631 & w52028;
assign w52030 = ~w51635 & ~w51638;
assign w52031 = ~w51604 & ~w52030;
assign w52032 = (w51626 & w52031) | (w51626 & w66903) | (w52031 & w66903);
assign w52033 = w51652 & ~w52028;
assign w52034 = ~w52022 & w52033;
assign w52035 = ~w51588 & w51614;
assign w52036 = ~w51604 & ~w51631;
assign w52037 = ~w52035 & w52036;
assign w52038 = ~w52034 & ~w52037;
assign w52039 = ~w51626 & ~w52038;
assign w52040 = w51587 & w51653;
assign w52041 = ~w52021 & ~w52040;
assign w52042 = ~w52032 & w52041;
assign w52043 = ~w52039 & w52042;
assign w52044 = ~w52027 & w52043;
assign w52045 = pi2727 & ~w52044;
assign w52046 = ~pi2727 & w52044;
assign w52047 = ~w52045 & ~w52046;
assign w52048 = ~w51479 & w51688;
assign w52049 = ~w51948 & ~w51952;
assign w52050 = (w51486 & ~w51948) | (w51486 & w66904) | (~w51948 & w66904);
assign w52051 = ~w52049 & w52050;
assign w52052 = ~w51466 & ~w51488;
assign w52053 = w51504 & ~w52052;
assign w52054 = w51498 & w51500;
assign w52055 = ~w51486 & ~w51526;
assign w52056 = w51959 & w52055;
assign w52057 = ~w52054 & w52056;
assign w52058 = ~w52053 & w52057;
assign w52059 = ~w52051 & ~w52058;
assign w52060 = (w51696 & ~w51523) | (w51696 & w66905) | (~w51523 & w66905);
assign w52061 = (pi2743 & w52059) | (pi2743 & w66906) | (w52059 & w66906);
assign w52062 = ~w52059 & w66907;
assign w52063 = ~w52061 & ~w52062;
assign w52064 = w51792 & w66908;
assign w52065 = w51726 & ~w52064;
assign w52066 = ~w51733 & w51752;
assign w52067 = ~w51970 & ~w52066;
assign w52068 = w51981 & w52067;
assign w52069 = w51752 & w51774;
assign w52070 = w51768 & ~w51792;
assign w52071 = ~w52069 & ~w52070;
assign w52072 = (w52071 & w52068) | (w52071 & w66909) | (w52068 & w66909);
assign w52073 = w51759 & ~w52072;
assign w52074 = ~w51974 & ~w52064;
assign w52075 = ~w51759 & ~w52074;
assign w52076 = ~w51726 & w52071;
assign w52077 = ~w52075 & w52076;
assign w52078 = w51794 & w52071;
assign w52079 = w51726 & ~w51974;
assign w52080 = ~w52078 & w52079;
assign w52081 = ~w52077 & ~w52080;
assign w52082 = ~w52073 & ~w52081;
assign w52083 = ~pi2736 & w52082;
assign w52084 = pi2736 & ~w52082;
assign w52085 = ~w52083 & ~w52084;
assign w52086 = w51871 & ~w51876;
assign w52087 = ~w51879 & ~w51914;
assign w52088 = ~w52006 & w52087;
assign w52089 = w51878 & w51892;
assign w52090 = ~w51905 & ~w52089;
assign w52091 = w52010 & w52087;
assign w52092 = w52090 & w52091;
assign w52093 = (~w52086 & w52088) | (~w52086 & w66910) | (w52088 & w66910);
assign w52094 = ~w52092 & w52093;
assign w52095 = ~w51900 & ~w52094;
assign w52096 = ~w51869 & ~w52090;
assign w52097 = ~w51900 & ~w52096;
assign w52098 = ~w51875 & ~w52010;
assign w52099 = ~w51913 & ~w52098;
assign w52100 = ~w52003 & ~w52099;
assign w52101 = (~w51880 & w51874) | (~w51880 & w66911) | (w51874 & w66911);
assign w52102 = w52090 & w52101;
assign w52103 = ~w52100 & w52102;
assign w52104 = ~w52097 & ~w52103;
assign w52105 = ~w52095 & ~w52104;
assign w52106 = ~pi2756 & w52105;
assign w52107 = pi2756 & ~w52105;
assign w52108 = ~w52106 & ~w52107;
assign w52109 = ~w51604 & w51611;
assign w52110 = w51610 & w51612;
assign w52111 = ~w51610 & ~w51612;
assign w52112 = ~w52110 & ~w52111;
assign w52113 = w51628 & ~w51656;
assign w52114 = (~w52113 & w52112) | (~w52113 & w64080) | (w52112 & w64080);
assign w52115 = ~w51607 & ~w52112;
assign w52116 = ~w52114 & w52115;
assign w52117 = (w51626 & w52116) | (w51626 & w66912) | (w52116 & w66912);
assign w52118 = ~w51626 & ~w51659;
assign w52119 = w52114 & w52118;
assign w52120 = ~w51630 & w51643;
assign w52121 = w51618 & w52120;
assign w52122 = ~w52109 & ~w52121;
assign w52123 = ~w52119 & w52122;
assign w52124 = ~w52117 & w52123;
assign w52125 = pi2744 & ~w52124;
assign w52126 = ~pi2744 & w52124;
assign w52127 = ~w52125 & ~w52126;
assign w52128 = ~w51383 & w51398;
assign w52129 = ~w51414 & ~w52128;
assign w52130 = ~w51438 & ~w52129;
assign w52131 = (w51395 & ~w51386) | (w51395 & w64081) | (~w51386 & w64081);
assign w52132 = ~w51370 & ~w51377;
assign w52133 = w51407 & ~w52132;
assign w52134 = w52131 & ~w52133;
assign w52135 = w51384 & w51396;
assign w52136 = ~w51377 & w51404;
assign w52137 = ~w51395 & ~w52135;
assign w52138 = ~w52136 & w52137;
assign w52139 = ~w52134 & ~w52138;
assign w52140 = ~w51385 & ~w51435;
assign w52141 = ~w51425 & w52140;
assign w52142 = ~w51388 & ~w52139;
assign w52143 = (w51395 & ~w51405) | (w51395 & w66913) | (~w51405 & w66913);
assign w52144 = ~w51397 & w52143;
assign w52145 = w51409 & ~w51430;
assign w52146 = ~w51395 & ~w52145;
assign w52147 = ~w52144 & ~w52146;
assign w52148 = ~w51414 & ~w51442;
assign w52149 = w51386 & ~w52148;
assign w52150 = w52140 & w66914;
assign w52151 = ~w52149 & w52150;
assign w52152 = ~w52147 & w52151;
assign w52153 = ~w51422 & ~w52152;
assign w52154 = (w52142 & w66915) | (w52142 & w66916) | (w66915 & w66916);
assign w52155 = ~w52153 & w52154;
assign w52156 = ~pi2737 & w52155;
assign w52157 = pi2737 & ~w52155;
assign w52158 = ~w52156 & ~w52157;
assign w52159 = ~pi6275 & pi9040;
assign w52160 = ~pi6144 & ~pi9040;
assign w52161 = ~w52159 & ~w52160;
assign w52162 = pi2710 & ~w52161;
assign w52163 = ~pi2710 & w52161;
assign w52164 = ~w52162 & ~w52163;
assign w52165 = ~pi5960 & pi9040;
assign w52166 = ~pi6032 & ~pi9040;
assign w52167 = ~w52165 & ~w52166;
assign w52168 = pi2705 & ~w52167;
assign w52169 = ~pi2705 & w52167;
assign w52170 = ~w52168 & ~w52169;
assign w52171 = ~w52164 & ~w52170;
assign w52172 = ~pi6241 & pi9040;
assign w52173 = ~pi6079 & ~pi9040;
assign w52174 = ~w52172 & ~w52173;
assign w52175 = pi2691 & ~w52174;
assign w52176 = ~pi2691 & w52174;
assign w52177 = ~w52175 & ~w52176;
assign w52178 = ~pi6042 & pi9040;
assign w52179 = ~pi6074 & ~pi9040;
assign w52180 = ~w52178 & ~w52179;
assign w52181 = pi2703 & ~w52180;
assign w52182 = ~pi2703 & w52180;
assign w52183 = ~w52181 & ~w52182;
assign w52184 = w52177 & w52183;
assign w52185 = ~pi6172 & pi9040;
assign w52186 = ~pi6086 & ~pi9040;
assign w52187 = ~w52185 & ~w52186;
assign w52188 = pi2683 & ~w52187;
assign w52189 = ~pi2683 & w52187;
assign w52190 = ~w52188 & ~w52189;
assign w52191 = w52184 & w52190;
assign w52192 = w52171 & w52191;
assign w52193 = ~w52177 & ~w52183;
assign w52194 = ~w52184 & ~w52193;
assign w52195 = ~w52164 & w52170;
assign w52196 = ~pi5991 & pi9040;
assign w52197 = ~pi6044 & ~pi9040;
assign w52198 = ~w52196 & ~w52197;
assign w52199 = pi2706 & ~w52198;
assign w52200 = ~pi2706 & w52198;
assign w52201 = ~w52199 & ~w52200;
assign w52202 = ~w52195 & w52201;
assign w52203 = w52164 & ~w52170;
assign w52204 = ~w52195 & ~w52203;
assign w52205 = ~w52202 & ~w52204;
assign w52206 = ~w52164 & w52183;
assign w52207 = w52164 & ~w52183;
assign w52208 = ~w52206 & ~w52207;
assign w52209 = w52170 & w52208;
assign w52210 = w52170 & w52183;
assign w52211 = w52164 & ~w52177;
assign w52212 = ~w52164 & w52177;
assign w52213 = ~w52211 & ~w52212;
assign w52214 = ~w52170 & ~w52213;
assign w52215 = w52170 & w52177;
assign w52216 = ~w52206 & ~w52215;
assign w52217 = (~w52210 & w52214) | (~w52210 & w64083) | (w52214 & w64083);
assign w52218 = (~w52205 & w52217) | (~w52205 & w66917) | (w52217 & w66917);
assign w52219 = w52194 & ~w52218;
assign w52220 = ~w52194 & ~w52205;
assign w52221 = ~w52190 & ~w52220;
assign w52222 = ~w52219 & w52221;
assign w52223 = ~w52170 & ~w52211;
assign w52224 = w52208 & ~w52223;
assign w52225 = w52201 & w52224;
assign w52226 = ~w52171 & w52201;
assign w52227 = ~w52224 & ~w52226;
assign w52228 = w52190 & ~w52225;
assign w52229 = ~w52227 & w52228;
assign w52230 = ~w52183 & w52202;
assign w52231 = w52213 & w52230;
assign w52232 = ~w52192 & ~w52231;
assign w52233 = ~w52229 & w52232;
assign w52234 = ~w52222 & w52233;
assign w52235 = ~pi2742 & w52234;
assign w52236 = pi2742 & ~w52234;
assign w52237 = ~w52235 & ~w52236;
assign w52238 = ~w51726 & ~w51790;
assign w52239 = ~w51775 & ~w52238;
assign w52240 = ~w51982 & ~w52239;
assign w52241 = (~w51726 & w51792) | (~w51726 & w66918) | (w51792 & w66918);
assign w52242 = ~w51748 & ~w51785;
assign w52243 = w51780 & w52242;
assign w52244 = w52241 & ~w52243;
assign w52245 = ~w51733 & ~w51785;
assign w52246 = ~w51968 & w52245;
assign w52247 = w51726 & ~w51985;
assign w52248 = ~w52246 & w52247;
assign w52249 = (w51759 & w52248) | (w51759 & w66919) | (w52248 & w66919);
assign w52250 = ~w51780 & w52241;
assign w52251 = w51747 & ~w51979;
assign w52252 = (w52251 & ~w52067) | (w52251 & w66920) | (~w52067 & w66920);
assign w52253 = w51760 & ~w51781;
assign w52254 = ~w52250 & w52253;
assign w52255 = ~w52252 & w52254;
assign w52256 = ~w52249 & ~w52255;
assign w52257 = ~w52240 & ~w52256;
assign w52258 = pi2749 & w52257;
assign w52259 = ~pi2749 & ~w52257;
assign w52260 = ~w52258 & ~w52259;
assign w52261 = ~w51605 & ~w51655;
assign w52262 = ~w51626 & ~w52261;
assign w52263 = (~w52028 & w51617) | (~w52028 & w66921) | (w51617 & w66921);
assign w52264 = ~w51629 & ~w51656;
assign w52265 = ~w51635 & w52264;
assign w52266 = ~w51626 & ~w52265;
assign w52267 = ~w52263 & ~w52266;
assign w52268 = ~w51604 & ~w52267;
assign w52269 = (~w51609 & w51640) | (~w51609 & w51610) | (w51640 & w51610);
assign w52270 = w52023 & ~w52269;
assign w52271 = w51650 & ~w51656;
assign w52272 = w51598 & w52271;
assign w52273 = ~w52021 & ~w52272;
assign w52274 = ~w52270 & w52273;
assign w52275 = w51626 & ~w52274;
assign w52276 = ~w51633 & ~w51661;
assign w52277 = ~w52262 & w52276;
assign w52278 = ~w52268 & ~w52275;
assign w52279 = (~pi2751 & ~w52278) | (~pi2751 & w66922) | (~w52278 & w66922);
assign w52280 = w52278 & w66923;
assign w52281 = ~w52279 & ~w52280;
assign w52282 = ~w52170 & ~w52183;
assign w52283 = ~w52210 & ~w52282;
assign w52284 = w52164 & w52283;
assign w52285 = ~w52195 & ~w52201;
assign w52286 = ~w52212 & w52285;
assign w52287 = ~w52284 & w52286;
assign w52288 = w52184 & w52287;
assign w52289 = w52193 & ~w52204;
assign w52290 = ~w52193 & w52204;
assign w52291 = ~w52289 & ~w52290;
assign w52292 = w52190 & ~w52202;
assign w52293 = ~w52291 & w52292;
assign w52294 = w52217 & ~w52285;
assign w52295 = ~w52217 & w66924;
assign w52296 = ~w52294 & ~w52295;
assign w52297 = ~w52190 & ~w52296;
assign w52298 = ~w52214 & ~w52289;
assign w52299 = w52225 & ~w52298;
assign w52300 = w52194 & ~w52203;
assign w52301 = w52190 & w52201;
assign w52302 = ~w52214 & w52301;
assign w52303 = ~w52300 & w52302;
assign w52304 = ~w52288 & ~w52293;
assign w52305 = ~w52299 & ~w52303;
assign w52306 = w52304 & w52305;
assign w52307 = ~w52297 & w52306;
assign w52308 = pi2733 & ~w52307;
assign w52309 = ~pi2733 & w52307;
assign w52310 = ~w52308 & ~w52309;
assign w52311 = ~w52298 & w52301;
assign w52312 = ~w52217 & w66925;
assign w52313 = ~w52201 & ~w52282;
assign w52314 = w52216 & w52313;
assign w52315 = ~w52312 & ~w52314;
assign w52316 = ~w52190 & ~w52315;
assign w52317 = w52191 & ~w52209;
assign w52318 = w52183 & w52212;
assign w52319 = ~w52190 & ~w52318;
assign w52320 = w52171 & w52183;
assign w52321 = ~w52215 & ~w52320;
assign w52322 = ~w52201 & ~w52319;
assign w52323 = ~w52321 & w52322;
assign w52324 = ~w52207 & ~w52319;
assign w52325 = w52201 & ~w52216;
assign w52326 = ~w52324 & w52325;
assign w52327 = ~w52311 & ~w52317;
assign w52328 = ~w52323 & ~w52326;
assign w52329 = w52327 & w52328;
assign w52330 = ~w52316 & w52329;
assign w52331 = pi2740 & ~w52330;
assign w52332 = ~pi2740 & w52330;
assign w52333 = ~w52331 & ~w52332;
assign w52334 = w52191 & w52203;
assign w52335 = w52164 & ~w52283;
assign w52336 = ~w52209 & ~w52335;
assign w52337 = w52201 & w52320;
assign w52338 = (~w52177 & ~w52336) | (~w52177 & w66926) | (~w52336 & w66926);
assign w52339 = ~w52201 & ~w52215;
assign w52340 = ~w52286 & w52339;
assign w52341 = ~w52338 & ~w52340;
assign w52342 = w52190 & ~w52341;
assign w52343 = w52226 & w52336;
assign w52344 = w52171 & w52193;
assign w52345 = ~w52287 & ~w52344;
assign w52346 = ~w52343 & w52345;
assign w52347 = ~w52190 & ~w52346;
assign w52348 = w52201 & w52212;
assign w52349 = w52336 & w66927;
assign w52350 = ~w52183 & ~w52201;
assign w52351 = w52215 & w52350;
assign w52352 = ~w52334 & ~w52351;
assign w52353 = ~w52349 & w52352;
assign w52354 = ~w52347 & w52353;
assign w52355 = (pi2746 & ~w52354) | (pi2746 & w66928) | (~w52354 & w66928);
assign w52356 = w52354 & w66929;
assign w52357 = ~w52355 & ~w52356;
assign w52358 = ~w51395 & ~w51427;
assign w52359 = w51364 & ~w51408;
assign w52360 = ~w52132 & w52359;
assign w52361 = (~w51395 & w52360) | (~w51395 & w66930) | (w52360 & w66930);
assign w52362 = ~w51442 & ~w51443;
assign w52363 = w52143 & ~w52362;
assign w52364 = ~w51387 & w52140;
assign w52365 = ~w52363 & w52364;
assign w52366 = (w51422 & ~w52365) | (w51422 & w66931) | (~w52365 & w66931);
assign w52367 = w51431 & ~w52360;
assign w52368 = ~w51425 & w51444;
assign w52369 = w52131 & w52368;
assign w52370 = ~w52367 & ~w52369;
assign w52371 = ~w51422 & ~w52370;
assign w52372 = w51412 & w51424;
assign w52373 = ~w51415 & ~w52358;
assign w52374 = ~w52372 & w52373;
assign w52375 = ~w52366 & w52374;
assign w52376 = ~w52371 & w52375;
assign w52377 = pi2752 & ~w52376;
assign w52378 = ~pi2752 & w52376;
assign w52379 = ~w52377 & ~w52378;
assign w52380 = w51869 & w51888;
assign w52381 = ~w51862 & ~w52380;
assign w52382 = w51900 & ~w52381;
assign w52383 = ~w51873 & ~w51912;
assign w52384 = w51852 & w51900;
assign w52385 = ~w52383 & w52384;
assign w52386 = ~w51872 & ~w52385;
assign w52387 = ~w51869 & ~w52386;
assign w52388 = ~w51907 & ~w51917;
assign w52389 = w51906 & w52388;
assign w52390 = w51881 & ~w52388;
assign w52391 = ~w51913 & ~w52089;
assign w52392 = ~w52389 & w52391;
assign w52393 = ~w52390 & w52392;
assign w52394 = ~w51900 & ~w52393;
assign w52395 = ~w51884 & ~w52387;
assign w52396 = ~w52382 & w52395;
assign w52397 = ~w52394 & w52396;
assign w52398 = pi2763 & ~w52397;
assign w52399 = ~pi2763 & w52397;
assign w52400 = ~w52398 & ~w52399;
assign w52401 = ~w51428 & w52362;
assign w52402 = w51395 & ~w52401;
assign w52403 = w51395 & ~w51399;
assign w52404 = w51396 & ~w52403;
assign w52405 = ~w52402 & ~w52404;
assign w52406 = ~w51422 & ~w52405;
assign w52407 = w51389 & w51395;
assign w52408 = w51371 & w51444;
assign w52409 = w51402 & ~w52408;
assign w52410 = ~w52407 & ~w52409;
assign w52411 = w51395 & w52132;
assign w52412 = ~w51364 & ~w52411;
assign w52413 = ~w51407 & ~w52412;
assign w52414 = w51384 & w51438;
assign w52415 = ~w51425 & ~w52135;
assign w52416 = ~w52414 & w52415;
assign w52417 = ~w52413 & w52416;
assign w52418 = w51422 & ~w52417;
assign w52419 = ~w52410 & ~w52418;
assign w52420 = ~w52406 & w52419;
assign w52421 = ~pi2774 & w52420;
assign w52422 = pi2774 & ~w52420;
assign w52423 = ~w52421 & ~w52422;
assign w52424 = ~pi6258 & pi9040;
assign w52425 = ~pi6379 & ~pi9040;
assign w52426 = ~w52424 & ~w52425;
assign w52427 = pi2738 & ~w52426;
assign w52428 = ~pi2738 & w52426;
assign w52429 = ~w52427 & ~w52428;
assign w52430 = ~pi6242 & pi9040;
assign w52431 = ~pi6384 & ~pi9040;
assign w52432 = ~w52430 & ~w52431;
assign w52433 = pi2754 & ~w52432;
assign w52434 = ~pi2754 & w52432;
assign w52435 = ~w52433 & ~w52434;
assign w52436 = ~w52429 & ~w52435;
assign w52437 = ~pi6279 & pi9040;
assign w52438 = ~pi6399 & ~pi9040;
assign w52439 = ~w52437 & ~w52438;
assign w52440 = pi2758 & ~w52439;
assign w52441 = ~pi2758 & w52439;
assign w52442 = ~w52440 & ~w52441;
assign w52443 = ~pi6228 & pi9040;
assign w52444 = ~pi6393 & ~pi9040;
assign w52445 = ~w52443 & ~w52444;
assign w52446 = pi2760 & ~w52445;
assign w52447 = ~pi2760 & w52445;
assign w52448 = ~w52446 & ~w52447;
assign w52449 = w52442 & ~w52448;
assign w52450 = w52436 & ~w52449;
assign w52451 = w52429 & w52435;
assign w52452 = ~w52436 & ~w52451;
assign w52453 = w52449 & w52452;
assign w52454 = ~w52450 & ~w52453;
assign w52455 = ~pi6248 & pi9040;
assign w52456 = ~pi6301 & ~pi9040;
assign w52457 = ~w52455 & ~w52456;
assign w52458 = pi2767 & ~w52457;
assign w52459 = ~pi2767 & w52457;
assign w52460 = ~w52458 & ~w52459;
assign w52461 = ~w52454 & w52460;
assign w52462 = ~pi6383 & pi9040;
assign w52463 = pi6387 & ~pi9040;
assign w52464 = ~w52462 & ~w52463;
assign w52465 = pi2765 & ~w52464;
assign w52466 = ~pi2765 & w52464;
assign w52467 = ~w52465 & ~w52466;
assign w52468 = w52435 & ~w52448;
assign w52469 = (~w52460 & ~w52468) | (~w52460 & w66932) | (~w52468 & w66932);
assign w52470 = ~w52442 & w52448;
assign w52471 = w52429 & ~w52435;
assign w52472 = w52470 & w52471;
assign w52473 = ~w52468 & ~w52472;
assign w52474 = w52469 & ~w52473;
assign w52475 = ~w52429 & w52448;
assign w52476 = ~w52468 & ~w52475;
assign w52477 = ~w52454 & w52476;
assign w52478 = ~w52442 & ~w52451;
assign w52479 = w52448 & w52460;
assign w52480 = w52435 & w52442;
assign w52481 = w52479 & ~w52480;
assign w52482 = ~w52478 & w52481;
assign w52483 = ~w52467 & ~w52482;
assign w52484 = ~w52474 & w52483;
assign w52485 = ~w52477 & w52484;
assign w52486 = ~w52442 & w52451;
assign w52487 = w52460 & ~w52486;
assign w52488 = w52429 & ~w52448;
assign w52489 = ~w52442 & w52488;
assign w52490 = ~w52487 & w52489;
assign w52491 = ~w52435 & ~w52442;
assign w52492 = ~w52475 & ~w52479;
assign w52493 = w52491 & ~w52492;
assign w52494 = w52442 & w52448;
assign w52495 = w52451 & w52494;
assign w52496 = w52467 & ~w52495;
assign w52497 = ~w52436 & ~w52475;
assign w52498 = ~w52494 & w52497;
assign w52499 = ~w52450 & ~w52460;
assign w52500 = ~w52498 & w52499;
assign w52501 = ~w52493 & w52496;
assign w52502 = ~w52490 & w52501;
assign w52503 = ~w52500 & w52502;
assign w52504 = ~w52485 & ~w52503;
assign w52505 = ~w52449 & ~w52470;
assign w52506 = w52435 & ~w52460;
assign w52507 = w52505 & w52506;
assign w52508 = ~w52461 & ~w52507;
assign w52509 = ~w52504 & w52508;
assign w52510 = ~pi2790 & w52509;
assign w52511 = pi2790 & ~w52509;
assign w52512 = ~w52510 & ~w52511;
assign w52513 = ~pi6385 & pi9040;
assign w52514 = ~pi6242 & ~pi9040;
assign w52515 = ~w52513 & ~w52514;
assign w52516 = pi2776 & ~w52515;
assign w52517 = ~pi2776 & w52515;
assign w52518 = ~w52516 & ~w52517;
assign w52519 = ~pi6181 & pi9040;
assign w52520 = ~pi6188 & ~pi9040;
assign w52521 = ~w52519 & ~w52520;
assign w52522 = pi2765 & ~w52521;
assign w52523 = ~pi2765 & w52521;
assign w52524 = ~w52522 & ~w52523;
assign w52525 = ~w52518 & w52524;
assign w52526 = ~pi6407 & pi9040;
assign w52527 = ~pi6302 & ~pi9040;
assign w52528 = ~w52526 & ~w52527;
assign w52529 = pi2738 & ~w52528;
assign w52530 = ~pi2738 & w52528;
assign w52531 = ~w52529 & ~w52530;
assign w52532 = ~pi6240 & pi9040;
assign w52533 = ~pi6231 & ~pi9040;
assign w52534 = ~w52532 & ~w52533;
assign w52535 = pi2780 & ~w52534;
assign w52536 = ~pi2780 & w52534;
assign w52537 = ~w52535 & ~w52536;
assign w52538 = w52531 & w52537;
assign w52539 = ~pi6366 & pi9040;
assign w52540 = ~pi6365 & ~pi9040;
assign w52541 = ~w52539 & ~w52540;
assign w52542 = pi2766 & ~w52541;
assign w52543 = ~pi2766 & w52541;
assign w52544 = ~w52542 & ~w52543;
assign w52545 = ~w52538 & ~w52544;
assign w52546 = ~w52538 & w64084;
assign w52547 = w52525 & w52546;
assign w52548 = ~pi6243 & pi9040;
assign w52549 = ~pi6248 & ~pi9040;
assign w52550 = ~w52548 & ~w52549;
assign w52551 = pi2779 & ~w52550;
assign w52552 = ~pi2779 & w52550;
assign w52553 = ~w52551 & ~w52552;
assign w52554 = ~w52524 & ~w52537;
assign w52555 = w52518 & w52554;
assign w52556 = w52545 & ~w52555;
assign w52557 = w52524 & ~w52531;
assign w52558 = w52518 & w52557;
assign w52559 = w52557 & w66933;
assign w52560 = ~w52531 & w52537;
assign w52561 = ~w52524 & w52560;
assign w52562 = (w52544 & ~w52560) | (w52544 & w66934) | (~w52560 & w66934);
assign w52563 = ~w52559 & w52562;
assign w52564 = ~w52556 & ~w52563;
assign w52565 = ~w52518 & ~w52537;
assign w52566 = w52531 & w52565;
assign w52567 = (w52544 & ~w52565) | (w52544 & w53412) | (~w52565 & w53412);
assign w52568 = w52525 & ~w52567;
assign w52569 = w52518 & w52537;
assign w52570 = w52524 & w52531;
assign w52571 = w52569 & w52570;
assign w52572 = ~w52568 & ~w52571;
assign w52573 = ~w52564 & w52572;
assign w52574 = ~w52553 & ~w52573;
assign w52575 = ~w52524 & ~w52531;
assign w52576 = ~w52565 & ~w52569;
assign w52577 = w52575 & ~w52576;
assign w52578 = w52518 & w52531;
assign w52579 = ~w52524 & w52578;
assign w52580 = w52525 & w52537;
assign w52581 = ~w52579 & ~w52580;
assign w52582 = ~w52538 & ~w52581;
assign w52583 = (w52544 & w52582) | (w52544 & w66935) | (w52582 & w66935);
assign w52584 = w52537 & w52579;
assign w52585 = ~w52544 & ~w52584;
assign w52586 = ~w52518 & w52575;
assign w52587 = ~w52558 & ~w52586;
assign w52588 = w52585 & w52587;
assign w52589 = w52557 & w52565;
assign w52590 = ~w52525 & w52531;
assign w52591 = ~w52537 & w52590;
assign w52592 = w52544 & ~w52589;
assign w52593 = w52581 & w52592;
assign w52594 = ~w52591 & w52593;
assign w52595 = w52553 & ~w52588;
assign w52596 = ~w52594 & w52595;
assign w52597 = ~w52547 & ~w52583;
assign w52598 = ~w52574 & w52597;
assign w52599 = ~w52596 & w52598;
assign w52600 = pi2791 & ~w52599;
assign w52601 = ~pi2791 & w52599;
assign w52602 = ~w52600 & ~w52601;
assign w52603 = ~w52475 & ~w52488;
assign w52604 = ~w52442 & w52603;
assign w52605 = w52603 & w64085;
assign w52606 = w52460 & ~w52605;
assign w52607 = w52471 & w52606;
assign w52608 = w52452 & ~w52494;
assign w52609 = (w52460 & w52505) | (w52460 & w66936) | (w52505 & w66936);
assign w52610 = ~w52608 & ~w52609;
assign w52611 = w52471 & w52494;
assign w52612 = w52480 & ~w52603;
assign w52613 = ~w52611 & ~w52612;
assign w52614 = ~w52604 & w52613;
assign w52615 = w52468 & ~w52614;
assign w52616 = w52467 & ~w52610;
assign w52617 = ~w52607 & w52616;
assign w52618 = ~w52615 & w52617;
assign w52619 = w52442 & ~w52476;
assign w52620 = w52449 & w52471;
assign w52621 = w52460 & ~w52620;
assign w52622 = (~w52460 & ~w52491) | (~w52460 & w64086) | (~w52491 & w64086);
assign w52623 = (w52476 & w52621) | (w52476 & w66937) | (w52621 & w66937);
assign w52624 = ~w52619 & ~w52623;
assign w52625 = ~w52454 & ~w52624;
assign w52626 = ~w52479 & ~w52489;
assign w52627 = w52435 & ~w52626;
assign w52628 = ~w52467 & ~w52472;
assign w52629 = ~w52627 & w52628;
assign w52630 = ~w52625 & w52629;
assign w52631 = ~w52618 & ~w52630;
assign w52632 = pi2798 & w52631;
assign w52633 = ~pi2798 & ~w52631;
assign w52634 = ~w52632 & ~w52633;
assign w52635 = ~pi6283 & pi9040;
assign w52636 = ~pi6177 & ~pi9040;
assign w52637 = ~w52635 & ~w52636;
assign w52638 = pi2762 & ~w52637;
assign w52639 = ~pi2762 & w52637;
assign w52640 = ~w52638 & ~w52639;
assign w52641 = ~pi6320 & pi9040;
assign w52642 = ~pi6274 & ~pi9040;
assign w52643 = ~w52641 & ~w52642;
assign w52644 = pi2773 & ~w52643;
assign w52645 = ~pi2773 & w52643;
assign w52646 = ~w52644 & ~w52645;
assign w52647 = w52640 & ~w52646;
assign w52648 = ~pi6537 & pi9040;
assign w52649 = ~pi6227 & ~pi9040;
assign w52650 = ~w52648 & ~w52649;
assign w52651 = pi2781 & ~w52650;
assign w52652 = ~pi2781 & w52650;
assign w52653 = ~w52651 & ~w52652;
assign w52654 = ~pi6262 & pi9040;
assign w52655 = ~pi6538 & ~pi9040;
assign w52656 = ~w52654 & ~w52655;
assign w52657 = pi2757 & ~w52656;
assign w52658 = ~pi2757 & w52656;
assign w52659 = ~w52657 & ~w52658;
assign w52660 = w52653 & ~w52659;
assign w52661 = w52647 & w52660;
assign w52662 = ~w52653 & w52659;
assign w52663 = ~w52646 & w52662;
assign w52664 = ~w52661 & ~w52663;
assign w52665 = ~pi6276 & pi9040;
assign w52666 = ~pi6303 & ~pi9040;
assign w52667 = ~w52665 & ~w52666;
assign w52668 = pi2782 & ~w52667;
assign w52669 = ~pi2782 & w52667;
assign w52670 = ~w52668 & ~w52669;
assign w52671 = w52640 & w52670;
assign w52672 = ~w52664 & w52671;
assign w52673 = ~pi6470 & pi9040;
assign w52674 = ~pi6247 & ~pi9040;
assign w52675 = ~w52673 & ~w52674;
assign w52676 = pi2777 & ~w52675;
assign w52677 = ~pi2777 & w52675;
assign w52678 = ~w52676 & ~w52677;
assign w52679 = ~w52672 & w52678;
assign w52680 = ~w52653 & ~w52670;
assign w52681 = w52640 & w52659;
assign w52682 = ~w52647 & w52680;
assign w52683 = ~w52681 & w52682;
assign w52684 = w52653 & w52670;
assign w52685 = ~w52640 & w52646;
assign w52686 = ~w52659 & ~w52685;
assign w52687 = ~w52647 & ~w52686;
assign w52688 = ~w52686 & w66938;
assign w52689 = w52664 & ~w52683;
assign w52690 = ~w52688 & w52689;
assign w52691 = ~w52679 & ~w52690;
assign w52692 = w52646 & ~w52662;
assign w52693 = w52681 & w52692;
assign w52694 = (~w52680 & ~w52692) | (~w52680 & w66939) | (~w52692 & w66939);
assign w52695 = (~w52694 & ~w52689) | (~w52694 & w66940) | (~w52689 & w66940);
assign w52696 = ~w52640 & ~w52659;
assign w52697 = ~w52692 & ~w52696;
assign w52698 = w52660 & w52685;
assign w52699 = ~w52697 & ~w52698;
assign w52700 = (w52678 & w52699) | (w52678 & w66941) | (w52699 & w66941);
assign w52701 = ~w52695 & w52700;
assign w52702 = ~w52661 & ~w52693;
assign w52703 = ~w52646 & w52653;
assign w52704 = ~w52640 & w52659;
assign w52705 = w52703 & w52704;
assign w52706 = w52702 & ~w52705;
assign w52707 = ~w52640 & ~w52646;
assign w52708 = ~w52670 & ~w52707;
assign w52709 = w52640 & ~w52653;
assign w52710 = w52708 & ~w52709;
assign w52711 = ~w52703 & w52704;
assign w52712 = w52710 & ~w52711;
assign w52713 = ~w52653 & w52696;
assign w52714 = ~w52708 & ~w52713;
assign w52715 = ~w52712 & ~w52714;
assign w52716 = ~w52646 & ~w52670;
assign w52717 = w52706 & w52716;
assign w52718 = ~w52715 & w52717;
assign w52719 = ~w52691 & ~w52701;
assign w52720 = ~w52718 & w52719;
assign w52721 = pi2787 & w52720;
assign w52722 = ~pi2787 & ~w52720;
assign w52723 = ~w52721 & ~w52722;
assign w52724 = w52435 & ~w52603;
assign w52725 = ~w52619 & w52622;
assign w52726 = ~w52724 & w52725;
assign w52727 = (w52613 & w52726) | (w52613 & w64087) | (w52726 & w64087);
assign w52728 = ~w52467 & ~w52727;
assign w52729 = (~w52622 & ~w52613) | (~w52622 & w64088) | (~w52613 & w64088);
assign w52730 = w52613 & w66942;
assign w52731 = w52467 & ~w52729;
assign w52732 = ~w52730 & w52731;
assign w52733 = ~w52470 & ~w52497;
assign w52734 = w52487 & ~w52733;
assign w52735 = w52491 & ~w52603;
assign w52736 = w52469 & ~w52735;
assign w52737 = ~w52735 & w66943;
assign w52738 = ~w52734 & ~w52737;
assign w52739 = w52475 & w52480;
assign w52740 = ~w52451 & w52469;
assign w52741 = ~w52507 & ~w52621;
assign w52742 = ~w52467 & ~w52739;
assign w52743 = (w52742 & ~w52741) | (w52742 & w66944) | (~w52741 & w66944);
assign w52744 = ~w52738 & w52743;
assign w52745 = w52436 & w52449;
assign w52746 = ~w52744 & w52745;
assign w52747 = ~w52728 & ~w52732;
assign w52748 = w52747 & w66945;
assign w52749 = (~pi2806 & ~w52747) | (~pi2806 & w66946) | (~w52747 & w66946);
assign w52750 = ~w52748 & ~w52749;
assign w52751 = ~pi6177 & pi9040;
assign w52752 = ~pi6246 & ~pi9040;
assign w52753 = ~w52751 & ~w52752;
assign w52754 = pi2753 & ~w52753;
assign w52755 = ~pi2753 & w52753;
assign w52756 = ~w52754 & ~w52755;
assign w52757 = ~pi6472 & pi9040;
assign w52758 = ~pi6373 & ~pi9040;
assign w52759 = ~w52757 & ~w52758;
assign w52760 = pi2775 & ~w52759;
assign w52761 = ~pi2775 & w52759;
assign w52762 = ~w52760 & ~w52761;
assign w52763 = ~pi6255 & pi9040;
assign w52764 = ~pi6310 & ~pi9040;
assign w52765 = ~w52763 & ~w52764;
assign w52766 = pi2778 & ~w52765;
assign w52767 = ~pi2778 & w52765;
assign w52768 = ~w52766 & ~w52767;
assign w52769 = w52762 & w52768;
assign w52770 = ~pi6245 & pi9040;
assign w52771 = ~pi6470 & ~pi9040;
assign w52772 = ~w52770 & ~w52771;
assign w52773 = pi2779 & ~w52772;
assign w52774 = ~pi2779 & w52772;
assign w52775 = ~w52773 & ~w52774;
assign w52776 = ~w52768 & w52775;
assign w52777 = ~pi6392 & pi9040;
assign w52778 = ~pi6269 & ~pi9040;
assign w52779 = ~w52777 & ~w52778;
assign w52780 = pi2741 & ~w52779;
assign w52781 = ~pi2741 & w52779;
assign w52782 = ~w52780 & ~w52781;
assign w52783 = ~pi6469 & pi9040;
assign w52784 = ~pi6262 & ~pi9040;
assign w52785 = ~w52783 & ~w52784;
assign w52786 = pi2780 & ~w52785;
assign w52787 = ~pi2780 & w52785;
assign w52788 = ~w52786 & ~w52787;
assign w52789 = w52782 & w52788;
assign w52790 = ~w52782 & ~w52788;
assign w52791 = ~w52789 & ~w52790;
assign w52792 = ~w52768 & w52791;
assign w52793 = ~w52775 & ~w52782;
assign w52794 = w52775 & w52782;
assign w52795 = ~w52793 & ~w52794;
assign w52796 = w52791 & w52795;
assign w52797 = w52762 & w52796;
assign w52798 = w52796 & w63332;
assign w52799 = (~w52776 & w52798) | (~w52776 & w63438) | (w52798 & w63438);
assign w52800 = ~w52791 & ~w52794;
assign w52801 = ~w52762 & ~w52788;
assign w52802 = w52794 & w52801;
assign w52803 = ~w52775 & ~w52801;
assign w52804 = ~w52802 & ~w52803;
assign w52805 = w52768 & ~w52804;
assign w52806 = w52800 & w52805;
assign w52807 = w52762 & w52790;
assign w52808 = w52776 & w52807;
assign w52809 = ~w52802 & ~w52808;
assign w52810 = ~w52806 & w52809;
assign w52811 = (w52769 & ~w52810) | (w52769 & w63439) | (~w52810 & w63439);
assign w52812 = ~w52775 & w52788;
assign w52813 = ~w52762 & ~w52782;
assign w52814 = w52812 & w52813;
assign w52815 = w52762 & ~w52775;
assign w52816 = (~w52788 & w52815) | (~w52788 & w64089) | (w52815 & w64089);
assign w52817 = ~w52776 & ~w52816;
assign w52818 = ~w52762 & ~w52768;
assign w52819 = w52817 & w52818;
assign w52820 = ~w52762 & w52768;
assign w52821 = ~w52801 & ~w52820;
assign w52822 = w52794 & ~w52821;
assign w52823 = ~w52808 & ~w52814;
assign w52824 = ~w52822 & w52823;
assign w52825 = (~w52756 & w52811) | (~w52756 & w64090) | (w52811 & w64090);
assign w52826 = w52782 & w52815;
assign w52827 = ~w52813 & ~w52826;
assign w52828 = w52792 & ~w52827;
assign w52829 = w52769 & w52793;
assign w52830 = w52776 & ~w52788;
assign w52831 = w52762 & w52789;
assign w52832 = w52788 & w52795;
assign w52833 = w52795 & w63440;
assign w52834 = ~w52831 & ~w52833;
assign w52835 = ~w52762 & w52775;
assign w52836 = ~w52815 & ~w52835;
assign w52837 = ~w52768 & ~w52812;
assign w52838 = w52836 & w52837;
assign w52839 = w52834 & ~w52838;
assign w52840 = w52795 & ~w52821;
assign w52841 = w52834 & w64091;
assign w52842 = (~w52829 & w52817) | (~w52829 & w66947) | (w52817 & w66947);
assign w52843 = ~w52841 & w52842;
assign w52844 = (w52756 & w52841) | (w52756 & w66948) | (w52841 & w66948);
assign w52845 = w52776 & w52831;
assign w52846 = w52768 & w52775;
assign w52847 = w52801 & w52846;
assign w52848 = ~w52845 & ~w52847;
assign w52849 = ~w52828 & w52848;
assign w52850 = ~w52844 & w52849;
assign w52851 = (~pi2795 & w52825) | (~pi2795 & w66949) | (w52825 & w66949);
assign w52852 = ~w52825 & w66950;
assign w52853 = ~w52851 & ~w52852;
assign w52854 = w52684 & w52696;
assign w52855 = w52647 & w52662;
assign w52856 = w52670 & ~w52855;
assign w52857 = ~w52661 & ~w52670;
assign w52858 = ~w52711 & w52857;
assign w52859 = ~w52856 & ~w52858;
assign w52860 = w52640 & ~w52660;
assign w52861 = w52692 & w52860;
assign w52862 = ~w52854 & ~w52861;
assign w52863 = ~w52859 & w66951;
assign w52864 = w52646 & w52670;
assign w52865 = ~w52659 & w52671;
assign w52866 = ~w52713 & ~w52865;
assign w52867 = ~w52864 & ~w52866;
assign w52868 = w52681 & w52716;
assign w52869 = ~w52678 & ~w52698;
assign w52870 = w52659 & ~w52855;
assign w52871 = ~w52699 & w66952;
assign w52872 = ~w52868 & w52869;
assign w52873 = ~w52867 & w52872;
assign w52874 = ~w52871 & w52873;
assign w52875 = ~w52863 & ~w52874;
assign w52876 = ~w52646 & w52688;
assign w52877 = w52713 & w52716;
assign w52878 = ~w52670 & w52861;
assign w52879 = w52660 & w52864;
assign w52880 = ~w52877 & ~w52879;
assign w52881 = ~w52878 & w52880;
assign w52882 = ~w52876 & w52881;
assign w52883 = ~w52875 & w52882;
assign w52884 = pi2803 & ~w52883;
assign w52885 = ~pi2803 & w52883;
assign w52886 = ~w52884 & ~w52885;
assign w52887 = w52662 & w52685;
assign w52888 = w52670 & ~w52887;
assign w52889 = ~w52660 & ~w52662;
assign w52890 = w52707 & w52889;
assign w52891 = w52888 & ~w52890;
assign w52892 = ~w52857 & ~w52891;
assign w52893 = w52716 & ~w52889;
assign w52894 = ~w52684 & ~w52865;
assign w52895 = ~w52660 & ~w52681;
assign w52896 = ~w52894 & w52895;
assign w52897 = w52708 & w52713;
assign w52898 = w52678 & ~w52893;
assign w52899 = ~w52897 & w52898;
assign w52900 = w52702 & ~w52896;
assign w52901 = w52899 & w52900;
assign w52902 = w52681 & w52684;
assign w52903 = ~w52855 & ~w52879;
assign w52904 = ~w52902 & w52903;
assign w52905 = w52869 & w52904;
assign w52906 = ~w52715 & w52905;
assign w52907 = ~w52901 & ~w52906;
assign w52908 = ~w52892 & ~w52907;
assign w52909 = ~pi2785 & w52908;
assign w52910 = pi2785 & ~w52908;
assign w52911 = ~w52909 & ~w52910;
assign w52912 = ~pi6227 & pi9040;
assign w52913 = ~pi6392 & ~pi9040;
assign w52914 = ~w52912 & ~w52913;
assign w52915 = pi2768 & ~w52914;
assign w52916 = ~pi2768 & w52914;
assign w52917 = ~w52915 & ~w52916;
assign w52918 = ~pi6244 & pi9040;
assign w52919 = ~pi6283 & ~pi9040;
assign w52920 = ~w52918 & ~w52919;
assign w52921 = pi2753 & ~w52920;
assign w52922 = ~pi2753 & w52920;
assign w52923 = ~w52921 & ~w52922;
assign w52924 = ~pi6538 & pi9040;
assign w52925 = ~pi6245 & ~pi9040;
assign w52926 = ~w52924 & ~w52925;
assign w52927 = pi2772 & ~w52926;
assign w52928 = ~pi2772 & w52926;
assign w52929 = ~w52927 & ~w52928;
assign w52930 = ~w52923 & w52929;
assign w52931 = ~pi6246 & pi9040;
assign w52932 = ~pi6320 & ~pi9040;
assign w52933 = ~w52931 & ~w52932;
assign w52934 = pi2741 & ~w52933;
assign w52935 = ~pi2741 & w52933;
assign w52936 = ~w52934 & ~w52935;
assign w52937 = w52930 & ~w52936;
assign w52938 = ~pi6373 & pi9040;
assign w52939 = ~pi6474 & ~pi9040;
assign w52940 = ~w52938 & ~w52939;
assign w52941 = pi2769 & ~w52940;
assign w52942 = ~pi2769 & w52940;
assign w52943 = ~w52941 & ~w52942;
assign w52944 = w52936 & ~w52943;
assign w52945 = w52923 & w52929;
assign w52946 = w52944 & w52945;
assign w52947 = ~w52936 & w52943;
assign w52948 = ~w52923 & ~w52947;
assign w52949 = ~pi6267 & pi9040;
assign w52950 = ~pi6276 & ~pi9040;
assign w52951 = ~w52949 & ~w52950;
assign w52952 = pi2759 & ~w52951;
assign w52953 = ~pi2759 & w52951;
assign w52954 = ~w52952 & ~w52953;
assign w52955 = w52929 & ~w52943;
assign w52956 = ~w52936 & w52955;
assign w52957 = w52923 & w52947;
assign w52958 = ~w52956 & ~w52957;
assign w52959 = ~w52948 & ~w52954;
assign w52960 = w52958 & w52959;
assign w52961 = ~w52937 & ~w52946;
assign w52962 = ~w52960 & w52961;
assign w52963 = ~w52917 & ~w52962;
assign w52964 = w52930 & w52947;
assign w52965 = ~w52936 & ~w52943;
assign w52966 = w52923 & w52965;
assign w52967 = w52917 & ~w52944;
assign w52968 = ~w52966 & w52967;
assign w52969 = w52917 & w52936;
assign w52970 = ~w52930 & w52969;
assign w52971 = w52948 & ~w52955;
assign w52972 = ~w52917 & ~w52971;
assign w52973 = ~w52968 & ~w52970;
assign w52974 = ~w52972 & w52973;
assign w52975 = (~w52917 & ~w52947) | (~w52917 & w66953) | (~w52947 & w66953);
assign w52976 = w52923 & ~w52929;
assign w52977 = ~w52975 & w52976;
assign w52978 = w52923 & w52943;
assign w52979 = w52969 & w52978;
assign w52980 = w52954 & ~w52964;
assign w52981 = ~w52979 & w52980;
assign w52982 = ~w52977 & w52981;
assign w52983 = ~w52974 & w52982;
assign w52984 = ~w52944 & ~w52947;
assign w52985 = w52945 & ~w52984;
assign w52986 = ~w52954 & ~w52985;
assign w52987 = w52930 & w52965;
assign w52988 = w52917 & ~w52955;
assign w52989 = w52948 & w52988;
assign w52990 = ~w52987 & ~w52989;
assign w52991 = w52986 & w52990;
assign w52992 = ~w52983 & ~w52991;
assign w52993 = ~w52963 & ~w52992;
assign w52994 = ~pi2789 & w52993;
assign w52995 = pi2789 & ~w52993;
assign w52996 = ~w52994 & ~w52995;
assign w52997 = w52812 & ~w52843;
assign w52998 = ~w52788 & ~w52795;
assign w52999 = ~w52814 & ~w52998;
assign w53000 = ~w52768 & ~w52999;
assign w53001 = ~w52791 & w52846;
assign w53002 = ~w52756 & ~w53001;
assign w53003 = ~w52797 & w53002;
assign w53004 = ~w53000 & w53003;
assign w53005 = w52756 & ~w52805;
assign w53006 = w52839 & w53005;
assign w53007 = ~w53004 & ~w53006;
assign w53008 = ~w52997 & ~w53007;
assign w53009 = pi2794 & w53008;
assign w53010 = ~pi2794 & ~w53008;
assign w53011 = ~w53009 & ~w53010;
assign w53012 = ~pi6188 & pi9040;
assign w53013 = ~pi6228 & ~pi9040;
assign w53014 = ~w53012 & ~w53013;
assign w53015 = pi2771 & ~w53014;
assign w53016 = ~pi2771 & w53014;
assign w53017 = ~w53015 & ~w53016;
assign w53018 = ~pi6384 & pi9040;
assign w53019 = ~pi6381 & ~pi9040;
assign w53020 = ~w53018 & ~w53019;
assign w53021 = pi2754 & ~w53020;
assign w53022 = ~pi2754 & w53020;
assign w53023 = ~w53021 & ~w53022;
assign w53024 = w53017 & w53023;
assign w53025 = ~pi6398 & pi9040;
assign w53026 = ~pi6279 & ~pi9040;
assign w53027 = ~w53025 & ~w53026;
assign w53028 = pi2761 & ~w53027;
assign w53029 = ~pi2761 & w53027;
assign w53030 = ~w53028 & ~w53029;
assign w53031 = ~pi6400 & pi9040;
assign w53032 = ~pi6243 & ~pi9040;
assign w53033 = ~w53031 & ~w53032;
assign w53034 = pi2764 & ~w53033;
assign w53035 = ~pi2764 & w53033;
assign w53036 = ~w53034 & ~w53035;
assign w53037 = ~w53030 & ~w53036;
assign w53038 = w53024 & w53037;
assign w53039 = ~pi6234 & pi9040;
assign w53040 = ~pi6385 & ~pi9040;
assign w53041 = ~w53039 & ~w53040;
assign w53042 = pi2755 & ~w53041;
assign w53043 = ~pi2755 & w53041;
assign w53044 = ~w53042 & ~w53043;
assign w53045 = w53036 & ~w53044;
assign w53046 = ~w53017 & ~w53023;
assign w53047 = w53045 & w53046;
assign w53048 = ~w53038 & ~w53047;
assign w53049 = ~w53023 & w53030;
assign w53050 = w53036 & w53049;
assign w53051 = ~w53036 & w53044;
assign w53052 = ~w53045 & ~w53051;
assign w53053 = ~w53023 & ~w53044;
assign w53054 = w53023 & ~w53030;
assign w53055 = ~w53049 & ~w53054;
assign w53056 = w53036 & w53055;
assign w53057 = (~w53053 & ~w53055) | (~w53053 & w63441) | (~w53055 & w63441);
assign w53058 = (~w53050 & ~w53057) | (~w53050 & w64092) | (~w53057 & w64092);
assign w53059 = ~w53048 & ~w53058;
assign w53060 = ~pi6387 & pi9040;
assign w53061 = ~pi6240 & ~pi9040;
assign w53062 = ~w53060 & ~w53061;
assign w53063 = pi2760 & ~w53062;
assign w53064 = ~pi2760 & w53062;
assign w53065 = ~w53063 & ~w53064;
assign w53066 = w53030 & ~w53044;
assign w53067 = w53036 & w53066;
assign w53068 = ~w53017 & ~w53055;
assign w53069 = ~w53030 & w53036;
assign w53070 = ~w53017 & w53069;
assign w53071 = w53017 & ~w53036;
assign w53072 = ~w53049 & w53071;
assign w53073 = ~w53067 & ~w53070;
assign w53074 = ~w53072 & w53073;
assign w53075 = ~w53068 & w53074;
assign w53076 = ~w53065 & ~w53075;
assign w53077 = w53051 & w53055;
assign w53078 = w53017 & w53067;
assign w53079 = ~w53036 & ~w53044;
assign w53080 = w53054 & w53079;
assign w53081 = ~w53023 & w53066;
assign w53082 = ~w53038 & w53065;
assign w53083 = ~w53070 & ~w53080;
assign w53084 = ~w53081 & w53083;
assign w53085 = ~w53077 & w53082;
assign w53086 = ~w53078 & w53085;
assign w53087 = w53084 & w53086;
assign w53088 = ~w53076 & ~w53087;
assign w53089 = ~w53024 & w53045;
assign w53090 = w53023 & ~w53037;
assign w53091 = (~w53044 & w53037) | (~w53044 & w53053) | (w53037 & w53053);
assign w53092 = w53030 & ~w53052;
assign w53093 = ~w53091 & ~w53092;
assign w53094 = w53089 & w53093;
assign w53095 = ~w53059 & ~w53094;
assign w53096 = ~w53088 & w53095;
assign w53097 = pi2807 & w53096;
assign w53098 = ~pi2807 & ~w53096;
assign w53099 = ~w53097 & ~w53098;
assign w53100 = w52481 & w52734;
assign w53101 = ~w52452 & w52736;
assign w53102 = w52475 & w52608;
assign w53103 = ~w52453 & w52496;
assign w53104 = ~w53102 & w53103;
assign w53105 = ~w53100 & w53104;
assign w53106 = ~w53101 & w53105;
assign w53107 = ~w52744 & ~w53106;
assign w53108 = ~pi2815 & w53107;
assign w53109 = pi2815 & ~w53107;
assign w53110 = ~w53108 & ~w53109;
assign w53111 = ~pi6302 & pi9040;
assign w53112 = ~pi6398 & ~pi9040;
assign w53113 = ~w53111 & ~w53112;
assign w53114 = pi2777 & ~w53113;
assign w53115 = ~pi2777 & w53113;
assign w53116 = ~w53114 & ~w53115;
assign w53117 = ~pi6379 & pi9040;
assign w53118 = ~pi6234 & ~pi9040;
assign w53119 = ~w53117 & ~w53118;
assign w53120 = pi2762 & ~w53119;
assign w53121 = ~pi2762 & w53119;
assign w53122 = ~w53120 & ~w53121;
assign w53123 = w53116 & w53122;
assign w53124 = ~pi6264 & pi9040;
assign w53125 = ~pi6366 & ~pi9040;
assign w53126 = ~w53124 & ~w53125;
assign w53127 = pi2748 & ~w53126;
assign w53128 = ~pi2748 & w53126;
assign w53129 = ~w53127 & ~w53128;
assign w53130 = ~w53123 & ~w53129;
assign w53131 = ~pi6231 & pi9040;
assign w53132 = ~pi6400 & ~pi9040;
assign w53133 = ~w53131 & ~w53132;
assign w53134 = pi2783 & ~w53133;
assign w53135 = ~pi2783 & w53133;
assign w53136 = ~w53134 & ~w53135;
assign w53137 = w53116 & w53136;
assign w53138 = w53130 & w53137;
assign w53139 = ~w53116 & w53136;
assign w53140 = w53116 & ~w53136;
assign w53141 = ~pi6301 & pi9040;
assign w53142 = ~pi6273 & ~pi9040;
assign w53143 = ~w53141 & ~w53142;
assign w53144 = pi2761 & ~w53143;
assign w53145 = ~pi2761 & w53143;
assign w53146 = ~w53144 & ~w53145;
assign w53147 = w53122 & ~w53146;
assign w53148 = ~w53122 & w53146;
assign w53149 = ~w53147 & ~w53148;
assign w53150 = ~w53140 & ~w53149;
assign w53151 = w53140 & w53149;
assign w53152 = ~w53150 & ~w53151;
assign w53153 = ~w53139 & w53152;
assign w53154 = ~w53122 & ~w53146;
assign w53155 = w53129 & ~w53154;
assign w53156 = w53116 & ~w53146;
assign w53157 = ~w53116 & ~w53136;
assign w53158 = w53146 & w53157;
assign w53159 = ~w53156 & ~w53158;
assign w53160 = w53155 & ~w53159;
assign w53161 = ~w53136 & ~w53146;
assign w53162 = w53155 & ~w53161;
assign w53163 = ~w53150 & ~w53162;
assign w53164 = w53122 & w53157;
assign w53165 = ~w53122 & w53139;
assign w53166 = ~w53164 & ~w53165;
assign w53167 = w53129 & ~w53166;
assign w53168 = ~w53160 & ~w53167;
assign w53169 = (~w53160 & w53168) | (~w53160 & w64093) | (w53168 & w64093);
assign w53170 = ~w53153 & ~w53169;
assign w53171 = ~w53116 & ~w53122;
assign w53172 = ~w53140 & ~w53147;
assign w53173 = ~w53139 & ~w53154;
assign w53174 = ~w53172 & ~w53173;
assign w53175 = ~w53171 & ~w53174;
assign w53176 = w53129 & w53161;
assign w53177 = ~w53139 & ~w53176;
assign w53178 = w53175 & ~w53177;
assign w53179 = w53116 & w53148;
assign w53180 = ~w53164 & ~w53179;
assign w53181 = w53130 & ~w53165;
assign w53182 = w53180 & w53181;
assign w53183 = ~pi6381 & pi9040;
assign w53184 = ~pi6181 & ~pi9040;
assign w53185 = ~w53183 & ~w53184;
assign w53186 = pi2764 & ~w53185;
assign w53187 = ~pi2764 & w53185;
assign w53188 = ~w53186 & ~w53187;
assign w53189 = (~w53188 & w53178) | (~w53188 & w64094) | (w53178 & w64094);
assign w53190 = w53122 & w53146;
assign w53191 = ~w53136 & w53190;
assign w53192 = ~w53116 & ~w53188;
assign w53193 = w53191 & ~w53192;
assign w53194 = ~w53129 & ~w53180;
assign w53195 = w53123 & ~w53163;
assign w53196 = w53129 & ~w53175;
assign w53197 = ~w53194 & ~w53195;
assign w53198 = (w53188 & ~w53197) | (w53188 & w66954) | (~w53197 & w66954);
assign w53199 = ~w53138 & ~w53193;
assign w53200 = ~w53189 & w53199;
assign w53201 = ~w53170 & w53200;
assign w53202 = (pi2784 & ~w53201) | (pi2784 & w66955) | (~w53201 & w66955);
assign w53203 = w53201 & w66956;
assign w53204 = ~w53202 & ~w53203;
assign w53205 = w53053 & w53069;
assign w53206 = w53024 & w53066;
assign w53207 = w53023 & w53044;
assign w53208 = w53037 & w53207;
assign w53209 = ~w53030 & w53044;
assign w53210 = ~w53023 & ~w53036;
assign w53211 = ~w53066 & w53210;
assign w53212 = ~w53209 & w53211;
assign w53213 = ~w53056 & ~w53212;
assign w53214 = w53036 & w53207;
assign w53215 = ~w53211 & ~w53214;
assign w53216 = w53030 & ~w53045;
assign w53217 = (~w53090 & ~w53215) | (~w53090 & w64095) | (~w53215 & w64095);
assign w53218 = ~w53017 & ~w53207;
assign w53219 = ~w53217 & w53218;
assign w53220 = (~w53208 & w53213) | (~w53208 & w64096) | (w53213 & w64096);
assign w53221 = ~w53219 & w53220;
assign w53222 = (~w53215 & w53213) | (~w53215 & w66957) | (w53213 & w66957);
assign w53223 = w53215 & w64097;
assign w53224 = ~w53047 & ~w53080;
assign w53225 = ~w53223 & w53224;
assign w53226 = ~w53222 & w53225;
assign w53227 = w53065 & ~w53226;
assign w53228 = ~w53205 & ~w53206;
assign w53229 = (w53228 & w53221) | (w53228 & w66958) | (w53221 & w66958);
assign w53230 = ~w53227 & w53229;
assign w53231 = pi2793 & w53230;
assign w53232 = ~pi2793 & ~w53230;
assign w53233 = ~w53231 & ~w53232;
assign w53234 = w52796 & w52818;
assign w53235 = (w52756 & ~w52810) | (w52756 & w66959) | (~w52810 & w66959);
assign w53236 = w52768 & w52791;
assign w53237 = w52812 & w53236;
assign w53238 = w52776 & ~w52801;
assign w53239 = ~w52790 & ~w53238;
assign w53240 = ~w52807 & ~w53239;
assign w53241 = w52815 & w64098;
assign w53242 = ~w52831 & ~w53241;
assign w53243 = (~w52756 & w53240) | (~w52756 & w64099) | (w53240 & w64099);
assign w53244 = ~w53237 & ~w53243;
assign w53245 = (w52762 & w52795) | (w52762 & w64100) | (w52795 & w64100);
assign w53246 = ~w52832 & w53245;
assign w53247 = ~w52791 & w64101;
assign w53248 = ~w52833 & ~w53247;
assign w53249 = ~w53246 & w53248;
assign w53250 = w52756 & ~w53249;
assign w53251 = ~w53244 & ~w53250;
assign w53252 = w52848 & ~w53234;
assign w53253 = ~w53251 & w53252;
assign w53254 = (pi2799 & ~w53253) | (pi2799 & w66960) | (~w53253 & w66960);
assign w53255 = w53253 & w66961;
assign w53256 = ~w53254 & ~w53255;
assign w53257 = w52789 & ~w52836;
assign w53258 = ~w52756 & w52800;
assign w53259 = ~w53257 & ~w53258;
assign w53260 = ~w52768 & ~w53259;
assign w53261 = ~w52762 & ~w53257;
assign w53262 = ~w53245 & ~w53261;
assign w53263 = w52834 & w53236;
assign w53264 = ~w53262 & ~w53263;
assign w53265 = ~w52756 & ~w53264;
assign w53266 = ~w53250 & ~w53260;
assign w53267 = ~w53265 & w53266;
assign w53268 = pi2788 & w53267;
assign w53269 = ~pi2788 & ~w53267;
assign w53270 = ~w53268 & ~w53269;
assign w53271 = ~w52518 & w52570;
assign w53272 = w52581 & ~w53271;
assign w53273 = w52545 & ~w53272;
assign w53274 = ~w52537 & w52570;
assign w53275 = ~w52524 & w52538;
assign w53276 = ~w52586 & ~w53275;
assign w53277 = (~w52544 & ~w53276) | (~w52544 & w66962) | (~w53276 & w66962);
assign w53278 = ~w52575 & ~w53274;
assign w53279 = ~w52561 & ~w52570;
assign w53280 = (w52544 & ~w53279) | (w52544 & w66963) | (~w53279 & w66963);
assign w53281 = w53278 & w53280;
assign w53282 = ~w52518 & w52560;
assign w53283 = ~w52584 & ~w53282;
assign w53284 = w52553 & ~w52559;
assign w53285 = w53283 & w53284;
assign w53286 = ~w53277 & w53285;
assign w53287 = ~w53281 & w53286;
assign w53288 = ~w52531 & w52569;
assign w53289 = ~w52546 & ~w53288;
assign w53290 = ~w52524 & ~w53289;
assign w53291 = w52569 & w52585;
assign w53292 = ~w52553 & ~w53290;
assign w53293 = ~w53291 & w53292;
assign w53294 = ~w52560 & ~w52569;
assign w53295 = ~w52579 & w53294;
assign w53296 = w52518 & ~w52531;
assign w53297 = w52553 & ~w53296;
assign w53298 = w52567 & ~w53297;
assign w53299 = w53295 & w53298;
assign w53300 = ~w53273 & ~w53299;
assign w53301 = (w53300 & w53287) | (w53300 & w66964) | (w53287 & w66964);
assign w53302 = pi2829 & w53301;
assign w53303 = ~pi2829 & ~w53301;
assign w53304 = ~w53302 & ~w53303;
assign w53305 = ~w53137 & ~w53161;
assign w53306 = ~w53156 & ~w53305;
assign w53307 = ~w53305 & w64102;
assign w53308 = (w53129 & w53307) | (w53129 & w66965) | (w53307 & w66965);
assign w53309 = w53139 & ~w53149;
assign w53310 = ~w53129 & w53140;
assign w53311 = ~w53309 & ~w53310;
assign w53312 = ~w53308 & w53311;
assign w53313 = w53188 & ~w53312;
assign w53314 = ~w53138 & ~w53162;
assign w53315 = w53146 & ~w53167;
assign w53316 = ~w53314 & ~w53315;
assign w53317 = w53146 & w53181;
assign w53318 = ~w53148 & ~w53166;
assign w53319 = w53151 & w53176;
assign w53320 = ~w53317 & ~w53318;
assign w53321 = ~w53319 & w53320;
assign w53322 = (~w53188 & ~w53321) | (~w53188 & w66966) | (~w53321 & w66966);
assign w53323 = ~w53313 & ~w53316;
assign w53324 = ~w53322 & w53323;
assign w53325 = ~pi2786 & w53324;
assign w53326 = pi2786 & ~w53324;
assign w53327 = ~w53325 & ~w53326;
assign w53328 = w53066 & w53210;
assign w53329 = (~w53051 & ~w53055) | (~w53051 & w66967) | (~w53055 & w66967);
assign w53330 = w53065 & ~w53209;
assign w53331 = ~w53329 & w53330;
assign w53332 = ~w53214 & ~w53328;
assign w53333 = ~w53331 & w53332;
assign w53334 = w53017 & ~w53333;
assign w53335 = w53037 & w53053;
assign w53336 = w53065 & ~w53214;
assign w53337 = (~w53335 & ~w53093) | (~w53335 & w66968) | (~w53093 & w66968);
assign w53338 = ~w53017 & ~w53337;
assign w53339 = w53036 & ~w53046;
assign w53340 = w53209 & w53339;
assign w53341 = ~w53052 & w64103;
assign w53342 = ~w53079 & ~w53081;
assign w53343 = ~w53017 & ~w53045;
assign w53344 = ~w53342 & ~w53343;
assign w53345 = w53048 & ~w53340;
assign w53346 = ~w53341 & w53345;
assign w53347 = ~w53344 & w53346;
assign w53348 = (~w53065 & ~w53346) | (~w53065 & w66969) | (~w53346 & w66969);
assign w53349 = ~w53059 & ~w53334;
assign w53350 = ~w53338 & ~w53348;
assign w53351 = w53349 & w53350;
assign w53352 = pi2804 & ~w53351;
assign w53353 = ~pi2804 & w53351;
assign w53354 = ~w53352 & ~w53353;
assign w53355 = w52917 & w52929;
assign w53356 = ~w52923 & ~w53355;
assign w53357 = w52936 & w52943;
assign w53358 = w52930 & w53357;
assign w53359 = ~w52917 & ~w52929;
assign w53360 = w52947 & w53359;
assign w53361 = ~w53358 & ~w53360;
assign w53362 = w53356 & ~w53361;
assign w53363 = w52976 & w52984;
assign w53364 = w52957 & w53355;
assign w53365 = ~w52945 & ~w52947;
assign w53366 = w52975 & ~w53365;
assign w53367 = w53361 & ~w53364;
assign w53368 = ~w53366 & w53367;
assign w53369 = ~w52917 & ~w52966;
assign w53370 = ~w52929 & w52936;
assign w53371 = w53369 & ~w53370;
assign w53372 = ~w52970 & ~w53363;
assign w53373 = (w53372 & ~w53368) | (w53372 & w66970) | (~w53368 & w66970);
assign w53374 = w52954 & ~w53373;
assign w53375 = ~w52978 & ~w52984;
assign w53376 = ~w52929 & w53375;
assign w53377 = (~w52954 & ~w53368) | (~w52954 & w66971) | (~w53368 & w66971);
assign w53378 = w52923 & w53370;
assign w53379 = ~w52987 & ~w53378;
assign w53380 = w52917 & ~w53379;
assign w53381 = ~w53362 & ~w53380;
assign w53382 = ~w53377 & w53381;
assign w53383 = ~w53374 & w53382;
assign w53384 = pi2792 & ~w53383;
assign w53385 = ~pi2792 & w53383;
assign w53386 = ~w53384 & ~w53385;
assign w53387 = ~w52661 & w66972;
assign w53388 = ~w52659 & w52707;
assign w53389 = w52888 & ~w53388;
assign w53390 = ~w52710 & ~w53387;
assign w53391 = ~w53389 & w53390;
assign w53392 = w52706 & ~w53391;
assign w53393 = ~w52678 & ~w53392;
assign w53394 = (w52864 & w52859) | (w52864 & w66973) | (w52859 & w66973);
assign w53395 = w52670 & ~w52709;
assign w53396 = ~w52663 & w53395;
assign w53397 = ~w52670 & w52687;
assign w53398 = w52678 & ~w52680;
assign w53399 = ~w53396 & w53398;
assign w53400 = ~w53397 & w53399;
assign w53401 = ~w52678 & ~w52710;
assign w53402 = w52692 & w52895;
assign w53403 = ~w53401 & w53402;
assign w53404 = ~w53400 & ~w53403;
assign w53405 = ~w53394 & w53404;
assign w53406 = ~w53393 & w53405;
assign w53407 = pi2801 & ~w53406;
assign w53408 = ~pi2801 & w53406;
assign w53409 = ~w53407 & ~w53408;
assign w53410 = w52525 & w52564;
assign w53411 = w52544 & w52586;
assign w53412 = ~w52531 & w52544;
assign w53413 = (~w53412 & w53290) | (~w53412 & w66974) | (w53290 & w66974);
assign w53414 = ~w52558 & ~w53274;
assign w53415 = w52544 & ~w53414;
assign w53416 = (~w52553 & w52587) | (~w52553 & w66975) | (w52587 & w66975);
assign w53417 = ~w53415 & w53416;
assign w53418 = ~w53413 & w53417;
assign w53419 = w52576 & ~w53278;
assign w53420 = w52524 & w52545;
assign w53421 = ~w52576 & w53420;
assign w53422 = ~w52590 & ~w53282;
assign w53423 = w52544 & ~w52554;
assign w53424 = ~w53422 & w53423;
assign w53425 = w52553 & ~w53419;
assign w53426 = ~w53421 & ~w53424;
assign w53427 = w53425 & w53426;
assign w53428 = ~w53418 & ~w53427;
assign w53429 = ~w53410 & ~w53411;
assign w53430 = ~w53428 & w53429;
assign w53431 = pi2814 & ~w53430;
assign w53432 = ~pi2814 & w53430;
assign w53433 = ~w53431 & ~w53432;
assign w53434 = w52917 & ~w52954;
assign w53435 = w52978 & w53370;
assign w53436 = w52944 & ~w52976;
assign w53437 = ~w52954 & ~w52964;
assign w53438 = ~w53436 & w53437;
assign w53439 = ~w53363 & w53438;
assign w53440 = ~w52929 & w53436;
assign w53441 = (~w52917 & ~w52958) | (~w52917 & w64104) | (~w52958 & w64104);
assign w53442 = ~w52930 & ~w52965;
assign w53443 = w52988 & ~w53442;
assign w53444 = w53361 & ~w53440;
assign w53445 = ~w53443 & w53444;
assign w53446 = ~w53441 & w53445;
assign w53447 = ~w52946 & ~w53435;
assign w53448 = (~w53446 & w66976) | (~w53446 & w66977) | (w66976 & w66977);
assign w53449 = ~w52923 & w53357;
assign w53450 = ~w52917 & ~w53449;
assign w53451 = w53361 & ~w53450;
assign w53452 = w53439 & w53451;
assign w53453 = ~w53448 & ~w53452;
assign w53454 = ~pi2796 & w53453;
assign w53455 = pi2796 & ~w53453;
assign w53456 = ~w53454 & ~w53455;
assign w53457 = ~w53306 & ~w53318;
assign w53458 = (w53129 & w53318) | (w53129 & w64106) | (w53318 & w64106);
assign w53459 = ~w53129 & ~w53152;
assign w53460 = ~w53458 & ~w53459;
assign w53461 = ~w53188 & ~w53460;
assign w53462 = ~w53129 & w53309;
assign w53463 = w53155 & ~w53174;
assign w53464 = w53457 & w53463;
assign w53465 = ~w53153 & ~w53464;
assign w53466 = w53188 & ~w53458;
assign w53467 = ~w53465 & w53466;
assign w53468 = (~w53462 & w53168) | (~w53462 & w66978) | (w53168 & w66978);
assign w53469 = ~w53461 & w53468;
assign w53470 = ~w53467 & w53469;
assign w53471 = pi2797 & ~w53470;
assign w53472 = ~pi2797 & w53470;
assign w53473 = ~w53471 & ~w53472;
assign w53474 = ~pi6310 & pi9040;
assign w53475 = ~pi6232 & ~pi9040;
assign w53476 = ~w53474 & ~w53475;
assign w53477 = pi2759 & ~w53476;
assign w53478 = ~pi2759 & w53476;
assign w53479 = ~w53477 & ~w53478;
assign w53480 = ~pi6303 & pi9040;
assign w53481 = ~pi6305 & ~pi9040;
assign w53482 = ~w53480 & ~w53481;
assign w53483 = pi2769 & ~w53482;
assign w53484 = ~pi2769 & w53482;
assign w53485 = ~w53483 & ~w53484;
assign w53486 = ~w53479 & ~w53485;
assign w53487 = ~pi6377 & pi9040;
assign w53488 = ~pi6537 & ~pi9040;
assign w53489 = ~w53487 & ~w53488;
assign w53490 = pi2781 & ~w53489;
assign w53491 = ~pi2781 & w53489;
assign w53492 = ~w53490 & ~w53491;
assign w53493 = ~w53479 & ~w53492;
assign w53494 = ~pi6247 & pi9040;
assign w53495 = ~pi6472 & ~pi9040;
assign w53496 = ~w53494 & ~w53495;
assign w53497 = pi2770 & ~w53496;
assign w53498 = ~pi2770 & w53496;
assign w53499 = ~w53497 & ~w53498;
assign w53500 = w53493 & w53499;
assign w53501 = ~w53479 & ~w53499;
assign w53502 = w53492 & w53501;
assign w53503 = ~w53500 & ~w53502;
assign w53504 = ~pi6269 & pi9040;
assign w53505 = ~pi6244 & ~pi9040;
assign w53506 = ~w53504 & ~w53505;
assign w53507 = pi2739 & ~w53506;
assign w53508 = ~pi2739 & w53506;
assign w53509 = ~w53507 & ~w53508;
assign w53510 = ~w53485 & ~w53499;
assign w53511 = w53479 & w53492;
assign w53512 = ~w53493 & ~w53511;
assign w53513 = ~w53479 & w53509;
assign w53514 = w53512 & ~w53513;
assign w53515 = w53512 & w64107;
assign w53516 = w53509 & ~w53515;
assign w53517 = w53503 & w53516;
assign w53518 = w53486 & w53517;
assign w53519 = ~pi6274 & pi9040;
assign w53520 = ~pi6299 & ~pi9040;
assign w53521 = ~w53519 & ~w53520;
assign w53522 = pi2757 & ~w53521;
assign w53523 = ~pi2757 & w53521;
assign w53524 = ~w53522 & ~w53523;
assign w53525 = w53485 & w53499;
assign w53526 = w53493 & ~w53525;
assign w53527 = ~w53479 & w53492;
assign w53528 = w53525 & w53527;
assign w53529 = ~w53485 & w53492;
assign w53530 = w53485 & ~w53492;
assign w53531 = ~w53529 & ~w53530;
assign w53532 = ~w53528 & w53531;
assign w53533 = w53509 & ~w53532;
assign w53534 = (~w53493 & ~w53532) | (~w53493 & w66979) | (~w53532 & w66979);
assign w53535 = ~w53533 & w53534;
assign w53536 = w53524 & ~w53526;
assign w53537 = ~w53535 & w53536;
assign w53538 = ~w53510 & ~w53527;
assign w53539 = w53509 & w53538;
assign w53540 = w53529 & w53539;
assign w53541 = ~w53510 & ~w53525;
assign w53542 = w53514 & ~w53541;
assign w53543 = ~w53485 & ~w53511;
assign w53544 = w53509 & ~w53543;
assign w53545 = w53502 & w53544;
assign w53546 = ~w53512 & w53541;
assign w53547 = ~w53542 & ~w53546;
assign w53548 = (~w53524 & ~w53547) | (~w53524 & w66980) | (~w53547 & w66980);
assign w53549 = ~w53518 & ~w53540;
assign w53550 = ~w53537 & ~w53548;
assign w53551 = w53549 & w53550;
assign w53552 = pi2809 & ~w53551;
assign w53553 = ~pi2809 & w53551;
assign w53554 = ~w53552 & ~w53553;
assign w53555 = ~w53068 & ~w53089;
assign w53556 = w53058 & w53555;
assign w53557 = w53090 & w53556;
assign w53558 = ~w53017 & ~w53342;
assign w53559 = ~w53328 & ~w53558;
assign w53560 = (w53065 & w53557) | (w53065 & w66981) | (w53557 & w66981);
assign w53561 = ~w53057 & w53343;
assign w53562 = (~w53072 & ~w53215) | (~w53072 & w66982) | (~w53215 & w66982);
assign w53563 = ~w53017 & ~w53058;
assign w53564 = ~w53065 & ~w53556;
assign w53565 = ~w53563 & w53564;
assign w53566 = (~w53561 & ~w53347) | (~w53561 & w64108) | (~w53347 & w64108);
assign w53567 = ~w53565 & w53566;
assign w53568 = w53567 & w66983;
assign w53569 = (pi2800 & ~w53567) | (pi2800 & w66984) | (~w53567 & w66984);
assign w53570 = ~w53568 & ~w53569;
assign w53571 = ~w52589 & ~w53280;
assign w53572 = ~w52553 & ~w53571;
assign w53573 = ~w53276 & w53295;
assign w53574 = ~w52578 & ~w53412;
assign w53575 = w52554 & ~w53574;
assign w53576 = w52557 & ~w53297;
assign w53577 = ~w53575 & ~w53576;
assign w53578 = ~w53573 & w53577;
assign w53579 = ~w52544 & ~w53578;
assign w53580 = ~w52524 & w52544;
assign w53581 = ~w53283 & w53580;
assign w53582 = ~w53280 & w53288;
assign w53583 = ~w53271 & ~w53575;
assign w53584 = ~w53582 & w53583;
assign w53585 = w52553 & ~w53584;
assign w53586 = ~w53579 & ~w53581;
assign w53587 = ~w53572 & w53586;
assign w53588 = w53587 & w66985;
assign w53589 = (pi2843 & ~w53587) | (pi2843 & w66986) | (~w53587 & w66986);
assign w53590 = ~w53588 & ~w53589;
assign w53591 = w52943 & w52945;
assign w53592 = w52917 & ~w53591;
assign w53593 = ~w53440 & w53592;
assign w53594 = ~w53450 & ~w53593;
assign w53595 = ~w52965 & ~w53356;
assign w53596 = w52929 & ~w52936;
assign w53597 = ~w53370 & ~w53596;
assign w53598 = ~w53595 & w53597;
assign w53599 = ~w52979 & w52986;
assign w53600 = ~w53598 & w53599;
assign w53601 = w52917 & ~w53375;
assign w53602 = ~w52929 & w52978;
assign w53603 = w53369 & ~w53602;
assign w53604 = ~w53601 & ~w53603;
assign w53605 = w52954 & ~w52987;
assign w53606 = ~w53604 & w53605;
assign w53607 = ~w53600 & ~w53606;
assign w53608 = ~w53594 & ~w53607;
assign w53609 = ~pi2810 & w53608;
assign w53610 = pi2810 & ~w53608;
assign w53611 = ~w53609 & ~w53610;
assign w53612 = w53516 & ~w53524;
assign w53613 = w53479 & w53499;
assign w53614 = ~w53485 & w53613;
assign w53615 = w53485 & w53493;
assign w53616 = w53503 & w63442;
assign w53617 = (~w53509 & ~w53531) | (~w53509 & w64109) | (~w53531 & w64109);
assign w53618 = w53616 & ~w53617;
assign w53619 = w53616 & w64110;
assign w53620 = ~w53502 & w53509;
assign w53621 = ~w53538 & w53620;
assign w53622 = ~w53619 & ~w53621;
assign w53623 = ~w53612 & ~w53622;
assign w53624 = ~w53616 & w53617;
assign w53625 = ~w53618 & ~w53624;
assign w53626 = ~w53509 & ~w53510;
assign w53627 = ~w53512 & w53626;
assign w53628 = w53524 & ~w53627;
assign w53629 = ~w53515 & w53628;
assign w53630 = (~w53629 & w53625) | (~w53629 & w66987) | (w53625 & w66987);
assign w53631 = ~w53545 & ~w53623;
assign w53632 = (pi2805 & ~w53631) | (pi2805 & w66988) | (~w53631 & w66988);
assign w53633 = w53631 & w66989;
assign w53634 = ~w53632 & ~w53633;
assign w53635 = ~w53486 & ~w53542;
assign w53636 = w53539 & ~w53635;
assign w53637 = ~w53512 & ~w53529;
assign w53638 = (~w53486 & w53512) | (~w53486 & w66990) | (w53512 & w66990);
assign w53639 = ~w53500 & ~w53524;
assign w53640 = ~w53638 & w53639;
assign w53641 = ~w53614 & ~w53640;
assign w53642 = ~w53509 & ~w53641;
assign w53643 = ~w53492 & ~w53509;
assign w53644 = (~w53643 & ~w53531) | (~w53643 & w66991) | (~w53531 & w66991);
assign w53645 = ~w53501 & ~w53613;
assign w53646 = ~w53644 & w53645;
assign w53647 = ~w53530 & ~w53613;
assign w53648 = ~w53511 & w53525;
assign w53649 = w53509 & ~w53647;
assign w53650 = ~w53648 & w53649;
assign w53651 = (~w53529 & ~w53649) | (~w53529 & w66992) | (~w53649 & w66992);
assign w53652 = w53501 & ~w53651;
assign w53653 = w53524 & ~w53528;
assign w53654 = ~w53646 & w53653;
assign w53655 = ~w53652 & w53654;
assign w53656 = w53493 & w53510;
assign w53657 = w53544 & ~w53637;
assign w53658 = ~w53524 & ~w53656;
assign w53659 = ~w53657 & w53658;
assign w53660 = ~w53655 & ~w53659;
assign w53661 = ~w53636 & ~w53642;
assign w53662 = ~w53660 & w53661;
assign w53663 = pi2816 & ~w53662;
assign w53664 = ~pi2816 & w53662;
assign w53665 = ~w53663 & ~w53664;
assign w53666 = ~w53486 & ~w53529;
assign w53667 = w53503 & w66993;
assign w53668 = ~w53486 & ~w53509;
assign w53669 = w53647 & w53668;
assign w53670 = ~w53650 & ~w53669;
assign w53671 = (~w53524 & ~w53670) | (~w53524 & w66994) | (~w53670 & w66994);
assign w53672 = w53525 & w53643;
assign w53673 = ~w53524 & ~w53672;
assign w53674 = ~w53509 & ~w53613;
assign w53675 = ~w53615 & w53674;
assign w53676 = (~w53675 & ~w53516) | (~w53675 & w66995) | (~w53516 & w66995);
assign w53677 = ~w53648 & ~w53676;
assign w53678 = ~w53673 & ~w53677;
assign w53679 = ~w53540 & ~w53671;
assign w53680 = ~w53678 & w53679;
assign w53681 = ~pi2811 & w53680;
assign w53682 = pi2811 & ~w53680;
assign w53683 = ~w53681 & ~w53682;
assign w53684 = w53130 & w53190;
assign w53685 = w53137 & w53154;
assign w53686 = (~w53129 & ~w53190) | (~w53129 & w66996) | (~w53190 & w66996);
assign w53687 = ~w53156 & ~w53172;
assign w53688 = (~w53685 & ~w53687) | (~w53685 & w66997) | (~w53687 & w66997);
assign w53689 = ~w53684 & w53688;
assign w53690 = w53188 & ~w53689;
assign w53691 = ~w53129 & w53307;
assign w53692 = (~w53130 & w53309) | (~w53130 & w66998) | (w53309 & w66998);
assign w53693 = w53688 & w53692;
assign w53694 = w53159 & w53686;
assign w53695 = ~w53122 & w53136;
assign w53696 = ~w53156 & w53695;
assign w53697 = ~w53160 & ~w53696;
assign w53698 = ~w53694 & w53697;
assign w53699 = ~w53188 & ~w53698;
assign w53700 = ~w53319 & ~w53691;
assign w53701 = ~w53693 & w53700;
assign w53702 = ~w53690 & w53701;
assign w53703 = ~w53699 & w53702;
assign w53704 = pi2808 & ~w53703;
assign w53705 = ~pi2808 & w53703;
assign w53706 = ~w53704 & ~w53705;
assign w53707 = ~pi6637 & pi9040;
assign w53708 = ~pi6491 & ~pi9040;
assign w53709 = ~w53707 & ~w53708;
assign w53710 = pi2844 & ~w53709;
assign w53711 = ~pi2844 & w53709;
assign w53712 = ~w53710 & ~w53711;
assign w53713 = ~pi6599 & pi9040;
assign w53714 = ~pi6485 & ~pi9040;
assign w53715 = ~w53713 & ~w53714;
assign w53716 = pi2802 & ~w53715;
assign w53717 = ~pi2802 & w53715;
assign w53718 = ~w53716 & ~w53717;
assign w53719 = ~w53712 & ~w53718;
assign w53720 = ~pi6416 & pi9040;
assign w53721 = ~pi6610 & ~pi9040;
assign w53722 = ~w53720 & ~w53721;
assign w53723 = pi2820 & ~w53722;
assign w53724 = ~pi2820 & w53722;
assign w53725 = ~w53723 & ~w53724;
assign w53726 = ~pi6404 & pi9040;
assign w53727 = ~pi6494 & ~pi9040;
assign w53728 = ~w53726 & ~w53727;
assign w53729 = pi2818 & ~w53728;
assign w53730 = ~pi2818 & w53728;
assign w53731 = ~w53729 & ~w53730;
assign w53732 = ~w53725 & w53731;
assign w53733 = w53719 & w53732;
assign w53734 = w53712 & ~w53725;
assign w53735 = ~w53718 & ~w53731;
assign w53736 = ~w53734 & w53735;
assign w53737 = w53718 & w53725;
assign w53738 = w53731 & w53737;
assign w53739 = ~w53736 & ~w53738;
assign w53740 = ~pi6598 & pi9040;
assign w53741 = ~pi6637 & ~pi9040;
assign w53742 = ~w53740 & ~w53741;
assign w53743 = pi2835 & ~w53742;
assign w53744 = ~pi2835 & w53742;
assign w53745 = ~w53743 & ~w53744;
assign w53746 = ~w53739 & ~w53745;
assign w53747 = ~w53712 & ~w53731;
assign w53748 = ~w53718 & ~w53725;
assign w53749 = ~w53737 & w53747;
assign w53750 = ~w53748 & w53749;
assign w53751 = w53712 & w53725;
assign w53752 = w53712 & w53718;
assign w53753 = ~w53719 & ~w53752;
assign w53754 = w53731 & w53753;
assign w53755 = w53753 & w64111;
assign w53756 = w53712 & ~w53731;
assign w53757 = ~w53736 & w53756;
assign w53758 = ~w53755 & ~w53757;
assign w53759 = w53745 & ~w53758;
assign w53760 = w53737 & w66999;
assign w53761 = w53731 & ~w53745;
assign w53762 = w53748 & w53761;
assign w53763 = ~w53760 & ~w53762;
assign w53764 = ~w53750 & w53763;
assign w53765 = ~w53759 & w53764;
assign w53766 = ~w53759 & w67000;
assign w53767 = ~pi6459 & pi9040;
assign w53768 = ~pi6614 & ~pi9040;
assign w53769 = ~w53767 & ~w53768;
assign w53770 = pi2839 & ~w53769;
assign w53771 = ~pi2839 & w53769;
assign w53772 = ~w53770 & ~w53771;
assign w53773 = ~w53766 & w53772;
assign w53774 = w53737 & w53747;
assign w53775 = ~w53745 & w53755;
assign w53776 = w53718 & w53731;
assign w53777 = ~w53756 & ~w53776;
assign w53778 = ~w53725 & ~w53745;
assign w53779 = ~w53777 & w53778;
assign w53780 = ~w53774 & ~w53779;
assign w53781 = ~w53775 & w53780;
assign w53782 = ~w53772 & ~w53781;
assign w53783 = w53731 & ~w53753;
assign w53784 = w53736 & ~w53750;
assign w53785 = w53745 & ~w53772;
assign w53786 = (w53785 & w53784) | (w53785 & w67001) | (w53784 & w67001);
assign w53787 = w53718 & w53745;
assign w53788 = w53734 & w53787;
assign w53789 = ~w53733 & ~w53788;
assign w53790 = ~w53786 & w53789;
assign w53791 = ~w53782 & w53790;
assign w53792 = ~w53773 & w53791;
assign w53793 = ~pi2861 & w53792;
assign w53794 = pi2861 & ~w53792;
assign w53795 = ~w53793 & ~w53794;
assign w53796 = ~w53739 & w53778;
assign w53797 = ~w53731 & ~w53745;
assign w53798 = ~w53753 & w53797;
assign w53799 = ~w53753 & w67002;
assign w53800 = w53725 & ~w53745;
assign w53801 = w53777 & w53800;
assign w53802 = ~w53732 & ~w53751;
assign w53803 = w53745 & ~w53802;
assign w53804 = ~w53754 & w53803;
assign w53805 = w53776 & w53778;
assign w53806 = ~w53712 & w53805;
assign w53807 = ~w53801 & ~w53806;
assign w53808 = ~w53799 & w53807;
assign w53809 = (w53772 & ~w53808) | (w53772 & w67003) | (~w53808 & w67003);
assign w53810 = w53725 & ~w53731;
assign w53811 = (w53745 & ~w53802) | (w53745 & w67004) | (~w53802 & w67004);
assign w53812 = w53731 & ~w53734;
assign w53813 = ~w53802 & ~w53812;
assign w53814 = ~w53745 & ~w53813;
assign w53815 = ~w53811 & ~w53814;
assign w53816 = ~w53734 & ~w53787;
assign w53817 = w53777 & ~w53816;
assign w53818 = w53763 & ~w53817;
assign w53819 = ~w53815 & w53818;
assign w53820 = ~w53772 & ~w53819;
assign w53821 = ~w53814 & w67005;
assign w53822 = w53748 & w53756;
assign w53823 = ~w53738 & ~w53822;
assign w53824 = w53745 & ~w53823;
assign w53825 = ~w53796 & ~w53824;
assign w53826 = ~w53821 & w53825;
assign w53827 = ~w53809 & w53826;
assign w53828 = ~w53820 & w53827;
assign w53829 = pi2857 & ~w53828;
assign w53830 = ~pi2857 & w53828;
assign w53831 = ~w53829 & ~w53830;
assign w53832 = ~pi6627 & pi9040;
assign w53833 = ~pi6619 & ~pi9040;
assign w53834 = ~w53832 & ~w53833;
assign w53835 = pi2821 & ~w53834;
assign w53836 = ~pi2821 & w53834;
assign w53837 = ~w53835 & ~w53836;
assign w53838 = ~pi6577 & pi9040;
assign w53839 = ~pi6598 & ~pi9040;
assign w53840 = ~w53838 & ~w53839;
assign w53841 = pi2842 & ~w53840;
assign w53842 = ~pi2842 & w53840;
assign w53843 = ~w53841 & ~w53842;
assign w53844 = ~pi6610 & pi9040;
assign w53845 = ~pi6604 & ~pi9040;
assign w53846 = ~w53844 & ~w53845;
assign w53847 = pi2813 & ~w53846;
assign w53848 = ~pi2813 & w53846;
assign w53849 = ~w53847 & ~w53848;
assign w53850 = ~w53843 & w53849;
assign w53851 = ~pi6555 & pi9040;
assign w53852 = ~pi6468 & ~pi9040;
assign w53853 = ~w53851 & ~w53852;
assign w53854 = pi2830 & ~w53853;
assign w53855 = ~pi2830 & w53853;
assign w53856 = ~w53854 & ~w53855;
assign w53857 = ~w53849 & ~w53856;
assign w53858 = ~w53850 & ~w53857;
assign w53859 = ~pi6481 & pi9040;
assign w53860 = ~pi6500 & ~pi9040;
assign w53861 = ~w53859 & ~w53860;
assign w53862 = pi2827 & ~w53861;
assign w53863 = ~pi2827 & w53861;
assign w53864 = ~w53862 & ~w53863;
assign w53865 = w53856 & ~w53864;
assign w53866 = w53843 & w53864;
assign w53867 = ~w53865 & ~w53866;
assign w53868 = ~w53858 & ~w53867;
assign w53869 = ~w53843 & ~w53849;
assign w53870 = ~w53864 & w53869;
assign w53871 = w53869 & w67006;
assign w53872 = w53843 & ~w53856;
assign w53873 = w53849 & ~w53864;
assign w53874 = w53872 & w53873;
assign w53875 = ~w53849 & w53865;
assign w53876 = ~w53874 & ~w53875;
assign w53877 = ~pi6419 & pi9040;
assign w53878 = ~pi6542 & ~pi9040;
assign w53879 = ~w53877 & ~w53878;
assign w53880 = pi2846 & ~w53879;
assign w53881 = ~pi2846 & w53879;
assign w53882 = ~w53880 & ~w53881;
assign w53883 = ~w53876 & ~w53882;
assign w53884 = w53843 & w53875;
assign w53885 = ~w53868 & ~w53871;
assign w53886 = ~w53884 & w53885;
assign w53887 = (w53837 & ~w53886) | (w53837 & w67007) | (~w53886 & w67007);
assign w53888 = w53843 & w53856;
assign w53889 = w53873 & w53888;
assign w53890 = ~w53849 & w53866;
assign w53891 = ~w53874 & ~w53890;
assign w53892 = ~w53857 & ~w53891;
assign w53893 = (~w53837 & ~w53869) | (~w53837 & w53902) | (~w53869 & w53902);
assign w53894 = ~w53889 & w53893;
assign w53895 = ~w53892 & w53894;
assign w53896 = (w53837 & ~w53866) | (w53837 & w67008) | (~w53866 & w67008);
assign w53897 = ~w53856 & w53864;
assign w53898 = ~w53850 & w53897;
assign w53899 = w53850 & ~w53897;
assign w53900 = ~w53898 & ~w53899;
assign w53901 = (w53882 & ~w53900) | (w53882 & w67009) | (~w53900 & w67009);
assign w53902 = ~w53837 & w53864;
assign w53903 = w53850 & ~w53856;
assign w53904 = w53902 & w53903;
assign w53905 = ~w53837 & ~w53849;
assign w53906 = w53872 & w53905;
assign w53907 = w53837 & ~w53864;
assign w53908 = w53850 & ~w53907;
assign w53909 = w53849 & w53864;
assign w53910 = w53856 & w53909;
assign w53911 = ~w53908 & ~w53910;
assign w53912 = ~w53843 & w53897;
assign w53913 = ~w53865 & ~w53888;
assign w53914 = ~w53912 & w53913;
assign w53915 = w53896 & w53914;
assign w53916 = ~w53911 & ~w53915;
assign w53917 = w53856 & w53902;
assign w53918 = ~w53906 & ~w53917;
assign w53919 = ~w53916 & w53918;
assign w53920 = ~w53882 & ~w53919;
assign w53921 = (~w53904 & w53895) | (~w53904 & w67010) | (w53895 & w67010);
assign w53922 = ~w53887 & w53921;
assign w53923 = ~w53920 & w53922;
assign w53924 = pi2852 & w53923;
assign w53925 = ~pi2852 & ~w53923;
assign w53926 = ~w53924 & ~w53925;
assign w53927 = ~w53753 & w53810;
assign w53928 = w53718 & ~w53731;
assign w53929 = ~w53800 & w53928;
assign w53930 = ~w53761 & ~w53929;
assign w53931 = ~w53712 & ~w53930;
assign w53932 = w53718 & ~w53803;
assign w53933 = w53734 & ~w53932;
assign w53934 = w53772 & ~w53927;
assign w53935 = ~w53931 & w53934;
assign w53936 = ~w53933 & w53935;
assign w53937 = w53712 & w53735;
assign w53938 = ~w53812 & ~w53937;
assign w53939 = w53745 & ~w53938;
assign w53940 = w53751 & w53776;
assign w53941 = ~w53772 & ~w53940;
assign w53942 = ~w53798 & w53941;
assign w53943 = ~w53939 & w53942;
assign w53944 = ~w53936 & ~w53943;
assign w53945 = ~w53806 & ~w53821;
assign w53946 = ~w53944 & w53945;
assign w53947 = ~pi2870 & ~w53946;
assign w53948 = pi2870 & w53946;
assign w53949 = ~w53947 & ~w53948;
assign w53950 = ~w53733 & ~w53805;
assign w53951 = w53778 & w53950;
assign w53952 = (w53718 & ~w53802) | (w53718 & w67011) | (~w53802 & w67011);
assign w53953 = w53781 & w53952;
assign w53954 = ~w53822 & ~w53951;
assign w53955 = (w53772 & w53953) | (w53772 & w67012) | (w53953 & w67012);
assign w53956 = ~w53774 & ~w53937;
assign w53957 = ~w53745 & ~w53956;
assign w53958 = (~w53772 & w53957) | (~w53772 & w67013) | (w53957 & w67013);
assign w53959 = ~w53765 & w53811;
assign w53960 = ~w53753 & w67014;
assign w53961 = w53735 & w53778;
assign w53962 = ~w53719 & ~w53735;
assign w53963 = w53785 & w53962;
assign w53964 = ~w53952 & w53963;
assign w53965 = ~w53960 & ~w53961;
assign w53966 = ~w53964 & w53965;
assign w53967 = ~w53958 & w53966;
assign w53968 = ~w53959 & w53967;
assign w53969 = (pi2869 & ~w53968) | (pi2869 & w67015) | (~w53968 & w67015);
assign w53970 = w53968 & w67016;
assign w53971 = ~w53969 & ~w53970;
assign w53972 = ~pi6604 & pi9040;
assign w53973 = ~pi6627 & ~pi9040;
assign w53974 = ~w53972 & ~w53973;
assign w53975 = pi2845 & ~w53974;
assign w53976 = ~pi2845 & w53974;
assign w53977 = ~w53975 & ~w53976;
assign w53978 = ~pi6468 & pi9040;
assign w53979 = ~pi6577 & ~pi9040;
assign w53980 = ~w53978 & ~w53979;
assign w53981 = pi2844 & ~w53980;
assign w53982 = ~pi2844 & w53980;
assign w53983 = ~w53981 & ~w53982;
assign w53984 = w53977 & w53983;
assign w53985 = ~pi6542 & pi9040;
assign w53986 = ~pi6465 & ~pi9040;
assign w53987 = ~w53985 & ~w53986;
assign w53988 = pi2826 & ~w53987;
assign w53989 = ~pi2826 & w53987;
assign w53990 = ~w53988 & ~w53989;
assign w53991 = ~pi6619 & pi9040;
assign w53992 = ~pi6484 & ~pi9040;
assign w53993 = ~w53991 & ~w53992;
assign w53994 = pi2841 & ~w53993;
assign w53995 = ~pi2841 & w53993;
assign w53996 = ~w53994 & ~w53995;
assign w53997 = w53990 & ~w53996;
assign w53998 = w53984 & w53997;
assign w53999 = ~pi6465 & pi9040;
assign w54000 = ~pi6481 & ~pi9040;
assign w54001 = ~w53999 & ~w54000;
assign w54002 = pi2818 & ~w54001;
assign w54003 = ~pi2818 & w54001;
assign w54004 = ~w54002 & ~w54003;
assign w54005 = w53984 & ~w53990;
assign w54006 = ~w53977 & w53997;
assign w54007 = ~w54005 & ~w54006;
assign w54008 = ~w53977 & ~w53983;
assign w54009 = ~w53984 & ~w54008;
assign w54010 = w54007 & ~w54009;
assign w54011 = ~w53977 & ~w53990;
assign w54012 = w53977 & ~w53983;
assign w54013 = ~w53990 & ~w53996;
assign w54014 = w54012 & w54013;
assign w54015 = ~pi6500 & pi9040;
assign w54016 = ~pi6555 & ~pi9040;
assign w54017 = ~w54015 & ~w54016;
assign w54018 = pi2828 & ~w54017;
assign w54019 = ~pi2828 & w54017;
assign w54020 = ~w54018 & ~w54019;
assign w54021 = (w54020 & w54010) | (w54020 & w64112) | (w54010 & w64112);
assign w54022 = ~w53977 & ~w53996;
assign w54023 = w53983 & w54022;
assign w54024 = (w54020 & ~w54022) | (w54020 & w54035) | (~w54022 & w54035);
assign w54025 = ~w54007 & ~w54024;
assign w54026 = w53990 & w54012;
assign w54027 = w54012 & w67017;
assign w54028 = ~w53998 & ~w54027;
assign w54029 = ~w54025 & w54028;
assign w54030 = ~w54021 & w54029;
assign w54031 = w54004 & ~w54030;
assign w54032 = ~w54012 & ~w54022;
assign w54033 = ~w53990 & ~w54020;
assign w54034 = ~w54032 & w54033;
assign w54035 = ~w53983 & w54020;
assign w54036 = w53997 & w54035;
assign w54037 = ~w53977 & w53990;
assign w54038 = w53984 & ~w53996;
assign w54039 = w53990 & w54008;
assign w54040 = ~w54038 & ~w54039;
assign w54041 = w54020 & ~w54040;
assign w54042 = w53996 & w54037;
assign w54043 = (w54042 & w54040) | (w54042 & w67018) | (w54040 & w67018);
assign w54044 = ~w54034 & ~w54036;
assign w54045 = ~w54043 & w54044;
assign w54046 = ~w54004 & ~w54045;
assign w54047 = ~w54009 & w54040;
assign w54048 = ~w54006 & w54020;
assign w54049 = ~w54047 & w67019;
assign w54050 = ~w53990 & w53996;
assign w54051 = w54008 & w54050;
assign w54052 = ~w54027 & ~w54051;
assign w54053 = w54020 & ~w54052;
assign w54054 = w53977 & ~w54020;
assign w54055 = w54050 & w54054;
assign w54056 = ~w53998 & ~w54055;
assign w54057 = ~w54053 & w54056;
assign w54058 = ~w54049 & w54057;
assign w54059 = ~w54046 & w54058;
assign w54060 = ~w54031 & w54059;
assign w54061 = pi2851 & ~w54060;
assign w54062 = ~pi2851 & w54060;
assign w54063 = ~w54061 & ~w54062;
assign w54064 = ~pi6613 & pi9040;
assign w54065 = ~pi6419 & ~pi9040;
assign w54066 = ~w54064 & ~w54065;
assign w54067 = pi2813 & ~w54066;
assign w54068 = ~pi2813 & w54066;
assign w54069 = ~w54067 & ~w54068;
assign w54070 = ~pi6480 & pi9040;
assign w54071 = ~pi6541 & ~pi9040;
assign w54072 = ~w54070 & ~w54071;
assign w54073 = pi2839 & ~w54072;
assign w54074 = ~pi2839 & w54072;
assign w54075 = ~w54073 & ~w54074;
assign w54076 = ~pi6494 & pi9040;
assign w54077 = ~pi6599 & ~pi9040;
assign w54078 = ~w54076 & ~w54077;
assign w54079 = pi2827 & ~w54078;
assign w54080 = ~pi2827 & w54078;
assign w54081 = ~w54079 & ~w54080;
assign w54082 = w54075 & ~w54081;
assign w54083 = ~w54075 & ~w54081;
assign w54084 = ~pi6408 & pi9040;
assign w54085 = ~pi6480 & ~pi9040;
assign w54086 = ~w54084 & ~w54085;
assign w54087 = pi2802 & ~w54086;
assign w54088 = ~pi2802 & w54086;
assign w54089 = ~w54087 & ~w54088;
assign w54090 = w54083 & w54089;
assign w54091 = ~w54081 & ~w54089;
assign w54092 = w54075 & w54091;
assign w54093 = ~w54090 & ~w54092;
assign w54094 = ~pi6541 & pi9040;
assign w54095 = ~pi6613 & ~pi9040;
assign w54096 = ~w54094 & ~w54095;
assign w54097 = pi2817 & ~w54096;
assign w54098 = ~pi2817 & w54096;
assign w54099 = ~w54097 & ~w54098;
assign w54100 = ~w54093 & w54099;
assign w54101 = ~pi6614 & pi9040;
assign w54102 = ~pi6416 & ~pi9040;
assign w54103 = ~w54101 & ~w54102;
assign w54104 = pi2840 & ~w54103;
assign w54105 = ~pi2840 & w54103;
assign w54106 = ~w54104 & ~w54105;
assign w54107 = ~w54089 & w54106;
assign w54108 = ~w54075 & w54081;
assign w54109 = ~w54089 & w54099;
assign w54110 = w54108 & w54109;
assign w54111 = w54075 & w54106;
assign w54112 = (~w54107 & w54110) | (~w54107 & w67020) | (w54110 & w67020);
assign w54113 = ~w54100 & ~w54112;
assign w54114 = w54089 & w54099;
assign w54115 = w54082 & w54114;
assign w54116 = ~w54106 & ~w54115;
assign w54117 = w54081 & w54089;
assign w54118 = ~w54099 & w54117;
assign w54119 = w54075 & ~w54099;
assign w54120 = ~w54082 & ~w54091;
assign w54121 = ~w54119 & ~w54120;
assign w54122 = ~w54118 & ~w54121;
assign w54123 = ~w54116 & ~w54122;
assign w54124 = w54075 & w54081;
assign w54125 = w54109 & w54124;
assign w54126 = ~w54089 & ~w54099;
assign w54127 = ~w54082 & ~w54108;
assign w54128 = w54126 & ~w54127;
assign w54129 = ~w54090 & ~w54125;
assign w54130 = ~w54128 & w54129;
assign w54131 = ~w54106 & ~w54130;
assign w54132 = ~w54123 & ~w54131;
assign w54133 = w54124 & w54126;
assign w54134 = w54089 & w54108;
assign w54135 = ~w54133 & ~w54134;
assign w54136 = ~w54106 & ~w54135;
assign w54137 = w54083 & w54126;
assign w54138 = ~w54110 & ~w54137;
assign w54139 = ~w54136 & w54138;
assign w54140 = ~w54075 & w54099;
assign w54141 = ~w54119 & ~w54140;
assign w54142 = ~w54089 & ~w54141;
assign w54143 = ~w54136 & w64113;
assign w54144 = w54132 & w54143;
assign w54145 = (~w54069 & w54144) | (~w54069 & w64114) | (w54144 & w64114);
assign w54146 = w54089 & ~w54106;
assign w54147 = ~w54069 & w54081;
assign w54148 = ~w54146 & ~w54147;
assign w54149 = ~w54107 & w54141;
assign w54150 = ~w54148 & w54149;
assign w54151 = ~w54109 & ~w54118;
assign w54152 = w54111 & ~w54151;
assign w54153 = (w54069 & ~w54139) | (w54069 & w67021) | (~w54139 & w67021);
assign w54154 = w54093 & w54138;
assign w54155 = ~w54091 & ~w54099;
assign w54156 = w54127 & w54155;
assign w54157 = w54106 & ~w54156;
assign w54158 = ~w54154 & w54157;
assign w54159 = ~w54150 & ~w54158;
assign w54160 = ~w54153 & w54159;
assign w54161 = ~w54145 & w67022;
assign w54162 = (~pi2848 & w54145) | (~pi2848 & w67023) | (w54145 & w67023);
assign w54163 = ~w54161 & ~w54162;
assign w54164 = ~w54122 & w67024;
assign w54165 = ~w54099 & ~w54135;
assign w54166 = w54113 & ~w54165;
assign w54167 = (w54069 & ~w54166) | (w54069 & w67025) | (~w54166 & w67025);
assign w54168 = ~w54091 & ~w54117;
assign w54169 = ~w54106 & ~w54168;
assign w54170 = w54083 & w54109;
assign w54171 = w54099 & w54106;
assign w54172 = w54075 & ~w54171;
assign w54173 = ~w54155 & w54172;
assign w54174 = ~w54169 & ~w54170;
assign w54175 = ~w54173 & w54174;
assign w54176 = ~w54107 & ~w54114;
assign w54177 = w54108 & ~w54176;
assign w54178 = w54083 & w67026;
assign w54179 = ~w54125 & ~w54177;
assign w54180 = ~w54178 & w54179;
assign w54181 = w54175 & w54180;
assign w54182 = ~w54069 & ~w54181;
assign w54183 = ~w54167 & ~w54182;
assign w54184 = pi2849 & ~w54183;
assign w54185 = ~pi2849 & w54183;
assign w54186 = ~w54184 & ~w54185;
assign w54187 = ~pi6501 & pi9040;
assign w54188 = ~pi6551 & ~pi9040;
assign w54189 = ~w54187 & ~w54188;
assign w54190 = pi2826 & ~w54189;
assign w54191 = ~pi2826 & w54189;
assign w54192 = ~w54190 & ~w54191;
assign w54193 = ~pi6409 & pi9040;
assign w54194 = ~pi6680 & ~pi9040;
assign w54195 = ~w54193 & ~w54194;
assign w54196 = pi2847 & ~w54195;
assign w54197 = ~pi2847 & w54195;
assign w54198 = ~w54196 & ~w54197;
assign w54199 = w54192 & w54198;
assign w54200 = ~pi6464 & pi9040;
assign w54201 = ~pi6463 & ~pi9040;
assign w54202 = ~w54200 & ~w54201;
assign w54203 = pi2825 & ~w54202;
assign w54204 = ~pi2825 & w54202;
assign w54205 = ~w54203 & ~w54204;
assign w54206 = ~pi6707 & pi9040;
assign w54207 = ~pi6501 & ~pi9040;
assign w54208 = ~w54206 & ~w54207;
assign w54209 = pi2824 & ~w54208;
assign w54210 = ~pi2824 & w54208;
assign w54211 = ~w54209 & ~w54210;
assign w54212 = ~w54205 & w54211;
assign w54213 = ~pi6504 & pi9040;
assign w54214 = ~pi6681 & ~pi9040;
assign w54215 = ~w54213 & ~w54214;
assign w54216 = pi2831 & ~w54215;
assign w54217 = ~pi2831 & w54215;
assign w54218 = ~w54216 & ~w54217;
assign w54219 = w54212 & ~w54218;
assign w54220 = ~w54211 & w54218;
assign w54221 = ~w54205 & w54220;
assign w54222 = ~w54219 & ~w54221;
assign w54223 = w54199 & ~w54222;
assign w54224 = ~pi6624 & pi9040;
assign w54225 = ~pi6506 & ~pi9040;
assign w54226 = ~w54224 & ~w54225;
assign w54227 = pi2845 & ~w54226;
assign w54228 = ~pi2845 & w54226;
assign w54229 = ~w54227 & ~w54228;
assign w54230 = w54205 & w54218;
assign w54231 = ~w54192 & ~w54211;
assign w54232 = ~w54199 & ~w54231;
assign w54233 = w54230 & w54232;
assign w54234 = w54192 & ~w54218;
assign w54235 = w54198 & w54205;
assign w54236 = w54198 & ~w54211;
assign w54237 = ~w54212 & ~w54236;
assign w54238 = w54205 & ~w54211;
assign w54239 = w54237 & ~w54238;
assign w54240 = ~w54235 & ~w54239;
assign w54241 = w54234 & ~w54240;
assign w54242 = ~w54192 & ~w54218;
assign w54243 = ~w54237 & w54242;
assign w54244 = ~w54233 & ~w54243;
assign w54245 = ~w54241 & w54244;
assign w54246 = w54229 & ~w54245;
assign w54247 = ~w54192 & w54218;
assign w54248 = ~w54205 & ~w54247;
assign w54249 = ~w54234 & ~w54248;
assign w54250 = w54198 & w54211;
assign w54251 = w54249 & w54250;
assign w54252 = w54192 & w54219;
assign w54253 = ~w54221 & ~w54252;
assign w54254 = ~w54251 & w54253;
assign w54255 = ~w54229 & ~w54254;
assign w54256 = ~w54198 & w54211;
assign w54257 = ~w54249 & w54256;
assign w54258 = ~w54234 & w54257;
assign w54259 = ~w54205 & w54218;
assign w54260 = w54229 & ~w54259;
assign w54261 = w54234 & w54238;
assign w54262 = ~w54231 & ~w54261;
assign w54263 = ~w54198 & ~w54260;
assign w54264 = ~w54262 & w54263;
assign w54265 = ~w54223 & ~w54264;
assign w54266 = ~w54258 & w54265;
assign w54267 = ~w54255 & w54266;
assign w54268 = ~w54246 & w54267;
assign w54269 = pi2858 & ~w54268;
assign w54270 = ~pi2858 & w54268;
assign w54271 = ~w54269 & ~w54270;
assign w54272 = ~w54008 & ~w54020;
assign w54273 = w54037 & w54272;
assign w54274 = (w54010 & w67027) | (w54010 & w67028) | (w67027 & w67028);
assign w54275 = w54007 & ~w54023;
assign w54276 = ~w54048 & ~w54275;
assign w54277 = w54052 & ~w54273;
assign w54278 = ~w54276 & w54277;
assign w54279 = (~w54004 & ~w54278) | (~w54004 & w67029) | (~w54278 & w67029);
assign w54280 = w53990 & ~w54020;
assign w54281 = ~w54013 & ~w54280;
assign w54282 = ~w54032 & w54281;
assign w54283 = ~w54024 & w54282;
assign w54284 = ~w54047 & w67030;
assign w54285 = ~w54030 & w54284;
assign w54286 = w53983 & w54011;
assign w54287 = ~w54039 & ~w54286;
assign w54288 = w54008 & w54013;
assign w54289 = ~w54005 & ~w54288;
assign w54290 = w54020 & ~w54289;
assign w54291 = ~w53996 & w54054;
assign w54292 = (~w54291 & w54287) | (~w54291 & w64115) | (w54287 & w64115);
assign w54293 = ~w54290 & w54292;
assign w54294 = (~w54283 & w54293) | (~w54283 & w67031) | (w54293 & w67031);
assign w54295 = ~w54285 & w54294;
assign w54296 = w54295 & w67032;
assign w54297 = (~pi2855 & ~w54295) | (~pi2855 & w67033) | (~w54295 & w67033);
assign w54298 = ~w54296 & ~w54297;
assign w54299 = ~pi6508 & pi9040;
assign w54300 = ~pi6498 & ~pi9040;
assign w54301 = ~w54299 & ~w54300;
assign w54302 = pi2812 & ~w54301;
assign w54303 = ~pi2812 & w54301;
assign w54304 = ~w54302 & ~w54303;
assign w54305 = ~pi6506 & pi9040;
assign w54306 = ~pi6602 & ~pi9040;
assign w54307 = ~w54305 & ~w54306;
assign w54308 = pi2824 & ~w54307;
assign w54309 = ~pi2824 & w54307;
assign w54310 = ~w54308 & ~w54309;
assign w54311 = w54304 & ~w54310;
assign w54312 = ~pi6483 & pi9040;
assign w54313 = ~pi6464 & ~pi9040;
assign w54314 = ~w54312 & ~w54313;
assign w54315 = pi2819 & ~w54314;
assign w54316 = ~pi2819 & w54314;
assign w54317 = ~w54315 & ~w54316;
assign w54318 = ~w54311 & ~w54317;
assign w54319 = ~w54304 & w54310;
assign w54320 = ~pi6460 & pi9040;
assign w54321 = ~pi6707 & ~pi9040;
assign w54322 = ~w54320 & ~w54321;
assign w54323 = pi2833 & ~w54322;
assign w54324 = ~pi2833 & w54322;
assign w54325 = ~w54323 & ~w54324;
assign w54326 = ~pi6495 & pi9040;
assign w54327 = ~pi6499 & ~pi9040;
assign w54328 = ~w54326 & ~w54327;
assign w54329 = pi2832 & ~w54328;
assign w54330 = ~pi2832 & w54328;
assign w54331 = ~w54329 & ~w54330;
assign w54332 = ~w54325 & ~w54331;
assign w54333 = ~w54319 & w54332;
assign w54334 = ~w54318 & ~w54333;
assign w54335 = ~pi6461 & pi9040;
assign w54336 = ~pi6502 & ~pi9040;
assign w54337 = ~w54335 & ~w54336;
assign w54338 = pi2831 & ~w54337;
assign w54339 = ~pi2831 & w54337;
assign w54340 = ~w54338 & ~w54339;
assign w54341 = w54304 & w54325;
assign w54342 = ~w54317 & ~w54341;
assign w54343 = ~w54304 & ~w54310;
assign w54344 = w54331 & w54343;
assign w54345 = w54342 & ~w54344;
assign w54346 = ~w54310 & w54331;
assign w54347 = w54310 & ~w54331;
assign w54348 = ~w54346 & ~w54347;
assign w54349 = w54304 & w54348;
assign w54350 = ~w54310 & ~w54317;
assign w54351 = ~w54304 & ~w54350;
assign w54352 = ~w54348 & w54351;
assign w54353 = ~w54349 & ~w54352;
assign w54354 = ~w54325 & ~w54353;
assign w54355 = w54325 & w54343;
assign w54356 = ~w54311 & ~w54355;
assign w54357 = w54345 & w54356;
assign w54358 = ~w54354 & w54357;
assign w54359 = ~w54334 & w54340;
assign w54360 = ~w54358 & w54359;
assign w54361 = w54304 & w54310;
assign w54362 = w54331 & w54361;
assign w54363 = w54317 & ~w54343;
assign w54364 = w54319 & w54325;
assign w54365 = w54348 & ~w54364;
assign w54366 = w54363 & w54365;
assign w54367 = (~w54362 & ~w54365) | (~w54362 & w67034) | (~w54365 & w67034);
assign w54368 = w54319 & ~w54325;
assign w54369 = ~w54355 & ~w54368;
assign w54370 = w54311 & w54332;
assign w54371 = w54317 & ~w54370;
assign w54372 = w54369 & w54371;
assign w54373 = ~w54345 & ~w54372;
assign w54374 = ~w54367 & w54373;
assign w54375 = ~w54331 & w54341;
assign w54376 = ~w54344 & w54369;
assign w54377 = w54369 & w67035;
assign w54378 = ~w54317 & ~w54340;
assign w54379 = (w54378 & ~w54348) | (w54378 & w67036) | (~w54348 & w67036);
assign w54380 = w54317 & w54325;
assign w54381 = w54340 & w54380;
assign w54382 = ~w54379 & ~w54381;
assign w54383 = w54377 & ~w54382;
assign w54384 = ~w54318 & ~w54340;
assign w54385 = ~w54377 & w54384;
assign w54386 = ~w54374 & w67037;
assign w54387 = ~w54360 & w54386;
assign w54388 = pi2866 & ~w54387;
assign w54389 = ~pi2866 & w54387;
assign w54390 = ~w54388 & ~w54389;
assign w54391 = ~w53889 & ~w53903;
assign w54392 = w53882 & ~w54391;
assign w54393 = w53843 & ~w53864;
assign w54394 = w53905 & ~w54393;
assign w54395 = ~w53884 & ~w54394;
assign w54396 = ~w53897 & ~w54393;
assign w54397 = ~w53882 & ~w54396;
assign w54398 = ~w54395 & w54397;
assign w54399 = ~w54392 & ~w54398;
assign w54400 = ~w53837 & ~w54399;
assign w54401 = w53882 & ~w54393;
assign w54402 = ~w53858 & ~w53865;
assign w54403 = w54401 & ~w54402;
assign w54404 = w53849 & ~w53882;
assign w54405 = ~w54396 & w54404;
assign w54406 = ~w53870 & ~w54405;
assign w54407 = ~w54403 & w54406;
assign w54408 = w53850 & w53917;
assign w54409 = w53856 & w53908;
assign w54410 = ~w53871 & ~w53882;
assign w54411 = w53891 & ~w54409;
assign w54412 = w54410 & w54411;
assign w54413 = w53865 & w53869;
assign w54414 = w53872 & w53891;
assign w54415 = w53882 & ~w54413;
assign w54416 = ~w54414 & w54415;
assign w54417 = ~w54412 & ~w54416;
assign w54418 = (~w54408 & w54407) | (~w54408 & w67038) | (w54407 & w67038);
assign w54419 = ~w54417 & w54418;
assign w54420 = ~w54400 & w54419;
assign w54421 = pi2874 & ~w54420;
assign w54422 = ~pi2874 & w54420;
assign w54423 = ~w54421 & ~w54422;
assign w54424 = ~pi6499 & pi9040;
assign w54425 = ~pi6698 & ~pi9040;
assign w54426 = ~w54424 & ~w54425;
assign w54427 = pi2846 & ~w54426;
assign w54428 = ~pi2846 & w54426;
assign w54429 = ~w54427 & ~w54428;
assign w54430 = ~pi6514 & pi9040;
assign w54431 = ~pi6460 & ~pi9040;
assign w54432 = ~w54430 & ~w54431;
assign w54433 = pi2830 & ~w54432;
assign w54434 = ~pi2830 & w54432;
assign w54435 = ~w54433 & ~w54434;
assign w54436 = ~w54429 & w54435;
assign w54437 = ~pi6745 & pi9040;
assign w54438 = ~pi6507 & ~pi9040;
assign w54439 = ~w54437 & ~w54438;
assign w54440 = pi2822 & ~w54439;
assign w54441 = ~pi2822 & w54439;
assign w54442 = ~w54440 & ~w54441;
assign w54443 = ~w54435 & w54442;
assign w54444 = ~pi6503 & pi9040;
assign w54445 = ~pi6495 & ~pi9040;
assign w54446 = ~w54444 & ~w54445;
assign w54447 = pi2836 & ~w54446;
assign w54448 = ~pi2836 & w54446;
assign w54449 = ~w54447 & ~w54448;
assign w54450 = w54443 & w54449;
assign w54451 = ~w54429 & ~w54442;
assign w54452 = w54429 & w54442;
assign w54453 = ~w54451 & ~w54452;
assign w54454 = ~pi6681 & pi9040;
assign w54455 = ~pi6603 & ~pi9040;
assign w54456 = ~w54454 & ~w54455;
assign w54457 = pi2823 & ~w54456;
assign w54458 = ~pi2823 & w54456;
assign w54459 = ~w54457 & ~w54458;
assign w54460 = w54435 & ~w54442;
assign w54461 = w54442 & ~w54449;
assign w54462 = ~w54459 & ~w54460;
assign w54463 = ~w54461 & w54462;
assign w54464 = w54453 & w54463;
assign w54465 = ~w54429 & w54449;
assign w54466 = ~w54442 & w54459;
assign w54467 = w54465 & w54466;
assign w54468 = ~w54450 & ~w54467;
assign w54469 = ~w54464 & w54468;
assign w54470 = w54436 & ~w54469;
assign w54471 = ~pi6405 & pi9040;
assign w54472 = ~pi6503 & ~pi9040;
assign w54473 = ~w54471 & ~w54472;
assign w54474 = pi2834 & ~w54473;
assign w54475 = ~pi2834 & w54473;
assign w54476 = ~w54474 & ~w54475;
assign w54477 = ~w54435 & ~w54453;
assign w54478 = ~w54429 & ~w54459;
assign w54479 = ~w54442 & w54478;
assign w54480 = ~w54477 & ~w54479;
assign w54481 = ~w54449 & ~w54480;
assign w54482 = ~w54435 & ~w54442;
assign w54483 = ~w54452 & w54459;
assign w54484 = ~w54482 & w54483;
assign w54485 = ~w54436 & w54484;
assign w54486 = ~w54443 & ~w54460;
assign w54487 = w54429 & w54449;
assign w54488 = w54486 & w54487;
assign w54489 = ~w54476 & ~w54488;
assign w54490 = ~w54485 & w54489;
assign w54491 = ~w54481 & w54490;
assign w54492 = w54429 & ~w54459;
assign w54493 = w54460 & w54492;
assign w54494 = w54476 & ~w54493;
assign w54495 = w54442 & w54459;
assign w54496 = w54435 & w54495;
assign w54497 = ~w54435 & ~w54459;
assign w54498 = ~w54429 & ~w54497;
assign w54499 = w54452 & ~w54459;
assign w54500 = w54452 & w54497;
assign w54501 = ~w54498 & ~w54500;
assign w54502 = w54449 & ~w54501;
assign w54503 = ~w54449 & ~w54492;
assign w54504 = ~w54498 & w54503;
assign w54505 = w54494 & ~w54496;
assign w54506 = ~w54504 & w54505;
assign w54507 = ~w54502 & w54506;
assign w54508 = ~w54491 & ~w54507;
assign w54509 = ~w54470 & ~w54508;
assign w54510 = ~pi2854 & w54509;
assign w54511 = pi2854 & ~w54509;
assign w54512 = ~w54510 & ~w54511;
assign w54513 = w54192 & w54211;
assign w54514 = ~w54242 & ~w54513;
assign w54515 = w54198 & ~w54220;
assign w54516 = w54514 & w54515;
assign w54517 = w54238 & w54242;
assign w54518 = w54222 & ~w54517;
assign w54519 = ~w54198 & ~w54518;
assign w54520 = w54230 & w54513;
assign w54521 = ~w54252 & ~w54520;
assign w54522 = w54229 & ~w54516;
assign w54523 = w54521 & w54522;
assign w54524 = ~w54519 & w54523;
assign w54525 = w54199 & w54221;
assign w54526 = ~w54205 & w54242;
assign w54527 = ~w54211 & w54526;
assign w54528 = w54211 & w54242;
assign w54529 = w54205 & w54528;
assign w54530 = ~w54229 & ~w54529;
assign w54531 = ~w54205 & w54247;
assign w54532 = ~w54198 & ~w54531;
assign w54533 = ~w54219 & ~w54514;
assign w54534 = ~w54532 & ~w54533;
assign w54535 = ~w54198 & ~w54514;
assign w54536 = ~w54534 & ~w54535;
assign w54537 = ~w54525 & ~w54527;
assign w54538 = w54530 & w54537;
assign w54539 = ~w54536 & w54538;
assign w54540 = ~w54524 & ~w54539;
assign w54541 = ~w54198 & ~w54252;
assign w54542 = w54230 & w54231;
assign w54543 = w54198 & ~w54542;
assign w54544 = w54211 & w54531;
assign w54545 = ~w54527 & w54543;
assign w54546 = ~w54544 & w54545;
assign w54547 = ~w54541 & ~w54546;
assign w54548 = ~w54540 & ~w54547;
assign w54549 = ~pi2860 & w54548;
assign w54550 = pi2860 & ~w54548;
assign w54551 = ~w54549 & ~w54550;
assign w54552 = ~pi6680 & pi9040;
assign w54553 = ~pi6421 & ~pi9040;
assign w54554 = ~w54552 & ~w54553;
assign w54555 = pi2837 & ~w54554;
assign w54556 = ~pi2837 & w54554;
assign w54557 = ~w54555 & ~w54556;
assign w54558 = ~pi6507 & pi9040;
assign w54559 = ~pi6508 & ~pi9040;
assign w54560 = ~w54558 & ~w54559;
assign w54561 = pi2822 & ~w54560;
assign w54562 = ~pi2822 & w54560;
assign w54563 = ~w54561 & ~w54562;
assign w54564 = w54557 & ~w54563;
assign w54565 = ~pi6421 & pi9040;
assign w54566 = ~pi6745 & ~pi9040;
assign w54567 = ~w54565 & ~w54566;
assign w54568 = pi2832 & ~w54567;
assign w54569 = ~pi2832 & w54567;
assign w54570 = ~w54568 & ~w54569;
assign w54571 = ~pi6602 & pi9040;
assign w54572 = ~pi6461 & ~pi9040;
assign w54573 = ~w54571 & ~w54572;
assign w54574 = pi2834 & ~w54573;
assign w54575 = ~pi2834 & w54573;
assign w54576 = ~w54574 & ~w54575;
assign w54577 = ~w54570 & ~w54576;
assign w54578 = ~w54563 & w54570;
assign w54579 = w54557 & w54576;
assign w54580 = w54578 & w54579;
assign w54581 = ~w54577 & ~w54580;
assign w54582 = w54564 & ~w54581;
assign w54583 = w54557 & ~w54570;
assign w54584 = ~w54576 & ~w54578;
assign w54585 = ~w54583 & w54584;
assign w54586 = ~pi6603 & pi9040;
assign w54587 = ~pi6405 & ~pi9040;
assign w54588 = ~w54586 & ~w54587;
assign w54589 = pi2838 & ~w54588;
assign w54590 = ~pi2838 & w54588;
assign w54591 = ~w54589 & ~w54590;
assign w54592 = w54585 & w54591;
assign w54593 = w54563 & ~w54570;
assign w54594 = w54579 & w54593;
assign w54595 = ~pi6502 & pi9040;
assign w54596 = ~pi6504 & ~pi9040;
assign w54597 = ~w54595 & ~w54596;
assign w54598 = pi2812 & ~w54597;
assign w54599 = ~pi2812 & w54597;
assign w54600 = ~w54598 & ~w54599;
assign w54601 = ~w54594 & ~w54600;
assign w54602 = ~w54582 & w54601;
assign w54603 = ~w54592 & w54602;
assign w54604 = w54570 & ~w54576;
assign w54605 = w54564 & w54604;
assign w54606 = (~w54591 & ~w54584) | (~w54591 & w67039) | (~w54584 & w67039);
assign w54607 = ~w54563 & w54576;
assign w54608 = ~w54570 & w54607;
assign w54609 = w54591 & ~w54608;
assign w54610 = ~w54576 & w54593;
assign w54611 = w54557 & w54610;
assign w54612 = w54609 & ~w54611;
assign w54613 = ~w54606 & ~w54612;
assign w54614 = ~w54578 & ~w54591;
assign w54615 = ~w54557 & w54576;
assign w54616 = ~w54614 & w54615;
assign w54617 = w54570 & w54576;
assign w54618 = w54563 & w54591;
assign w54619 = w54617 & w54618;
assign w54620 = w54600 & ~w54605;
assign w54621 = ~w54619 & w54620;
assign w54622 = ~w54616 & w54621;
assign w54623 = ~w54613 & w54622;
assign w54624 = ~w54603 & ~w54623;
assign w54625 = ~w54557 & ~w54570;
assign w54626 = w54607 & ~w54625;
assign w54627 = ~w54584 & ~w54600;
assign w54628 = ~w54626 & w54627;
assign w54629 = w54557 & ~w54576;
assign w54630 = ~w54563 & w54629;
assign w54631 = ~w54594 & ~w54630;
assign w54632 = ~w54628 & w54631;
assign w54633 = ~w54591 & ~w54632;
assign w54634 = ~w54624 & ~w54633;
assign w54635 = ~pi2853 & w54634;
assign w54636 = pi2853 & ~w54634;
assign w54637 = ~w54635 & ~w54636;
assign w54638 = w54435 & w54453;
assign w54639 = (w54459 & w54453) | (w54459 & w67040) | (w54453 & w67040);
assign w54640 = ~w54638 & w54639;
assign w54641 = w54461 & w54640;
assign w54642 = ~w54435 & w54467;
assign w54643 = w54435 & ~w54449;
assign w54644 = ~w54442 & ~w54459;
assign w54645 = w54643 & w54644;
assign w54646 = w54487 & w54497;
assign w54647 = w54429 & w54643;
assign w54648 = ~w54429 & ~w54435;
assign w54649 = ~w54644 & w54648;
assign w54650 = ~w54647 & ~w54649;
assign w54651 = w54476 & w54650;
assign w54652 = w54469 & w54651;
assign w54653 = w54499 & ~w54643;
assign w54654 = w54483 & w67041;
assign w54655 = ~w54476 & ~w54654;
assign w54656 = w54429 & w54459;
assign w54657 = w54482 & w54656;
assign w54658 = ~w54443 & w54478;
assign w54659 = ~w54657 & ~w54658;
assign w54660 = ~w54449 & ~w54659;
assign w54661 = w54465 & w54495;
assign w54662 = ~w54479 & ~w54661;
assign w54663 = w54435 & ~w54662;
assign w54664 = ~w54653 & ~w54660;
assign w54665 = w54664 & w67042;
assign w54666 = ~w54652 & ~w54665;
assign w54667 = ~w54645 & ~w54646;
assign w54668 = ~w54642 & w54667;
assign w54669 = ~w54641 & w54668;
assign w54670 = ~w54666 & w54669;
assign w54671 = pi2850 & ~w54670;
assign w54672 = ~pi2850 & w54670;
assign w54673 = ~w54671 & ~w54672;
assign w54674 = w53915 & ~w54401;
assign w54675 = ~w53843 & w53865;
assign w54676 = ~w53892 & ~w54675;
assign w54677 = w53857 & w53864;
assign w54678 = ~w53910 & ~w54677;
assign w54679 = ~w53902 & ~w54394;
assign w54680 = w54678 & ~w54679;
assign w54681 = w53896 & ~w54678;
assign w54682 = ~w54680 & ~w54681;
assign w54683 = w54676 & w54682;
assign w54684 = w53882 & ~w54683;
assign w54685 = w53888 & w54404;
assign w54686 = ~w53868 & ~w54685;
assign w54687 = ~w53837 & ~w54686;
assign w54688 = ~w53904 & ~w54398;
assign w54689 = ~w54674 & ~w54687;
assign w54690 = w54688 & w54689;
assign w54691 = ~w54684 & w54690;
assign w54692 = pi2893 & ~w54691;
assign w54693 = ~pi2893 & w54691;
assign w54694 = ~w54692 & ~w54693;
assign w54695 = w54106 & ~w54114;
assign w54696 = ~w54127 & w54695;
assign w54697 = ~w54106 & w54156;
assign w54698 = ~w54125 & w54171;
assign w54699 = w54127 & w54698;
assign w54700 = ~w54170 & ~w54696;
assign w54701 = ~w54697 & w54700;
assign w54702 = (~w54069 & ~w54701) | (~w54069 & w67043) | (~w54701 & w67043);
assign w54703 = w54099 & w54134;
assign w54704 = ~w54125 & ~w54703;
assign w54705 = ~w54123 & w54704;
assign w54706 = ~w54175 & ~w54705;
assign w54707 = (~w54124 & w54141) | (~w54124 & w64116) | (w54141 & w64116);
assign w54708 = (~w54106 & ~w54707) | (~w54106 & w67044) | (~w54707 & w67044);
assign w54709 = ~w54157 & ~w54708;
assign w54710 = ~w54115 & w54704;
assign w54711 = ~w54709 & w54710;
assign w54712 = w54069 & ~w54711;
assign w54713 = ~w54702 & ~w54706;
assign w54714 = w54713 & w67045;
assign w54715 = (pi2856 & ~w54713) | (pi2856 & w67046) | (~w54713 & w67046);
assign w54716 = ~w54714 & ~w54715;
assign w54717 = ~w54449 & ~w54452;
assign w54718 = ~w54499 & ~w54717;
assign w54719 = w54486 & ~w54718;
assign w54720 = ~w54496 & ~w54647;
assign w54721 = w54719 & ~w54720;
assign w54722 = w54460 & w54465;
assign w54723 = (~w54450 & w54718) | (~w54450 & w67047) | (w54718 & w67047);
assign w54724 = ~w54453 & w67048;
assign w54725 = ~w54722 & ~w54724;
assign w54726 = w54655 & w54725;
assign w54727 = w54723 & w54726;
assign w54728 = w54463 & w54723;
assign w54729 = w54494 & ~w54640;
assign w54730 = ~w54728 & w54729;
assign w54731 = ~w54727 & ~w54730;
assign w54732 = ~w54721 & ~w54731;
assign w54733 = ~pi2865 & w54732;
assign w54734 = pi2865 & ~w54732;
assign w54735 = ~w54733 & ~w54734;
assign w54736 = ~w54261 & ~w54520;
assign w54737 = ~w54527 & w54736;
assign w54738 = ~w54198 & ~w54737;
assign w54739 = ~w54218 & ~w54235;
assign w54740 = ~w54232 & w54739;
assign w54741 = w54236 & ~w54242;
assign w54742 = w54249 & w54741;
assign w54743 = ~w54231 & ~w54236;
assign w54744 = w54259 & w54743;
assign w54745 = ~w54740 & ~w54744;
assign w54746 = w54530 & w54745;
assign w54747 = ~w54742 & w54746;
assign w54748 = ~w54212 & w54247;
assign w54749 = ~w54252 & ~w54748;
assign w54750 = ~w54198 & ~w54749;
assign w54751 = w54242 & w54250;
assign w54752 = w54229 & ~w54751;
assign w54753 = ~w54525 & w54752;
assign w54754 = w54736 & w54753;
assign w54755 = ~w54750 & w54754;
assign w54756 = ~w54747 & ~w54755;
assign w54757 = ~w54230 & w54250;
assign w54758 = ~w54248 & w54757;
assign w54759 = ~w54738 & ~w54758;
assign w54760 = ~w54756 & w54759;
assign w54761 = pi2875 & ~w54760;
assign w54762 = ~pi2875 & w54760;
assign w54763 = ~w54761 & ~w54762;
assign w54764 = (~w54722 & w54650) | (~w54722 & w67049) | (w54650 & w67049);
assign w54765 = ~w54459 & ~w54764;
assign w54766 = w54461 & w54656;
assign w54767 = (w54766 & ~w54650) | (w54766 & w67050) | (~w54650 & w67050);
assign w54768 = ~w54435 & w54644;
assign w54769 = ~w54661 & ~w54722;
assign w54770 = ~w54768 & w54769;
assign w54771 = w54720 & w54770;
assign w54772 = ~w54476 & ~w54771;
assign w54773 = ~w54429 & ~w54486;
assign w54774 = ~w54657 & ~w54773;
assign w54775 = (~w54449 & w54773) | (~w54449 & w67051) | (w54773 & w67051);
assign w54776 = ~w54501 & ~w54503;
assign w54777 = w54774 & w54776;
assign w54778 = ~w54654 & ~w54775;
assign w54779 = ~w54777 & w54778;
assign w54780 = w54476 & ~w54779;
assign w54781 = ~w54646 & ~w54767;
assign w54782 = ~w54765 & w54781;
assign w54783 = ~w54772 & w54782;
assign w54784 = ~w54780 & w54783;
assign w54785 = pi2864 & ~w54784;
assign w54786 = ~pi2864 & w54784;
assign w54787 = ~w54785 & ~w54786;
assign w54788 = w54332 & w54343;
assign w54789 = w54325 & w54347;
assign w54790 = ~w54788 & ~w54789;
assign w54791 = w54317 & ~w54790;
assign w54792 = w54325 & w54331;
assign w54793 = w54343 & ~w54792;
assign w54794 = w54340 & ~w54793;
assign w54795 = ~w54366 & w54794;
assign w54796 = ~w54791 & ~w54795;
assign w54797 = ~w54317 & ~w54343;
assign w54798 = ~w54365 & w54797;
assign w54799 = ~w54796 & ~w54798;
assign w54800 = ~w54317 & w54319;
assign w54801 = ~w54311 & ~w54800;
assign w54802 = ~w54332 & ~w54792;
assign w54803 = ~w54364 & w54802;
assign w54804 = w54801 & ~w54803;
assign w54805 = ~w54801 & w54802;
assign w54806 = ~w54340 & ~w54804;
assign w54807 = ~w54805 & w54806;
assign w54808 = ~w54799 & ~w54807;
assign w54809 = ~pi2876 & w54808;
assign w54810 = pi2876 & ~w54808;
assign w54811 = ~w54809 & ~w54810;
assign w54812 = ~w54020 & w54287;
assign w54813 = w54012 & w54050;
assign w54814 = w54012 & w53997;
assign w54815 = w53984 & ~w53997;
assign w54816 = ~w54281 & w54815;
assign w54817 = ~w54813 & ~w54814;
assign w54818 = ~w54816 & w54817;
assign w54819 = w53977 & w54818;
assign w54820 = w54812 & ~w54819;
assign w54821 = (~w54004 & w54047) | (~w54004 & w67052) | (w54047 & w67052);
assign w54822 = ~w54051 & ~w54814;
assign w54823 = w54020 & ~w54822;
assign w54824 = ~w54287 & w67053;
assign w54825 = ~w54823 & ~w54824;
assign w54826 = ~w54821 & w54825;
assign w54827 = ~w54820 & ~w54826;
assign w54828 = ~w53983 & ~w54026;
assign w54829 = ~w54047 & w67054;
assign w54830 = w54287 & w67055;
assign w54831 = w54818 & ~w54830;
assign w54832 = ~w54829 & w54831;
assign w54833 = w54004 & ~w54832;
assign w54834 = ~w54827 & ~w54833;
assign w54835 = pi2862 & w54834;
assign w54836 = ~pi2862 & ~w54834;
assign w54837 = ~w54835 & ~w54836;
assign w54838 = w54570 & w54629;
assign w54839 = w54629 & w67056;
assign w54840 = ~w54563 & ~w54591;
assign w54841 = ~w54563 & w54625;
assign w54842 = ~w54838 & ~w54841;
assign w54843 = w54840 & w54842;
assign w54844 = w54842 & w67057;
assign w54845 = ~w54839 & ~w54844;
assign w54846 = w54557 & w54591;
assign w54847 = ~w54576 & ~w54846;
assign w54848 = ~w54845 & w54847;
assign w54849 = ~w54578 & ~w54593;
assign w54850 = ~w54617 & ~w54849;
assign w54851 = ~w54849 & w67058;
assign w54852 = w54604 & w54840;
assign w54853 = ~w54600 & ~w54852;
assign w54854 = w54578 & w54591;
assign w54855 = ~w54614 & ~w54854;
assign w54856 = w54579 & ~w54855;
assign w54857 = ~w54851 & w54853;
assign w54858 = ~w54856 & w54857;
assign w54859 = w54845 & w54858;
assign w54860 = w54618 & ~w54629;
assign w54861 = ~w54606 & ~w54840;
assign w54862 = ~w54581 & ~w54861;
assign w54863 = w54615 & w54849;
assign w54864 = w54600 & ~w54860;
assign w54865 = ~w54863 & w54864;
assign w54866 = ~w54862 & w54865;
assign w54867 = ~w54859 & ~w54866;
assign w54868 = ~w54557 & w54563;
assign w54869 = ~w54564 & ~w54868;
assign w54870 = ~w54583 & ~w54615;
assign w54871 = ~w54869 & ~w54870;
assign w54872 = w54609 & w54871;
assign w54873 = ~w54848 & ~w54872;
assign w54874 = ~w54867 & w54873;
assign w54875 = pi2863 & ~w54874;
assign w54876 = ~pi2863 & w54874;
assign w54877 = ~w54875 & ~w54876;
assign w54878 = ~w54361 & w54792;
assign w54879 = ~w54341 & ~w54346;
assign w54880 = w54340 & ~w54347;
assign w54881 = w54317 & ~w54879;
assign w54882 = ~w54880 & w54881;
assign w54883 = ~w54878 & ~w54882;
assign w54884 = ~w54340 & ~w54350;
assign w54885 = w54878 & w54884;
assign w54886 = ~w54883 & ~w54885;
assign w54887 = w54340 & w54373;
assign w54888 = ~w54304 & ~w54331;
assign w54889 = w54310 & w54332;
assign w54890 = ~w54888 & ~w54889;
assign w54891 = ~w54340 & ~w54890;
assign w54892 = w54376 & w54891;
assign w54893 = w54378 & ~w54888;
assign w54894 = w54879 & w54893;
assign w54895 = ~w54892 & ~w54894;
assign w54896 = ~w54886 & w54895;
assign w54897 = ~w54887 & w54896;
assign w54898 = pi2884 & ~w54897;
assign w54899 = ~pi2884 & w54897;
assign w54900 = ~w54898 & ~w54899;
assign w54901 = (~w54788 & ~w54353) | (~w54788 & w67059) | (~w54353 & w67059);
assign w54902 = ~w54340 & ~w54901;
assign w54903 = w54342 & ~w54356;
assign w54904 = w54331 & w54364;
assign w54905 = ~w54903 & ~w54904;
assign w54906 = ~w54354 & w54905;
assign w54907 = w54340 & ~w54906;
assign w54908 = ~w54343 & ~w54888;
assign w54909 = ~w54355 & ~w54908;
assign w54910 = (~w54340 & w54909) | (~w54340 & w67060) | (w54909 & w67060);
assign w54911 = ~w54375 & ~w54910;
assign w54912 = ~w54317 & ~w54911;
assign w54913 = ~w54310 & w54380;
assign w54914 = w54353 & w54913;
assign w54915 = ~w54902 & ~w54914;
assign w54916 = ~w54907 & ~w54912;
assign w54917 = (~pi2883 & ~w54916) | (~pi2883 & w67061) | (~w54916 & w67061);
assign w54918 = w54916 & w67062;
assign w54919 = ~w54917 & ~w54918;
assign w54920 = ~w54012 & w54050;
assign w54921 = ~w53997 & w54032;
assign w54922 = w54272 & ~w54921;
assign w54923 = w54024 & ~w54026;
assign w54924 = ~w54922 & ~w54923;
assign w54925 = ~w54920 & ~w54924;
assign w54926 = ~w54004 & ~w54925;
assign w54927 = ~w54014 & ~w54920;
assign w54928 = ~w54047 & w67063;
assign w54929 = (~w54814 & w54289) | (~w54814 & w67064) | (w54289 & w67064);
assign w54930 = ~w54020 & ~w54929;
assign w54931 = ~w53998 & ~w54813;
assign w54932 = ~w54273 & w54931;
assign w54933 = ~w54041 & w54932;
assign w54934 = w54004 & ~w54933;
assign w54935 = ~w54928 & ~w54930;
assign w54936 = ~w54934 & w54935;
assign w54937 = ~w54926 & w54936;
assign w54938 = ~pi2871 & w54937;
assign w54939 = pi2871 & ~w54937;
assign w54940 = ~w54938 & ~w54939;
assign w54941 = w54140 & w54168;
assign w54942 = ~w54082 & ~w54169;
assign w54943 = w54124 & ~w54176;
assign w54944 = ~w54941 & ~w54943;
assign w54945 = (w54132 & w67065) | (w54132 & w67066) | (w67065 & w67066);
assign w54946 = w54069 & ~w54132;
assign w54947 = ~w54082 & w54146;
assign w54948 = ~w54141 & w54947;
assign w54949 = (~w54948 & ~w54158) | (~w54948 & w67067) | (~w54158 & w67067);
assign w54950 = ~w54946 & w54949;
assign w54951 = w54950 & w67068;
assign w54952 = (~pi2859 & ~w54950) | (~pi2859 & w67069) | (~w54950 & w67069);
assign w54953 = ~w54951 & ~w54952;
assign w54954 = ~w54528 & w54737;
assign w54955 = w54235 & ~w54954;
assign w54956 = ~w54238 & ~w54748;
assign w54957 = ~w54220 & ~w54956;
assign w54958 = ~w54542 & w54741;
assign w54959 = w54229 & ~w54958;
assign w54960 = ~w54257 & w54959;
assign w54961 = ~w54957 & w54960;
assign w54962 = ~w54526 & w54543;
assign w54963 = w54192 & w54220;
assign w54964 = w54532 & ~w54963;
assign w54965 = ~w54962 & ~w54964;
assign w54966 = ~w54229 & ~w54544;
assign w54967 = w54521 & w54966;
assign w54968 = ~w54965 & w54967;
assign w54969 = ~w54961 & ~w54968;
assign w54970 = ~w54192 & ~w54198;
assign w54971 = w54957 & w54970;
assign w54972 = ~w54955 & ~w54971;
assign w54973 = ~w54969 & w54972;
assign w54974 = ~pi2877 & w54973;
assign w54975 = pi2877 & ~w54973;
assign w54976 = ~w54974 & ~w54975;
assign w54977 = w54591 & ~w54600;
assign w54978 = w54617 & w54868;
assign w54979 = ~w54605 & ~w54610;
assign w54980 = ~w54863 & w54979;
assign w54981 = ~w54594 & ~w54978;
assign w54982 = (w54981 & w54980) | (w54981 & w67070) | (w54980 & w67070);
assign w54983 = ~w54977 & ~w54982;
assign w54984 = w54600 & ~w54842;
assign w54985 = w54601 & ~w54604;
assign w54986 = w54980 & w54985;
assign w54987 = ~w54984 & ~w54986;
assign w54988 = w54591 & ~w54987;
assign w54989 = w54593 & w67071;
assign w54990 = ~w54839 & ~w54989;
assign w54991 = (w54600 & w54843) | (w54600 & w67072) | (w54843 & w67072);
assign w54992 = ~w54557 & w54604;
assign w54993 = w54853 & w54992;
assign w54994 = ~w54991 & ~w54993;
assign w54995 = ~w54983 & w54994;
assign w54996 = ~w54988 & w54995;
assign w54997 = pi2867 & ~w54996;
assign w54998 = ~pi2867 & w54996;
assign w54999 = ~w54997 & ~w54998;
assign w55000 = w53914 & w54394;
assign w55001 = ~w53875 & ~w53912;
assign w55002 = w53837 & ~w55001;
assign w55003 = ~w53903 & ~w53909;
assign w55004 = (~w53902 & w55002) | (~w53902 & w67073) | (w55002 & w67073);
assign w55005 = ~w53882 & ~w55004;
assign w55006 = w53850 & w53864;
assign w55007 = w53837 & ~w53849;
assign w55008 = w53856 & w54393;
assign w55009 = ~w55007 & w55008;
assign w55010 = ~w53866 & ~w53907;
assign w55011 = w53857 & ~w55010;
assign w55012 = w53882 & ~w55006;
assign w55013 = ~w55009 & w55012;
assign w55014 = ~w55011 & w55013;
assign w55015 = ~w55005 & ~w55014;
assign w55016 = ~w54676 & w55007;
assign w55017 = ~w53837 & w53873;
assign w55018 = ~w54401 & w55017;
assign w55019 = ~w55000 & ~w55018;
assign w55020 = ~w55016 & w55019;
assign w55021 = ~w55015 & w55020;
assign w55022 = ~pi2898 & ~w55021;
assign w55023 = pi2898 & w55021;
assign w55024 = ~w55022 & ~w55023;
assign w55025 = w54604 & w54614;
assign w55026 = w54600 & w54850;
assign w55027 = ~w54989 & ~w55026;
assign w55028 = w54591 & ~w55027;
assign w55029 = w54617 & w54846;
assign w55030 = w54576 & w54591;
assign w55031 = ~w54593 & ~w55030;
assign w55032 = ~w54870 & w55031;
assign w55033 = w54600 & ~w55032;
assign w55034 = w54847 & w54869;
assign w55035 = ~w54580 & ~w54619;
assign w55036 = ~w54841 & w55035;
assign w55037 = w54601 & ~w55034;
assign w55038 = w55036 & w55037;
assign w55039 = ~w55033 & ~w55038;
assign w55040 = ~w55025 & ~w55029;
assign w55041 = ~w55028 & w55040;
assign w55042 = ~w55039 & w55041;
assign w55043 = pi2889 & ~w55042;
assign w55044 = ~pi2889 & w55042;
assign w55045 = ~w55043 & ~w55044;
assign w55046 = ~pi6671 & pi9040;
assign w55047 = ~pi6732 & ~pi9040;
assign w55048 = ~w55046 & ~w55047;
assign w55049 = pi2911 & ~w55048;
assign w55050 = ~pi2911 & w55048;
assign w55051 = ~w55049 & ~w55050;
assign w55052 = ~pi6676 & pi9040;
assign w55053 = ~pi6839 & ~pi9040;
assign w55054 = ~w55052 & ~w55053;
assign w55055 = pi2905 & ~w55054;
assign w55056 = ~pi2905 & w55054;
assign w55057 = ~w55055 & ~w55056;
assign w55058 = ~pi6668 & pi9040;
assign w55059 = ~pi6794 & ~pi9040;
assign w55060 = ~w55058 & ~w55059;
assign w55061 = pi2881 & ~w55060;
assign w55062 = ~pi2881 & w55060;
assign w55063 = ~w55061 & ~w55062;
assign w55064 = w55057 & w55063;
assign w55065 = ~pi6684 & pi9040;
assign w55066 = ~pi6806 & ~pi9040;
assign w55067 = ~w55065 & ~w55066;
assign w55068 = pi2908 & ~w55067;
assign w55069 = ~pi2908 & w55067;
assign w55070 = ~w55068 & ~w55069;
assign w55071 = w55064 & w55070;
assign w55072 = ~w55051 & w55071;
assign w55073 = ~w55051 & ~w55070;
assign w55074 = w55057 & w55073;
assign w55075 = ~w55057 & ~w55063;
assign w55076 = w55051 & ~w55070;
assign w55077 = w55075 & w55076;
assign w55078 = ~w55057 & w55070;
assign w55079 = ~w55051 & w55070;
assign w55080 = ~w55064 & ~w55075;
assign w55081 = ~w55079 & w55080;
assign w55082 = w55080 & w64118;
assign w55083 = ~w55077 & ~w55082;
assign w55084 = ~w55082 & w67074;
assign w55085 = ~pi6737 & pi9040;
assign w55086 = ~pi6655 & ~pi9040;
assign w55087 = ~w55085 & ~w55086;
assign w55088 = pi2900 & ~w55087;
assign w55089 = ~pi2900 & w55087;
assign w55090 = ~w55088 & ~w55089;
assign w55091 = w55063 & w55073;
assign w55092 = w55090 & ~w55091;
assign w55093 = ~w55084 & w55092;
assign w55094 = ~w55051 & w55063;
assign w55095 = ~w55064 & ~w55094;
assign w55096 = ~w55057 & w55090;
assign w55097 = ~w55076 & ~w55096;
assign w55098 = ~w55095 & ~w55097;
assign w55099 = ~w55063 & ~w55073;
assign w55100 = ~w55078 & w55099;
assign w55101 = w55063 & w55070;
assign w55102 = ~w55090 & ~w55094;
assign w55103 = ~w55101 & w55102;
assign w55104 = ~w55100 & w55103;
assign w55105 = ~pi6663 & pi9040;
assign w55106 = ~pi6811 & ~pi9040;
assign w55107 = ~w55105 & ~w55106;
assign w55108 = pi2901 & ~w55107;
assign w55109 = ~pi2901 & w55107;
assign w55110 = ~w55108 & ~w55109;
assign w55111 = (~w55110 & w55104) | (~w55110 & w67075) | (w55104 & w67075);
assign w55112 = ~w55063 & w55070;
assign w55113 = ~w55079 & ~w55090;
assign w55114 = w55112 & w55113;
assign w55115 = w55075 & w55079;
assign w55116 = ~w55071 & ~w55115;
assign w55117 = w55090 & ~w55116;
assign w55118 = w55063 & ~w55084;
assign w55119 = ~w55070 & w55090;
assign w55120 = w55095 & w55119;
assign w55121 = w55057 & w55112;
assign w55122 = ~w55091 & ~w55121;
assign w55123 = ~w55090 & ~w55122;
assign w55124 = ~w55117 & ~w55120;
assign w55125 = ~w55123 & w55124;
assign w55126 = (w55110 & ~w55125) | (w55110 & w67076) | (~w55125 & w67076);
assign w55127 = ~w55072 & ~w55114;
assign w55128 = ~w55111 & w55127;
assign w55129 = ~w55093 & w55128;
assign w55130 = ~w55126 & w55129;
assign w55131 = pi2921 & ~w55130;
assign w55132 = ~pi2921 & w55130;
assign w55133 = ~w55131 & ~w55132;
assign w55134 = w55076 & w55080;
assign w55135 = w55113 & ~w55134;
assign w55136 = w55090 & ~w55134;
assign w55137 = w55073 & w55075;
assign w55138 = ~w55121 & ~w55137;
assign w55139 = w55136 & w55138;
assign w55140 = w55110 & ~w55135;
assign w55141 = ~w55139 & w55140;
assign w55142 = (~w55091 & w55116) | (~w55091 & w67077) | (w55116 & w67077);
assign w55143 = w55083 & w55142;
assign w55144 = ~w55110 & ~w55143;
assign w55145 = ~w55118 & w55136;
assign w55146 = w55051 & w55070;
assign w55147 = w55075 & w55146;
assign w55148 = w55057 & ~w55110;
assign w55149 = ~w55101 & w55148;
assign w55150 = ~w55134 & w55149;
assign w55151 = ~w55090 & ~w55147;
assign w55152 = ~w55150 & w55151;
assign w55153 = ~w55145 & ~w55152;
assign w55154 = ~w55141 & ~w55144;
assign w55155 = ~w55153 & w55154;
assign w55156 = ~pi2926 & w55155;
assign w55157 = pi2926 & ~w55155;
assign w55158 = ~w55156 & ~w55157;
assign w55159 = ~pi6738 & pi9040;
assign w55160 = ~pi6765 & ~pi9040;
assign w55161 = ~w55159 & ~w55160;
assign w55162 = pi2903 & ~w55161;
assign w55163 = ~pi2903 & w55161;
assign w55164 = ~w55162 & ~w55163;
assign w55165 = ~pi6987 & pi9040;
assign w55166 = ~pi6736 & ~pi9040;
assign w55167 = ~w55165 & ~w55166;
assign w55168 = pi2897 & ~w55167;
assign w55169 = ~pi2897 & w55167;
assign w55170 = ~w55168 & ~w55169;
assign w55171 = w55164 & ~w55170;
assign w55172 = ~pi6727 & pi9040;
assign w55173 = ~pi6722 & ~pi9040;
assign w55174 = ~w55172 & ~w55173;
assign w55175 = pi2872 & ~w55174;
assign w55176 = ~pi2872 & w55174;
assign w55177 = ~w55175 & ~w55176;
assign w55178 = w55171 & ~w55177;
assign w55179 = w55164 & w55170;
assign w55180 = ~pi6667 & pi9040;
assign w55181 = ~pi6809 & ~pi9040;
assign w55182 = ~w55180 & ~w55181;
assign w55183 = pi2895 & ~w55182;
assign w55184 = ~pi2895 & w55182;
assign w55185 = ~w55183 & ~w55184;
assign w55186 = w55177 & ~w55185;
assign w55187 = w55179 & w55186;
assign w55188 = ~w55178 & ~w55187;
assign w55189 = ~pi6765 & pi9040;
assign w55190 = ~pi6674 & ~pi9040;
assign w55191 = ~w55189 & ~w55190;
assign w55192 = pi2878 & ~w55191;
assign w55193 = ~pi2878 & w55191;
assign w55194 = ~w55192 & ~w55193;
assign w55195 = ~w55188 & ~w55194;
assign w55196 = ~w55177 & w55185;
assign w55197 = ~w55170 & ~w55196;
assign w55198 = w55164 & ~w55185;
assign w55199 = w55197 & ~w55198;
assign w55200 = w55197 & w67078;
assign w55201 = ~pi6735 & pi9040;
assign w55202 = ~pi6766 & ~pi9040;
assign w55203 = ~w55201 & ~w55202;
assign w55204 = pi2890 & ~w55203;
assign w55205 = ~pi2890 & w55203;
assign w55206 = ~w55204 & ~w55205;
assign w55207 = w55170 & w55185;
assign w55208 = w55177 & w55194;
assign w55209 = w55207 & w55208;
assign w55210 = ~w55164 & w55170;
assign w55211 = w55194 & w55210;
assign w55212 = ~w55170 & w55186;
assign w55213 = w55186 & w67079;
assign w55214 = w55194 & ~w55213;
assign w55215 = ~w55177 & ~w55185;
assign w55216 = w55170 & w55215;
assign w55217 = ~w55212 & ~w55216;
assign w55218 = w55214 & ~w55217;
assign w55219 = ~w55186 & ~w55196;
assign w55220 = w55179 & ~w55219;
assign w55221 = w55164 & w55194;
assign w55222 = ~w55164 & w55177;
assign w55223 = ~w55221 & ~w55222;
assign w55224 = (~w55170 & ~w55171) | (~w55170 & w67080) | (~w55171 & w67080);
assign w55225 = w55223 & w55224;
assign w55226 = ~w55220 & ~w55225;
assign w55227 = w55196 & w55226;
assign w55228 = w55206 & ~w55209;
assign w55229 = ~w55211 & w55228;
assign w55230 = ~w55200 & w55229;
assign w55231 = ~w55218 & w55230;
assign w55232 = ~w55227 & w55231;
assign w55233 = w55170 & w55196;
assign w55234 = (~w55194 & ~w55196) | (~w55194 & w67081) | (~w55196 & w67081);
assign w55235 = ~w55177 & w55198;
assign w55236 = w55234 & ~w55235;
assign w55237 = ~w55197 & w55236;
assign w55238 = w55171 & w55215;
assign w55239 = w55194 & w55199;
assign w55240 = ~w55206 & ~w55238;
assign w55241 = ~w55220 & w55240;
assign w55242 = ~w55239 & w55241;
assign w55243 = ~w55237 & w55242;
assign w55244 = (~w55195 & w55232) | (~w55195 & w67082) | (w55232 & w67082);
assign w55245 = pi2918 & w55244;
assign w55246 = ~pi2918 & ~w55244;
assign w55247 = ~w55245 & ~w55246;
assign w55248 = ~pi6774 & pi9040;
assign w55249 = ~pi6896 & ~pi9040;
assign w55250 = ~w55248 & ~w55249;
assign w55251 = pi2880 & ~w55250;
assign w55252 = ~pi2880 & w55250;
assign w55253 = ~w55251 & ~w55252;
assign w55254 = ~pi6896 & pi9040;
assign w55255 = ~pi6730 & ~pi9040;
assign w55256 = ~w55254 & ~w55255;
assign w55257 = pi2899 & ~w55256;
assign w55258 = ~pi2899 & w55256;
assign w55259 = ~w55257 & ~w55258;
assign w55260 = w55253 & ~w55259;
assign w55261 = ~pi6634 & pi9040;
assign w55262 = ~pi6661 & ~pi9040;
assign w55263 = ~w55261 & ~w55262;
assign w55264 = pi2886 & ~w55263;
assign w55265 = ~pi2886 & w55263;
assign w55266 = ~w55264 & ~w55265;
assign w55267 = w55260 & ~w55266;
assign w55268 = ~w55253 & w55259;
assign w55269 = ~pi6632 & pi9040;
assign w55270 = ~pi6735 & ~pi9040;
assign w55271 = ~w55269 & ~w55270;
assign w55272 = pi2881 & ~w55271;
assign w55273 = ~pi2881 & w55271;
assign w55274 = ~w55272 & ~w55273;
assign w55275 = ~w55266 & w55274;
assign w55276 = w55268 & w55275;
assign w55277 = ~w55267 & ~w55276;
assign w55278 = ~pi6658 & pi9040;
assign w55279 = ~pi6853 & ~pi9040;
assign w55280 = ~w55278 & ~w55279;
assign w55281 = pi2909 & ~w55280;
assign w55282 = ~pi2909 & w55280;
assign w55283 = ~w55281 & ~w55282;
assign w55284 = w55274 & w55283;
assign w55285 = ~pi6807 & pi9040;
assign w55286 = ~pi6721 & ~pi9040;
assign w55287 = ~w55285 & ~w55286;
assign w55288 = pi2908 & ~w55287;
assign w55289 = ~pi2908 & w55287;
assign w55290 = ~w55288 & ~w55289;
assign w55291 = ~w55284 & w55290;
assign w55292 = ~w55277 & ~w55291;
assign w55293 = ~w55253 & w55274;
assign w55294 = ~w55266 & ~w55293;
assign w55295 = w55259 & ~w55266;
assign w55296 = ~w55293 & ~w55295;
assign w55297 = ~w55259 & w55274;
assign w55298 = w55253 & ~w55274;
assign w55299 = ~w55297 & ~w55298;
assign w55300 = ~w55296 & w55299;
assign w55301 = ~w55283 & w55300;
assign w55302 = ~w55283 & ~w55297;
assign w55303 = w55266 & ~w55274;
assign w55304 = w55253 & w55303;
assign w55305 = (w55302 & ~w55277) | (w55302 & w67083) | (~w55277 & w67083);
assign w55306 = ~w55301 & ~w55305;
assign w55307 = w55294 & ~w55306;
assign w55308 = ~w55253 & w55266;
assign w55309 = ~w55303 & ~w55308;
assign w55310 = ~w55294 & w55309;
assign w55311 = ~w55276 & ~w55283;
assign w55312 = w55310 & w55311;
assign w55313 = ~w55253 & ~w55274;
assign w55314 = ~w55259 & ~w55283;
assign w55315 = w55313 & w55314;
assign w55316 = w55259 & w55313;
assign w55317 = w55313 & w67084;
assign w55318 = ~w55315 & ~w55317;
assign w55319 = ~w55259 & ~w55284;
assign w55320 = ~w55309 & ~w55319;
assign w55321 = ~w55313 & ~w55320;
assign w55322 = w55318 & ~w55321;
assign w55323 = w55290 & ~w55312;
assign w55324 = ~w55322 & w55323;
assign w55325 = w55259 & w55283;
assign w55326 = ~w55300 & w55325;
assign w55327 = ~w55310 & w55314;
assign w55328 = ~w55290 & ~w55326;
assign w55329 = ~w55327 & w55328;
assign w55330 = ~w55324 & ~w55329;
assign w55331 = ~w55292 & ~w55307;
assign w55332 = ~w55330 & w55331;
assign w55333 = pi2929 & ~w55332;
assign w55334 = ~pi2929 & w55332;
assign w55335 = ~w55333 & ~w55334;
assign w55336 = w55308 & w55325;
assign w55337 = w55283 & ~w55299;
assign w55338 = w55302 & ~w55304;
assign w55339 = (~w55268 & w55299) | (~w55268 & w67085) | (w55299 & w67085);
assign w55340 = ~w55338 & w55339;
assign w55341 = ~w55260 & ~w55268;
assign w55342 = w55294 & w55341;
assign w55343 = ~w55253 & w55342;
assign w55344 = w55260 & w55275;
assign w55345 = ~w55336 & ~w55344;
assign w55346 = ~w55317 & w55345;
assign w55347 = ~w55343 & w55346;
assign w55348 = (~w55290 & ~w55347) | (~w55290 & w67086) | (~w55347 & w67086);
assign w55349 = w55295 & w55337;
assign w55350 = ~w55266 & ~w55283;
assign w55351 = ~w55341 & w55350;
assign w55352 = ~w55299 & w67087;
assign w55353 = w55259 & w55310;
assign w55354 = w55266 & w55315;
assign w55355 = ~w55351 & ~w55354;
assign w55356 = ~w55352 & w55355;
assign w55357 = (w55290 & ~w55356) | (w55290 & w67088) | (~w55356 & w67088);
assign w55358 = ~w55275 & w55283;
assign w55359 = ~w55253 & ~w55266;
assign w55360 = w55303 & w55260;
assign w55361 = ~w55359 & ~w55360;
assign w55362 = w55358 & ~w55361;
assign w55363 = ~w55353 & ~w55362;
assign w55364 = ~w55325 & ~w55361;
assign w55365 = ~w55363 & w55364;
assign w55366 = ~w55348 & ~w55349;
assign w55367 = ~w55357 & ~w55365;
assign w55368 = w55366 & w55367;
assign w55369 = pi2923 & ~w55368;
assign w55370 = ~pi2923 & w55368;
assign w55371 = ~w55369 & ~w55370;
assign w55372 = ~pi6726 & pi9040;
assign w55373 = ~pi6670 & ~pi9040;
assign w55374 = ~w55372 & ~w55373;
assign w55375 = pi2868 & ~w55374;
assign w55376 = ~pi2868 & w55374;
assign w55377 = ~w55375 & ~w55376;
assign w55378 = ~pi6739 & pi9040;
assign w55379 = ~pi6801 & ~pi9040;
assign w55380 = ~w55378 & ~w55379;
assign w55381 = pi2879 & ~w55380;
assign w55382 = ~pi2879 & w55380;
assign w55383 = ~w55381 & ~w55382;
assign w55384 = ~w55377 & ~w55383;
assign w55385 = ~pi6828 & pi9040;
assign w55386 = ~pi6699 & ~pi9040;
assign w55387 = ~w55385 & ~w55386;
assign w55388 = pi2901 & ~w55387;
assign w55389 = ~pi2901 & w55387;
assign w55390 = ~w55388 & ~w55389;
assign w55391 = w55383 & w55390;
assign w55392 = w55377 & w55391;
assign w55393 = ~w55384 & ~w55392;
assign w55394 = ~pi6662 & pi9040;
assign w55395 = ~pi6671 & ~pi9040;
assign w55396 = ~w55394 & ~w55395;
assign w55397 = pi2905 & ~w55396;
assign w55398 = ~pi2905 & w55396;
assign w55399 = ~w55397 & ~w55398;
assign w55400 = ~w55390 & w55399;
assign w55401 = ~w55391 & ~w55400;
assign w55402 = ~w55377 & w55399;
assign w55403 = w55390 & w55402;
assign w55404 = ~w55377 & w55383;
assign w55405 = ~pi6660 & pi9040;
assign w55406 = ~pi6769 & ~pi9040;
assign w55407 = ~w55405 & ~w55406;
assign w55408 = pi2894 & ~w55407;
assign w55409 = ~pi2894 & w55407;
assign w55410 = ~w55408 & ~w55409;
assign w55411 = ~w55404 & ~w55410;
assign w55412 = ~w55403 & ~w55411;
assign w55413 = ~w55401 & w55412;
assign w55414 = ~pi6672 & pi9040;
assign w55415 = ~pi6668 & ~pi9040;
assign w55416 = ~w55414 & ~w55415;
assign w55417 = pi2904 & ~w55416;
assign w55418 = ~pi2904 & w55416;
assign w55419 = ~w55417 & ~w55418;
assign w55420 = ~w55390 & ~w55410;
assign w55421 = w55384 & w55420;
assign w55422 = w55390 & ~w55410;
assign w55423 = ~w55383 & w55399;
assign w55424 = w55383 & ~w55399;
assign w55425 = ~w55423 & ~w55424;
assign w55426 = w55377 & w55425;
assign w55427 = w55425 & w63443;
assign w55428 = ~w55421 & ~w55427;
assign w55429 = w55410 & ~w55424;
assign w55430 = ~w55393 & ~w55429;
assign w55431 = w55428 & w55430;
assign w55432 = w55383 & w55410;
assign w55433 = ~w55390 & w55432;
assign w55434 = ~w55403 & ~w55433;
assign w55435 = ~w55425 & ~w55434;
assign w55436 = w55377 & ~w55399;
assign w55437 = w55390 & ~w55436;
assign w55438 = w55377 & ~w55390;
assign w55439 = (w55410 & w55437) | (w55410 & w67089) | (w55437 & w67089);
assign w55440 = w55377 & w55400;
assign w55441 = (~w55410 & ~w55402) | (~w55410 & w55420) | (~w55402 & w55420);
assign w55442 = ~w55440 & w55441;
assign w55443 = ~w55439 & ~w55442;
assign w55444 = ~w55435 & ~w55443;
assign w55445 = ~w55431 & w55444;
assign w55446 = ~w55419 & ~w55445;
assign w55447 = w55425 & w55437;
assign w55448 = w55410 & ~w55440;
assign w55449 = ~w55447 & w55448;
assign w55450 = w55377 & w55401;
assign w55451 = ~w55410 & ~w55450;
assign w55452 = ~w55413 & w55451;
assign w55453 = w55419 & ~w55449;
assign w55454 = ~w55452 & w55453;
assign w55455 = w55390 & w55410;
assign w55456 = ~w55377 & ~w55455;
assign w55457 = w55435 & w55456;
assign w55458 = ~w55399 & w55421;
assign w55459 = (~w55458 & ~w55413) | (~w55458 & w67090) | (~w55413 & w67090);
assign w55460 = ~w55457 & w55459;
assign w55461 = ~w55454 & w55460;
assign w55462 = ~w55446 & w55461;
assign w55463 = pi2920 & ~w55462;
assign w55464 = ~pi2920 & w55462;
assign w55465 = ~w55463 & ~w55464;
assign w55466 = ~pi6800 & pi9040;
assign w55467 = ~pi6734 & ~pi9040;
assign w55468 = ~w55466 & ~w55467;
assign w55469 = pi2904 & ~w55468;
assign w55470 = ~pi2904 & w55468;
assign w55471 = ~w55469 & ~w55470;
assign w55472 = ~pi6801 & pi9040;
assign w55473 = ~pi6828 & ~pi9040;
assign w55474 = ~w55472 & ~w55473;
assign w55475 = pi2885 & ~w55474;
assign w55476 = ~pi2885 & w55474;
assign w55477 = ~w55475 & ~w55476;
assign w55478 = w55471 & ~w55477;
assign w55479 = ~pi6699 & pi9040;
assign w55480 = ~pi6662 & ~pi9040;
assign w55481 = ~w55479 & ~w55480;
assign w55482 = pi2879 & ~w55481;
assign w55483 = ~pi2879 & w55481;
assign w55484 = ~w55482 & ~w55483;
assign w55485 = ~pi6669 & pi9040;
assign w55486 = ~pi6800 & ~pi9040;
assign w55487 = ~w55485 & ~w55486;
assign w55488 = pi2887 & ~w55487;
assign w55489 = ~pi2887 & w55487;
assign w55490 = ~w55488 & ~w55489;
assign w55491 = ~w55484 & ~w55490;
assign w55492 = ~pi6655 & pi9040;
assign w55493 = ~pi6663 & ~pi9040;
assign w55494 = ~w55492 & ~w55493;
assign w55495 = pi2902 & ~w55494;
assign w55496 = ~pi2902 & w55494;
assign w55497 = ~w55495 & ~w55496;
assign w55498 = ~w55484 & w55497;
assign w55499 = ~w55491 & ~w55498;
assign w55500 = w55478 & ~w55499;
assign w55501 = w55484 & ~w55490;
assign w55502 = ~w55484 & w55490;
assign w55503 = ~w55501 & ~w55502;
assign w55504 = ~w55477 & w55490;
assign w55505 = w55471 & ~w55491;
assign w55506 = ~w55504 & w55505;
assign w55507 = w55503 & w55506;
assign w55508 = ~w55500 & ~w55507;
assign w55509 = ~w55471 & ~w55498;
assign w55510 = w55504 & w55509;
assign w55511 = ~w55471 & w55477;
assign w55512 = w55491 & w55511;
assign w55513 = ~w55506 & ~w55512;
assign w55514 = ~w55497 & ~w55513;
assign w55515 = ~pi6740 & pi9040;
assign w55516 = ~pi6669 & ~pi9040;
assign w55517 = ~w55515 & ~w55516;
assign w55518 = pi2888 & ~w55517;
assign w55519 = ~pi2888 & w55517;
assign w55520 = ~w55518 & ~w55519;
assign w55521 = ~w55510 & ~w55520;
assign w55522 = w55508 & w55521;
assign w55523 = ~w55514 & w55522;
assign w55524 = ~w55471 & ~w55484;
assign w55525 = w55471 & w55484;
assign w55526 = ~w55524 & ~w55525;
assign w55527 = w55490 & w55526;
assign w55528 = w55471 & w55477;
assign w55529 = w55502 & w55528;
assign w55530 = ~w55497 & ~w55529;
assign w55531 = w55527 & w55530;
assign w55532 = w55471 & w55497;
assign w55533 = ~w55501 & w55532;
assign w55534 = ~w55507 & w67091;
assign w55535 = w55477 & ~w55490;
assign w55536 = ~w55504 & ~w55535;
assign w55537 = w55524 & w55536;
assign w55538 = w55520 & ~w55537;
assign w55539 = ~w55531 & w55538;
assign w55540 = ~w55534 & w55539;
assign w55541 = w55497 & ~w55512;
assign w55542 = ~w55503 & w55511;
assign w55543 = ~w55491 & ~w55542;
assign w55544 = w55541 & ~w55543;
assign w55545 = ~w55478 & ~w55511;
assign w55546 = w55484 & ~w55497;
assign w55547 = w55545 & w55546;
assign w55548 = ~w55544 & ~w55547;
assign w55549 = (w55548 & w55523) | (w55548 & w67092) | (w55523 & w67092);
assign w55550 = pi2914 & ~w55549;
assign w55551 = ~pi2914 & w55549;
assign w55552 = ~w55550 & ~w55551;
assign w55553 = ~pi6853 & pi9040;
assign w55554 = ~pi6632 & ~pi9040;
assign w55555 = ~w55553 & ~w55554;
assign w55556 = pi2892 & ~w55555;
assign w55557 = ~pi2892 & w55555;
assign w55558 = ~w55556 & ~w55557;
assign w55559 = ~pi6731 & pi9040;
assign w55560 = ~pi6866 & ~pi9040;
assign w55561 = ~w55559 & ~w55560;
assign w55562 = pi2891 & ~w55561;
assign w55563 = ~pi2891 & w55561;
assign w55564 = ~w55562 & ~w55563;
assign w55565 = ~pi6866 & pi9040;
assign w55566 = ~pi6673 & ~pi9040;
assign w55567 = ~w55565 & ~w55566;
assign w55568 = pi2872 & ~w55567;
assign w55569 = ~pi2872 & w55567;
assign w55570 = ~w55568 & ~w55569;
assign w55571 = w55564 & ~w55570;
assign w55572 = ~pi6763 & pi9040;
assign w55573 = ~pi6664 & ~pi9040;
assign w55574 = ~w55572 & ~w55573;
assign w55575 = pi2907 & ~w55574;
assign w55576 = ~pi2907 & w55574;
assign w55577 = ~w55575 & ~w55576;
assign w55578 = w55570 & w55577;
assign w55579 = ~w55571 & ~w55578;
assign w55580 = ~pi6673 & pi9040;
assign w55581 = ~pi6738 & ~pi9040;
assign w55582 = ~w55580 & ~w55581;
assign w55583 = pi2896 & ~w55582;
assign w55584 = ~pi2896 & w55582;
assign w55585 = ~w55583 & ~w55584;
assign w55586 = ~w55564 & w55585;
assign w55587 = ~w55570 & ~w55577;
assign w55588 = ~w55578 & ~w55587;
assign w55589 = ~w55564 & w55570;
assign w55590 = ~w55571 & ~w55589;
assign w55591 = w55588 & ~w55590;
assign w55592 = w55558 & w55591;
assign w55593 = ~w55571 & w55588;
assign w55594 = ~w55592 & ~w55593;
assign w55595 = (w55585 & w55592) | (w55585 & w63333) | (w55592 & w63333);
assign w55596 = (~w55592 & w63444) | (~w55592 & w63445) | (w63444 & w63445);
assign w55597 = ~w55596 & w64119;
assign w55598 = ~w55577 & ~w55586;
assign w55599 = w55564 & ~w55585;
assign w55600 = w55558 & w55570;
assign w55601 = ~w55599 & ~w55600;
assign w55602 = ~w55598 & ~w55601;
assign w55603 = ~w55558 & w55587;
assign w55604 = ~w55602 & ~w55603;
assign w55605 = ~w55558 & w55590;
assign w55606 = w55604 & w55605;
assign w55607 = w55558 & w55577;
assign w55608 = ~w55558 & ~w55570;
assign w55609 = w55579 & ~w55608;
assign w55610 = ~w55558 & w55564;
assign w55611 = ~w55585 & ~w55610;
assign w55612 = ~w55607 & w55611;
assign w55613 = ~w55609 & w55612;
assign w55614 = ~w55606 & ~w55613;
assign w55615 = ~w55597 & w55614;
assign w55616 = ~pi6809 & pi9040;
assign w55617 = ~pi6658 & ~pi9040;
assign w55618 = ~w55616 & ~w55617;
assign w55619 = pi2897 & ~w55618;
assign w55620 = ~pi2897 & w55618;
assign w55621 = ~w55619 & ~w55620;
assign w55622 = ~w55615 & ~w55621;
assign w55623 = ~w55564 & w55588;
assign w55624 = w55564 & ~w55588;
assign w55625 = ~w55623 & ~w55624;
assign w55626 = w55558 & ~w55625;
assign w55627 = w55564 & w55577;
assign w55628 = ~w55589 & ~w55627;
assign w55629 = ~w55585 & ~w55628;
assign w55630 = ~w55625 & w64120;
assign w55631 = w55577 & ~w55585;
assign w55632 = ~w55599 & ~w55631;
assign w55633 = w55609 & w55632;
assign w55634 = ~w55586 & ~w55587;
assign w55635 = ~w55558 & ~w55590;
assign w55636 = ~w55634 & w55635;
assign w55637 = ~w55633 & ~w55636;
assign w55638 = w55577 & w55599;
assign w55639 = (w55621 & ~w55637) | (w55621 & w67093) | (~w55637 & w67093);
assign w55640 = ~w55558 & ~w55577;
assign w55641 = w55564 & w55640;
assign w55642 = w55585 & w55641;
assign w55643 = w55608 & w55631;
assign w55644 = ~w55564 & ~w55640;
assign w55645 = w55640 & w63446;
assign w55646 = ~w55644 & ~w55645;
assign w55647 = w55585 & ~w55646;
assign w55648 = w55590 & ~w55607;
assign w55649 = ~w55608 & ~w55640;
assign w55650 = w55648 & w55649;
assign w55651 = w55647 & w55650;
assign w55652 = ~w55642 & ~w55643;
assign w55653 = ~w55630 & w55652;
assign w55654 = ~w55651 & w55653;
assign w55655 = ~w55639 & w55654;
assign w55656 = ~w55622 & w55655;
assign w55657 = pi2924 & ~w55656;
assign w55658 = ~pi2924 & w55656;
assign w55659 = ~w55657 & ~w55658;
assign w55660 = ~pi6769 & pi9040;
assign w55661 = ~pi6676 & ~pi9040;
assign w55662 = ~w55660 & ~w55661;
assign w55663 = pi2882 & ~w55662;
assign w55664 = ~pi2882 & w55662;
assign w55665 = ~w55663 & ~w55664;
assign w55666 = ~pi6732 & pi9040;
assign w55667 = ~pi6684 & ~pi9040;
assign w55668 = ~w55666 & ~w55667;
assign w55669 = pi2910 & ~w55668;
assign w55670 = ~pi2910 & w55668;
assign w55671 = ~w55669 & ~w55670;
assign w55672 = ~pi6839 & pi9040;
assign w55673 = ~pi6737 & ~pi9040;
assign w55674 = ~w55672 & ~w55673;
assign w55675 = pi2888 & ~w55674;
assign w55676 = ~pi2888 & w55674;
assign w55677 = ~w55675 & ~w55676;
assign w55678 = ~w55671 & w55677;
assign w55679 = ~pi6670 & pi9040;
assign w55680 = ~pi6672 & ~pi9040;
assign w55681 = ~w55679 & ~w55680;
assign w55682 = pi2887 & ~w55681;
assign w55683 = ~pi2887 & w55681;
assign w55684 = ~w55682 & ~w55683;
assign w55685 = ~pi6806 & pi9040;
assign w55686 = ~pi6726 & ~pi9040;
assign w55687 = ~w55685 & ~w55686;
assign w55688 = pi2907 & ~w55687;
assign w55689 = ~pi2907 & w55687;
assign w55690 = ~w55688 & ~w55689;
assign w55691 = w55684 & ~w55690;
assign w55692 = w55678 & w55691;
assign w55693 = ~w55665 & w55692;
assign w55694 = ~pi6706 & pi9040;
assign w55695 = ~pi6739 & ~pi9040;
assign w55696 = ~w55694 & ~w55695;
assign w55697 = pi2891 & ~w55696;
assign w55698 = ~pi2891 & w55696;
assign w55699 = ~w55697 & ~w55698;
assign w55700 = ~w55684 & ~w55690;
assign w55701 = w55671 & w55700;
assign w55702 = w55700 & w67094;
assign w55703 = ~w55684 & w55690;
assign w55704 = ~w55677 & w55703;
assign w55705 = ~w55702 & ~w55704;
assign w55706 = w55665 & ~w55705;
assign w55707 = w55684 & w55690;
assign w55708 = w55671 & w55690;
assign w55709 = w55671 & ~w55677;
assign w55710 = ~w55678 & ~w55709;
assign w55711 = ~w55708 & ~w55710;
assign w55712 = ~w55707 & ~w55711;
assign w55713 = ~w55665 & ~w55712;
assign w55714 = w55677 & w55684;
assign w55715 = ~w55671 & ~w55690;
assign w55716 = ~w55708 & ~w55715;
assign w55717 = w55714 & ~w55716;
assign w55718 = ~w55706 & ~w55717;
assign w55719 = ~w55713 & w55718;
assign w55720 = ~w55699 & ~w55719;
assign w55721 = w55707 & w55709;
assign w55722 = ~w55702 & ~w55721;
assign w55723 = w55700 & w55710;
assign w55724 = w55684 & w55709;
assign w55725 = ~w55723 & ~w55724;
assign w55726 = w55703 & ~w55710;
assign w55727 = (~w55726 & w55725) | (~w55726 & w67095) | (w55725 & w67095);
assign w55728 = w55665 & ~w55727;
assign w55729 = ~w55678 & ~w55691;
assign w55730 = w55665 & ~w55692;
assign w55731 = ~w55729 & w55730;
assign w55732 = ~w55665 & ~w55684;
assign w55733 = w55710 & w55732;
assign w55734 = ~w55721 & ~w55733;
assign w55735 = ~w55731 & w55734;
assign w55736 = (~w55693 & w55735) | (~w55693 & w67096) | (w55735 & w67096);
assign w55737 = ~w55728 & w55736;
assign w55738 = ~w55720 & w55737;
assign w55739 = pi2912 & ~w55738;
assign w55740 = ~pi2912 & w55738;
assign w55741 = ~w55739 & ~w55740;
assign w55742 = ~w55211 & ~w55238;
assign w55743 = ~w55223 & ~w55742;
assign w55744 = ~w55171 & w55208;
assign w55745 = w55177 & w55185;
assign w55746 = ~w55170 & w55745;
assign w55747 = ~w55194 & ~w55746;
assign w55748 = ~w55179 & ~w55196;
assign w55749 = w55234 & ~w55748;
assign w55750 = ~w55207 & ~w55219;
assign w55751 = ~w55219 & w67097;
assign w55752 = ~w55749 & ~w55751;
assign w55753 = ~w55210 & w55747;
assign w55754 = w55752 & w55753;
assign w55755 = w55171 & w55745;
assign w55756 = ~w55164 & ~w55194;
assign w55757 = w55196 & w55756;
assign w55758 = ~w55755 & ~w55757;
assign w55759 = w55225 & ~w55758;
assign w55760 = w55210 & w55219;
assign w55761 = w55206 & ~w55744;
assign w55762 = ~w55760 & w55761;
assign w55763 = ~w55759 & w55762;
assign w55764 = ~w55754 & w55763;
assign w55765 = w55221 & w55233;
assign w55766 = ~w55206 & w55758;
assign w55767 = ~w55765 & w55766;
assign w55768 = w55752 & w55767;
assign w55769 = ~w55764 & ~w55768;
assign w55770 = ~w55743 & ~w55769;
assign w55771 = pi2934 & w55770;
assign w55772 = ~pi2934 & ~w55770;
assign w55773 = ~w55771 & ~w55772;
assign w55774 = w55207 & w55222;
assign w55775 = ~w55187 & ~w55774;
assign w55776 = ~w55171 & ~w55215;
assign w55777 = ~w55198 & ~w55776;
assign w55778 = ~w55197 & w55777;
assign w55779 = ~w55212 & w55775;
assign w55780 = ~w55778 & w55779;
assign w55781 = ~w55747 & ~w55755;
assign w55782 = ~w55194 & ~w55780;
assign w55783 = (~w55206 & ~w55780) | (~w55206 & w67098) | (~w55780 & w67098);
assign w55784 = ~w55782 & w55783;
assign w55785 = w55194 & ~w55777;
assign w55786 = ~w55236 & ~w55785;
assign w55787 = w55206 & ~w55213;
assign w55788 = w55758 & w55775;
assign w55789 = w55787 & w55788;
assign w55790 = ~w55786 & w55789;
assign w55791 = ~w55784 & ~w55790;
assign w55792 = pi2951 & w55791;
assign w55793 = ~pi2951 & ~w55791;
assign w55794 = ~w55792 & ~w55793;
assign w55795 = w55073 & ~w55090;
assign w55796 = ~w55080 & ~w55795;
assign w55797 = ~w55081 & ~w55796;
assign w55798 = w55071 & w55113;
assign w55799 = ~w55057 & ~w55101;
assign w55800 = ~w55075 & ~w55146;
assign w55801 = ~w55078 & ~w55800;
assign w55802 = w55092 & ~w55801;
assign w55803 = ~w55799 & w55802;
assign w55804 = ~w55147 & ~w55798;
assign w55805 = ~w55797 & w55804;
assign w55806 = ~w55803 & w55805;
assign w55807 = w55110 & ~w55806;
assign w55808 = ~w55090 & ~w55134;
assign w55809 = w55078 & w55094;
assign w55810 = w55090 & ~w55809;
assign w55811 = ~w55077 & w55810;
assign w55812 = ~w55808 & ~w55811;
assign w55813 = ~w55072 & ~w55090;
assign w55814 = ~w55081 & ~w55115;
assign w55815 = w55813 & w55814;
assign w55816 = ~w55110 & ~w55802;
assign w55817 = ~w55815 & w55816;
assign w55818 = ~w55812 & ~w55817;
assign w55819 = ~w55807 & w55818;
assign w55820 = pi2935 & ~w55819;
assign w55821 = ~pi2935 & w55819;
assign w55822 = ~w55820 & ~w55821;
assign w55823 = w55577 & ~w55637;
assign w55824 = ~w55591 & ~w55600;
assign w55825 = w55594 & ~w55824;
assign w55826 = w55611 & ~w55644;
assign w55827 = w55621 & ~w55826;
assign w55828 = ~w55647 & w55827;
assign w55829 = ~w55825 & w55828;
assign w55830 = w55585 & w55624;
assign w55831 = ~w55585 & ~w55627;
assign w55832 = w55648 & w55831;
assign w55833 = ~w55592 & ~w55621;
assign w55834 = ~w55830 & ~w55832;
assign w55835 = w55833 & w55834;
assign w55836 = (~w55823 & w55829) | (~w55823 & w67099) | (w55829 & w67099);
assign w55837 = pi2925 & w55836;
assign w55838 = ~pi2925 & ~w55836;
assign w55839 = ~w55837 & ~w55838;
assign w55840 = ~w55383 & ~w55402;
assign w55841 = ~w55390 & w55840;
assign w55842 = ~w55392 & ~w55841;
assign w55843 = ~w55410 & ~w55842;
assign w55844 = w55390 & w55423;
assign w55845 = w55423 & w64121;
assign w55846 = w55400 & ~w55840;
assign w55847 = (w55410 & w55846) | (w55410 & w64122) | (w55846 & w64122);
assign w55848 = ~w55384 & w55390;
assign w55849 = ~w55377 & ~w55425;
assign w55850 = ~w55426 & ~w55849;
assign w55851 = ~w55848 & ~w55850;
assign w55852 = ~w55850 & w64123;
assign w55853 = ~w55431 & ~w55847;
assign w55854 = ~w55852 & w55853;
assign w55855 = w55419 & ~w55843;
assign w55856 = w55854 & w55855;
assign w55857 = ~w55846 & w67100;
assign w55858 = ~w55851 & w55857;
assign w55859 = ~w55377 & ~w55401;
assign w55860 = (~w55410 & w55859) | (~w55410 & w67101) | (w55859 & w67101);
assign w55861 = w55424 & w55438;
assign w55862 = ~w55419 & ~w55861;
assign w55863 = ~w55860 & w55862;
assign w55864 = w55384 & w55447;
assign w55865 = w55402 & w55432;
assign w55866 = ~w55864 & ~w55865;
assign w55867 = (~w55856 & w67190) | (~w55856 & w67191) | (w67190 & w67191);
assign w55868 = (w55856 & w67192) | (w55856 & w67193) | (w67192 & w67193);
assign w55869 = ~w55867 & ~w55868;
assign w55870 = ~w55422 & ~w55433;
assign w55871 = ~w55399 & ~w55870;
assign w55872 = w55402 & w55455;
assign w55873 = ~w55871 & ~w55872;
assign w55874 = ~w55851 & w55873;
assign w55875 = w55419 & ~w55874;
assign w55876 = ~w55392 & ~w55420;
assign w55877 = w55425 & ~w55876;
assign w55878 = ~w55390 & ~w55423;
assign w55879 = w55412 & ~w55878;
assign w55880 = ~w55877 & ~w55879;
assign w55881 = ~w55419 & ~w55880;
assign w55882 = ~w55457 & ~w55881;
assign w55883 = ~w55875 & w55882;
assign w55884 = ~pi2916 & w55883;
assign w55885 = pi2916 & ~w55883;
assign w55886 = ~w55884 & ~w55885;
assign w55887 = (w55283 & w55267) | (w55283 & w67102) | (w55267 & w67102);
assign w55888 = ~w55309 & w55341;
assign w55889 = ~w55887 & ~w55888;
assign w55890 = ~w55301 & w55889;
assign w55891 = w55290 & ~w55890;
assign w55892 = w55303 & w55341;
assign w55893 = ~w55283 & ~w55892;
assign w55894 = w55266 & w55274;
assign w55895 = w55341 & w55894;
assign w55896 = w55283 & ~w55317;
assign w55897 = ~w55895 & w55896;
assign w55898 = ~w55893 & ~w55897;
assign w55899 = ~w55299 & w55361;
assign w55900 = w55889 & w55899;
assign w55901 = w55363 & ~w55900;
assign w55902 = ~w55290 & ~w55901;
assign w55903 = ~w55891 & ~w55898;
assign w55904 = ~w55902 & w55903;
assign w55905 = pi2950 & w55904;
assign w55906 = ~pi2950 & ~w55904;
assign w55907 = ~w55905 & ~w55906;
assign w55908 = ~w55503 & ~w55528;
assign w55909 = ~w55497 & ~w55908;
assign w55910 = w55526 & w55536;
assign w55911 = ~w55524 & w55536;
assign w55912 = ~w55908 & ~w55911;
assign w55913 = w55497 & ~w55912;
assign w55914 = w55524 & w55913;
assign w55915 = ~w55512 & ~w55520;
assign w55916 = ~w55910 & w55915;
assign w55917 = ~w55909 & w55916;
assign w55918 = ~w55914 & w55917;
assign w55919 = w55502 & w55511;
assign w55920 = ~w55497 & w55919;
assign w55921 = ~w55502 & ~w55526;
assign w55922 = w55541 & w55921;
assign w55923 = w55526 & ~w55536;
assign w55924 = w55520 & ~w55920;
assign w55925 = ~w55923 & w55924;
assign w55926 = ~w55922 & w55925;
assign w55927 = ~w55918 & ~w55926;
assign w55928 = ~pi2915 & w55927;
assign w55929 = pi2915 & ~w55927;
assign w55930 = ~w55928 & ~w55929;
assign w55931 = ~w55588 & w55831;
assign w55932 = ~w55650 & ~w55931;
assign w55933 = ~w55558 & ~w55593;
assign w55934 = w55932 & w55933;
assign w55935 = (w55621 & w55934) | (w55621 & w67103) | (w55934 & w67103);
assign w55936 = (w55621 & w55932) | (w55621 & w67104) | (w55932 & w67104);
assign w55937 = ~w55595 & w55932;
assign w55938 = ~w55936 & ~w55937;
assign w55939 = ~w55935 & ~w55938;
assign w55940 = ~pi2917 & w55939;
assign w55941 = pi2917 & ~w55939;
assign w55942 = ~w55940 & ~w55941;
assign w55943 = ~w55316 & ~w55344;
assign w55944 = w55283 & ~w55943;
assign w55945 = ~w55895 & ~w55944;
assign w55946 = (w55290 & ~w55945) | (w55290 & w67105) | (~w55945 & w67105);
assign w55947 = w55260 & w55358;
assign w55948 = ~w55253 & ~w55283;
assign w55949 = ~w55350 & ~w55359;
assign w55950 = w55274 & ~w55948;
assign w55951 = ~w55949 & w55950;
assign w55952 = ~w55342 & ~w55947;
assign w55953 = ~w55951 & w55952;
assign w55954 = w55318 & w55953;
assign w55955 = ~w55290 & ~w55954;
assign w55956 = (~w55283 & w55343) | (~w55283 & w67106) | (w55343 & w67106);
assign w55957 = ~w55336 & ~w55349;
assign w55958 = ~w55956 & w55957;
assign w55959 = ~w55946 & w55958;
assign w55960 = ~w55955 & w55959;
assign w55961 = pi2939 & ~w55960;
assign w55962 = ~pi2939 & w55960;
assign w55963 = ~w55961 & ~w55962;
assign w55964 = w55383 & ~w55436;
assign w55965 = ~w55456 & ~w55964;
assign w55966 = ~w55420 & ~w55423;
assign w55967 = w55456 & w55966;
assign w55968 = w55419 & ~w55965;
assign w55969 = ~w55967 & w55968;
assign w55970 = (w55439 & ~w55853) | (w55439 & w67107) | (~w55853 & w67107);
assign w55971 = ~w55437 & w64125;
assign w55972 = (w55410 & w55971) | (w55410 & w67108) | (w55971 & w67108);
assign w55973 = w55404 & w55422;
assign w55974 = ~w55404 & w55420;
assign w55975 = ~w55425 & w55974;
assign w55976 = ~w55973 & ~w55975;
assign w55977 = ~w55864 & w55976;
assign w55978 = (~w55419 & ~w55977) | (~w55419 & w67109) | (~w55977 & w67109);
assign w55979 = w55428 & ~w55969;
assign w55980 = ~w55978 & w55979;
assign w55981 = ~w55970 & w55980;
assign w55982 = ~pi2919 & ~w55981;
assign w55983 = pi2919 & w55981;
assign w55984 = ~w55982 & ~w55983;
assign w55985 = ~w55602 & w64126;
assign w55986 = ~w55625 & w55985;
assign w55987 = ~w55645 & ~w55651;
assign w55988 = ~w55986 & w55987;
assign w55989 = (w55621 & ~w55988) | (w55621 & w64127) | (~w55988 & w64127);
assign w55990 = w55629 & ~w55649;
assign w55991 = w55609 & w55621;
assign w55992 = w55599 & w55600;
assign w55993 = ~w55570 & w55577;
assign w55994 = w55586 & w55993;
assign w55995 = ~w55992 & ~w55994;
assign w55996 = ~w55991 & ~w55995;
assign w55997 = ~w55604 & ~w55621;
assign w55998 = ~w55642 & ~w55990;
assign w55999 = ~w55996 & w55998;
assign w56000 = ~w55997 & w55999;
assign w56001 = ~w55989 & w67110;
assign w56002 = (~pi2932 & w55989) | (~pi2932 & w67111) | (w55989 & w67111);
assign w56003 = ~w56001 & ~w56002;
assign w56004 = (~w55064 & w55809) | (~w55064 & w67112) | (w55809 & w67112);
assign w56005 = w55057 & w55119;
assign w56006 = w55800 & ~w56005;
assign w56007 = ~w56004 & w56006;
assign w56008 = ~w55147 & ~w56007;
assign w56009 = w55110 & ~w56008;
assign w56010 = ~w55096 & ~w55136;
assign w56011 = ~w55115 & ~w56010;
assign w56012 = ~w55079 & ~w55138;
assign w56013 = ~w55090 & ~w55809;
assign w56014 = ~w56012 & w56013;
assign w56015 = ~w56011 & ~w56014;
assign w56016 = ~w55074 & ~w55078;
assign w56017 = w55051 & ~w55063;
assign w56018 = w56016 & ~w56017;
assign w56019 = ~w55813 & w56018;
assign w56020 = ~w55075 & w55090;
assign w56021 = ~w56016 & ~w56020;
assign w56022 = ~w55110 & ~w56021;
assign w56023 = ~w56019 & w56022;
assign w56024 = ~w56009 & ~w56023;
assign w56025 = ~w56015 & w56024;
assign w56026 = pi2955 & w56025;
assign w56027 = ~pi2955 & ~w56025;
assign w56028 = ~w56026 & ~w56027;
assign w56029 = ~pi6664 & pi9040;
assign w56030 = ~pi6634 & ~pi9040;
assign w56031 = ~w56029 & ~w56030;
assign w56032 = pi2899 & ~w56031;
assign w56033 = ~pi2899 & w56031;
assign w56034 = ~w56032 & ~w56033;
assign w56035 = ~pi6799 & pi9040;
assign w56036 = ~pi6731 & ~pi9040;
assign w56037 = ~w56035 & ~w56036;
assign w56038 = pi2890 & ~w56037;
assign w56039 = ~pi2890 & w56037;
assign w56040 = ~w56038 & ~w56039;
assign w56041 = ~w56034 & ~w56040;
assign w56042 = ~pi6722 & pi9040;
assign w56043 = ~pi6667 & ~pi9040;
assign w56044 = ~w56042 & ~w56043;
assign w56045 = pi2895 & ~w56044;
assign w56046 = ~pi2895 & w56044;
assign w56047 = ~w56045 & ~w56046;
assign w56048 = ~pi6766 & pi9040;
assign w56049 = ~pi6987 & ~pi9040;
assign w56050 = ~w56048 & ~w56049;
assign w56051 = pi2906 & ~w56050;
assign w56052 = ~pi2906 & w56050;
assign w56053 = ~w56051 & ~w56052;
assign w56054 = w56047 & w56053;
assign w56055 = ~pi6730 & pi9040;
assign w56056 = ~pi6763 & ~pi9040;
assign w56057 = ~w56055 & ~w56056;
assign w56058 = pi2880 & ~w56057;
assign w56059 = ~pi2880 & w56057;
assign w56060 = ~w56058 & ~w56059;
assign w56061 = w56054 & w56060;
assign w56062 = w56041 & w56061;
assign w56063 = ~pi6721 & pi9040;
assign w56064 = ~pi6799 & ~pi9040;
assign w56065 = ~w56063 & ~w56064;
assign w56066 = pi2873 & ~w56065;
assign w56067 = ~pi2873 & w56065;
assign w56068 = ~w56066 & ~w56067;
assign w56069 = ~w56047 & ~w56053;
assign w56070 = w56041 & w56069;
assign w56071 = w56034 & ~w56047;
assign w56072 = w56034 & ~w56040;
assign w56073 = w56053 & w56072;
assign w56074 = ~w56034 & w56047;
assign w56075 = w56040 & w56074;
assign w56076 = ~w56073 & ~w56075;
assign w56077 = ~w56071 & w56076;
assign w56078 = w56060 & ~w56077;
assign w56079 = w56053 & w56071;
assign w56080 = ~w56070 & ~w56079;
assign w56081 = ~w56078 & w56080;
assign w56082 = w56068 & ~w56081;
assign w56083 = ~w56040 & w56068;
assign w56084 = w56034 & w56040;
assign w56085 = ~w56041 & ~w56084;
assign w56086 = ~w56083 & w56085;
assign w56087 = ~w56054 & ~w56069;
assign w56088 = ~w56073 & w56087;
assign w56089 = ~w56086 & ~w56088;
assign w56090 = w56086 & w56087;
assign w56091 = ~w56060 & ~w56089;
assign w56092 = ~w56090 & w56091;
assign w56093 = w56060 & ~w56068;
assign w56094 = ~w56041 & w56093;
assign w56095 = w56077 & w56094;
assign w56096 = ~w56062 & ~w56095;
assign w56097 = ~w56092 & w56096;
assign w56098 = ~w56082 & w56097;
assign w56099 = pi2942 & ~w56098;
assign w56100 = ~pi2942 & w56098;
assign w56101 = ~w56099 & ~w56100;
assign w56102 = w55471 & w55490;
assign w56103 = ~w55471 & ~w55490;
assign w56104 = ~w56102 & ~w56103;
assign w56105 = ~w55477 & ~w56104;
assign w56106 = ~w56104 & w67113;
assign w56107 = w55497 & ~w56106;
assign w56108 = w55484 & w55511;
assign w56109 = ~w55497 & ~w56108;
assign w56110 = ~w55484 & ~w55545;
assign w56111 = w55484 & w56103;
assign w56112 = ~w56102 & ~w56111;
assign w56113 = ~w56110 & w56112;
assign w56114 = w56109 & ~w56113;
assign w56115 = w55526 & w67114;
assign w56116 = w55525 & w55535;
assign w56117 = ~w56115 & ~w56116;
assign w56118 = (w56117 & w56114) | (w56117 & w67115) | (w56114 & w67115);
assign w56119 = w55520 & ~w56118;
assign w56120 = ~w55520 & ~w56105;
assign w56121 = w56117 & w56120;
assign w56122 = w55541 & ~w56121;
assign w56123 = ~w55512 & ~w56106;
assign w56124 = ~w55520 & ~w56123;
assign w56125 = ~w55497 & w56117;
assign w56126 = ~w56124 & w56125;
assign w56127 = ~w56122 & ~w56126;
assign w56128 = ~w56119 & ~w56127;
assign w56129 = ~pi2928 & w56128;
assign w56130 = pi2928 & ~w56128;
assign w56131 = ~w56129 & ~w56130;
assign w56132 = w56069 & ~w56072;
assign w56133 = ~w56073 & ~w56132;
assign w56134 = w56060 & w56068;
assign w56135 = ~w56133 & w56134;
assign w56136 = w56083 & w56133;
assign w56137 = ~w56071 & ~w56074;
assign w56138 = w56085 & w56137;
assign w56139 = ~w56133 & ~w56138;
assign w56140 = w56076 & ~w56139;
assign w56141 = (~w56068 & w56139) | (~w56068 & w67116) | (w56139 & w67116);
assign w56142 = w56034 & ~w56068;
assign w56143 = w56040 & w56053;
assign w56144 = ~w56047 & w56143;
assign w56145 = ~w56142 & w56144;
assign w56146 = ~w56136 & ~w56145;
assign w56147 = ~w56141 & w56146;
assign w56148 = ~w56060 & ~w56147;
assign w56149 = w56069 & w56086;
assign w56150 = ~w56068 & ~w56069;
assign w56151 = ~w56085 & w56150;
assign w56152 = ~w56149 & ~w56151;
assign w56153 = w56060 & ~w56152;
assign w56154 = ~w56053 & w56068;
assign w56155 = w56138 & w56154;
assign w56156 = ~w56134 & ~w56142;
assign w56157 = w56047 & w56143;
assign w56158 = ~w56156 & w56157;
assign w56159 = ~w56135 & ~w56158;
assign w56160 = ~w56155 & w56159;
assign w56161 = ~w56153 & w56160;
assign w56162 = ~w56148 & w56161;
assign w56163 = pi2940 & ~w56162;
assign w56164 = ~pi2940 & w56162;
assign w56165 = ~w56163 & ~w56164;
assign w56166 = w55665 & w55701;
assign w56167 = w55699 & ~w56166;
assign w56168 = ~w55677 & w55684;
assign w56169 = w55665 & w55677;
assign w56170 = ~w56168 & ~w56169;
assign w56171 = w55708 & w56170;
assign w56172 = ~w55707 & ~w55714;
assign w56173 = w55716 & ~w56172;
assign w56174 = (w55665 & w56173) | (w55665 & w67117) | (w56173 & w67117);
assign w56175 = ~w55665 & ~w55690;
assign w56176 = w56168 & w56175;
assign w56177 = ~w56171 & ~w56176;
assign w56178 = ~w56174 & w56177;
assign w56179 = ~w56167 & ~w56178;
assign w56180 = ~w55671 & ~w55684;
assign w56181 = w55690 & w56180;
assign w56182 = ~w55691 & ~w56181;
assign w56183 = w55713 & ~w56182;
assign w56184 = w55677 & ~w55684;
assign w56185 = ~w56168 & ~w56184;
assign w56186 = (~w55700 & w56185) | (~w55700 & w67118) | (w56185 & w67118);
assign w56187 = w55665 & w56186;
assign w56188 = ~w55707 & w56185;
assign w56189 = w56187 & ~w56188;
assign w56190 = (~w55707 & ~w56185) | (~w55707 & w67119) | (~w56185 & w67119);
assign w56191 = (~w55665 & ~w55714) | (~w55665 & w56175) | (~w55714 & w56175);
assign w56192 = ~w56190 & w56191;
assign w56193 = w55722 & ~w56181;
assign w56194 = ~w56192 & w56193;
assign w56195 = ~w56189 & w56194;
assign w56196 = w55699 & ~w56195;
assign w56197 = ~w56179 & ~w56183;
assign w56198 = ~w56196 & w56197;
assign w56199 = pi2933 & ~w56198;
assign w56200 = ~pi2933 & w56198;
assign w56201 = ~w56199 & ~w56200;
assign w56202 = w55179 & w55185;
assign w56203 = w55214 & ~w56202;
assign w56204 = ~w55747 & ~w56203;
assign w56205 = ~w55164 & w55215;
assign w56206 = ~w55209 & ~w56205;
assign w56207 = w55226 & w56206;
assign w56208 = ~w55206 & ~w56207;
assign w56209 = w55194 & w55750;
assign w56210 = ~w55210 & ~w55216;
assign w56211 = w55747 & ~w56210;
assign w56212 = ~w55751 & w56211;
assign w56213 = ~w55238 & ~w56209;
assign w56214 = ~w56212 & w56213;
assign w56215 = w55206 & ~w56214;
assign w56216 = ~w56204 & ~w56208;
assign w56217 = ~w56215 & w56216;
assign w56218 = ~pi2958 & w56217;
assign w56219 = pi2958 & ~w56217;
assign w56220 = ~w56218 & ~w56219;
assign w56221 = ~w56041 & ~w56143;
assign w56222 = w56041 & w56053;
assign w56223 = ~w56221 & ~w56222;
assign w56224 = w56134 & ~w56223;
assign w56225 = (~w56061 & ~w56140) | (~w56061 & w67120) | (~w56140 & w67120);
assign w56226 = ~w56084 & ~w56225;
assign w56227 = ~w56040 & ~w56047;
assign w56228 = ~w56068 & ~w56227;
assign w56229 = ~w56074 & ~w56143;
assign w56230 = w56228 & w56229;
assign w56231 = ~w56139 & ~w56230;
assign w56232 = ~w56060 & ~w56231;
assign w56233 = ~w56034 & w56054;
assign w56234 = ~w56060 & ~w56233;
assign w56235 = ~w56221 & w56228;
assign w56236 = ~w56234 & w56235;
assign w56237 = ~w56071 & ~w56234;
assign w56238 = w56068 & ~w56229;
assign w56239 = ~w56237 & w56238;
assign w56240 = ~w56236 & ~w56239;
assign w56241 = ~w56232 & w56240;
assign w56242 = ~w56226 & w56241;
assign w56243 = pi2943 & ~w56242;
assign w56244 = ~pi2943 & w56242;
assign w56245 = ~w56243 & ~w56244;
assign w56246 = ~w55678 & ~w56172;
assign w56247 = ~w56181 & ~w56246;
assign w56248 = (w55665 & w56246) | (w55665 & w67121) | (w56246 & w67121);
assign w56249 = w55716 & w56188;
assign w56250 = ~w55707 & w56169;
assign w56251 = ~w56180 & w56250;
assign w56252 = w55665 & ~w55714;
assign w56253 = w55690 & ~w55710;
assign w56254 = ~w56252 & w56253;
assign w56255 = ~w56176 & ~w56251;
assign w56256 = w55725 & w56255;
assign w56257 = ~w56254 & w56256;
assign w56258 = ~w55716 & w56191;
assign w56259 = w56256 & w64128;
assign w56260 = ~w56248 & ~w56249;
assign w56261 = (w55699 & w56259) | (w55699 & w67122) | (w56259 & w67122);
assign w56262 = ~w55671 & w56170;
assign w56263 = ~w56191 & w56262;
assign w56264 = (~w56263 & w56257) | (~w56263 & w67123) | (w56257 & w67123);
assign w56265 = ~w56261 & w56264;
assign w56266 = pi2922 & w56265;
assign w56267 = ~pi2922 & ~w56265;
assign w56268 = ~w56266 & ~w56267;
assign w56269 = w56061 & w56072;
assign w56270 = w56040 & ~w56137;
assign w56271 = ~w56034 & ~w56068;
assign w56272 = (~w56040 & w56137) | (~w56040 & w64129) | (w56137 & w64129);
assign w56273 = ~w56270 & ~w56272;
assign w56274 = ~w56228 & ~w56273;
assign w56275 = ~w56068 & ~w56138;
assign w56276 = ~w56270 & w56275;
assign w56277 = ~w56274 & ~w56276;
assign w56278 = ~w56060 & ~w56222;
assign w56279 = ~w56277 & w56278;
assign w56280 = ~w56053 & w56273;
assign w56281 = ~w56223 & w56271;
assign w56282 = ~w56280 & ~w56281;
assign w56283 = w56060 & ~w56282;
assign w56284 = ~w56047 & w56222;
assign w56285 = w56053 & w56075;
assign w56286 = ~w56284 & ~w56285;
assign w56287 = w56068 & ~w56286;
assign w56288 = ~w56068 & w56144;
assign w56289 = ~w56269 & ~w56288;
assign w56290 = ~w56287 & w56289;
assign w56291 = ~w56279 & w56290;
assign w56292 = w56291 & w67124;
assign w56293 = (~pi2927 & ~w56291) | (~pi2927 & w67125) | (~w56291 & w67125);
assign w56294 = ~w56292 & ~w56293;
assign w56295 = w55497 & ~w55919;
assign w56296 = w55504 & w55525;
assign w56297 = w56109 & ~w56296;
assign w56298 = ~w56295 & ~w56297;
assign w56299 = ~w55525 & ~w55532;
assign w56300 = ~w55912 & ~w56299;
assign w56301 = ~w55477 & ~w55484;
assign w56302 = w56104 & w56301;
assign w56303 = w55530 & ~w56302;
assign w56304 = w55503 & w56303;
assign w56305 = ~w55520 & ~w55542;
assign w56306 = ~w56300 & w56305;
assign w56307 = ~w56304 & w56306;
assign w56308 = ~w56111 & w56303;
assign w56309 = ~w55913 & ~w56308;
assign w56310 = w55520 & ~w56116;
assign w56311 = ~w56309 & w56310;
assign w56312 = ~w56307 & ~w56311;
assign w56313 = ~w56312 & w67126;
assign w56314 = (pi2931 & w56312) | (pi2931 & w67127) | (w56312 & w67127);
assign w56315 = ~w56313 & ~w56314;
assign w56316 = w55665 & ~w55715;
assign w56317 = w56184 & ~w56316;
assign w56318 = ~w56187 & ~w56317;
assign w56319 = ~w55699 & ~w56318;
assign w56320 = w55699 & w55700;
assign w56321 = ~w56181 & ~w56320;
assign w56322 = ~w55677 & ~w56321;
assign w56323 = ~w55721 & ~w56322;
assign w56324 = w55665 & ~w56323;
assign w56325 = ~w55665 & w55710;
assign w56326 = ~w56176 & ~w56325;
assign w56327 = ~w56186 & ~w56326;
assign w56328 = ~w55677 & ~w55732;
assign w56329 = ~w55724 & w56328;
assign w56330 = w55699 & ~w55700;
assign w56331 = ~w56329 & w56330;
assign w56332 = w56247 & w56331;
assign w56333 = ~w56327 & ~w56332;
assign w56334 = ~w56324 & w56333;
assign w56335 = ~w56319 & w56334;
assign w56336 = ~pi2948 & ~w56335;
assign w56337 = pi2948 & w56335;
assign w56338 = ~w56336 & ~w56337;
assign w56339 = ~pi6909 & pi9040;
assign w56340 = ~pi6864 & ~pi9040;
assign w56341 = ~w56339 & ~w56340;
assign w56342 = pi2956 & ~w56341;
assign w56343 = ~pi2956 & w56341;
assign w56344 = ~w56342 & ~w56343;
assign w56345 = ~pi7018 & pi9040;
assign w56346 = ~pi6879 & ~pi9040;
assign w56347 = ~w56345 & ~w56346;
assign w56348 = pi2970 & ~w56347;
assign w56349 = ~pi2970 & w56347;
assign w56350 = ~w56348 & ~w56349;
assign w56351 = w56344 & ~w56350;
assign w56352 = ~w56344 & w56350;
assign w56353 = ~w56351 & ~w56352;
assign w56354 = ~pi6936 & pi9040;
assign w56355 = ~pi6913 & ~pi9040;
assign w56356 = ~w56354 & ~w56355;
assign w56357 = pi2936 & ~w56356;
assign w56358 = ~pi2936 & w56356;
assign w56359 = ~w56357 & ~w56358;
assign w56360 = w56353 & w56359;
assign w56361 = ~pi6999 & pi9040;
assign w56362 = ~pi7028 & ~pi9040;
assign w56363 = ~w56361 & ~w56362;
assign w56364 = pi2953 & ~w56363;
assign w56365 = ~pi2953 & w56363;
assign w56366 = ~w56364 & ~w56365;
assign w56367 = ~w56344 & ~w56366;
assign w56368 = ~w56350 & ~w56366;
assign w56369 = w56350 & w56366;
assign w56370 = ~w56368 & ~w56369;
assign w56371 = ~w56359 & ~w56367;
assign w56372 = ~w56370 & w56371;
assign w56373 = ~w56360 & ~w56372;
assign w56374 = ~pi7080 & pi9040;
assign w56375 = ~pi6884 & ~pi9040;
assign w56376 = ~w56374 & ~w56375;
assign w56377 = pi2949 & ~w56376;
assign w56378 = ~pi2949 & w56376;
assign w56379 = ~w56377 & ~w56378;
assign w56380 = ~w56373 & ~w56379;
assign w56381 = w56350 & w56379;
assign w56382 = w56350 & ~w56359;
assign w56383 = ~w56381 & ~w56382;
assign w56384 = w56367 & ~w56383;
assign w56385 = w56359 & w56366;
assign w56386 = w56353 & w56385;
assign w56387 = ~w56384 & ~w56386;
assign w56388 = ~pi6868 & pi9040;
assign w56389 = pi6999 & ~pi9040;
assign w56390 = ~w56388 & ~w56389;
assign w56391 = pi2961 & ~w56390;
assign w56392 = ~pi2961 & w56390;
assign w56393 = ~w56391 & ~w56392;
assign w56394 = (w56393 & w56380) | (w56393 & w67128) | (w56380 & w67128);
assign w56395 = w56344 & w56359;
assign w56396 = ~w56344 & ~w56359;
assign w56397 = ~w56395 & ~w56396;
assign w56398 = w56368 & ~w56397;
assign w56399 = w56350 & ~w56366;
assign w56400 = w56395 & w56399;
assign w56401 = ~w56379 & ~w56400;
assign w56402 = w56359 & w56370;
assign w56403 = w56401 & w56402;
assign w56404 = ~w56372 & w56381;
assign w56405 = w56387 & w56404;
assign w56406 = ~w56398 & ~w56403;
assign w56407 = ~w56405 & w56406;
assign w56408 = ~w56393 & ~w56407;
assign w56409 = ~w56359 & ~w56366;
assign w56410 = w56351 & w56409;
assign w56411 = w56379 & ~w56410;
assign w56412 = ~w56385 & ~w56409;
assign w56413 = w56351 & w56412;
assign w56414 = ~w56409 & ~w56413;
assign w56415 = w56411 & ~w56414;
assign w56416 = w56366 & ~w56379;
assign w56417 = w56353 & w56416;
assign w56418 = ~w56415 & ~w56417;
assign w56419 = ~w56394 & w56418;
assign w56420 = ~w56408 & w56419;
assign w56421 = ~pi3189 & ~w56420;
assign w56422 = pi3189 & w56420;
assign w56423 = ~w56421 & ~w56422;
assign w56424 = ~pi7011 & pi9040;
assign w56425 = ~pi6889 & ~pi9040;
assign w56426 = ~w56424 & ~w56425;
assign w56427 = pi2972 & ~w56426;
assign w56428 = ~pi2972 & w56426;
assign w56429 = ~w56427 & ~w56428;
assign w56430 = ~pi6874 & pi9040;
assign w56431 = ~pi7063 & ~pi9040;
assign w56432 = ~w56430 & ~w56431;
assign w56433 = pi2969 & ~w56432;
assign w56434 = ~pi2969 & w56432;
assign w56435 = ~w56433 & ~w56434;
assign w56436 = ~w56429 & ~w56435;
assign w56437 = ~pi6989 & pi9040;
assign w56438 = ~pi6872 & ~pi9040;
assign w56439 = ~w56437 & ~w56438;
assign w56440 = pi2961 & ~w56439;
assign w56441 = ~pi2961 & w56439;
assign w56442 = ~w56440 & ~w56441;
assign w56443 = ~pi7028 & pi9040;
assign w56444 = ~pi6895 & ~pi9040;
assign w56445 = ~w56443 & ~w56444;
assign w56446 = pi2945 & ~w56445;
assign w56447 = ~pi2945 & w56445;
assign w56448 = ~w56446 & ~w56447;
assign w56449 = ~pi7020 & pi9040;
assign w56450 = ~pi6860 & ~pi9040;
assign w56451 = ~w56449 & ~w56450;
assign w56452 = pi2936 & ~w56451;
assign w56453 = ~pi2936 & w56451;
assign w56454 = ~w56452 & ~w56453;
assign w56455 = w56448 & ~w56454;
assign w56456 = ~w56429 & w56455;
assign w56457 = ~w56442 & w56456;
assign w56458 = ~w56435 & w56442;
assign w56459 = (w56448 & ~w56436) | (w56448 & w56455) | (~w56436 & w56455);
assign w56460 = w56458 & ~w56459;
assign w56461 = w56435 & ~w56442;
assign w56462 = ~w56429 & ~w56448;
assign w56463 = w56461 & w56462;
assign w56464 = ~w56460 & ~w56463;
assign w56465 = ~w56429 & w56454;
assign w56466 = w56429 & ~w56454;
assign w56467 = ~w56465 & ~w56466;
assign w56468 = ~w56448 & ~w56467;
assign w56469 = ~w56464 & w56468;
assign w56470 = ~w56457 & ~w56469;
assign w56471 = w56436 & ~w56470;
assign w56472 = ~w56458 & ~w56461;
assign w56473 = ~w56448 & ~w56454;
assign w56474 = ~pi6860 & pi9040;
assign w56475 = ~pi7018 & ~pi9040;
assign w56476 = ~w56474 & ~w56475;
assign w56477 = pi2967 & ~w56476;
assign w56478 = ~pi2967 & w56476;
assign w56479 = ~w56477 & ~w56478;
assign w56480 = w56435 & ~w56454;
assign w56481 = ~w56465 & ~w56480;
assign w56482 = w56461 & w56481;
assign w56483 = w56458 & ~w56465;
assign w56484 = ~w56458 & w56465;
assign w56485 = ~w56483 & ~w56484;
assign w56486 = w56448 & ~w56485;
assign w56487 = (w56479 & ~w56472) | (w56479 & w67129) | (~w56472 & w67129);
assign w56488 = ~w56482 & w56487;
assign w56489 = ~w56486 & w56488;
assign w56490 = ~w56442 & w56466;
assign w56491 = w56466 & w67130;
assign w56492 = w56435 & w56442;
assign w56493 = w56448 & ~w56492;
assign w56494 = ~w56462 & w56467;
assign w56495 = ~w56493 & w56494;
assign w56496 = ~w56479 & ~w56491;
assign w56497 = ~w56495 & w56496;
assign w56498 = w56464 & w56497;
assign w56499 = ~w56436 & ~w56472;
assign w56500 = w56448 & ~w56467;
assign w56501 = w56499 & w56500;
assign w56502 = (~w56501 & w56498) | (~w56501 & w67131) | (w56498 & w67131);
assign w56503 = ~w56471 & w56502;
assign w56504 = pi3191 & ~w56503;
assign w56505 = ~pi3191 & w56503;
assign w56506 = ~w56504 & ~w56505;
assign w56507 = ~pi6895 & pi9040;
assign w56508 = ~pi6922 & ~pi9040;
assign w56509 = ~w56507 & ~w56508;
assign w56510 = pi2938 & ~w56509;
assign w56511 = ~pi2938 & w56509;
assign w56512 = ~w56510 & ~w56511;
assign w56513 = ~pi7016 & pi9040;
assign w56514 = ~pi6870 & ~pi9040;
assign w56515 = ~w56513 & ~w56514;
assign w56516 = pi2962 & ~w56515;
assign w56517 = ~pi2962 & w56515;
assign w56518 = ~w56516 & ~w56517;
assign w56519 = ~pi6927 & pi9040;
assign w56520 = ~pi7013 & ~pi9040;
assign w56521 = ~w56519 & ~w56520;
assign w56522 = pi2953 & ~w56521;
assign w56523 = ~pi2953 & w56521;
assign w56524 = ~w56522 & ~w56523;
assign w56525 = w56518 & ~w56524;
assign w56526 = ~pi6870 & pi9040;
assign w56527 = ~pi7011 & ~pi9040;
assign w56528 = ~w56526 & ~w56527;
assign w56529 = pi2957 & ~w56528;
assign w56530 = ~pi2957 & w56528;
assign w56531 = ~w56529 & ~w56530;
assign w56532 = ~w56525 & ~w56531;
assign w56533 = w56512 & w56524;
assign w56534 = w56518 & w56533;
assign w56535 = w56512 & ~w56518;
assign w56536 = ~pi6913 & pi9040;
assign w56537 = ~pi6915 & ~pi9040;
assign w56538 = ~w56536 & ~w56537;
assign w56539 = pi2954 & ~w56538;
assign w56540 = ~pi2954 & w56538;
assign w56541 = ~w56539 & ~w56540;
assign w56542 = (~w56524 & w56535) | (~w56524 & w64130) | (w56535 & w64130);
assign w56543 = ~w56534 & ~w56542;
assign w56544 = w56532 & ~w56543;
assign w56545 = ~w56512 & w56544;
assign w56546 = w56518 & ~w56541;
assign w56547 = ~w56512 & ~w56546;
assign w56548 = ~w56518 & w56541;
assign w56549 = w56524 & ~w56548;
assign w56550 = ~w56548 & w64131;
assign w56551 = ~w56532 & w56547;
assign w56552 = ~w56550 & w56551;
assign w56553 = ~pi6872 & pi9040;
assign w56554 = ~pi6927 & ~pi9040;
assign w56555 = ~w56553 & ~w56554;
assign w56556 = pi2970 & ~w56555;
assign w56557 = ~pi2970 & w56555;
assign w56558 = ~w56556 & ~w56557;
assign w56559 = ~w56518 & ~w56541;
assign w56560 = w56524 & w56531;
assign w56561 = w56559 & w56560;
assign w56562 = w56512 & w56531;
assign w56563 = w56546 & w56562;
assign w56564 = ~w56512 & w56518;
assign w56565 = ~w56535 & ~w56564;
assign w56566 = ~w56531 & ~w56565;
assign w56567 = w56541 & w56566;
assign w56568 = ~w56565 & w63447;
assign w56569 = w56533 & w56546;
assign w56570 = ~w56568 & ~w56569;
assign w56571 = ~w56558 & ~w56561;
assign w56572 = ~w56563 & w56571;
assign w56573 = ~w56552 & w56572;
assign w56574 = w56573 & w67132;
assign w56575 = ~w56512 & ~w56524;
assign w56576 = ~w56533 & ~w56575;
assign w56577 = w56559 & w56576;
assign w56578 = w56570 & ~w56577;
assign w56579 = w56552 & ~w56578;
assign w56580 = w56546 & w56575;
assign w56581 = w56531 & ~w56580;
assign w56582 = w56535 & w56541;
assign w56583 = ~w56550 & ~w56582;
assign w56584 = w56581 & w56583;
assign w56585 = w56547 & ~w56548;
assign w56586 = ~w56535 & ~w56576;
assign w56587 = ~w56582 & ~w56585;
assign w56588 = (~w56531 & ~w56587) | (~w56531 & w64132) | (~w56587 & w64132);
assign w56589 = ~w56584 & ~w56588;
assign w56590 = (w56558 & w56578) | (w56558 & w64133) | (w56578 & w64133);
assign w56591 = ~w56589 & w56590;
assign w56592 = ~w56512 & w56541;
assign w56593 = w56518 & ~w56592;
assign w56594 = ~w56524 & w56548;
assign w56595 = ~w56593 & ~w56594;
assign w56596 = w56581 & w56586;
assign w56597 = ~w56595 & w56596;
assign w56598 = ~w56545 & ~w56597;
assign w56599 = (w56598 & w56591) | (w56598 & w67133) | (w56591 & w67133);
assign w56600 = pi3192 & ~w56599;
assign w56601 = ~pi3192 & w56599;
assign w56602 = ~w56600 & ~w56601;
assign w56603 = ~w56353 & ~w56366;
assign w56604 = ~w56350 & w56359;
assign w56605 = ~w56382 & ~w56604;
assign w56606 = ~w56368 & w56605;
assign w56607 = ~w56603 & ~w56606;
assign w56608 = w56351 & w56366;
assign w56609 = ~w56379 & ~w56608;
assign w56610 = ~w56607 & w56609;
assign w56611 = w56605 & w67134;
assign w56612 = w56379 & ~w56611;
assign w56613 = ~w56610 & ~w56612;
assign w56614 = w56344 & ~w56399;
assign w56615 = w56607 & w56614;
assign w56616 = (~w56400 & ~w56607) | (~w56400 & w67135) | (~w56607 & w67135);
assign w56617 = (~w56393 & w56613) | (~w56393 & w67136) | (w56613 & w67136);
assign w56618 = w56605 & ~w56614;
assign w56619 = w56393 & ~w56618;
assign w56620 = (w56411 & w56615) | (w56411 & w67137) | (w56615 & w67137);
assign w56621 = ~w56410 & ~w56611;
assign w56622 = w56393 & ~w56621;
assign w56623 = (w56401 & ~w56607) | (w56401 & w67138) | (~w56607 & w67138);
assign w56624 = ~w56622 & w56623;
assign w56625 = ~w56620 & ~w56624;
assign w56626 = ~w56617 & ~w56625;
assign w56627 = ~pi3242 & w56626;
assign w56628 = pi3242 & ~w56626;
assign w56629 = ~w56627 & ~w56628;
assign w56630 = ~pi6889 & pi9040;
assign w56631 = pi6868 & ~pi9040;
assign w56632 = ~w56630 & ~w56631;
assign w56633 = pi2962 & ~w56632;
assign w56634 = ~pi2962 & w56632;
assign w56635 = ~w56633 & ~w56634;
assign w56636 = ~pi7063 & pi9040;
assign w56637 = ~pi6878 & ~pi9040;
assign w56638 = ~w56636 & ~w56637;
assign w56639 = pi2941 & ~w56638;
assign w56640 = ~pi2941 & w56638;
assign w56641 = ~w56639 & ~w56640;
assign w56642 = ~pi6879 & pi9040;
assign w56643 = ~pi6989 & ~pi9040;
assign w56644 = ~w56642 & ~w56643;
assign w56645 = pi2975 & ~w56644;
assign w56646 = ~pi2975 & w56644;
assign w56647 = ~w56645 & ~w56646;
assign w56648 = ~pi7048 & pi9040;
assign w56649 = ~pi7080 & ~pi9040;
assign w56650 = ~w56648 & ~w56649;
assign w56651 = pi2966 & ~w56650;
assign w56652 = ~pi2966 & w56650;
assign w56653 = ~w56651 & ~w56652;
assign w56654 = ~w56647 & ~w56653;
assign w56655 = ~pi6878 & pi9040;
assign w56656 = ~pi6909 & ~pi9040;
assign w56657 = ~w56655 & ~w56656;
assign w56658 = pi2947 & ~w56657;
assign w56659 = ~pi2947 & w56657;
assign w56660 = ~w56658 & ~w56659;
assign w56661 = w56654 & w56660;
assign w56662 = ~pi6915 & pi9040;
assign w56663 = ~pi7020 & ~pi9040;
assign w56664 = ~w56662 & ~w56663;
assign w56665 = pi2954 & ~w56664;
assign w56666 = ~pi2954 & w56664;
assign w56667 = ~w56665 & ~w56666;
assign w56668 = w56653 & w56667;
assign w56669 = ~w56660 & w56668;
assign w56670 = ~w56641 & ~w56661;
assign w56671 = ~w56669 & w56670;
assign w56672 = w56660 & w56667;
assign w56673 = ~w56660 & ~w56667;
assign w56674 = ~w56672 & ~w56673;
assign w56675 = w56653 & ~w56667;
assign w56676 = w56647 & ~w56660;
assign w56677 = w56675 & w56676;
assign w56678 = ~w56674 & ~w56677;
assign w56679 = (w56641 & ~w56678) | (w56641 & w64134) | (~w56678 & w64134);
assign w56680 = ~w56653 & ~w56660;
assign w56681 = w56647 & ~w56653;
assign w56682 = ~w56667 & w56681;
assign w56683 = ~w56680 & ~w56682;
assign w56684 = w56679 & w56683;
assign w56685 = ~w56647 & w56672;
assign w56686 = w56660 & ~w56667;
assign w56687 = w56653 & w56686;
assign w56688 = w56647 & w56687;
assign w56689 = ~w56685 & ~w56688;
assign w56690 = (w56689 & w56684) | (w56689 & w67139) | (w56684 & w67139);
assign w56691 = w56635 & ~w56690;
assign w56692 = ~w56673 & ~w56681;
assign w56693 = ~w56641 & ~w56680;
assign w56694 = ~w56672 & ~w56693;
assign w56695 = ~w56692 & ~w56694;
assign w56696 = w56641 & ~w56686;
assign w56697 = (~w56647 & w56680) | (~w56647 & w67140) | (w56680 & w67140);
assign w56698 = ~w56696 & w56697;
assign w56699 = (~w56635 & w56695) | (~w56635 & w67141) | (w56695 & w67141);
assign w56700 = ~w56647 & w56653;
assign w56701 = ~w56641 & ~w56700;
assign w56702 = ~w56681 & w56701;
assign w56703 = w56701 & w67142;
assign w56704 = w56647 & w56668;
assign w56705 = ~w56661 & ~w56704;
assign w56706 = w56641 & w56705;
assign w56707 = w56654 & w56667;
assign w56708 = w56673 & w56681;
assign w56709 = ~w56688 & ~w56708;
assign w56710 = ~w56707 & w56709;
assign w56711 = w56706 & ~w56710;
assign w56712 = w56672 & w56700;
assign w56713 = ~w56703 & ~w56712;
assign w56714 = ~w56699 & w56713;
assign w56715 = ~w56711 & w56714;
assign w56716 = ~w56691 & w56715;
assign w56717 = ~pi3186 & w56716;
assign w56718 = pi3186 & ~w56716;
assign w56719 = ~w56717 & ~w56718;
assign w56720 = ~w56369 & w56397;
assign w56721 = w56373 & w56720;
assign w56722 = ~w56379 & ~w56412;
assign w56723 = ~w56344 & w56385;
assign w56724 = w56379 & ~w56723;
assign w56725 = w56604 & w56724;
assign w56726 = ~w56722 & ~w56725;
assign w56727 = w56398 & w56726;
assign w56728 = w56350 & ~w56379;
assign w56729 = ~w56369 & ~w56723;
assign w56730 = ~w56728 & ~w56729;
assign w56731 = ~w56393 & ~w56730;
assign w56732 = ~w56721 & w56731;
assign w56733 = ~w56727 & w56732;
assign w56734 = w56370 & w56396;
assign w56735 = w56344 & w56728;
assign w56736 = w56393 & ~w56400;
assign w56737 = ~w56410 & ~w56735;
assign w56738 = w56736 & w56737;
assign w56739 = ~w56734 & w56738;
assign w56740 = w56726 & w56739;
assign w56741 = ~w56733 & ~w56740;
assign w56742 = ~pi3185 & w56741;
assign w56743 = pi3185 & ~w56741;
assign w56744 = ~w56742 & ~w56743;
assign w56745 = ~pi7000 & pi9040;
assign w56746 = ~pi7073 & ~pi9040;
assign w56747 = ~w56745 & ~w56746;
assign w56748 = pi2974 & ~w56747;
assign w56749 = ~pi2974 & w56747;
assign w56750 = ~w56748 & ~w56749;
assign w56751 = ~pi6977 & pi9040;
assign w56752 = ~pi6997 & ~pi9040;
assign w56753 = ~w56751 & ~w56752;
assign w56754 = pi2972 & ~w56753;
assign w56755 = ~pi2972 & w56753;
assign w56756 = ~w56754 & ~w56755;
assign w56757 = w56750 & w56756;
assign w56758 = ~pi6995 & pi9040;
assign w56759 = ~pi7098 & ~pi9040;
assign w56760 = ~w56758 & ~w56759;
assign w56761 = pi2967 & ~w56760;
assign w56762 = ~pi2967 & w56760;
assign w56763 = ~w56761 & ~w56762;
assign w56764 = ~pi7167 & pi9040;
assign w56765 = ~pi6964 & ~pi9040;
assign w56766 = ~w56764 & ~w56765;
assign w56767 = pi2930 & ~w56766;
assign w56768 = ~pi2930 & w56766;
assign w56769 = ~w56767 & ~w56768;
assign w56770 = ~w56763 & ~w56769;
assign w56771 = ~pi7073 & pi9040;
assign w56772 = ~pi6963 & ~pi9040;
assign w56773 = ~w56771 & ~w56772;
assign w56774 = pi2968 & ~w56773;
assign w56775 = ~pi2968 & w56773;
assign w56776 = ~w56774 & ~w56775;
assign w56777 = w56750 & w56776;
assign w56778 = w56770 & w56777;
assign w56779 = w56763 & w56769;
assign w56780 = ~w56770 & ~w56779;
assign w56781 = ~w56750 & ~w56763;
assign w56782 = w56780 & ~w56781;
assign w56783 = w56756 & ~w56769;
assign w56784 = ~w56776 & ~w56783;
assign w56785 = w56782 & w56784;
assign w56786 = ~w56778 & ~w56785;
assign w56787 = w56757 & ~w56786;
assign w56788 = ~pi7098 & pi9040;
assign w56789 = ~pi6861 & ~pi9040;
assign w56790 = ~w56788 & ~w56789;
assign w56791 = pi2946 & ~w56790;
assign w56792 = ~pi2946 & w56790;
assign w56793 = ~w56791 & ~w56792;
assign w56794 = w56750 & w56763;
assign w56795 = ~w56756 & ~w56780;
assign w56796 = w56756 & w56780;
assign w56797 = ~w56795 & ~w56796;
assign w56798 = w56794 & w56797;
assign w56799 = ~w56756 & ~w56763;
assign w56800 = w56756 & w56763;
assign w56801 = ~w56799 & ~w56800;
assign w56802 = ~w56794 & ~w56801;
assign w56803 = ~w56776 & ~w56780;
assign w56804 = ~w56802 & w56803;
assign w56805 = (~w56750 & w56804) | (~w56750 & w67143) | (w56804 & w67143);
assign w56806 = w56780 & ~w56801;
assign w56807 = w56776 & w56806;
assign w56808 = ~w56798 & ~w56807;
assign w56809 = (~w56793 & ~w56808) | (~w56793 & w67144) | (~w56808 & w67144);
assign w56810 = w56763 & ~w56776;
assign w56811 = w56783 & w56810;
assign w56812 = ~w56756 & ~w56776;
assign w56813 = ~w56763 & ~w56812;
assign w56814 = ~w56756 & w56769;
assign w56815 = w56810 & w56814;
assign w56816 = ~w56813 & ~w56815;
assign w56817 = w56750 & ~w56816;
assign w56818 = ~w56750 & ~w56810;
assign w56819 = ~w56813 & w56818;
assign w56820 = w56769 & w56776;
assign w56821 = w56756 & w56820;
assign w56822 = ~w56811 & ~w56821;
assign w56823 = ~w56819 & w56822;
assign w56824 = ~w56817 & w56823;
assign w56825 = w56793 & ~w56824;
assign w56826 = ~w56787 & ~w56825;
assign w56827 = ~w56809 & w56826;
assign w56828 = pi3244 & w56827;
assign w56829 = ~pi3244 & ~w56827;
assign w56830 = ~w56828 & ~w56829;
assign w56831 = w56769 & ~w56801;
assign w56832 = w56776 & ~w56831;
assign w56833 = ~w56750 & ~w56784;
assign w56834 = ~w56832 & w56833;
assign w56835 = w56794 & w56812;
assign w56836 = ~w56816 & ~w56818;
assign w56837 = ~w56797 & w56836;
assign w56838 = ~w56769 & w56837;
assign w56839 = ~w56800 & w56818;
assign w56840 = ~w56776 & ~w56814;
assign w56841 = ~w56782 & ~w56840;
assign w56842 = w56839 & ~w56841;
assign w56843 = w56777 & w56796;
assign w56844 = ~w56793 & ~w56804;
assign w56845 = ~w56843 & w56844;
assign w56846 = ~w56842 & w56845;
assign w56847 = w56750 & w56814;
assign w56848 = ~w56769 & w56812;
assign w56849 = w56802 & ~w56848;
assign w56850 = w56793 & ~w56847;
assign w56851 = ~w56849 & w56850;
assign w56852 = w56786 & w56851;
assign w56853 = ~w56846 & ~w56852;
assign w56854 = ~w56834 & ~w56835;
assign w56855 = ~w56838 & w56854;
assign w56856 = (pi3190 & w56853) | (pi3190 & w67145) | (w56853 & w67145);
assign w56857 = ~w56853 & w67146;
assign w56858 = ~w56856 & ~w56857;
assign w56859 = ~pi7025 & pi9040;
assign w56860 = ~pi6911 & ~pi9040;
assign w56861 = ~w56859 & ~w56860;
assign w56862 = pi2973 & ~w56861;
assign w56863 = ~pi2973 & w56861;
assign w56864 = ~w56862 & ~w56863;
assign w56865 = ~pi6861 & pi9040;
assign w56866 = ~pi7134 & ~pi9040;
assign w56867 = ~w56865 & ~w56866;
assign w56868 = pi2944 & ~w56867;
assign w56869 = ~pi2944 & w56867;
assign w56870 = ~w56868 & ~w56869;
assign w56871 = ~w56864 & w56870;
assign w56872 = ~pi7022 & pi9040;
assign w56873 = ~pi6995 & ~pi9040;
assign w56874 = ~w56872 & ~w56873;
assign w56875 = pi2964 & ~w56874;
assign w56876 = ~pi2964 & w56874;
assign w56877 = ~w56875 & ~w56876;
assign w56878 = w56871 & ~w56877;
assign w56879 = ~pi7010 & pi9040;
assign w56880 = ~pi6977 & ~pi9040;
assign w56881 = ~w56879 & ~w56880;
assign w56882 = pi2947 & ~w56881;
assign w56883 = ~pi2947 & w56881;
assign w56884 = ~w56882 & ~w56883;
assign w56885 = w56871 & w67147;
assign w56886 = ~pi6964 & pi9040;
assign w56887 = ~pi7025 & ~pi9040;
assign w56888 = ~w56886 & ~w56887;
assign w56889 = pi2963 & ~w56888;
assign w56890 = ~pi2963 & w56888;
assign w56891 = ~w56889 & ~w56890;
assign w56892 = ~w56885 & w56891;
assign w56893 = ~w56864 & ~w56884;
assign w56894 = ~w56864 & w56884;
assign w56895 = ~w56870 & w56877;
assign w56896 = w56894 & w56895;
assign w56897 = ~w56893 & ~w56896;
assign w56898 = ~pi6918 & pi9040;
assign w56899 = pi6885 & ~pi9040;
assign w56900 = ~w56898 & ~w56899;
assign w56901 = pi2966 & ~w56900;
assign w56902 = ~pi2966 & w56900;
assign w56903 = ~w56901 & ~w56902;
assign w56904 = ~w56897 & w56903;
assign w56905 = ~w56891 & ~w56904;
assign w56906 = ~w56892 & ~w56905;
assign w56907 = w56870 & ~w56884;
assign w56908 = ~w56864 & ~w56907;
assign w56909 = ~w56870 & w56884;
assign w56910 = w56864 & ~w56877;
assign w56911 = w56909 & w56910;
assign w56912 = w56891 & w56911;
assign w56913 = ~w56877 & ~w56891;
assign w56914 = w56870 & w56884;
assign w56915 = ~w56870 & ~w56884;
assign w56916 = ~w56871 & ~w56915;
assign w56917 = ~w56914 & w56916;
assign w56918 = w56913 & ~w56917;
assign w56919 = ~w56912 & ~w56918;
assign w56920 = ~w56908 & ~w56919;
assign w56921 = ~w56877 & w56915;
assign w56922 = w56864 & w56921;
assign w56923 = ~w56870 & ~w56891;
assign w56924 = ~w56864 & w56923;
assign w56925 = w56877 & ~w56893;
assign w56926 = w56891 & w56914;
assign w56927 = ~w56915 & ~w56924;
assign w56928 = w56925 & ~w56926;
assign w56929 = w56927 & w56928;
assign w56930 = ~w56864 & w56915;
assign w56931 = w56864 & w56914;
assign w56932 = (w56891 & ~w56915) | (w56891 & w56946) | (~w56915 & w56946);
assign w56933 = ~w56931 & w56932;
assign w56934 = ~w56891 & ~w56894;
assign w56935 = w56877 & ~w56884;
assign w56936 = w56870 & w56935;
assign w56937 = w56934 & ~w56936;
assign w56938 = ~w56933 & ~w56937;
assign w56939 = ~w56870 & ~w56925;
assign w56940 = w56938 & w56939;
assign w56941 = ~w56903 & ~w56922;
assign w56942 = ~w56929 & w56941;
assign w56943 = ~w56940 & w56942;
assign w56944 = w56877 & ~w56909;
assign w56945 = ~w56907 & ~w56944;
assign w56946 = w56864 & w56891;
assign w56947 = ~w56945 & w56946;
assign w56948 = w56903 & ~w56911;
assign w56949 = ~w56878 & w56948;
assign w56950 = ~w56947 & w56949;
assign w56951 = ~w56943 & ~w56950;
assign w56952 = ~w56906 & ~w56920;
assign w56953 = ~w56951 & w56952;
assign w56954 = pi3237 & ~w56953;
assign w56955 = ~pi3237 & w56953;
assign w56956 = ~w56954 & ~w56955;
assign w56957 = ~w56653 & w56673;
assign w56958 = (~w56635 & ~w56705) | (~w56635 & w67148) | (~w56705 & w67148);
assign w56959 = w56686 & w56700;
assign w56960 = ~w56708 & ~w56959;
assign w56961 = ~w56958 & w56960;
assign w56962 = w56641 & ~w56961;
assign w56963 = w56674 & ~w56700;
assign w56964 = w56678 & ~w56702;
assign w56965 = ~w56963 & ~w56964;
assign w56966 = ~w56673 & ~w56682;
assign w56967 = w56706 & w56966;
assign w56968 = ~w56965 & ~w56967;
assign w56969 = w56635 & ~w56968;
assign w56970 = ~w56674 & w56700;
assign w56971 = ~w56963 & ~w56970;
assign w56972 = w56635 & ~w56681;
assign w56973 = ~w56641 & ~w56972;
assign w56974 = ~w56971 & w56973;
assign w56975 = ~w56962 & ~w56974;
assign w56976 = ~w56969 & w56975;
assign w56977 = pi3261 & ~w56976;
assign w56978 = ~pi3261 & w56976;
assign w56979 = ~w56977 & ~w56978;
assign w56980 = w56560 & w56592;
assign w56981 = w56533 & w56559;
assign w56982 = w56541 & ~w56564;
assign w56983 = w56583 & w56982;
assign w56984 = w56524 & w56564;
assign w56985 = ~w56531 & ~w56984;
assign w56986 = ~w56983 & w56985;
assign w56987 = ~w56546 & ~w56549;
assign w56988 = ~w56594 & w56987;
assign w56989 = w56987 & w64135;
assign w56990 = ~w56542 & ~w56550;
assign w56991 = w56531 & w56990;
assign w56992 = ~w56989 & ~w56991;
assign w56993 = ~w56986 & w56992;
assign w56994 = ~w56558 & ~w56981;
assign w56995 = ~w56993 & w56994;
assign w56996 = w56982 & w56991;
assign w56997 = (w56558 & w56543) | (w56558 & w67149) | (w56543 & w67149);
assign w56998 = w56578 & w56997;
assign w56999 = ~w56996 & w56998;
assign w57000 = ~w56995 & ~w56999;
assign w57001 = ~w56580 & ~w56980;
assign w57002 = ~w57000 & w67150;
assign w57003 = (~pi3193 & w57000) | (~pi3193 & w67151) | (w57000 & w67151);
assign w57004 = ~w57002 & ~w57003;
assign w57005 = ~pi7134 & pi9040;
assign w57006 = ~pi6937 & ~pi9040;
assign w57007 = ~w57005 & ~w57006;
assign w57008 = pi2946 & ~w57007;
assign w57009 = ~pi2946 & w57007;
assign w57010 = ~w57008 & ~w57009;
assign w57011 = ~pi6991 & pi9040;
assign w57012 = ~pi7010 & ~pi9040;
assign w57013 = ~w57011 & ~w57012;
assign w57014 = pi2971 & ~w57013;
assign w57015 = ~pi2971 & w57013;
assign w57016 = ~w57014 & ~w57015;
assign w57017 = ~w57010 & w57016;
assign w57018 = ~pi6885 & pi9040;
assign w57019 = ~pi6991 & ~pi9040;
assign w57020 = ~w57018 & ~w57019;
assign w57021 = pi2930 & ~w57020;
assign w57022 = ~pi2930 & w57020;
assign w57023 = ~w57021 & ~w57022;
assign w57024 = ~pi6917 & pi9040;
assign w57025 = ~pi7001 & ~pi9040;
assign w57026 = ~w57024 & ~w57025;
assign w57027 = pi2959 & ~w57026;
assign w57028 = ~pi2959 & w57026;
assign w57029 = ~w57027 & ~w57028;
assign w57030 = ~w57023 & ~w57029;
assign w57031 = w57017 & w57030;
assign w57032 = w57010 & w57016;
assign w57033 = ~pi6970 & pi9040;
assign w57034 = ~pi6897 & ~pi9040;
assign w57035 = ~w57033 & ~w57034;
assign w57036 = pi2960 & ~w57035;
assign w57037 = ~pi2960 & w57035;
assign w57038 = ~w57036 & ~w57037;
assign w57039 = w57023 & ~w57038;
assign w57040 = w57032 & w57039;
assign w57041 = ~pi7001 & pi9040;
assign w57042 = ~pi6905 & ~pi9040;
assign w57043 = ~w57041 & ~w57042;
assign w57044 = pi2952 & ~w57043;
assign w57045 = ~pi2952 & w57043;
assign w57046 = ~w57044 & ~w57045;
assign w57047 = ~w57040 & ~w57046;
assign w57048 = ~w57010 & w57038;
assign w57049 = ~w57023 & w57048;
assign w57050 = ~w57016 & ~w57038;
assign w57051 = ~w57023 & w57050;
assign w57052 = w57050 & w67152;
assign w57053 = w57010 & w57023;
assign w57054 = ~w57049 & ~w57053;
assign w57055 = ~w57052 & w57054;
assign w57056 = ~w57048 & ~w57050;
assign w57057 = w57054 & w67153;
assign w57058 = ~w57040 & w57046;
assign w57059 = ~w57057 & w57058;
assign w57060 = (~w57029 & ~w57055) | (~w57029 & w67154) | (~w57055 & w67154);
assign w57061 = ~w57059 & w57060;
assign w57062 = ~w57010 & ~w57023;
assign w57063 = w57010 & w57038;
assign w57064 = ~w57010 & ~w57038;
assign w57065 = w57023 & w57064;
assign w57066 = w57064 & w63448;
assign w57067 = (w57029 & ~w57063) | (w57029 & w67155) | (~w57063 & w67155);
assign w57068 = ~w57066 & w57067;
assign w57069 = ~w57048 & ~w57062;
assign w57070 = ~w57040 & w57069;
assign w57071 = w57068 & w57070;
assign w57072 = w57023 & w57029;
assign w57073 = ~w57023 & ~w57032;
assign w57074 = ~w57072 & ~w57073;
assign w57075 = w57063 & ~w57074;
assign w57076 = w57016 & ~w57023;
assign w57077 = w57048 & w57076;
assign w57078 = w57046 & ~w57077;
assign w57079 = ~w57075 & w57078;
assign w57080 = ~w57071 & w57079;
assign w57081 = ~w57063 & ~w57064;
assign w57082 = w57076 & ~w57081;
assign w57083 = w57029 & w57057;
assign w57084 = w57047 & ~w57082;
assign w57085 = ~w57083 & w57084;
assign w57086 = ~w57080 & ~w57085;
assign w57087 = ~w57031 & ~w57061;
assign w57088 = ~w57086 & w57087;
assign w57089 = pi3187 & ~w57088;
assign w57090 = ~pi3187 & w57088;
assign w57091 = ~w57089 & ~w57090;
assign w57092 = w56674 & w56681;
assign w57093 = w56673 & w56654;
assign w57094 = ~w56669 & ~w57093;
assign w57095 = (~w56701 & ~w57094) | (~w56701 & w67156) | (~w57094 & w67156);
assign w57096 = ~w57092 & ~w57095;
assign w57097 = w56635 & ~w57096;
assign w57098 = ~w56688 & ~w57092;
assign w57099 = w56679 & ~w57098;
assign w57100 = ~w56687 & ~w56707;
assign w57101 = w56641 & ~w57100;
assign w57102 = (~w56674 & w57101) | (~w56674 & w67157) | (w57101 & w67157);
assign w57103 = ~w56641 & ~w56707;
assign w57104 = ~w56669 & w57103;
assign w57105 = ~w56679 & ~w57104;
assign w57106 = ~w56641 & ~w56653;
assign w57107 = w56672 & w57106;
assign w57108 = ~w56661 & ~w57107;
assign w57109 = w56709 & w57108;
assign w57110 = ~w57105 & w57109;
assign w57111 = ~w56635 & ~w57110;
assign w57112 = ~w57099 & ~w57102;
assign w57113 = ~w57097 & w57112;
assign w57114 = ~w57111 & w57113;
assign w57115 = pi3241 & ~w57114;
assign w57116 = ~pi3241 & w57114;
assign w57117 = ~w57115 & ~w57116;
assign w57118 = w56369 & ~w56397;
assign w57119 = (~w56396 & ~w56370) | (~w56396 & w67158) | (~w56370 & w67158);
assign w57120 = w56381 & ~w57119;
assign w57121 = w56367 & ~w56605;
assign w57122 = w56722 & ~w57121;
assign w57123 = ~w56413 & ~w57118;
assign w57124 = ~w57122 & w57123;
assign w57125 = (w56393 & ~w57124) | (w56393 & w67159) | (~w57124 & w67159);
assign w57126 = ~w56359 & w56615;
assign w57127 = ~w56352 & w56409;
assign w57128 = w56724 & ~w57127;
assign w57129 = w56605 & w67160;
assign w57130 = w56401 & ~w57121;
assign w57131 = ~w57129 & w57130;
assign w57132 = ~w57128 & ~w57131;
assign w57133 = ~w57126 & ~w57132;
assign w57134 = ~w56393 & ~w57133;
assign w57135 = w56368 & w56395;
assign w57136 = w56379 & ~w57135;
assign w57137 = w56352 & w56385;
assign w57138 = w56609 & ~w57137;
assign w57139 = ~w57136 & ~w57138;
assign w57140 = ~w57125 & ~w57139;
assign w57141 = ~w57134 & w67161;
assign w57142 = (pi3249 & w57134) | (pi3249 & w67162) | (w57134 & w67162);
assign w57143 = ~w57141 & ~w57142;
assign w57144 = w57016 & ~w57029;
assign w57145 = ~w57062 & ~w57144;
assign w57146 = ~w57053 & ~w57145;
assign w57147 = ~w57016 & w57038;
assign w57148 = w57030 & w57147;
assign w57149 = w57023 & w57048;
assign w57150 = w57048 & w64136;
assign w57151 = ~w57066 & ~w57148;
assign w57152 = ~w57150 & w57151;
assign w57153 = w57146 & ~w57152;
assign w57154 = ~w57017 & w57072;
assign w57155 = w57053 & w57147;
assign w57156 = ~w57029 & ~w57081;
assign w57157 = w57146 & w57156;
assign w57158 = ~w57154 & ~w57155;
assign w57159 = ~w57052 & w57158;
assign w57160 = ~w57157 & w57159;
assign w57161 = w57046 & ~w57160;
assign w57162 = w57029 & ~w57032;
assign w57163 = ~w57023 & w57038;
assign w57164 = ~w57029 & w57032;
assign w57165 = ~w57162 & w57163;
assign w57166 = ~w57164 & w57165;
assign w57167 = ~w57039 & ~w57049;
assign w57168 = ~w57016 & ~w57167;
assign w57169 = ~w57163 & w57164;
assign w57170 = ~w57150 & ~w57169;
assign w57171 = ~w57166 & w57170;
assign w57172 = ~w57168 & w57171;
assign w57173 = ~w57046 & ~w57172;
assign w57174 = w57064 & w57076;
assign w57175 = ~w57053 & ~w57174;
assign w57176 = w57162 & ~w57175;
assign w57177 = ~w57153 & ~w57176;
assign w57178 = ~w57161 & w57177;
assign w57179 = ~w57173 & w57178;
assign w57180 = pi3243 & w57179;
assign w57181 = ~pi3243 & ~w57179;
assign w57182 = ~w57180 & ~w57181;
assign w57183 = w56757 & w56770;
assign w57184 = ~w56750 & w56806;
assign w57185 = ~w57183 & ~w57184;
assign w57186 = ~w56776 & ~w57185;
assign w57187 = ~w56750 & w56800;
assign w57188 = ~w56821 & ~w57187;
assign w57189 = ~w56848 & ~w57183;
assign w57190 = w57188 & w57189;
assign w57191 = ~w56793 & ~w57190;
assign w57192 = w56793 & ~w56800;
assign w57193 = ~w56781 & ~w56794;
assign w57194 = w56820 & w57193;
assign w57195 = ~w57192 & w57194;
assign w57196 = w56797 & w56839;
assign w57197 = w56794 & w56807;
assign w57198 = ~w56837 & ~w57196;
assign w57199 = (w56793 & ~w57198) | (w56793 & w67163) | (~w57198 & w67163);
assign w57200 = ~w56835 & ~w57195;
assign w57201 = ~w57191 & w57200;
assign w57202 = ~w57186 & w57201;
assign w57203 = ~w57199 & w57202;
assign w57204 = pi3260 & w57203;
assign w57205 = ~pi3260 & ~w57203;
assign w57206 = ~w57204 & ~w57205;
assign w57207 = w56776 & w56797;
assign w57208 = ~w56783 & ~w56800;
assign w57209 = ~w56750 & ~w56814;
assign w57210 = w57208 & w57209;
assign w57211 = w56756 & ~w56810;
assign w57212 = ~w56780 & ~w56812;
assign w57213 = ~w57211 & w57212;
assign w57214 = ~w57210 & ~w57213;
assign w57215 = ~w57188 & ~w57214;
assign w57216 = w56750 & w56840;
assign w57217 = w57208 & w57216;
assign w57218 = w56793 & ~w56811;
assign w57219 = ~w57217 & w57218;
assign w57220 = ~w57207 & w57219;
assign w57221 = ~w57215 & w57220;
assign w57222 = ~w56793 & ~w56847;
assign w57223 = ~w57183 & w57222;
assign w57224 = ~w57197 & w57223;
assign w57225 = w57214 & w57224;
assign w57226 = ~w57221 & ~w57225;
assign w57227 = ~pi3245 & w57226;
assign w57228 = pi3245 & ~w57226;
assign w57229 = ~w57227 & ~w57228;
assign w57230 = (~w56676 & ~w57103) | (~w56676 & w67164) | (~w57103 & w67164);
assign w57231 = ~w56675 & ~w57230;
assign w57232 = ~w57101 & ~w57231;
assign w57233 = ~w56635 & ~w57232;
assign w57234 = ~w56686 & ~w56700;
assign w57235 = w56641 & ~w56675;
assign w57236 = ~w57234 & w57235;
assign w57237 = ~w56677 & ~w57107;
assign w57238 = ~w56712 & w57237;
assign w57239 = (w56635 & ~w57238) | (w56635 & w67165) | (~w57238 & w67165);
assign w57240 = ~w56700 & ~w57094;
assign w57241 = ~w56959 & ~w57240;
assign w57242 = ~w56641 & ~w57241;
assign w57243 = ~w56692 & w56696;
assign w57244 = ~w56971 & w57243;
assign w57245 = ~w57239 & ~w57244;
assign w57246 = ~w57242 & w57245;
assign w57247 = ~w57233 & w57246;
assign w57248 = pi3328 & w57247;
assign w57249 = ~pi3328 & ~w57247;
assign w57250 = ~w57248 & ~w57249;
assign w57251 = ~w56531 & ~w56550;
assign w57252 = w56547 & w57251;
assign w57253 = ~w56576 & w56982;
assign w57254 = w56531 & w56564;
assign w57255 = w56564 & w56560;
assign w57256 = ~w57253 & ~w57255;
assign w57257 = ~w57252 & w57256;
assign w57258 = w56558 & ~w57257;
assign w57259 = ~w56575 & w56990;
assign w57260 = ~w56531 & w56565;
assign w57261 = ~w57259 & w57260;
assign w57262 = w56565 & ~w56575;
assign w57263 = ~w56581 & ~w57262;
assign w57264 = ~w56988 & w57263;
assign w57265 = ~w57253 & w67166;
assign w57266 = w56991 & w57265;
assign w57267 = ~w57264 & ~w57266;
assign w57268 = ~w56558 & ~w57267;
assign w57269 = ~w56989 & ~w57261;
assign w57270 = ~w57258 & w57269;
assign w57271 = ~w57268 & w57270;
assign w57272 = pi3236 & w57271;
assign w57273 = ~pi3236 & ~w57271;
assign w57274 = ~w57272 & ~w57273;
assign w57275 = ~w57029 & ~w57149;
assign w57276 = w57152 & ~w57275;
assign w57277 = ~w57065 & ~w57077;
assign w57278 = ~w57052 & w57277;
assign w57279 = (~w57046 & w57276) | (~w57046 & w64137) | (w57276 & w64137);
assign w57280 = ~w57040 & ~w57155;
assign w57281 = w57016 & w57038;
assign w57282 = ~w57051 & ~w57281;
assign w57283 = w57068 & ~w57282;
assign w57284 = w57030 & w57056;
assign w57285 = w57152 & ~w57284;
assign w57286 = (w57046 & ~w57285) | (w57046 & w67167) | (~w57285 & w67167);
assign w57287 = ~w57279 & w57280;
assign w57288 = w57278 & w57280;
assign w57289 = w57029 & ~w57046;
assign w57290 = ~w57288 & w57289;
assign w57291 = (~w57290 & ~w57287) | (~w57290 & w67168) | (~w57287 & w67168);
assign w57292 = pi3262 & w57291;
assign w57293 = ~pi3262 & ~w57291;
assign w57294 = ~w57292 & ~w57293;
assign w57295 = ~w56582 & ~w57254;
assign w57296 = w56595 & ~w57295;
assign w57297 = ~w56524 & w56592;
assign w57298 = ~w56561 & ~w57297;
assign w57299 = ~w56577 & w57298;
assign w57300 = ~w57296 & w57299;
assign w57301 = w56558 & ~w57300;
assign w57302 = ~w56595 & ~w57251;
assign w57303 = w56987 & w67169;
assign w57304 = ~w57302 & ~w57303;
assign w57305 = ~w56558 & ~w57304;
assign w57306 = w56546 & ~w57302;
assign w57307 = (w57306 & w56993) | (w57306 & w67170) | (w56993 & w67170);
assign w57308 = ~w56579 & ~w57301;
assign w57309 = ~w57305 & w57308;
assign w57310 = w57309 & w67171;
assign w57311 = (pi3231 & ~w57309) | (pi3231 & w67172) | (~w57309 & w67172);
assign w57312 = ~w57310 & ~w57311;
assign w57313 = ~w56877 & ~w56884;
assign w57314 = w56864 & ~w56870;
assign w57315 = ~w56871 & ~w57314;
assign w57316 = w57313 & w57315;
assign w57317 = w56871 & w56935;
assign w57318 = w56891 & ~w57317;
assign w57319 = ~w57316 & w57318;
assign w57320 = ~w56891 & ~w56911;
assign w57321 = ~w57319 & ~w57320;
assign w57322 = w56924 & w56935;
assign w57323 = w56933 & w57315;
assign w57324 = w56913 & ~w57315;
assign w57325 = w56877 & w56931;
assign w57326 = ~w56903 & ~w57325;
assign w57327 = ~w56911 & ~w57322;
assign w57328 = ~w57324 & w57327;
assign w57329 = w57328 & w67173;
assign w57330 = ~w56884 & w57314;
assign w57331 = w57314 & w56935;
assign w57332 = ~w56877 & w56930;
assign w57333 = w56903 & ~w57331;
assign w57334 = ~w57332 & w57333;
assign w57335 = w56895 & w56946;
assign w57336 = ~w56885 & ~w57335;
assign w57337 = ~w56938 & w57336;
assign w57338 = w57334 & w57337;
assign w57339 = ~w57329 & ~w57338;
assign w57340 = ~w57321 & ~w57339;
assign w57341 = ~pi3173 & w57340;
assign w57342 = pi3173 & ~w57340;
assign w57343 = ~w57341 & ~w57342;
assign w57344 = w56435 & w56456;
assign w57345 = ~w56435 & w56466;
assign w57346 = ~w56442 & w56454;
assign w57347 = ~w56429 & ~w57346;
assign w57348 = (w56448 & ~w56481) | (w56448 & w64138) | (~w56481 & w64138);
assign w57349 = w56461 & w56465;
assign w57350 = ~w56435 & ~w56442;
assign w57351 = w56467 & w57350;
assign w57352 = ~w57349 & ~w57351;
assign w57353 = w56454 & w57348;
assign w57354 = w57352 & w57353;
assign w57355 = ~w57347 & w57354;
assign w57356 = w56442 & w56465;
assign w57357 = ~w56442 & w56481;
assign w57358 = ~w57356 & ~w57357;
assign w57359 = ~w57348 & ~w57358;
assign w57360 = ~w56429 & ~w56454;
assign w57361 = w56492 & w57360;
assign w57362 = w56479 & ~w57345;
assign w57363 = ~w57361 & w57362;
assign w57364 = ~w57359 & w57363;
assign w57365 = ~w57355 & w57364;
assign w57366 = ~w56435 & w56454;
assign w57367 = ~w57347 & ~w57366;
assign w57368 = w56459 & ~w57367;
assign w57369 = w56442 & ~w56448;
assign w57370 = w56429 & w57369;
assign w57371 = ~w56490 & ~w57370;
assign w57372 = w56435 & ~w57371;
assign w57373 = w56462 & w57346;
assign w57374 = ~w56479 & ~w57373;
assign w57375 = ~w57368 & w57374;
assign w57376 = ~w57372 & w57375;
assign w57377 = ~w56469 & ~w57344;
assign w57378 = (w57377 & w57365) | (w57377 & w67174) | (w57365 & w67174);
assign w57379 = pi3323 & ~w57378;
assign w57380 = ~pi3323 & w57378;
assign w57381 = ~w57379 & ~w57380;
assign w57382 = ~pi6867 & pi9040;
assign w57383 = ~pi6970 & ~pi9040;
assign w57384 = ~w57382 & ~w57383;
assign w57385 = pi2952 & ~w57384;
assign w57386 = ~pi2952 & w57384;
assign w57387 = ~w57385 & ~w57386;
assign w57388 = ~pi6905 & pi9040;
assign w57389 = ~pi6867 & ~pi9040;
assign w57390 = ~w57388 & ~w57389;
assign w57391 = pi2973 & ~w57390;
assign w57392 = ~pi2973 & w57390;
assign w57393 = ~w57391 & ~w57392;
assign w57394 = ~w57387 & ~w57393;
assign w57395 = ~pi6971 & pi9040;
assign w57396 = ~pi6917 & ~pi9040;
assign w57397 = ~w57395 & ~w57396;
assign w57398 = pi2960 & ~w57397;
assign w57399 = ~pi2960 & w57397;
assign w57400 = ~w57398 & ~w57399;
assign w57401 = ~pi6998 & pi9040;
assign w57402 = ~pi7022 & ~pi9040;
assign w57403 = ~w57401 & ~w57402;
assign w57404 = pi2965 & ~w57403;
assign w57405 = ~pi2965 & w57403;
assign w57406 = ~w57404 & ~w57405;
assign w57407 = w57400 & w57406;
assign w57408 = ~pi6963 & pi9040;
assign w57409 = pi6918 & ~pi9040;
assign w57410 = ~w57408 & ~w57409;
assign w57411 = pi2944 & ~w57410;
assign w57412 = ~pi2944 & w57410;
assign w57413 = ~w57411 & ~w57412;
assign w57414 = w57407 & w57413;
assign w57415 = w57394 & w57414;
assign w57416 = ~w57400 & ~w57406;
assign w57417 = ~w57407 & ~w57416;
assign w57418 = ~pi6997 & pi9040;
assign w57419 = ~pi6971 & ~pi9040;
assign w57420 = ~w57418 & ~w57419;
assign w57421 = pi2937 & ~w57420;
assign w57422 = ~pi2937 & w57420;
assign w57423 = ~w57421 & ~w57422;
assign w57424 = ~w57387 & w57423;
assign w57425 = w57387 & w57393;
assign w57426 = ~w57394 & ~w57425;
assign w57427 = ~w57424 & w57426;
assign w57428 = ~w57393 & w57400;
assign w57429 = ~w57387 & w57406;
assign w57430 = ~w57428 & ~w57429;
assign w57431 = ~w57394 & ~w57430;
assign w57432 = ~w57427 & ~w57431;
assign w57433 = w57417 & ~w57432;
assign w57434 = ~w57417 & ~w57427;
assign w57435 = ~w57413 & ~w57434;
assign w57436 = ~w57433 & w57435;
assign w57437 = w57393 & ~w57400;
assign w57438 = ~w57431 & ~w57437;
assign w57439 = w57413 & w57423;
assign w57440 = ~w57438 & w57439;
assign w57441 = w57413 & ~w57423;
assign w57442 = ~w57387 & ~w57400;
assign w57443 = ~w57437 & ~w57442;
assign w57444 = w57430 & w57441;
assign w57445 = w57443 & w57444;
assign w57446 = ~w57393 & w57406;
assign w57447 = w57393 & ~w57406;
assign w57448 = ~w57446 & ~w57447;
assign w57449 = w57423 & ~w57443;
assign w57450 = w57448 & w57449;
assign w57451 = ~w57415 & ~w57445;
assign w57452 = ~w57450 & w57451;
assign w57453 = ~w57440 & w57452;
assign w57454 = ~w57436 & w57453;
assign w57455 = ~pi3264 & w57454;
assign w57456 = pi3264 & ~w57454;
assign w57457 = ~w57455 & ~w57456;
assign w57458 = w57416 & ~w57426;
assign w57459 = ~w57431 & ~w57458;
assign w57460 = ~w57423 & ~w57459;
assign w57461 = w57387 & w57406;
assign w57462 = ~w57400 & w57461;
assign w57463 = ~w57424 & ~w57462;
assign w57464 = ~w57394 & w57423;
assign w57465 = ~w57407 & ~w57429;
assign w57466 = w57464 & ~w57465;
assign w57467 = w57426 & w64139;
assign w57468 = ~w57416 & w57423;
assign w57469 = ~w57426 & ~w57468;
assign w57470 = (w57469 & w57459) | (w57469 & w63449) | (w57459 & w63449);
assign w57471 = ~w57466 & ~w57467;
assign w57472 = ~w57470 & w57471;
assign w57473 = ~w57470 & w64140;
assign w57474 = (~w57413 & w57473) | (~w57413 & w67175) | (w57473 & w67175);
assign w57475 = w57413 & ~w57472;
assign w57476 = w57387 & ~w57393;
assign w57477 = ~w57446 & ~w57476;
assign w57478 = w57387 & w57400;
assign w57479 = w57393 & ~w57442;
assign w57480 = ~w57478 & w57479;
assign w57481 = ~w57423 & w57477;
assign w57482 = ~w57480 & w57481;
assign w57483 = w57461 & w57482;
assign w57484 = ~w57387 & ~w57448;
assign w57485 = ~w57467 & ~w57484;
assign w57486 = ~w57442 & w57464;
assign w57487 = ~w57485 & w57486;
assign w57488 = ~w57483 & ~w57487;
assign w57489 = ~w57475 & w57488;
assign w57490 = (pi3331 & ~w57489) | (pi3331 & w67176) | (~w57489 & w67176);
assign w57491 = w57489 & w67177;
assign w57492 = ~w57490 & ~w57491;
assign w57493 = w56458 & w56495;
assign w57494 = w56455 & w57350;
assign w57495 = w56466 & w56492;
assign w57496 = ~w56436 & ~w57495;
assign w57497 = w57369 & ~w57496;
assign w57498 = ~w56442 & w57345;
assign w57499 = ~w56429 & ~w56492;
assign w57500 = w56448 & ~w57499;
assign w57501 = ~w56480 & ~w57366;
assign w57502 = ~w57346 & ~w57501;
assign w57503 = w57500 & ~w57502;
assign w57504 = w56442 & ~w56454;
assign w57505 = w56435 & ~w57504;
assign w57506 = w57347 & w57505;
assign w57507 = w56479 & ~w57498;
assign w57508 = ~w57506 & w57507;
assign w57509 = ~w57497 & ~w57503;
assign w57510 = w57508 & w57509;
assign w57511 = w56472 & w57360;
assign w57512 = ~w56455 & ~w57360;
assign w57513 = w56499 & w57512;
assign w57514 = w56442 & w56448;
assign w57515 = ~w56481 & w57514;
assign w57516 = w57374 & ~w57511;
assign w57517 = ~w57515 & w57516;
assign w57518 = ~w57513 & w57517;
assign w57519 = ~w57510 & ~w57518;
assign w57520 = ~w57493 & ~w57494;
assign w57521 = ~w57519 & w57520;
assign w57522 = pi3271 & w57521;
assign w57523 = ~pi3271 & ~w57521;
assign w57524 = ~w57522 & ~w57523;
assign w57525 = w56907 & w56910;
assign w57526 = w56891 & w57525;
assign w57527 = w56923 & w56893;
assign w57528 = w56871 & w56892;
assign w57529 = w56913 & w56914;
assign w57530 = ~w56877 & ~w56923;
assign w57531 = w56916 & w57530;
assign w57532 = ~w57527 & ~w57529;
assign w57533 = ~w57531 & w57532;
assign w57534 = w57334 & w57533;
assign w57535 = ~w57528 & w57534;
assign w57536 = w56907 & ~w56910;
assign w57537 = w57320 & ~w57536;
assign w57538 = w56892 & ~w57330;
assign w57539 = ~w57537 & ~w57538;
assign w57540 = ~w56896 & w57326;
assign w57541 = ~w57539 & w57540;
assign w57542 = ~w57535 & ~w57541;
assign w57543 = ~w56896 & ~w57325;
assign w57544 = ~w57332 & w57543;
assign w57545 = ~w56891 & ~w57544;
assign w57546 = ~w57335 & ~w57526;
assign w57547 = ~w57545 & w57546;
assign w57548 = ~w57542 & w57547;
assign w57549 = pi3247 & ~w57548;
assign w57550 = ~pi3247 & w57548;
assign w57551 = ~w57549 & ~w57550;
assign w57552 = (~w56923 & ~w56934) | (~w56923 & w67178) | (~w56934 & w67178);
assign w57553 = w56864 & ~w56944;
assign w57554 = ~w57552 & w57553;
assign w57555 = w56935 & w57315;
assign w57556 = ~w56896 & ~w56903;
assign w57557 = ~w57555 & w57556;
assign w57558 = ~w57554 & w57557;
assign w57559 = ~w56921 & w57318;
assign w57560 = w57552 & ~w57559;
assign w57561 = w56948 & ~w57525;
assign w57562 = ~w57325 & w57561;
assign w57563 = ~w57560 & w57562;
assign w57564 = ~w56878 & ~w56894;
assign w57565 = ~w56903 & ~w57564;
assign w57566 = ~w57331 & w57543;
assign w57567 = ~w57565 & w57566;
assign w57568 = w56891 & ~w57567;
assign w57569 = ~w56891 & w57555;
assign w57570 = (~w57569 & w57563) | (~w57569 & w67179) | (w57563 & w67179);
assign w57571 = ~w57568 & w57570;
assign w57572 = ~pi3248 & w57571;
assign w57573 = pi3248 & ~w57571;
assign w57574 = ~w57572 & ~w57573;
assign w57575 = w57429 & w57479;
assign w57576 = w57424 & w57428;
assign w57577 = (~w57428 & ~w57479) | (~w57428 & w64141) | (~w57479 & w64141);
assign w57578 = (~w57576 & ~w57577) | (~w57576 & w67180) | (~w57577 & w67180);
assign w57579 = ~w57406 & ~w57578;
assign w57580 = ~w57423 & ~w57461;
assign w57581 = ~w57477 & w57580;
assign w57582 = ~w57575 & ~w57581;
assign w57583 = ~w57579 & w57582;
assign w57584 = w57413 & ~w57583;
assign w57585 = ~w57423 & w57462;
assign w57586 = w57394 & w57416;
assign w57587 = ~w57482 & ~w57586;
assign w57588 = w57423 & w57446;
assign w57589 = w57578 & w57588;
assign w57590 = (w57587 & w67181) | (w57587 & w67182) | (w67181 & w67182);
assign w57591 = ~w57589 & w57590;
assign w57592 = ~w57584 & w57591;
assign w57593 = ~pi3350 & w57592;
assign w57594 = pi3350 & ~w57592;
assign w57595 = ~w57593 & ~w57594;
assign w57596 = w57502 & w57512;
assign w57597 = ~w57349 & ~w57495;
assign w57598 = ~w56457 & w57597;
assign w57599 = ~w57596 & w57598;
assign w57600 = w56479 & ~w57599;
assign w57601 = w57348 & ~w57498;
assign w57602 = w56435 & w57504;
assign w57603 = ~w56448 & ~w57602;
assign w57604 = w57352 & w57603;
assign w57605 = ~w57601 & ~w57604;
assign w57606 = ~w57500 & w57504;
assign w57607 = ~w56491 & ~w57606;
assign w57608 = ~w57354 & w57607;
assign w57609 = ~w56479 & ~w57608;
assign w57610 = ~w57600 & ~w57605;
assign w57611 = ~w57609 & w57610;
assign w57612 = pi3349 & w57611;
assign w57613 = ~pi3349 & ~w57611;
assign w57614 = ~w57612 & ~w57613;
assign w57615 = w57414 & ~w57425;
assign w57616 = w57406 & w57428;
assign w57617 = ~w57413 & ~w57616;
assign w57618 = ~w57428 & ~w57461;
assign w57619 = ~w57423 & ~w57442;
assign w57620 = w57618 & w57619;
assign w57621 = (~w57620 & w57459) | (~w57620 & w67183) | (w57459 & w67183);
assign w57622 = w57617 & ~w57621;
assign w57623 = ~w57437 & ~w57617;
assign w57624 = w57423 & ~w57623;
assign w57625 = w57387 & ~w57406;
assign w57626 = w57441 & ~w57625;
assign w57627 = ~w57624 & ~w57626;
assign w57628 = ~w57618 & ~w57627;
assign w57629 = w57439 & ~w57485;
assign w57630 = ~w57423 & w57616;
assign w57631 = ~w57615 & ~w57630;
assign w57632 = ~w57629 & w57631;
assign w57633 = ~w57622 & w57632;
assign w57634 = ~w57628 & w57633;
assign w57635 = pi3329 & ~w57634;
assign w57636 = ~pi3329 & w57634;
assign w57637 = ~w57635 & ~w57636;
assign w57638 = ~w57068 & ~w57275;
assign w57639 = w57029 & ~w57167;
assign w57640 = w57010 & ~w57029;
assign w57641 = ~w57039 & w57640;
assign w57642 = ~w57281 & w57641;
assign w57643 = ~w57174 & ~w57642;
assign w57644 = ~w57639 & w57643;
assign w57645 = w57046 & ~w57644;
assign w57646 = ~w57076 & w57146;
assign w57647 = ~w57072 & ~w57076;
assign w57648 = w57063 & ~w57647;
assign w57649 = ~w57040 & ~w57051;
assign w57650 = ~w57648 & w57649;
assign w57651 = ~w57646 & w57650;
assign w57652 = ~w57046 & ~w57651;
assign w57653 = ~w57638 & ~w57645;
assign w57654 = ~w57652 & w57653;
assign w57655 = ~pi3273 & w57654;
assign w57656 = pi3273 & ~w57654;
assign w57657 = ~w57655 & ~w57656;
assign w57658 = ~pi7135 & pi9040;
assign w57659 = ~pi7117 & ~pi9040;
assign w57660 = ~w57658 & ~w57659;
assign w57661 = pi3267 & ~w57660;
assign w57662 = ~pi3267 & w57660;
assign w57663 = ~w57661 & ~w57662;
assign w57664 = ~pi7177 & pi9040;
assign w57665 = ~pi7143 & ~pi9040;
assign w57666 = ~w57664 & ~w57665;
assign w57667 = pi3325 & ~w57666;
assign w57668 = ~pi3325 & w57666;
assign w57669 = ~w57667 & ~w57668;
assign w57670 = w57663 & w57669;
assign w57671 = ~pi7153 & pi9040;
assign w57672 = ~pi7156 & ~pi9040;
assign w57673 = ~w57671 & ~w57672;
assign w57674 = pi3403 & ~w57673;
assign w57675 = ~pi3403 & w57673;
assign w57676 = ~w57674 & ~w57675;
assign w57677 = w57669 & w57676;
assign w57678 = ~pi7248 & pi9040;
assign w57679 = ~pi7148 & ~pi9040;
assign w57680 = ~w57678 & ~w57679;
assign w57681 = pi3272 & ~w57680;
assign w57682 = ~pi3272 & w57680;
assign w57683 = ~w57681 & ~w57682;
assign w57684 = ~w57677 & ~w57683;
assign w57685 = w57670 & w57684;
assign w57686 = ~w57663 & w57683;
assign w57687 = ~w57669 & w57676;
assign w57688 = w57686 & w57687;
assign w57689 = ~w57685 & ~w57688;
assign w57690 = ~w57663 & ~w57683;
assign w57691 = ~w57669 & ~w57676;
assign w57692 = w57686 & ~w57691;
assign w57693 = w57663 & ~w57683;
assign w57694 = ~w57669 & ~w57683;
assign w57695 = ~w57693 & ~w57694;
assign w57696 = ~w57692 & w57695;
assign w57697 = w57663 & w57676;
assign w57698 = ~w57663 & ~w57676;
assign w57699 = ~w57697 & ~w57698;
assign w57700 = ~w57688 & w57699;
assign w57701 = ~w57696 & ~w57700;
assign w57702 = w57684 & w57695;
assign w57703 = (~w57702 & w57701) | (~w57702 & w64143) | (w57701 & w64143);
assign w57704 = (w57689 & ~w57703) | (w57689 & w67184) | (~w57703 & w67184);
assign w57705 = ~pi7141 & pi9040;
assign w57706 = ~pi7150 & ~pi9040;
assign w57707 = ~w57705 & ~w57706;
assign w57708 = pi3269 & ~w57707;
assign w57709 = ~pi3269 & w57707;
assign w57710 = ~w57708 & ~w57709;
assign w57711 = ~w57704 & w57710;
assign w57712 = ~pi7117 & pi9040;
assign w57713 = ~pi7294 & ~pi9040;
assign w57714 = ~w57712 & ~w57713;
assign w57715 = pi3347 & ~w57714;
assign w57716 = ~pi3347 & w57714;
assign w57717 = ~w57715 & ~w57716;
assign w57718 = ~w57663 & ~w57710;
assign w57719 = w57687 & w57718;
assign w57720 = w57669 & w57683;
assign w57721 = ~w57697 & w57710;
assign w57722 = w57720 & ~w57721;
assign w57723 = w57663 & ~w57676;
assign w57724 = ~w57669 & w57683;
assign w57725 = w57663 & w57724;
assign w57726 = (w57710 & ~w57724) | (w57710 & w64144) | (~w57724 & w64144);
assign w57727 = w57723 & ~w57726;
assign w57728 = ~w57669 & ~w57697;
assign w57729 = ~w57683 & w57710;
assign w57730 = ~w57670 & w57729;
assign w57731 = ~w57728 & w57730;
assign w57732 = ~w57719 & ~w57722;
assign w57733 = w57732 & w64145;
assign w57734 = ~w57717 & ~w57733;
assign w57735 = w57676 & ~w57683;
assign w57736 = w57670 & w57735;
assign w57737 = ~w57727 & ~w57736;
assign w57738 = w57676 & w57686;
assign w57739 = ~w57724 & ~w57735;
assign w57740 = w57663 & w57710;
assign w57741 = ~w57739 & w57740;
assign w57742 = w57683 & w57723;
assign w57743 = w57710 & ~w57742;
assign w57744 = w57718 & w57724;
assign w57745 = w57669 & ~w57686;
assign w57746 = w57699 & w57745;
assign w57747 = ~w57744 & ~w57746;
assign w57748 = ~w57743 & ~w57747;
assign w57749 = w57694 & ~w57699;
assign w57750 = ~w57738 & ~w57741;
assign w57751 = ~w57749 & w57750;
assign w57752 = ~w57748 & w57751;
assign w57753 = ~w57737 & w57752;
assign w57754 = w57752 & w64146;
assign w57755 = ~w57669 & w57710;
assign w57756 = w57683 & w57755;
assign w57757 = ~w57723 & ~w57756;
assign w57758 = ~w57727 & ~w57757;
assign w57759 = ~w57683 & ~w57710;
assign w57760 = ~w57699 & w57759;
assign w57761 = w57677 & w57686;
assign w57762 = ~w57760 & ~w57761;
assign w57763 = ~w57758 & w57762;
assign w57764 = w57717 & ~w57763;
assign w57765 = ~w57734 & ~w57764;
assign w57766 = ~w57754 & w57765;
assign w57767 = w57766 & w67185;
assign w57768 = (~pi3762 & ~w57766) | (~pi3762 & w67186) | (~w57766 & w67186);
assign w57769 = ~w57767 & ~w57768;
assign w57770 = ~pi7136 & pi9040;
assign w57771 = ~pi7161 & ~pi9040;
assign w57772 = ~w57770 & ~w57771;
assign w57773 = pi3270 & ~w57772;
assign w57774 = ~pi3270 & w57772;
assign w57775 = ~w57773 & ~w57774;
assign w57776 = ~pi7137 & pi9040;
assign w57777 = ~pi7232 & ~pi9040;
assign w57778 = ~w57776 & ~w57777;
assign w57779 = pi3268 & ~w57778;
assign w57780 = ~pi3268 & w57778;
assign w57781 = ~w57779 & ~w57780;
assign w57782 = w57775 & ~w57781;
assign w57783 = ~pi7294 & pi9040;
assign w57784 = ~pi7137 & ~pi9040;
assign w57785 = ~w57783 & ~w57784;
assign w57786 = pi3357 & ~w57785;
assign w57787 = ~pi3357 & w57785;
assign w57788 = ~w57786 & ~w57787;
assign w57789 = ~w57782 & w57788;
assign w57790 = ~pi7146 & pi9040;
assign w57791 = ~pi7142 & ~pi9040;
assign w57792 = ~w57790 & ~w57791;
assign w57793 = pi3310 & ~w57792;
assign w57794 = ~pi3310 & w57792;
assign w57795 = ~w57793 & ~w57794;
assign w57796 = w57775 & w57795;
assign w57797 = ~w57789 & ~w57796;
assign w57798 = ~w57775 & w57788;
assign w57799 = ~w57796 & ~w57798;
assign w57800 = w57781 & ~w57799;
assign w57801 = ~w57797 & ~w57800;
assign w57802 = ~pi7101 & pi9040;
assign w57803 = ~pi7285 & ~pi9040;
assign w57804 = ~w57802 & ~w57803;
assign w57805 = pi3348 & ~w57804;
assign w57806 = ~pi3348 & w57804;
assign w57807 = ~w57805 & ~w57806;
assign w57808 = ~w57801 & ~w57807;
assign w57809 = ~w57781 & w57788;
assign w57810 = ~w57775 & ~w57795;
assign w57811 = ~w57809 & w57810;
assign w57812 = ~w57796 & ~w57811;
assign w57813 = w57808 & ~w57812;
assign w57814 = ~w57781 & ~w57795;
assign w57815 = ~w57807 & w57814;
assign w57816 = w57775 & w57788;
assign w57817 = w57795 & ~w57816;
assign w57818 = ~w57775 & w57781;
assign w57819 = ~w57782 & ~w57818;
assign w57820 = w57817 & w57819;
assign w57821 = (w57775 & w57820) | (w57775 & w63450) | (w57820 & w63450);
assign w57822 = ~w57775 & ~w57788;
assign w57823 = w57781 & w57795;
assign w57824 = ~w57814 & ~w57823;
assign w57825 = w57822 & w57824;
assign w57826 = ~w57788 & w57796;
assign w57827 = ~w57795 & w57816;
assign w57828 = ~w57826 & ~w57827;
assign w57829 = w57775 & w57828;
assign w57830 = (w57807 & w57825) | (w57807 & w63451) | (w57825 & w63451);
assign w57831 = ~w57829 & w57830;
assign w57832 = w57789 & w57831;
assign w57833 = ~w57821 & ~w57825;
assign w57834 = ~w57832 & w57833;
assign w57835 = ~pi7156 & pi9040;
assign w57836 = ~pi7164 & ~pi9040;
assign w57837 = ~w57835 & ~w57836;
assign w57838 = pi3404 & ~w57837;
assign w57839 = ~pi3404 & w57837;
assign w57840 = ~w57838 & ~w57839;
assign w57841 = (w57840 & ~w57834) | (w57840 & w64147) | (~w57834 & w64147);
assign w57842 = w57795 & w57807;
assign w57843 = w57809 & w57842;
assign w57844 = w57822 & w57823;
assign w57845 = ~w57808 & ~w57831;
assign w57846 = w57775 & ~w57809;
assign w57847 = w57814 & w57846;
assign w57848 = ~w57843 & ~w57847;
assign w57849 = (~w57845 & w64149) | (~w57845 & w64150) | (w64149 & w64150);
assign w57850 = ~w57841 & w64151;
assign w57851 = (pi3763 & w57841) | (pi3763 & w64152) | (w57841 & w64152);
assign w57852 = ~w57850 & ~w57851;
assign w57853 = w57788 & ~w57807;
assign w57854 = ~w57819 & w57853;
assign w57855 = w57822 & w57842;
assign w57856 = w57788 & w57814;
assign w57857 = ~w57855 & ~w57856;
assign w57858 = ~w57821 & w57857;
assign w57859 = (~w57798 & w57821) | (~w57798 & w64153) | (w57821 & w64153);
assign w57860 = ~w57854 & ~w57859;
assign w57861 = ~w57840 & ~w57860;
assign w57862 = (~w57781 & ~w57817) | (~w57781 & w63452) | (~w57817 & w63452);
assign w57863 = ~w57800 & ~w57862;
assign w57864 = ~w57807 & w57863;
assign w57865 = ~w57795 & w57822;
assign w57866 = w57807 & ~w57865;
assign w57867 = ~w57863 & w57866;
assign w57868 = w57858 & w57867;
assign w57869 = (w57840 & w57868) | (w57840 & w64154) | (w57868 & w64154);
assign w57870 = w57807 & ~w57840;
assign w57871 = ~w57816 & w57870;
assign w57872 = (~w57871 & w57863) | (~w57871 & w63453) | (w57863 & w63453);
assign w57873 = w57819 & ~w57872;
assign w57874 = ~w57795 & w57798;
assign w57875 = ~w57846 & ~w57874;
assign w57876 = w57815 & w57875;
assign w57877 = ~w57873 & ~w57876;
assign w57878 = ~w57861 & w57877;
assign w57879 = w57878 & w63454;
assign w57880 = (pi3783 & ~w57878) | (pi3783 & w63455) | (~w57878 & w63455);
assign w57881 = ~w57879 & ~w57880;
assign w57882 = ~pi7164 & pi9040;
assign w57883 = ~pi7159 & ~pi9040;
assign w57884 = ~w57882 & ~w57883;
assign w57885 = pi3404 & ~w57884;
assign w57886 = ~pi3404 & w57884;
assign w57887 = ~w57885 & ~w57886;
assign w57888 = ~pi7250 & pi9040;
assign w57889 = ~pi7153 & ~pi9040;
assign w57890 = ~w57888 & ~w57889;
assign w57891 = pi3309 & ~w57890;
assign w57892 = ~pi3309 & w57890;
assign w57893 = ~w57891 & ~w57892;
assign w57894 = ~w57887 & ~w57893;
assign w57895 = w57887 & w57893;
assign w57896 = ~w57894 & ~w57895;
assign w57897 = ~pi7285 & pi9040;
assign w57898 = ~pi7250 & ~pi9040;
assign w57899 = ~w57897 & ~w57898;
assign w57900 = pi3358 & ~w57899;
assign w57901 = ~pi3358 & w57899;
assign w57902 = ~w57900 & ~w57901;
assign w57903 = ~pi7148 & pi9040;
assign w57904 = ~pi7141 & ~pi9040;
assign w57905 = ~w57903 & ~w57904;
assign w57906 = pi3272 & ~w57905;
assign w57907 = ~pi3272 & w57905;
assign w57908 = ~w57906 & ~w57907;
assign w57909 = ~w57902 & w57908;
assign w57910 = ~pi7158 & pi9040;
assign w57911 = ~pi7177 & ~pi9040;
assign w57912 = ~w57910 & ~w57911;
assign w57913 = pi3310 & ~w57912;
assign w57914 = ~pi3310 & w57912;
assign w57915 = ~w57913 & ~w57914;
assign w57916 = w57908 & w57915;
assign w57917 = ~w57909 & ~w57916;
assign w57918 = ~pi7232 & pi9040;
assign w57919 = ~pi7101 & ~pi9040;
assign w57920 = ~w57918 & ~w57919;
assign w57921 = pi3267 & ~w57920;
assign w57922 = ~pi3267 & w57920;
assign w57923 = ~w57921 & ~w57922;
assign w57924 = ~w57917 & ~w57923;
assign w57925 = ~w57902 & w57915;
assign w57926 = ~w57924 & ~w57925;
assign w57927 = ~w57896 & ~w57926;
assign w57928 = ~w57887 & ~w57915;
assign w57929 = w57893 & ~w57908;
assign w57930 = w57928 & w57929;
assign w57931 = w57902 & ~w57930;
assign w57932 = ~w57908 & ~w57915;
assign w57933 = ~w57887 & w57893;
assign w57934 = ~w57916 & ~w57932;
assign w57935 = w57933 & w57934;
assign w57936 = ~w57932 & ~w57935;
assign w57937 = w57931 & ~w57936;
assign w57938 = w57908 & w57928;
assign w57939 = w57928 & w64155;
assign w57940 = w57894 & w57932;
assign w57941 = ~w57939 & ~w57940;
assign w57942 = w57887 & w57902;
assign w57943 = w57893 & ~w57915;
assign w57944 = ~w57893 & w57916;
assign w57945 = ~w57943 & ~w57944;
assign w57946 = w57942 & ~w57945;
assign w57947 = ~w57893 & ~w57915;
assign w57948 = w57887 & w57947;
assign w57949 = ~w57887 & ~w57908;
assign w57950 = w57887 & w57908;
assign w57951 = ~w57949 & ~w57950;
assign w57952 = w57915 & w57951;
assign w57953 = ~w57948 & ~w57952;
assign w57954 = w57909 & ~w57953;
assign w57955 = w57923 & w57941;
assign w57956 = ~w57946 & w57955;
assign w57957 = ~w57954 & w57956;
assign w57958 = ~w57909 & w57948;
assign w57959 = ~w57908 & w57915;
assign w57960 = w57887 & w57959;
assign w57961 = ~w57930 & ~w57960;
assign w57962 = ~w57902 & ~w57961;
assign w57963 = ~w57923 & ~w57958;
assign w57964 = ~w57962 & w57963;
assign w57965 = ~w57957 & ~w57964;
assign w57966 = ~w57927 & ~w57937;
assign w57967 = ~w57965 & w57966;
assign w57968 = pi3710 & ~w57967;
assign w57969 = ~pi3710 & w57967;
assign w57970 = ~w57968 & ~w57969;
assign w57971 = ~w57807 & ~w57828;
assign w57972 = ~w57855 & ~w57971;
assign w57973 = ~w57781 & ~w57972;
assign w57974 = w57807 & ~w57875;
assign w57975 = w57816 & w57823;
assign w57976 = w57795 & w57798;
assign w57977 = ~w57865 & ~w57976;
assign w57978 = ~w57807 & ~w57977;
assign w57979 = ~w57840 & ~w57975;
assign w57980 = ~w57974 & w57979;
assign w57981 = ~w57978 & w57980;
assign w57982 = w57807 & ~w57809;
assign w57983 = w57775 & ~w57853;
assign w57984 = ~w57982 & w57983;
assign w57985 = w57798 & w57823;
assign w57986 = w57840 & ~w57985;
assign w57987 = ~w57825 & w57986;
assign w57988 = w57857 & ~w57984;
assign w57989 = w57987 & w57988;
assign w57990 = ~w57981 & ~w57989;
assign w57991 = ~w57973 & ~w57990;
assign w57992 = pi3781 & w57991;
assign w57993 = ~pi3781 & ~w57991;
assign w57994 = ~w57992 & ~w57993;
assign w57995 = w57943 & w57950;
assign w57996 = ~w57923 & ~w57995;
assign w57997 = ~w57887 & w57959;
assign w57998 = ~w57893 & w57997;
assign w57999 = w57902 & ~w57938;
assign w58000 = w57951 & w63456;
assign w58001 = ~w57902 & ~w57995;
assign w58002 = ~w58000 & w58001;
assign w58003 = (~w57999 & ~w58002) | (~w57999 & w64156) | (~w58002 & w64156);
assign w58004 = ~w57933 & ~w57948;
assign w58005 = ~w57934 & ~w58004;
assign w58006 = w57996 & ~w57998;
assign w58007 = ~w58005 & w58006;
assign w58008 = ~w58003 & w58007;
assign w58009 = w57947 & w57950;
assign w58010 = ~w57941 & ~w58003;
assign w58011 = w57929 & w57961;
assign w58012 = ~w57894 & ~w57942;
assign w58013 = w57915 & ~w57949;
assign w58014 = ~w58012 & w58013;
assign w58015 = w57923 & ~w58009;
assign w58016 = ~w58014 & w58015;
assign w58017 = ~w58011 & w58016;
assign w58018 = ~w58010 & w58017;
assign w58019 = ~w58008 & ~w58018;
assign w58020 = ~pi3761 & w58019;
assign w58021 = pi3761 & ~w58019;
assign w58022 = ~w58020 & ~w58021;
assign w58023 = ~pi7169 & pi9040;
assign w58024 = ~pi7292 & ~pi9040;
assign w58025 = ~w58023 & ~w58024;
assign w58026 = pi3347 & ~w58025;
assign w58027 = ~pi3347 & w58025;
assign w58028 = ~w58026 & ~w58027;
assign w58029 = ~pi7157 & pi9040;
assign w58030 = ~pi7233 & ~pi9040;
assign w58031 = ~w58029 & ~w58030;
assign w58032 = pi3332 & ~w58031;
assign w58033 = ~pi3332 & w58031;
assign w58034 = ~w58032 & ~w58033;
assign w58035 = ~w58028 & ~w58034;
assign w58036 = ~pi7272 & pi9040;
assign w58037 = ~pi7147 & ~pi9040;
assign w58038 = ~w58036 & ~w58037;
assign w58039 = pi3266 & ~w58038;
assign w58040 = ~pi3266 & w58038;
assign w58041 = ~w58039 & ~w58040;
assign w58042 = ~pi7218 & pi9040;
assign w58043 = ~pi7224 & ~pi9040;
assign w58044 = ~w58042 & ~w58043;
assign w58045 = pi3325 & ~w58044;
assign w58046 = ~pi3325 & w58044;
assign w58047 = ~w58045 & ~w58046;
assign w58048 = w58041 & ~w58047;
assign w58049 = w58035 & ~w58048;
assign w58050 = ~w58041 & w58047;
assign w58051 = w58034 & w58041;
assign w58052 = ~w58050 & ~w58051;
assign w58053 = ~w58048 & ~w58050;
assign w58054 = w58028 & w58053;
assign w58055 = ~w58028 & ~w58053;
assign w58056 = ~w58054 & ~w58055;
assign w58057 = w58034 & ~w58056;
assign w58058 = (~w58049 & w58056) | (~w58049 & w63335) | (w58056 & w63335);
assign w58059 = ~pi7118 & pi9040;
assign w58060 = ~pi7235 & ~pi9040;
assign w58061 = ~w58059 & ~w58060;
assign w58062 = pi3405 & ~w58061;
assign w58063 = ~pi3405 & w58061;
assign w58064 = ~w58062 & ~w58063;
assign w58065 = ~w58058 & ~w58064;
assign w58066 = ~w58034 & ~w58041;
assign w58067 = ~w58028 & w58064;
assign w58068 = ~w58066 & w58067;
assign w58069 = w58053 & w58068;
assign w58070 = ~w58035 & ~w58069;
assign w58071 = w58028 & w58047;
assign w58072 = w58052 & ~w58071;
assign w58073 = w58028 & w58064;
assign w58074 = ~w58034 & ~w58047;
assign w58075 = w58034 & w58047;
assign w58076 = ~w58074 & ~w58075;
assign w58077 = ~w58035 & w58076;
assign w58078 = (w58050 & ~w58076) | (w58050 & w63457) | (~w58076 & w63457);
assign w58079 = w58073 & w58078;
assign w58080 = w58028 & w58041;
assign w58081 = ~w58034 & w58064;
assign w58082 = ~w58074 & ~w58081;
assign w58083 = w58080 & ~w58082;
assign w58084 = (~w58083 & w58070) | (~w58083 & w63336) | (w58070 & w63336);
assign w58085 = ~w58079 & w58084;
assign w58086 = ~w58065 & w58085;
assign w58087 = ~pi7293 & pi9040;
assign w58088 = ~pi7155 & ~pi9040;
assign w58089 = ~w58087 & ~w58088;
assign w58090 = pi3324 & ~w58089;
assign w58091 = ~pi3324 & w58089;
assign w58092 = ~w58090 & ~w58091;
assign w58093 = ~w58086 & ~w58092;
assign w58094 = ~w58047 & w58069;
assign w58095 = w58051 & ~w58056;
assign w58096 = w58047 & w58066;
assign w58097 = (~w58096 & w58056) | (~w58096 & w63458) | (w58056 & w63458);
assign w58098 = ~w58064 & ~w58097;
assign w58099 = w58073 & w58074;
assign w58100 = ~w58047 & ~w58064;
assign w58101 = w58028 & ~w58064;
assign w58102 = ~w58048 & ~w58101;
assign w58103 = ~w58100 & ~w58102;
assign w58104 = ~w58051 & w58068;
assign w58105 = ~w58047 & ~w58080;
assign w58106 = ~w58103 & ~w58104;
assign w58107 = (w58106 & ~w58058) | (w58106 & w64157) | (~w58058 & w64157);
assign w58108 = w58092 & ~w58107;
assign w58109 = ~w58094 & ~w58099;
assign w58110 = ~w58098 & w58109;
assign w58111 = ~w58093 & w58110;
assign w58112 = w58111 & w63459;
assign w58113 = (pi3759 & ~w58111) | (pi3759 & w63460) | (~w58111 & w63460);
assign w58114 = ~w58112 & ~w58113;
assign w58115 = w57789 & ~w57824;
assign w58116 = ~w57807 & w57819;
assign w58117 = ~w57775 & w58116;
assign w58118 = w57782 & w57842;
assign w58119 = w57840 & ~w58118;
assign w58120 = ~w58115 & w58119;
assign w58121 = ~w57876 & w58120;
assign w58122 = ~w58117 & w58121;
assign w58123 = w57782 & w57795;
assign w58124 = ~w57844 & ~w57874;
assign w58125 = (~w57807 & ~w58124) | (~w57807 & w64158) | (~w58124 & w64158);
assign w58126 = ~w57840 & ~w57847;
assign w58127 = ~w58125 & w58126;
assign w58128 = ~w58122 & ~w58127;
assign w58129 = ~w57820 & ~w57827;
assign w58130 = w57870 & ~w58129;
assign w58131 = w58116 & w58129;
assign w58132 = ~w57820 & w57982;
assign w58133 = (w58132 & w57832) | (w58132 & w64159) | (w57832 & w64159);
assign w58134 = ~w58130 & ~w58131;
assign w58135 = ~w58128 & w58134;
assign w58136 = w58135 & w64160;
assign w58137 = (~pi3778 & ~w58135) | (~pi3778 & w64161) | (~w58135 & w64161);
assign w58138 = ~w58136 & ~w58137;
assign w58139 = w58047 & w58104;
assign w58140 = w58053 & w58073;
assign w58141 = ~w58028 & ~w58041;
assign w58142 = ~w58080 & ~w58141;
assign w58143 = ~w58053 & w58142;
assign w58144 = w58034 & w58143;
assign w58145 = ~w58092 & ~w58140;
assign w58146 = ~w58144 & w58145;
assign w58147 = w58035 & w58100;
assign w58148 = w58066 & w58071;
assign w58149 = w58092 & ~w58148;
assign w58150 = ~w58067 & ~w58101;
assign w58151 = ~w58072 & ~w58150;
assign w58152 = w58074 & w58080;
assign w58153 = ~w58069 & ~w58152;
assign w58154 = ~w58151 & w58153;
assign w58155 = w58064 & ~w58154;
assign w58156 = w58041 & w58047;
assign w58157 = ~w58101 & ~w58156;
assign w58158 = w58034 & ~w58157;
assign w58159 = ~w58147 & w58149;
assign w58160 = ~w58158 & w58159;
assign w58161 = (~w58146 & w58155) | (~w58146 & w64162) | (w58155 & w64162);
assign w58162 = w58047 & ~w58066;
assign w58163 = ~w58064 & ~w58092;
assign w58164 = ~w58142 & w58163;
assign w58165 = ~w58162 & w58164;
assign w58166 = ~w58139 & ~w58165;
assign w58167 = ~w58161 & w58166;
assign w58168 = pi3776 & w58167;
assign w58169 = ~pi3776 & ~w58167;
assign w58170 = ~w58168 & ~w58169;
assign w58171 = ~w57663 & w57739;
assign w58172 = (~w57710 & w58171) | (~w57710 & w64163) | (w58171 & w64163);
assign w58173 = w57684 & ~w57728;
assign w58174 = w57683 & ~w57692;
assign w58175 = w57726 & w58174;
assign w58176 = ~w57761 & ~w58173;
assign w58177 = ~w58175 & w58176;
assign w58178 = (w57717 & ~w58177) | (w57717 & w64164) | (~w58177 & w64164);
assign w58179 = w57717 & ~w57735;
assign w58180 = ~w57676 & ~w57694;
assign w58181 = ~w57720 & w58180;
assign w58182 = ~w57677 & w57710;
assign w58183 = ~w57738 & w58182;
assign w58184 = ~w58179 & w58183;
assign w58185 = ~w58181 & w58184;
assign w58186 = ~w57689 & w57748;
assign w58187 = w57676 & ~w57740;
assign w58188 = w57745 & w58187;
assign w58189 = (~w57717 & w58188) | (~w57717 & w64165) | (w58188 & w64165);
assign w58190 = ~w58185 & ~w58189;
assign w58191 = ~w58186 & w58190;
assign w58192 = ~w58178 & w58191;
assign w58193 = (pi3849 & ~w58192) | (pi3849 & w64166) | (~w58192 & w64166);
assign w58194 = w58192 & w64167;
assign w58195 = ~w58193 & ~w58194;
assign w58196 = ~pi7154 & pi9040;
assign w58197 = ~pi7246 & ~pi9040;
assign w58198 = ~w58196 & ~w58197;
assign w58199 = pi3326 & ~w58198;
assign w58200 = ~pi3326 & w58198;
assign w58201 = ~w58199 & ~w58200;
assign w58202 = ~pi7159 & pi9040;
assign w58203 = ~pi7165 & ~pi9040;
assign w58204 = ~w58202 & ~w58203;
assign w58205 = pi3357 & ~w58204;
assign w58206 = ~pi3357 & w58204;
assign w58207 = ~w58205 & ~w58206;
assign w58208 = w58201 & ~w58207;
assign w58209 = ~pi7142 & pi9040;
assign w58210 = ~pi7248 & ~pi9040;
assign w58211 = ~w58209 & ~w58210;
assign w58212 = pi3360 & ~w58211;
assign w58213 = ~pi3360 & w58211;
assign w58214 = ~w58212 & ~w58213;
assign w58215 = w58208 & w58214;
assign w58216 = ~pi7161 & pi9040;
assign w58217 = ~pi7154 & ~pi9040;
assign w58218 = ~w58216 & ~w58217;
assign w58219 = pi3422 & ~w58218;
assign w58220 = ~pi3422 & w58218;
assign w58221 = ~w58219 & ~w58220;
assign w58222 = w58207 & ~w58221;
assign w58223 = w58201 & ~w58214;
assign w58224 = ~w58201 & w58214;
assign w58225 = ~w58223 & ~w58224;
assign w58226 = w58222 & ~w58225;
assign w58227 = ~w58215 & ~w58226;
assign w58228 = ~pi7144 & pi9040;
assign w58229 = ~pi7146 & ~pi9040;
assign w58230 = ~w58228 & ~w58229;
assign w58231 = pi3314 & ~w58230;
assign w58232 = ~pi3314 & w58230;
assign w58233 = ~w58231 & ~w58232;
assign w58234 = ~w58227 & w58233;
assign w58235 = ~pi7150 & pi9040;
assign w58236 = ~pi7136 & ~pi9040;
assign w58237 = ~w58235 & ~w58236;
assign w58238 = pi3270 & ~w58237;
assign w58239 = ~pi3270 & w58237;
assign w58240 = ~w58238 & ~w58239;
assign w58241 = ~w58221 & w58223;
assign w58242 = w58207 & w58221;
assign w58243 = ~w58201 & w58242;
assign w58244 = (~w58233 & ~w58242) | (~w58233 & w64168) | (~w58242 & w64168);
assign w58245 = w58207 & ~w58214;
assign w58246 = ~w58221 & w58245;
assign w58247 = w58244 & ~w58246;
assign w58248 = ~w58207 & w58221;
assign w58249 = ~w58222 & ~w58248;
assign w58250 = ~w58201 & ~w58214;
assign w58251 = ~w58201 & ~w58221;
assign w58252 = ~w58250 & ~w58251;
assign w58253 = ~w58249 & w58252;
assign w58254 = ~w58243 & ~w58253;
assign w58255 = ~w58253 & w63461;
assign w58256 = (~w58247 & w58255) | (~w58247 & w64169) | (w58255 & w64169);
assign w58257 = w58214 & ~w58221;
assign w58258 = ~w58201 & ~w58207;
assign w58259 = w58257 & w58258;
assign w58260 = w58208 & w63462;
assign w58261 = ~w58259 & ~w58260;
assign w58262 = ~w58233 & ~w58251;
assign w58263 = w58222 & w58262;
assign w58264 = ~w58241 & ~w58263;
assign w58265 = w58261 & w58264;
assign w58266 = ~w58256 & w58265;
assign w58267 = ~w58240 & ~w58266;
assign w58268 = (w58257 & w58226) | (w58257 & w64170) | (w58226 & w64170);
assign w58269 = ~w58245 & ~w58248;
assign w58270 = w58250 & w58269;
assign w58271 = ~w58243 & ~w58270;
assign w58272 = (w58233 & w58270) | (w58233 & w64171) | (w58270 & w64171);
assign w58273 = ~w58268 & ~w58272;
assign w58274 = w58240 & ~w58273;
assign w58275 = w58224 & w58248;
assign w58276 = ~w58214 & w58221;
assign w58277 = w58240 & w58276;
assign w58278 = ~w58275 & ~w58277;
assign w58279 = ~w58233 & ~w58278;
assign w58280 = ~w58234 & ~w58279;
assign w58281 = ~w58274 & w58280;
assign w58282 = ~w58267 & w58281;
assign w58283 = ~pi3800 & w58282;
assign w58284 = pi3800 & ~w58282;
assign w58285 = ~w58283 & ~w58284;
assign w58286 = ~w58214 & ~w58233;
assign w58287 = w58251 & w58286;
assign w58288 = w58201 & w58233;
assign w58289 = ~w58263 & ~w58288;
assign w58290 = w58207 & w58223;
assign w58291 = w58233 & ~w58241;
assign w58292 = w58254 & w58291;
assign w58293 = ~w58241 & ~w58243;
assign w58294 = ~w58233 & ~w58293;
assign w58295 = ~w58260 & ~w58290;
assign w58296 = ~w58294 & w58295;
assign w58297 = ~w58292 & w58296;
assign w58298 = ~w58257 & ~w58258;
assign w58299 = w58262 & ~w58298;
assign w58300 = ~w58287 & ~w58299;
assign w58301 = (w58297 & w64172) | (w58297 & w64173) | (w64172 & w64173);
assign w58302 = w58221 & w58290;
assign w58303 = w58240 & ~w58297;
assign w58304 = ~w58246 & w58261;
assign w58305 = w58291 & ~w58304;
assign w58306 = w58224 & w58262;
assign w58307 = ~w58302 & ~w58306;
assign w58308 = ~w58305 & w58307;
assign w58309 = ~w58303 & w58308;
assign w58310 = w58309 & w64174;
assign w58311 = (pi3843 & ~w58309) | (pi3843 & w64175) | (~w58309 & w64175);
assign w58312 = ~w58310 & ~w58311;
assign w58313 = w57722 & w57723;
assign w58314 = (w57717 & w57753) | (w57717 & w63464) | (w57753 & w63464);
assign w58315 = ~w57717 & ~w57752;
assign w58316 = w57698 & w57729;
assign w58317 = ~w57728 & w58179;
assign w58318 = w57743 & w58317;
assign w58319 = ~w58313 & ~w58316;
assign w58320 = ~w58318 & w58319;
assign w58321 = ~w58315 & w58320;
assign w58322 = ~w58314 & w58321;
assign w58323 = pi3809 & ~w58322;
assign w58324 = ~pi3809 & w58322;
assign w58325 = ~w58323 & ~w58324;
assign w58326 = ~pi7229 & pi9040;
assign w58327 = ~pi7138 & ~pi9040;
assign w58328 = ~w58326 & ~w58327;
assign w58329 = pi3326 & ~w58328;
assign w58330 = ~pi3326 & w58328;
assign w58331 = ~w58329 & ~w58330;
assign w58332 = ~pi7145 & pi9040;
assign w58333 = ~pi7426 & ~pi9040;
assign w58334 = ~w58332 & ~w58333;
assign w58335 = pi3387 & ~w58334;
assign w58336 = ~pi3387 & w58334;
assign w58337 = ~w58335 & ~w58336;
assign w58338 = w58331 & w58337;
assign w58339 = ~pi7235 & pi9040;
assign w58340 = ~pi7230 & ~pi9040;
assign w58341 = ~w58339 & ~w58340;
assign w58342 = pi3351 & ~w58341;
assign w58343 = ~pi3351 & w58341;
assign w58344 = ~w58342 & ~w58343;
assign w58345 = ~pi7147 & pi9040;
assign w58346 = ~pi7423 & ~pi9040;
assign w58347 = ~w58345 & ~w58346;
assign w58348 = pi3311 & ~w58347;
assign w58349 = ~pi3311 & w58347;
assign w58350 = ~w58348 & ~w58349;
assign w58351 = ~w58344 & ~w58350;
assign w58352 = ~w58344 & w58350;
assign w58353 = ~pi7423 & pi9040;
assign w58354 = ~pi7234 & ~pi9040;
assign w58355 = ~w58353 & ~w58354;
assign w58356 = pi3353 & ~w58355;
assign w58357 = ~pi3353 & w58355;
assign w58358 = ~w58356 & ~w58357;
assign w58359 = w58352 & ~w58358;
assign w58360 = w58344 & ~w58350;
assign w58361 = w58331 & w58360;
assign w58362 = w58360 & w58365;
assign w58363 = ~w58359 & ~w58362;
assign w58364 = w58331 & w58350;
assign w58365 = w58331 & ~w58358;
assign w58366 = ~w58337 & ~w58344;
assign w58367 = ~w58364 & w58366;
assign w58368 = ~w58365 & w58367;
assign w58369 = w58363 & ~w58368;
assign w58370 = w58351 & w58369;
assign w58371 = ~w58352 & ~w58360;
assign w58372 = ~w58331 & ~w58371;
assign w58373 = (w58350 & w58371) | (w58350 & w58364) | (w58371 & w58364);
assign w58374 = (w58371 & w64176) | (w58371 & w64177) | (w64176 & w64177);
assign w58375 = (~w58338 & w58370) | (~w58338 & w63465) | (w58370 & w63465);
assign w58376 = w58344 & ~w58358;
assign w58377 = ~w58331 & w58350;
assign w58378 = w58376 & ~w58377;
assign w58379 = ~w58361 & ~w58378;
assign w58380 = w58337 & w58344;
assign w58381 = w58379 & w58380;
assign w58382 = w58369 & ~w58381;
assign w58383 = ~w58331 & w58360;
assign w58384 = w58360 & w63337;
assign w58385 = ~w58350 & ~w58358;
assign w58386 = ~w58331 & w58385;
assign w58387 = w58385 & w63338;
assign w58388 = ~w58384 & ~w58387;
assign w58389 = w58337 & ~w58344;
assign w58390 = ~w58358 & ~w58389;
assign w58391 = w58373 & w58390;
assign w58392 = ~w58331 & ~w58337;
assign w58393 = w58351 & w58392;
assign w58394 = w58352 & w58365;
assign w58395 = w58337 & ~w58394;
assign w58396 = w58352 & w58395;
assign w58397 = w58338 & w58385;
assign w58398 = ~w58393 & ~w58397;
assign w58399 = w58388 & w58398;
assign w58400 = ~w58391 & w58399;
assign w58401 = ~w58396 & w58400;
assign w58402 = w58382 & w58401;
assign w58403 = ~pi7138 & pi9040;
assign w58404 = ~pi7118 & ~pi9040;
assign w58405 = ~w58403 & ~w58404;
assign w58406 = pi3422 & ~w58405;
assign w58407 = ~pi3422 & w58405;
assign w58408 = ~w58406 & ~w58407;
assign w58409 = (w58408 & w58402) | (w58408 & w63466) | (w58402 & w63466);
assign w58410 = w58338 & ~w58363;
assign w58411 = w58408 & ~w58410;
assign w58412 = ~w58382 & ~w58411;
assign w58413 = w58344 & w58364;
assign w58414 = ~w58372 & ~w58413;
assign w58415 = ~w58337 & ~w58358;
assign w58416 = ~w58414 & w58415;
assign w58417 = ~w58412 & ~w58416;
assign w58418 = (pi3764 & w58409) | (pi3764 & w64178) | (w58409 & w64178);
assign w58419 = ~w58409 & w64179;
assign w58420 = ~w58418 & ~w58419;
assign w58421 = ~w58034 & ~w58064;
assign w58422 = w58143 & w58421;
assign w58423 = (~w58055 & w58056) | (~w58055 & w63467) | (w58056 & w63467);
assign w58424 = ~w58064 & ~w58423;
assign w58425 = ~w58079 & w58153;
assign w58426 = (w58092 & w58424) | (w58092 & w64180) | (w58424 & w64180);
assign w58427 = w58047 & ~w58421;
assign w58428 = ~w58150 & w58427;
assign w58429 = ~w58097 & w58428;
assign w58430 = w58053 & ~w58076;
assign w58431 = (~w58092 & w58151) | (~w58092 & w64181) | (w58151 & w64181);
assign w58432 = ~w58099 & ~w58422;
assign w58433 = ~w58431 & w58432;
assign w58434 = ~w58429 & w58433;
assign w58435 = ~w58426 & w58434;
assign w58436 = ~pi3824 & w58435;
assign w58437 = pi3824 & ~w58435;
assign w58438 = ~w58436 & ~w58437;
assign w58439 = ~w57928 & ~w57951;
assign w58440 = ~w57951 & w64182;
assign w58441 = ~w57930 & ~w58440;
assign w58442 = ~w57923 & ~w58441;
assign w58443 = w58002 & ~w58442;
assign w58444 = ~w57893 & ~w57951;
assign w58445 = w57996 & ~w58444;
assign w58446 = ~w58000 & w58445;
assign w58447 = w57931 & ~w58446;
assign w58448 = ~w58443 & ~w58447;
assign w58449 = w57902 & ~w58440;
assign w58450 = w58004 & ~w58439;
assign w58451 = ~w57902 & ~w57915;
assign w58452 = ~w57902 & ~w57933;
assign w58453 = ~w58451 & ~w58452;
assign w58454 = ~w58450 & ~w58453;
assign w58455 = ~w57995 & ~w58000;
assign w58456 = (w58455 & w58454) | (w58455 & w64183) | (w58454 & w64183);
assign w58457 = w57923 & ~w58456;
assign w58458 = ~w58448 & ~w58457;
assign w58459 = ~pi3771 & w58458;
assign w58460 = pi3771 & ~w58458;
assign w58461 = ~w58459 & ~w58460;
assign w58462 = w58053 & ~w58080;
assign w58463 = w58163 & w58462;
assign w58464 = w58077 & ~w58142;
assign w58465 = ~w58048 & ~w58092;
assign w58466 = ~w58078 & w58465;
assign w58467 = ~w58163 & ~w58466;
assign w58468 = ~w58464 & ~w58467;
assign w58469 = w58081 & w58462;
assign w58470 = w58149 & ~w58469;
assign w58471 = ~w58057 & w58470;
assign w58472 = ~w58468 & ~w58471;
assign w58473 = ~w58035 & ~w58064;
assign w58474 = w58156 & w58473;
assign w58475 = ~w58095 & w58474;
assign w58476 = ~w58463 & ~w58475;
assign w58477 = ~w58472 & w58476;
assign w58478 = pi3810 & ~w58477;
assign w58479 = ~pi3810 & w58477;
assign w58480 = ~w58478 & ~w58479;
assign w58481 = ~pi7224 & pi9040;
assign w58482 = ~pi7157 & ~pi9040;
assign w58483 = ~w58481 & ~w58482;
assign w58484 = pi3266 & ~w58483;
assign w58485 = ~pi3266 & w58483;
assign w58486 = ~w58484 & ~w58485;
assign w58487 = ~pi7228 & pi9040;
assign w58488 = ~pi7166 & ~pi9040;
assign w58489 = ~w58487 & ~w58488;
assign w58490 = pi3359 & ~w58489;
assign w58491 = ~pi3359 & w58489;
assign w58492 = ~w58490 & ~w58491;
assign w58493 = ~w58486 & w58492;
assign w58494 = ~pi7426 & pi9040;
assign w58495 = ~pi7169 & ~pi9040;
assign w58496 = ~w58494 & ~w58495;
assign w58497 = pi3324 & ~w58496;
assign w58498 = ~pi3324 & w58496;
assign w58499 = ~w58497 & ~w58498;
assign w58500 = w58493 & ~w58499;
assign w58501 = ~pi7234 & pi9040;
assign w58502 = ~pi7151 & ~pi9040;
assign w58503 = ~w58501 & ~w58502;
assign w58504 = pi3356 & ~w58503;
assign w58505 = ~pi3356 & w58503;
assign w58506 = ~w58504 & ~w58505;
assign w58507 = w58493 & w58544;
assign w58508 = w58486 & w58506;
assign w58509 = ~w58486 & ~w58506;
assign w58510 = ~w58508 & ~w58509;
assign w58511 = w58499 & ~w58510;
assign w58512 = ~w58499 & ~w58506;
assign w58513 = w58486 & w58492;
assign w58514 = w58512 & w58513;
assign w58515 = ~pi7140 & pi9040;
assign w58516 = ~pi7218 & ~pi9040;
assign w58517 = ~w58515 & ~w58516;
assign w58518 = pi3327 & ~w58517;
assign w58519 = ~pi3327 & w58517;
assign w58520 = ~w58518 & ~w58519;
assign w58521 = (w58520 & w58511) | (w58520 & w64184) | (w58511 & w64184);
assign w58522 = w58499 & w58520;
assign w58523 = w58499 & ~w58506;
assign w58524 = ~w58508 & ~w58523;
assign w58525 = ~w58522 & ~w58524;
assign w58526 = w58499 & ~w58525;
assign w58527 = ~w58492 & w58526;
assign w58528 = ~w58492 & w58512;
assign w58529 = ~w58499 & w58508;
assign w58530 = ~w58528 & ~w58529;
assign w58531 = ~w58520 & ~w58530;
assign w58532 = ~pi7151 & pi9040;
assign w58533 = ~pi7160 & ~pi9040;
assign w58534 = ~w58532 & ~w58533;
assign w58535 = pi3346 & ~w58534;
assign w58536 = ~pi3346 & w58534;
assign w58537 = ~w58535 & ~w58536;
assign w58538 = ~w58507 & w58537;
assign w58539 = ~w58531 & w58538;
assign w58540 = ~w58521 & w58539;
assign w58541 = w58513 & w58523;
assign w58542 = ~w58537 & ~w58541;
assign w58543 = w58520 & ~w58530;
assign w58544 = ~w58499 & w58506;
assign w58545 = w58493 & ~w58523;
assign w58546 = ~w58544 & w58545;
assign w58547 = w58542 & ~w58546;
assign w58548 = ~w58543 & w58547;
assign w58549 = (~w58548 & ~w58540) | (~w58548 & w64185) | (~w58540 & w64185);
assign w58550 = ~w58486 & ~w58492;
assign w58551 = w58523 & w58550;
assign w58552 = ~w58499 & ~w58509;
assign w58553 = ~w58551 & ~w58552;
assign w58554 = ~w58486 & w58553;
assign w58555 = w58486 & ~w58499;
assign w58556 = ~w58537 & ~w58555;
assign w58557 = ~w58554 & w58556;
assign w58558 = ~w58500 & ~w58541;
assign w58559 = ~w58557 & w58558;
assign w58560 = ~w58520 & ~w58559;
assign w58561 = ~w58549 & ~w58560;
assign w58562 = ~pi3779 & w58561;
assign w58563 = pi3779 & ~w58561;
assign w58564 = ~w58562 & ~w58563;
assign w58565 = w58379 & w64186;
assign w58566 = ~w58393 & ~w58413;
assign w58567 = w58358 & ~w58566;
assign w58568 = (w58408 & w58371) | (w58408 & w63468) | (w58371 & w63468);
assign w58569 = ~w58567 & w58568;
assign w58570 = w58337 & w58358;
assign w58571 = w58360 & w58570;
assign w58572 = w58331 & ~w58344;
assign w58573 = w58337 & ~w58572;
assign w58574 = ~w58360 & ~w58377;
assign w58575 = w58573 & w58574;
assign w58576 = ~w58394 & ~w58571;
assign w58577 = ~w58575 & w58576;
assign w58578 = ~w58352 & ~w58386;
assign w58579 = w58337 & w58578;
assign w58580 = w58577 & w58579;
assign w58581 = w58569 & ~w58580;
assign w58582 = w58358 & w58377;
assign w58583 = ~w58572 & ~w58582;
assign w58584 = ~w58337 & ~w58583;
assign w58585 = w58388 & ~w58408;
assign w58586 = ~w58584 & w58585;
assign w58587 = w58577 & w58586;
assign w58588 = ~w58581 & ~w58587;
assign w58589 = ~w58359 & w58573;
assign w58590 = ~w58578 & w58589;
assign w58591 = ~w58362 & ~w58590;
assign w58592 = ~w58380 & ~w58591;
assign w58593 = ~w58565 & ~w58592;
assign w58594 = ~w58588 & w58593;
assign w58595 = pi3760 & ~w58594;
assign w58596 = ~pi3760 & w58594;
assign w58597 = ~w58595 & ~w58596;
assign w58598 = w57677 & w57759;
assign w58599 = w57690 & w57755;
assign w58600 = ~w57688 & ~w57736;
assign w58601 = ~w57742 & ~w58598;
assign w58602 = ~w58599 & w58601;
assign w58603 = w58600 & w58602;
assign w58604 = w57717 & ~w58603;
assign w58605 = w57691 & w57693;
assign w58606 = (~w57717 & w57696) | (~w57717 & w64187) | (w57696 & w64187);
assign w58607 = ~w57701 & w58171;
assign w58608 = w57710 & ~w58606;
assign w58609 = ~w58607 & w58608;
assign w58610 = w57693 & ~w57717;
assign w58611 = ~w57710 & ~w58610;
assign w58612 = ~w57701 & w58611;
assign w58613 = ~w58609 & ~w58612;
assign w58614 = ~w58604 & ~w58613;
assign w58615 = ~pi3867 & ~w58614;
assign w58616 = pi3867 & w58614;
assign w58617 = ~w58615 & ~w58616;
assign w58618 = ~w58233 & w58268;
assign w58619 = w58269 & ~w58293;
assign w58620 = ~w58249 & ~w58252;
assign w58621 = (~w58233 & ~w58208) | (~w58233 & w58286) | (~w58208 & w58286);
assign w58622 = ~w58302 & w58621;
assign w58623 = ~w58620 & w58622;
assign w58624 = ~w58619 & w58623;
assign w58625 = w58221 & w58245;
assign w58626 = ~w58208 & ~w58625;
assign w58627 = w58249 & w58626;
assign w58628 = (~w58240 & w58627) | (~w58240 & w64188) | (w58627 & w64188);
assign w58629 = ~w58624 & w58628;
assign w58630 = ~w58225 & w58248;
assign w58631 = w58201 & w58248;
assign w58632 = ~w58207 & ~w58631;
assign w58633 = ~w58627 & w64189;
assign w58634 = ~w58263 & ~w58270;
assign w58635 = w58286 & ~w58634;
assign w58636 = w58242 & ~w58288;
assign w58637 = w58225 & w58636;
assign w58638 = ~w58630 & ~w58637;
assign w58639 = ~w58635 & w58638;
assign w58640 = (w58240 & ~w58639) | (w58240 & w64190) | (~w58639 & w64190);
assign w58641 = w58223 & w58248;
assign w58642 = ~w58259 & ~w58641;
assign w58643 = w58233 & ~w58642;
assign w58644 = ~w58618 & ~w58643;
assign w58645 = ~w58629 & w58644;
assign w58646 = (pi3864 & ~w58645) | (pi3864 & w64191) | (~w58645 & w64191);
assign w58647 = w58645 & w64192;
assign w58648 = ~w58646 & ~w58647;
assign w58649 = w58358 & w58371;
assign w58650 = w58371 & w64193;
assign w58651 = ~w58383 & w58395;
assign w58652 = ~w58376 & w58377;
assign w58653 = ~w58337 & ~w58652;
assign w58654 = ~w58362 & w58653;
assign w58655 = ~w58651 & ~w58654;
assign w58656 = ~w58650 & ~w58655;
assign w58657 = (w58408 & w58655) | (w58408 & w64194) | (w58655 & w64194);
assign w58658 = ~w58401 & ~w58408;
assign w58659 = ~w58387 & ~w58650;
assign w58660 = ~w58337 & ~w58659;
assign w58661 = ~w58565 & ~w58571;
assign w58662 = ~w58660 & w58661;
assign w58663 = ~w58657 & w58662;
assign w58664 = ~w58658 & w58663;
assign w58665 = pi3767 & ~w58664;
assign w58666 = ~pi3767 & w58664;
assign w58667 = ~w58665 & ~w58666;
assign w58668 = ~pi7162 & pi9040;
assign w58669 = ~pi7140 & ~pi9040;
assign w58670 = ~w58668 & ~w58669;
assign w58671 = pi3346 & ~w58670;
assign w58672 = ~pi3346 & w58670;
assign w58673 = ~w58671 & ~w58672;
assign w58674 = ~pi7231 & pi9040;
assign w58675 = ~pi7236 & ~pi9040;
assign w58676 = ~w58674 & ~w58675;
assign w58677 = pi3351 & ~w58676;
assign w58678 = ~pi3351 & w58676;
assign w58679 = ~w58677 & ~w58678;
assign w58680 = ~w58673 & w58679;
assign w58681 = ~pi7236 & pi9040;
assign w58682 = ~pi7229 & ~pi9040;
assign w58683 = ~w58681 & ~w58682;
assign w58684 = pi3356 & ~w58683;
assign w58685 = ~pi3356 & w58683;
assign w58686 = ~w58684 & ~w58685;
assign w58687 = ~pi7155 & pi9040;
assign w58688 = ~pi7162 & ~pi9040;
assign w58689 = ~w58687 & ~w58688;
assign w58690 = pi3330 & ~w58689;
assign w58691 = ~pi3330 & w58689;
assign w58692 = ~w58690 & ~w58691;
assign w58693 = w58686 & w58692;
assign w58694 = w58680 & w58693;
assign w58695 = ~pi7166 & pi9040;
assign w58696 = ~pi7085 & ~pi9040;
assign w58697 = ~w58695 & ~w58696;
assign w58698 = pi3311 & ~w58697;
assign w58699 = ~pi3311 & w58697;
assign w58700 = ~w58698 & ~w58699;
assign w58701 = ~pi7160 & pi9040;
assign w58702 = ~pi7228 & ~pi9040;
assign w58703 = ~w58701 & ~w58702;
assign w58704 = pi3265 & ~w58703;
assign w58705 = ~pi3265 & w58703;
assign w58706 = ~w58704 & ~w58705;
assign w58707 = ~w58679 & ~w58706;
assign w58708 = ~w58673 & ~w58692;
assign w58709 = w58673 & w58692;
assign w58710 = w58707 & ~w58708;
assign w58711 = ~w58709 & w58710;
assign w58712 = ~w58673 & ~w58679;
assign w58713 = w58686 & w58706;
assign w58714 = w58712 & ~w58713;
assign w58715 = w58673 & ~w58686;
assign w58716 = w58673 & ~w58679;
assign w58717 = ~w58680 & ~w58716;
assign w58718 = (~w58715 & w58717) | (~w58715 & w64195) | (w58717 & w64195);
assign w58719 = w58673 & w58679;
assign w58720 = ~w58715 & ~w58719;
assign w58721 = w58679 & w58715;
assign w58722 = ~w58720 & ~w58721;
assign w58723 = ~w58718 & ~w58722;
assign w58724 = ~w58692 & ~w58714;
assign w58725 = ~w58723 & w58724;
assign w58726 = ~w58694 & w58700;
assign w58727 = ~w58711 & w58726;
assign w58728 = ~w58725 & w58727;
assign w58729 = ~w58686 & ~w58692;
assign w58730 = w58712 & w58729;
assign w58731 = w58706 & w58723;
assign w58732 = ~w58700 & ~w58730;
assign w58733 = ~w58731 & w58732;
assign w58734 = ~w58728 & ~w58733;
assign w58735 = ~w58686 & w58709;
assign w58736 = w58692 & w58712;
assign w58737 = ~w58700 & ~w58736;
assign w58738 = w58718 & w58737;
assign w58739 = ~w58735 & ~w58738;
assign w58740 = ~w58706 & ~w58739;
assign w58741 = w58692 & w58706;
assign w58742 = ~w58693 & ~w58729;
assign w58743 = w58680 & ~w58706;
assign w58744 = ~w58742 & w58743;
assign w58745 = w58708 & w58713;
assign w58746 = w58716 & ~w58742;
assign w58747 = ~w58745 & ~w58746;
assign w58748 = w58717 & w58742;
assign w58749 = ~w58744 & ~w58748;
assign w58750 = w58747 & w58749;
assign w58751 = ~w58715 & w58741;
assign w58752 = ~w58750 & w58751;
assign w58753 = ~w58740 & ~w58752;
assign w58754 = ~w58734 & w58753;
assign w58755 = pi3789 & ~w58754;
assign w58756 = ~pi3789 & w58754;
assign w58757 = ~w58755 & ~w58756;
assign w58758 = ~w57895 & ~w57928;
assign w58759 = ~w57908 & ~w58758;
assign w58760 = ~w57944 & ~w58759;
assign w58761 = ~w58759 & w63469;
assign w58762 = w57947 & w57951;
assign w58763 = w58001 & ~w58762;
assign w58764 = ~w57997 & w58763;
assign w58765 = w57895 & w57959;
assign w58766 = (~w58765 & w58764) | (~w58765 & w63470) | (w58764 & w63470);
assign w58767 = w57887 & w57944;
assign w58768 = ~w58453 & ~w58767;
assign w58769 = w57902 & ~w57939;
assign w58770 = ~w58768 & ~w58769;
assign w58771 = w57887 & ~w58451;
assign w58772 = w58760 & w58771;
assign w58773 = (~w57935 & ~w58763) | (~w57935 & w64196) | (~w58763 & w64196);
assign w58774 = ~w58772 & w58773;
assign w58775 = ~w57923 & ~w58774;
assign w58776 = (~w58770 & w58766) | (~w58770 & w64197) | (w58766 & w64197);
assign w58777 = ~w58775 & w58776;
assign w58778 = ~pi3770 & w58777;
assign w58779 = pi3770 & ~w58777;
assign w58780 = ~w58778 & ~w58779;
assign w58781 = w58493 & w58512;
assign w58782 = ~w58499 & ~w58537;
assign w58783 = w58499 & w58537;
assign w58784 = w58492 & ~w58783;
assign w58785 = w58486 & ~w58782;
assign w58786 = ~w58784 & w58785;
assign w58787 = ~w58781 & ~w58786;
assign w58788 = w58520 & ~w58787;
assign w58789 = ~w58486 & ~w58520;
assign w58790 = ~w58492 & w58506;
assign w58791 = ~w58544 & ~w58790;
assign w58792 = w58789 & ~w58791;
assign w58793 = w58522 & w58545;
assign w58794 = w58499 & w58506;
assign w58795 = w58510 & ~w58794;
assign w58796 = w58510 & w64198;
assign w58797 = w58492 & w58525;
assign w58798 = ~w58792 & ~w58793;
assign w58799 = ~w58796 & w58798;
assign w58800 = (~w58537 & ~w58799) | (~w58537 & w64199) | (~w58799 & w64199);
assign w58801 = ~w58492 & w58511;
assign w58802 = ~w58513 & ~w58550;
assign w58803 = ~w58499 & ~w58802;
assign w58804 = ~w58546 & ~w58803;
assign w58805 = ~w58520 & ~w58804;
assign w58806 = ~w58801 & ~w58805;
assign w58807 = w58537 & ~w58806;
assign w58808 = ~w58788 & ~w58800;
assign w58809 = ~w58807 & w58808;
assign w58810 = pi3847 & w58809;
assign w58811 = ~pi3847 & ~w58809;
assign w58812 = ~w58810 & ~w58811;
assign w58813 = w58693 & w58707;
assign w58814 = w58686 & w58712;
assign w58815 = ~w58709 & ~w58814;
assign w58816 = ~w58706 & ~w58815;
assign w58817 = w58679 & w58708;
assign w58818 = ~w58736 & ~w58817;
assign w58819 = w58716 & w58729;
assign w58820 = (w58706 & ~w58818) | (w58706 & w64200) | (~w58818 & w64200);
assign w58821 = w58693 & ~w58719;
assign w58822 = ~w58816 & ~w58821;
assign w58823 = ~w58820 & w58822;
assign w58824 = w58700 & ~w58823;
assign w58825 = ~w58735 & ~w58814;
assign w58826 = w58818 & w58825;
assign w58827 = ~w58700 & ~w58722;
assign w58828 = w58826 & w58827;
assign w58829 = w58721 & w58741;
assign w58830 = ~w58692 & ~w58706;
assign w58831 = ~w58741 & ~w58830;
assign w58832 = ~w58720 & ~w58831;
assign w58833 = ~w58680 & w58706;
assign w58834 = ~w58743 & ~w58833;
assign w58835 = w58686 & ~w58719;
assign w58836 = ~w58741 & w58835;
assign w58837 = ~w58834 & w58836;
assign w58838 = ~w58832 & ~w58837;
assign w58839 = ~w58700 & ~w58838;
assign w58840 = ~w58813 & ~w58829;
assign w58841 = (w58840 & ~w58828) | (w58840 & w64201) | (~w58828 & w64201);
assign w58842 = ~w58839 & w58841;
assign w58843 = ~w58824 & w58842;
assign w58844 = pi3780 & ~w58843;
assign w58845 = ~pi3780 & w58843;
assign w58846 = ~w58844 & ~w58845;
assign w58847 = w58693 & w58719;
assign w58848 = (~w58706 & w58828) | (~w58706 & w64202) | (w58828 & w64202);
assign w58849 = ~w58706 & ~w58729;
assign w58850 = w58717 & w58849;
assign w58851 = w58741 & w58826;
assign w58852 = w58729 & ~w58834;
assign w58853 = ~w58819 & ~w58850;
assign w58854 = ~w58852 & w58853;
assign w58855 = ~w58851 & w58854;
assign w58856 = w58700 & ~w58855;
assign w58857 = ~w58747 & w58820;
assign w58858 = ~w58700 & ~w58743;
assign w58859 = ~w58850 & w58858;
assign w58860 = ~w58826 & w58859;
assign w58861 = ~w58857 & ~w58860;
assign w58862 = ~w58848 & w58861;
assign w58863 = ~w58856 & w58862;
assign w58864 = pi3844 & ~w58863;
assign w58865 = ~pi3844 & w58863;
assign w58866 = ~w58864 & ~w58865;
assign w58867 = ~w58700 & ~w58750;
assign w58868 = w58708 & w64203;
assign w58869 = ~w58722 & ~w58868;
assign w58870 = (~w58706 & w58722) | (~w58706 & w64204) | (w58722 & w64204);
assign w58871 = w58692 & w58814;
assign w58872 = ~w58870 & ~w58871;
assign w58873 = w58700 & ~w58872;
assign w58874 = w58700 & ~w58712;
assign w58875 = w58869 & w58874;
assign w58876 = w58679 & ~w58686;
assign w58877 = w58692 & w58876;
assign w58878 = ~w58730 & ~w58877;
assign w58879 = ~w58875 & w58878;
assign w58880 = w58706 & ~w58879;
assign w58881 = ~w58867 & ~w58873;
assign w58882 = ~w58880 & w58881;
assign w58883 = ~pi3857 & w58882;
assign w58884 = pi3857 & ~w58882;
assign w58885 = ~w58883 & ~w58884;
assign w58886 = w58570 & ~w58656;
assign w58887 = (~w58392 & w58567) | (~w58392 & w63471) | (w58567 & w63471);
assign w58888 = w58649 & ~w58887;
assign w58889 = w58350 & ~w58389;
assign w58890 = ~w58378 & w58889;
assign w58891 = ~w58582 & w58890;
assign w58892 = (~w58408 & ~w58591) | (~w58408 & w64205) | (~w58591 & w64205);
assign w58893 = ~w58337 & w58379;
assign w58894 = w58408 & ~w58589;
assign w58895 = ~w58893 & w58894;
assign w58896 = ~w58888 & ~w58895;
assign w58897 = ~w58892 & w58896;
assign w58898 = (pi3841 & ~w58897) | (pi3841 & w64206) | (~w58897 & w64206);
assign w58899 = w58897 & w64207;
assign w58900 = ~w58898 & ~w58899;
assign w58901 = ~w58544 & ~w58550;
assign w58902 = w58790 & w58901;
assign w58903 = ~w58541 & ~w58902;
assign w58904 = ~w58508 & ~w58537;
assign w58905 = ~w58790 & w58904;
assign w58906 = ~w58553 & w58905;
assign w58907 = w58903 & ~w58906;
assign w58908 = ~w58520 & ~w58907;
assign w58909 = ~w58790 & ~w58901;
assign w58910 = w58789 & ~w58909;
assign w58911 = w58486 & w58528;
assign w58912 = ~w58789 & w58909;
assign w58913 = w58903 & ~w58911;
assign w58914 = ~w58910 & ~w58912;
assign w58915 = w58913 & w58914;
assign w58916 = w58537 & ~w58915;
assign w58917 = w58782 & ~w58789;
assign w58918 = w58790 & w58917;
assign w58919 = w58520 & ~w58552;
assign w58920 = w58542 & w58919;
assign w58921 = ~w58801 & w58920;
assign w58922 = ~w58918 & ~w58921;
assign w58923 = ~w58908 & w58922;
assign w58924 = ~w58916 & w58923;
assign w58925 = pi3856 & ~w58924;
assign w58926 = ~pi3856 & w58924;
assign w58927 = ~w58925 & ~w58926;
assign w58928 = (w58233 & ~w58245) | (w58233 & w64208) | (~w58245 & w64208);
assign w58929 = w58620 & w58928;
assign w58930 = ~w58631 & w58928;
assign w58931 = ~w58626 & w58930;
assign w58932 = ~w58263 & ~w58275;
assign w58933 = ~w58302 & w58932;
assign w58934 = (w58240 & ~w58933) | (w58240 & w64209) | (~w58933 & w64209);
assign w58935 = w58244 & ~w58269;
assign w58936 = ~w58930 & ~w58935;
assign w58937 = w58224 & ~w58248;
assign w58938 = ~w58936 & ~w58937;
assign w58939 = ~w58240 & ~w58938;
assign w58940 = ~w58271 & w58627;
assign w58941 = (~w58233 & w58940) | (~w58233 & w64210) | (w58940 & w64210);
assign w58942 = ~w58929 & ~w58934;
assign w58943 = ~w58939 & ~w58941;
assign w58944 = w58942 & w58943;
assign w58945 = pi3921 & ~w58944;
assign w58946 = ~pi3921 & w58944;
assign w58947 = ~w58945 & ~w58946;
assign w58948 = w58520 & w58795;
assign w58949 = ~w58781 & ~w58948;
assign w58950 = w58537 & ~w58949;
assign w58951 = w58492 & w58794;
assign w58952 = ~w58508 & ~w58951;
assign w58953 = w58526 & ~w58952;
assign w58954 = w58520 & w58555;
assign w58955 = ~w58794 & ~w58802;
assign w58956 = ~w58954 & w58955;
assign w58957 = ~w58953 & ~w58956;
assign w58958 = ~w58537 & ~w58957;
assign w58959 = ~w58509 & ~w58790;
assign w58960 = w58783 & ~w58959;
assign w58961 = ~w58520 & ~w58529;
assign w58962 = ~w58960 & w58961;
assign w58963 = w58520 & ~w58951;
assign w58964 = ~w58911 & w58963;
assign w58965 = ~w58962 & ~w58964;
assign w58966 = ~w58950 & ~w58965;
assign w58967 = ~w58958 & w58966;
assign w58968 = ~pi3917 & w58967;
assign w58969 = pi3917 & ~w58967;
assign w58970 = ~w58968 & ~w58969;
assign w58971 = ~pi7386 & pi9040;
assign w58972 = ~pi7431 & ~pi9040;
assign w58973 = ~w58971 & ~w58972;
assign w58974 = pi3782 & ~w58973;
assign w58975 = ~pi3782 & w58973;
assign w58976 = ~w58974 & ~w58975;
assign w58977 = ~pi7454 & pi9040;
assign w58978 = ~pi7425 & ~pi9040;
assign w58979 = ~w58977 & ~w58978;
assign w58980 = pi3895 & ~w58979;
assign w58981 = ~pi3895 & w58979;
assign w58982 = ~w58980 & ~w58981;
assign w58983 = ~w58976 & ~w58982;
assign w58984 = ~pi7431 & pi9040;
assign w58985 = ~pi7568 & ~pi9040;
assign w58986 = ~w58984 & ~w58985;
assign w58987 = pi3866 & ~w58986;
assign w58988 = ~pi3866 & w58986;
assign w58989 = ~w58987 & ~w58988;
assign w58990 = ~pi7453 & pi9040;
assign w58991 = ~pi7461 & ~pi9040;
assign w58992 = ~w58990 & ~w58991;
assign w58993 = pi3929 & ~w58992;
assign w58994 = ~pi3929 & w58992;
assign w58995 = ~w58993 & ~w58994;
assign w58996 = ~w58989 & ~w58995;
assign w58997 = ~pi7534 & pi9040;
assign w58998 = ~pi7385 & ~pi9040;
assign w58999 = ~w58997 & ~w58998;
assign w59000 = pi3912 & ~w58999;
assign w59001 = ~pi3912 & w58999;
assign w59002 = ~w59000 & ~w59001;
assign w59003 = w58996 & ~w59002;
assign w59004 = w58983 & w59003;
assign w59005 = ~pi7449 & pi9040;
assign w59006 = ~pi7534 & ~pi9040;
assign w59007 = ~w59005 & ~w59006;
assign w59008 = pi3936 & ~w59007;
assign w59009 = ~pi3936 & w59007;
assign w59010 = ~w59008 & ~w59009;
assign w59011 = ~w58989 & ~w59002;
assign w59012 = ~w58976 & w58995;
assign w59013 = ~w59011 & w59012;
assign w59014 = w58989 & w58995;
assign w59015 = w58976 & ~w59014;
assign w59016 = ~w58982 & ~w59013;
assign w59017 = ~w59015 & w59016;
assign w59018 = w58995 & w59002;
assign w59019 = w58976 & w59018;
assign w59020 = ~w58976 & w58989;
assign w59021 = w58976 & ~w58989;
assign w59022 = ~w59020 & ~w59021;
assign w59023 = w58976 & w59003;
assign w59024 = ~w58976 & w59002;
assign w59025 = w58996 & ~w59024;
assign w59026 = w58995 & ~w59002;
assign w59027 = ~w58995 & w59002;
assign w59028 = w58989 & ~w59027;
assign w59029 = ~w59026 & w59028;
assign w59030 = ~w59025 & ~w59029;
assign w59031 = ~w59023 & ~w59030;
assign w59032 = ~w59030 & w64211;
assign w59033 = w58982 & ~w59019;
assign w59034 = ~w59032 & w59033;
assign w59035 = ~w58982 & w59002;
assign w59036 = ~w59022 & w59035;
assign w59037 = w59010 & ~w59036;
assign w59038 = ~w59017 & w59037;
assign w59039 = ~w59034 & w59038;
assign w59040 = ~w58996 & ~w59002;
assign w59041 = w58982 & ~w59020;
assign w59042 = w59040 & w59041;
assign w59043 = ~w59036 & ~w59042;
assign w59044 = ~w58976 & ~w58995;
assign w59045 = ~w58982 & w58989;
assign w59046 = w59044 & w59045;
assign w59047 = w58976 & w59014;
assign w59048 = w59014 & w64212;
assign w59049 = ~w59046 & ~w59048;
assign w59050 = w58989 & w59027;
assign w59051 = w58982 & ~w58989;
assign w59052 = ~w59050 & ~w59051;
assign w59053 = ~w58976 & ~w59052;
assign w59054 = w59043 & w59049;
assign w59055 = (~w59010 & ~w59054) | (~w59010 & w64213) | (~w59054 & w64213);
assign w59056 = ~w59043 & w59053;
assign w59057 = w58996 & w59024;
assign w59058 = ~w59047 & ~w59057;
assign w59059 = w58982 & ~w59058;
assign w59060 = ~w59004 & ~w59059;
assign w59061 = ~w59056 & w59060;
assign w59062 = ~w59055 & w59061;
assign w59063 = ~w59039 & w59062;
assign w59064 = pi5202 & ~w59063;
assign w59065 = ~pi5202 & w59063;
assign w59066 = ~w59064 & ~w59065;
assign w59067 = ~pi7424 & pi9040;
assign w59068 = ~pi7410 & ~pi9040;
assign w59069 = ~w59067 & ~w59068;
assign w59070 = pi3892 & ~w59069;
assign w59071 = ~pi3892 & w59069;
assign w59072 = ~w59070 & ~w59071;
assign w59073 = ~pi7413 & pi9040;
assign w59074 = ~pi7383 & ~pi9040;
assign w59075 = ~w59073 & ~w59074;
assign w59076 = pi3862 & ~w59075;
assign w59077 = ~pi3862 & w59075;
assign w59078 = ~w59076 & ~w59077;
assign w59079 = w59072 & w59078;
assign w59080 = ~pi7417 & pi9040;
assign w59081 = ~pi7444 & ~pi9040;
assign w59082 = ~w59080 & ~w59081;
assign w59083 = pi3845 & ~w59082;
assign w59084 = ~pi3845 & w59082;
assign w59085 = ~w59083 & ~w59084;
assign w59086 = w59079 & ~w59085;
assign w59087 = ~w59072 & ~w59085;
assign w59088 = ~w59078 & w59087;
assign w59089 = ~w59086 & ~w59088;
assign w59090 = ~pi7412 & pi9040;
assign w59091 = ~pi7369 & ~pi9040;
assign w59092 = ~w59090 & ~w59091;
assign w59093 = pi3839 & ~w59092;
assign w59094 = ~pi3839 & w59092;
assign w59095 = ~w59093 & ~w59094;
assign w59096 = ~w59089 & ~w59095;
assign w59097 = ~pi7518 & pi9040;
assign w59098 = ~pi7450 & ~pi9040;
assign w59099 = ~w59097 & ~w59098;
assign w59100 = pi3931 & ~w59099;
assign w59101 = ~pi3931 & w59099;
assign w59102 = ~w59100 & ~w59101;
assign w59103 = w59085 & ~w59102;
assign w59104 = w59072 & ~w59078;
assign w59105 = ~w59103 & ~w59104;
assign w59106 = ~w59078 & w59103;
assign w59107 = (w59095 & ~w59103) | (w59095 & w64214) | (~w59103 & w64214);
assign w59108 = ~w59072 & w59095;
assign w59109 = ~w59107 & ~w59108;
assign w59110 = ~w59105 & ~w59109;
assign w59111 = ~pi7383 & pi9040;
assign w59112 = ~pi7412 & ~pi9040;
assign w59113 = ~w59111 & ~w59112;
assign w59114 = pi3863 & ~w59113;
assign w59115 = ~pi3863 & w59113;
assign w59116 = ~w59114 & ~w59115;
assign w59117 = ~w59072 & w59078;
assign w59118 = w59085 & w59117;
assign w59119 = w59117 & w59123;
assign w59120 = w59116 & ~w59119;
assign w59121 = ~w59096 & w59120;
assign w59122 = ~w59110 & w59121;
assign w59123 = w59085 & w59102;
assign w59124 = ~w59079 & w59095;
assign w59125 = w59123 & ~w59124;
assign w59126 = w59104 & ~w59107;
assign w59127 = w59078 & ~w59102;
assign w59128 = ~w59072 & ~w59095;
assign w59129 = w59127 & w59128;
assign w59130 = ~w59116 & ~w59129;
assign w59131 = ~w59125 & w59130;
assign w59132 = ~w59126 & w59131;
assign w59133 = w59072 & ~w59095;
assign w59134 = w59106 & w59133;
assign w59135 = w59087 & w59102;
assign w59136 = w59079 & w64215;
assign w59137 = ~w59135 & ~w59136;
assign w59138 = ~w59116 & ~w59137;
assign w59139 = ~w59078 & w59102;
assign w59140 = ~w59085 & w59139;
assign w59141 = w59078 & w59102;
assign w59142 = ~w59118 & ~w59141;
assign w59143 = ~w59140 & w59142;
assign w59144 = (~w59105 & ~w59142) | (~w59105 & w64216) | (~w59142 & w64216);
assign w59145 = ~w59127 & ~w59139;
assign w59146 = w59087 & w59145;
assign w59147 = ~w59138 & ~w59146;
assign w59148 = ~w59144 & w59147;
assign w59149 = w59095 & ~w59148;
assign w59150 = (~w59134 & w59122) | (~w59134 & w64217) | (w59122 & w64217);
assign w59151 = ~w59149 & w59150;
assign w59152 = pi5217 & ~w59151;
assign w59153 = ~pi5217 & w59151;
assign w59154 = ~w59152 & ~w59153;
assign w59155 = ~pi7511 & pi9040;
assign w59156 = ~pi7446 & ~pi9040;
assign w59157 = ~w59155 & ~w59156;
assign w59158 = pi3842 & ~w59157;
assign w59159 = ~pi3842 & w59157;
assign w59160 = ~w59158 & ~w59159;
assign w59161 = ~pi7522 & pi9040;
assign w59162 = ~pi7439 & ~pi9040;
assign w59163 = ~w59161 & ~w59162;
assign w59164 = pi3851 & ~w59163;
assign w59165 = ~pi3851 & w59163;
assign w59166 = ~w59164 & ~w59165;
assign w59167 = ~w59160 & ~w59166;
assign w59168 = ~pi7591 & pi9040;
assign w59169 = ~pi7421 & ~pi9040;
assign w59170 = ~w59168 & ~w59169;
assign w59171 = pi3865 & ~w59170;
assign w59172 = ~pi3865 & w59170;
assign w59173 = ~w59171 & ~w59172;
assign w59174 = ~w59166 & w59173;
assign w59175 = ~w59167 & ~w59174;
assign w59176 = ~pi7466 & pi9040;
assign w59177 = ~pi7422 & ~pi9040;
assign w59178 = ~w59176 & ~w59177;
assign w59179 = pi3958 & ~w59178;
assign w59180 = ~pi3958 & w59178;
assign w59181 = ~w59179 & ~w59180;
assign w59182 = ~w59173 & w59181;
assign w59183 = ~pi7421 & pi9040;
assign w59184 = ~pi7521 & ~pi9040;
assign w59185 = ~w59183 & ~w59184;
assign w59186 = pi3930 & ~w59185;
assign w59187 = ~pi3930 & w59185;
assign w59188 = ~w59186 & ~w59187;
assign w59189 = w59160 & ~w59188;
assign w59190 = w59181 & w59189;
assign w59191 = ~pi7434 & pi9040;
assign w59192 = ~pi7511 & ~pi9040;
assign w59193 = ~w59191 & ~w59192;
assign w59194 = pi3940 & ~w59193;
assign w59195 = ~pi3940 & w59193;
assign w59196 = ~w59194 & ~w59195;
assign w59197 = ~w59173 & ~w59188;
assign w59198 = w59173 & w59188;
assign w59199 = ~w59197 & ~w59198;
assign w59200 = ~w59160 & ~w59199;
assign w59201 = ~w59160 & ~w59188;
assign w59202 = w59181 & w59201;
assign w59203 = ~w59196 & ~w59202;
assign w59204 = ~w59200 & w59203;
assign w59205 = ~w59182 & ~w59190;
assign w59206 = ~w59204 & w59205;
assign w59207 = ~w59175 & ~w59206;
assign w59208 = ~w59160 & w59181;
assign w59209 = ~w59173 & w59188;
assign w59210 = w59208 & w59209;
assign w59211 = ~w59160 & w59198;
assign w59212 = (~w59166 & ~w59198) | (~w59166 & w64218) | (~w59198 & w64218);
assign w59213 = w59173 & ~w59181;
assign w59214 = ~w59212 & w59213;
assign w59215 = ~w59173 & ~w59189;
assign w59216 = w59160 & w59188;
assign w59217 = ~w59201 & ~w59216;
assign w59218 = ~w59182 & w59217;
assign w59219 = w59166 & ~w59218;
assign w59220 = ~w59215 & w59219;
assign w59221 = ~w59181 & w59197;
assign w59222 = w59160 & w59209;
assign w59223 = ~w59221 & ~w59222;
assign w59224 = ~w59166 & ~w59223;
assign w59225 = w59196 & ~w59210;
assign w59226 = ~w59214 & w59225;
assign w59227 = ~w59224 & w59226;
assign w59228 = ~w59220 & w59227;
assign w59229 = w59189 & w64219;
assign w59230 = ~w59196 & ~w59229;
assign w59231 = w59166 & ~w59223;
assign w59232 = w59181 & w59200;
assign w59233 = w59230 & ~w59231;
assign w59234 = ~w59232 & w59233;
assign w59235 = ~w59228 & ~w59234;
assign w59236 = ~w59207 & ~w59235;
assign w59237 = ~pi5280 & w59236;
assign w59238 = pi5280 & ~w59236;
assign w59239 = ~w59237 & ~w59238;
assign w59240 = ~pi7462 & pi9040;
assign w59241 = ~pi7386 & ~pi9040;
assign w59242 = ~w59240 & ~w59241;
assign w59243 = pi3936 & ~w59242;
assign w59244 = ~pi3936 & w59242;
assign w59245 = ~w59243 & ~w59244;
assign w59246 = ~pi7450 & pi9040;
assign w59247 = ~pi7424 & ~pi9040;
assign w59248 = ~w59246 & ~w59247;
assign w59249 = pi3853 & ~w59248;
assign w59250 = ~pi3853 & w59248;
assign w59251 = ~w59249 & ~w59250;
assign w59252 = ~w59245 & ~w59251;
assign w59253 = w59245 & w59251;
assign w59254 = ~w59252 & ~w59253;
assign w59255 = ~pi7444 & pi9040;
assign w59256 = ~pi7409 & ~pi9040;
assign w59257 = ~w59255 & ~w59256;
assign w59258 = pi3929 & ~w59257;
assign w59259 = ~pi3929 & w59257;
assign w59260 = ~w59258 & ~w59259;
assign w59261 = ~w59254 & w59260;
assign w59262 = ~pi7409 & pi9040;
assign w59263 = ~pi7433 & ~pi9040;
assign w59264 = ~w59262 & ~w59263;
assign w59265 = pi3875 & ~w59264;
assign w59266 = ~pi3875 & w59264;
assign w59267 = ~w59265 & ~w59266;
assign w59268 = ~w59261 & ~w59267;
assign w59269 = ~pi7410 & pi9040;
assign w59270 = ~pi7518 & ~pi9040;
assign w59271 = ~w59269 & ~w59270;
assign w59272 = pi3845 & ~w59271;
assign w59273 = ~pi3845 & w59271;
assign w59274 = ~w59272 & ~w59273;
assign w59275 = ~w59245 & w59274;
assign w59276 = w59251 & ~w59260;
assign w59277 = w59275 & w59276;
assign w59278 = w59267 & ~w59277;
assign w59279 = ~w59251 & w59260;
assign w59280 = w59245 & w59260;
assign w59281 = ~w59245 & w59276;
assign w59282 = ~w59280 & ~w59281;
assign w59283 = ~w59281 & w63472;
assign w59284 = ~w59279 & w59283;
assign w59285 = w59278 & ~w59284;
assign w59286 = ~w59268 & ~w59285;
assign w59287 = ~w59260 & w59267;
assign w59288 = w59274 & ~w59287;
assign w59289 = ~w59254 & w59288;
assign w59290 = ~pi7429 & pi9040;
assign w59291 = ~pi7411 & ~pi9040;
assign w59292 = ~w59290 & ~w59291;
assign w59293 = pi3892 & ~w59292;
assign w59294 = ~pi3892 & w59292;
assign w59295 = ~w59293 & ~w59294;
assign w59296 = (~w59267 & w59281) | (~w59267 & w63473) | (w59281 & w63473);
assign w59297 = ~w59274 & w59296;
assign w59298 = ~w59251 & ~w59260;
assign w59299 = w59245 & ~w59274;
assign w59300 = w59245 & w59267;
assign w59301 = ~w59299 & ~w59300;
assign w59302 = w59298 & ~w59301;
assign w59303 = ~w59289 & ~w59295;
assign w59304 = ~w59302 & w59303;
assign w59305 = ~w59297 & w59304;
assign w59306 = ~w59260 & ~w59274;
assign w59307 = w59252 & w59306;
assign w59308 = w59260 & ~w59274;
assign w59309 = ~w59267 & ~w59308;
assign w59310 = ~w59275 & ~w59299;
assign w59311 = w59260 & ~w59310;
assign w59312 = w59245 & w59274;
assign w59313 = w59298 & w59312;
assign w59314 = (w59309 & w59311) | (w59309 & w63474) | (w59311 & w63474);
assign w59315 = w59251 & w59260;
assign w59316 = ~w59298 & ~w59308;
assign w59317 = ~w59315 & w59316;
assign w59318 = w59300 & w59317;
assign w59319 = ~w59277 & w59295;
assign w59320 = ~w59307 & w59319;
assign w59321 = ~w59318 & w59320;
assign w59322 = ~w59314 & w59321;
assign w59323 = ~w59305 & ~w59322;
assign w59324 = ~w59286 & ~w59323;
assign w59325 = ~pi5307 & w59324;
assign w59326 = pi5307 & ~w59324;
assign w59327 = ~w59325 & ~w59326;
assign w59328 = ~pi7415 & pi9040;
assign w59329 = ~pi7434 & ~pi9040;
assign w59330 = ~w59328 & ~w59329;
assign w59331 = pi3863 & ~w59330;
assign w59332 = ~pi3863 & w59330;
assign w59333 = ~w59331 & ~w59332;
assign w59334 = ~pi7440 & pi9040;
assign w59335 = ~pi7591 & ~pi9040;
assign w59336 = ~w59334 & ~w59335;
assign w59337 = pi3989 & ~w59336;
assign w59338 = ~pi3989 & w59336;
assign w59339 = ~w59337 & ~w59338;
assign w59340 = ~w59333 & w59339;
assign w59341 = ~pi7396 & pi9040;
assign w59342 = ~pi7379 & ~pi9040;
assign w59343 = ~w59341 & ~w59342;
assign w59344 = pi3842 & ~w59343;
assign w59345 = ~pi3842 & w59343;
assign w59346 = ~w59344 & ~w59345;
assign w59347 = ~pi7521 & pi9040;
assign w59348 = ~pi7440 & ~pi9040;
assign w59349 = ~w59347 & ~w59348;
assign w59350 = pi3931 & ~w59349;
assign w59351 = ~pi3931 & w59349;
assign w59352 = ~w59350 & ~w59351;
assign w59353 = ~w59346 & ~w59352;
assign w59354 = ~pi7436 & pi9040;
assign w59355 = ~pi7414 & ~pi9040;
assign w59356 = ~w59354 & ~w59355;
assign w59357 = pi3935 & ~w59356;
assign w59358 = ~pi3935 & w59356;
assign w59359 = ~w59357 & ~w59358;
assign w59360 = w59353 & w59359;
assign w59361 = w59340 & w59360;
assign w59362 = ~w59352 & ~w59359;
assign w59363 = w59333 & w59362;
assign w59364 = w59339 & w59363;
assign w59365 = ~w59333 & ~w59359;
assign w59366 = w59352 & ~w59365;
assign w59367 = w59339 & w59346;
assign w59368 = ~w59366 & w59367;
assign w59369 = ~pi7575 & pi9040;
assign w59370 = ~pi7430 & ~pi9040;
assign w59371 = ~w59369 & ~w59370;
assign w59372 = pi3865 & ~w59371;
assign w59373 = ~pi3865 & w59371;
assign w59374 = ~w59372 & ~w59373;
assign w59375 = w59340 & w59352;
assign w59376 = (~w59346 & w59375) | (~w59346 & w63475) | (w59375 & w63475);
assign w59377 = w59333 & ~w59339;
assign w59378 = w59352 & w59377;
assign w59379 = ~w59376 & ~w59378;
assign w59380 = (w59333 & w59376) | (w59333 & w64220) | (w59376 & w64220);
assign w59381 = ~w59346 & ~w59359;
assign w59382 = ~w59333 & ~w59352;
assign w59383 = ~w59376 & ~w59382;
assign w59384 = ~w59381 & ~w59383;
assign w59385 = ~w59368 & w59374;
assign w59386 = ~w59380 & w59385;
assign w59387 = ~w59384 & w59386;
assign w59388 = w59346 & w59352;
assign w59389 = ~w59353 & ~w59388;
assign w59390 = ~w59333 & w59389;
assign w59391 = w59389 & w64221;
assign w59392 = w59333 & w59346;
assign w59393 = w59339 & ~w59359;
assign w59394 = w59392 & w59393;
assign w59395 = w59333 & w59360;
assign w59396 = ~w59365 & ~w59395;
assign w59397 = ~w59333 & ~w59346;
assign w59398 = w59389 & ~w59397;
assign w59399 = ~w59339 & ~w59398;
assign w59400 = ~w59396 & w59399;
assign w59401 = w59346 & w59363;
assign w59402 = w59352 & w59359;
assign w59403 = ~w59392 & ~w59397;
assign w59404 = w59339 & w59402;
assign w59405 = w59403 & w59404;
assign w59406 = ~w59401 & ~w59405;
assign w59407 = ~w59374 & ~w59394;
assign w59408 = ~w59391 & w59407;
assign w59409 = w59406 & w59408;
assign w59410 = ~w59400 & w59409;
assign w59411 = ~w59387 & ~w59410;
assign w59412 = ~w59389 & ~w59392;
assign w59413 = ~w59339 & w59412;
assign w59414 = ~w59359 & ~w59388;
assign w59415 = ~w59402 & ~w59403;
assign w59416 = ~w59414 & w59415;
assign w59417 = ~w59413 & ~w59416;
assign w59418 = w59346 & w59359;
assign w59419 = ~w59381 & ~w59418;
assign w59420 = ~w59339 & ~w59419;
assign w59421 = w59417 & w59420;
assign w59422 = ~w59361 & ~w59364;
assign w59423 = ~w59421 & w59422;
assign w59424 = ~w59411 & w59423;
assign w59425 = ~pi5238 & ~w59424;
assign w59426 = pi5238 & w59424;
assign w59427 = ~w59425 & ~w59426;
assign w59428 = ~pi7446 & pi9040;
assign w59429 = ~pi7415 & ~pi9040;
assign w59430 = ~w59428 & ~w59429;
assign w59431 = pi3943 & ~w59430;
assign w59432 = ~pi3943 & w59430;
assign w59433 = ~w59431 & ~w59432;
assign w59434 = ~pi7397 & pi9040;
assign w59435 = ~pi7537 & ~pi9040;
assign w59436 = ~w59434 & ~w59435;
assign w59437 = pi3939 & ~w59436;
assign w59438 = ~pi3939 & w59436;
assign w59439 = ~w59437 & ~w59438;
assign w59440 = ~w59433 & w59439;
assign w59441 = ~pi7519 & pi9040;
assign w59442 = ~pi7528 & ~pi9040;
assign w59443 = ~w59441 & ~w59442;
assign w59444 = pi3840 & ~w59443;
assign w59445 = ~pi3840 & w59443;
assign w59446 = ~w59444 & ~w59445;
assign w59447 = ~pi7460 & pi9040;
assign w59448 = ~pi7456 & ~pi9040;
assign w59449 = ~w59447 & ~w59448;
assign w59450 = pi3915 & ~w59449;
assign w59451 = ~pi3915 & w59449;
assign w59452 = ~w59450 & ~w59451;
assign w59453 = ~w59446 & ~w59452;
assign w59454 = ~pi7537 & pi9040;
assign w59455 = ~pi7522 & ~pi9040;
assign w59456 = ~w59454 & ~w59455;
assign w59457 = pi3960 & ~w59456;
assign w59458 = ~pi3960 & w59456;
assign w59459 = ~w59457 & ~w59458;
assign w59460 = ~w59433 & ~w59459;
assign w59461 = w59453 & w59460;
assign w59462 = w59446 & ~w59452;
assign w59463 = w59459 & w59462;
assign w59464 = ~w59461 & ~w59463;
assign w59465 = w59440 & ~w59464;
assign w59466 = ~w59433 & w59452;
assign w59467 = (~w59439 & w59463) | (~w59439 & w64222) | (w59463 & w64222);
assign w59468 = w59433 & w59453;
assign w59469 = w59453 & w64223;
assign w59470 = ~pi7439 & pi9040;
assign w59471 = ~pi7397 & ~pi9040;
assign w59472 = ~w59470 & ~w59471;
assign w59473 = pi3870 & ~w59472;
assign w59474 = ~pi3870 & w59472;
assign w59475 = ~w59473 & ~w59474;
assign w59476 = ~w59469 & ~w59475;
assign w59477 = w59446 & w59452;
assign w59478 = w59459 & ~w59477;
assign w59479 = ~w59446 & w59452;
assign w59480 = ~w59459 & ~w59479;
assign w59481 = ~w59478 & ~w59480;
assign w59482 = w59433 & w59481;
assign w59483 = w59433 & ~w59459;
assign w59484 = w59462 & w59483;
assign w59485 = (~w59484 & ~w59481) | (~w59484 & w64224) | (~w59481 & w64224);
assign w59486 = w59433 & w59439;
assign w59487 = w59462 & w59486;
assign w59488 = w59433 & ~w59446;
assign w59489 = ~w59433 & w59446;
assign w59490 = ~w59488 & ~w59489;
assign w59491 = ~w59439 & ~w59459;
assign w59492 = ~w59490 & w59491;
assign w59493 = ~w59487 & ~w59492;
assign w59494 = ~w59485 & ~w59493;
assign w59495 = ~w59459 & w59489;
assign w59496 = w59489 & w59551;
assign w59497 = w59439 & w59459;
assign w59498 = w59488 & w59497;
assign w59499 = w59477 & w59486;
assign w59500 = w59440 & w59453;
assign w59501 = ~w59461 & ~w59498;
assign w59502 = ~w59499 & ~w59500;
assign w59503 = w59501 & w59502;
assign w59504 = ~w59496 & w59503;
assign w59505 = ~w59467 & w59476;
assign w59506 = w59504 & w59505;
assign w59507 = ~w59494 & w59506;
assign w59508 = ~w59433 & ~w59439;
assign w59509 = w59453 & w59508;
assign w59510 = w59459 & w59509;
assign w59511 = w59440 & w59479;
assign w59512 = w59475 & ~w59511;
assign w59513 = ~w59510 & w59512;
assign w59514 = ~w59482 & w59513;
assign w59515 = w59493 & w59514;
assign w59516 = (~w59465 & w59507) | (~w59465 & w64225) | (w59507 & w64225);
assign w59517 = pi5216 & ~w59516;
assign w59518 = ~pi5216 & w59516;
assign w59519 = ~w59517 & ~w59518;
assign w59520 = w59011 & w59012;
assign w59521 = w59022 & w59027;
assign w59522 = ~w58989 & w59018;
assign w59523 = (w58982 & w59521) | (w58982 & w64226) | (w59521 & w64226);
assign w59524 = ~w59023 & w59049;
assign w59525 = ~w59523 & w59524;
assign w59526 = ~w59520 & w59525;
assign w59527 = w59010 & ~w59526;
assign w59528 = ~w59010 & ~w59013;
assign w59529 = ~w59022 & w59026;
assign w59530 = w59528 & w59529;
assign w59531 = w58982 & w58995;
assign w59532 = w59024 & w59531;
assign w59533 = ~w59521 & w59528;
assign w59534 = w59010 & ~w59025;
assign w59535 = ~w59047 & w59534;
assign w59536 = ~w58982 & ~w59533;
assign w59537 = ~w59535 & w59536;
assign w59538 = w58982 & ~w59010;
assign w59539 = w59031 & w59538;
assign w59540 = w58989 & ~w59024;
assign w59541 = w59044 & w59540;
assign w59542 = ~w59532 & ~w59541;
assign w59543 = ~w59530 & w59542;
assign w59544 = ~w59537 & w59543;
assign w59545 = ~w59539 & w59544;
assign w59546 = (pi5191 & ~w59545) | (pi5191 & w64227) | (~w59545 & w64227);
assign w59547 = w59545 & w64228;
assign w59548 = ~w59546 & ~w59547;
assign w59549 = w59439 & w59452;
assign w59550 = w59475 & ~w59549;
assign w59551 = w59452 & ~w59459;
assign w59552 = w59488 & w59551;
assign w59553 = ~w59495 & ~w59552;
assign w59554 = ~w59550 & ~w59553;
assign w59555 = w59462 & ~w59483;
assign w59556 = ~w59552 & ~w59555;
assign w59557 = ~w59439 & ~w59556;
assign w59558 = ~w59459 & ~w59462;
assign w59559 = ~w59479 & ~w59558;
assign w59560 = w59433 & ~w59439;
assign w59561 = (w59560 & w59558) | (w59560 & w64229) | (w59558 & w64229);
assign w59562 = ~w59557 & ~w59561;
assign w59563 = w59480 & ~w59562;
assign w59564 = ~w59481 & w59508;
assign w59565 = w59486 & w59559;
assign w59566 = ~w59475 & ~w59564;
assign w59567 = ~w59565 & w59566;
assign w59568 = w59453 & w59483;
assign w59569 = w59433 & ~w59453;
assign w59570 = ~w59549 & ~w59569;
assign w59571 = w59478 & ~w59570;
assign w59572 = ~w59439 & ~w59483;
assign w59573 = w59481 & w59572;
assign w59574 = w59475 & ~w59500;
assign w59575 = ~w59568 & w59574;
assign w59576 = ~w59571 & w59575;
assign w59577 = ~w59573 & w59576;
assign w59578 = ~w59567 & ~w59577;
assign w59579 = ~w59554 & ~w59563;
assign w59580 = ~w59578 & w59579;
assign w59581 = pi5350 & ~w59580;
assign w59582 = ~pi5350 & w59580;
assign w59583 = ~w59581 & ~w59582;
assign w59584 = ~pi7461 & pi9040;
assign w59585 = ~pi7429 & ~pi9040;
assign w59586 = ~w59584 & ~w59585;
assign w59587 = pi3912 & ~w59586;
assign w59588 = ~pi3912 & w59586;
assign w59589 = ~w59587 & ~w59588;
assign w59590 = ~pi7425 & pi9040;
assign w59591 = ~pi7376 & ~pi9040;
assign w59592 = ~w59590 & ~w59591;
assign w59593 = pi3915 & ~w59592;
assign w59594 = ~pi3915 & w59592;
assign w59595 = ~w59593 & ~w59594;
assign w59596 = ~w59589 & w59595;
assign w59597 = ~pi7411 & pi9040;
assign w59598 = ~pi7453 & ~pi9040;
assign w59599 = ~w59597 & ~w59598;
assign w59600 = pi3870 & ~w59599;
assign w59601 = ~pi3870 & w59599;
assign w59602 = ~w59600 & ~w59601;
assign w59603 = ~pi7376 & pi9040;
assign w59604 = ~pi7589 & ~pi9040;
assign w59605 = ~w59603 & ~w59604;
assign w59606 = pi3972 & ~w59605;
assign w59607 = ~pi3972 & w59605;
assign w59608 = ~w59606 & ~w59607;
assign w59609 = w59602 & w59608;
assign w59610 = w59596 & w59609;
assign w59611 = ~w59589 & ~w59595;
assign w59612 = ~w59602 & w59608;
assign w59613 = w59611 & w59612;
assign w59614 = ~w59610 & ~w59613;
assign w59615 = ~pi7568 & pi9040;
assign w59616 = ~pi7462 & ~pi9040;
assign w59617 = ~w59615 & ~w59616;
assign w59618 = pi3861 & ~w59617;
assign w59619 = ~pi3861 & w59617;
assign w59620 = ~w59618 & ~w59619;
assign w59621 = ~w59614 & w59620;
assign w59622 = w59595 & w59602;
assign w59623 = w59589 & w59620;
assign w59624 = w59622 & w59623;
assign w59625 = w59595 & ~w59608;
assign w59626 = w59589 & w59625;
assign w59627 = w59589 & ~w59595;
assign w59628 = ~w59596 & ~w59627;
assign w59629 = w59612 & ~w59628;
assign w59630 = ~w59595 & ~w59602;
assign w59631 = ~w59611 & ~w59630;
assign w59632 = ~w59609 & ~w59631;
assign w59633 = ~w59629 & ~w59632;
assign w59634 = w59620 & ~w59633;
assign w59635 = w59602 & w59627;
assign w59636 = ~w59602 & w59625;
assign w59637 = ~w59635 & ~w59636;
assign w59638 = ~w59620 & ~w59637;
assign w59639 = ~w59610 & ~w59624;
assign w59640 = ~w59626 & w59639;
assign w59641 = ~w59638 & w59640;
assign w59642 = ~w59634 & w59641;
assign w59643 = ~pi7385 & pi9040;
assign w59644 = ~pi7427 & ~pi9040;
assign w59645 = ~w59643 & ~w59644;
assign w59646 = pi3866 & ~w59645;
assign w59647 = ~pi3866 & w59645;
assign w59648 = ~w59646 & ~w59647;
assign w59649 = w59609 & ~w59620;
assign w59650 = w59589 & w59608;
assign w59651 = w59589 & ~w59602;
assign w59652 = w59602 & ~w59627;
assign w59653 = ~w59651 & ~w59652;
assign w59654 = (~w59650 & w59652) | (~w59650 & w64230) | (w59652 & w64230);
assign w59655 = (w59620 & ~w59652) | (w59620 & w64231) | (~w59652 & w64231);
assign w59656 = w59654 & w59655;
assign w59657 = ~w59649 & ~w59656;
assign w59658 = ~w59595 & ~w59657;
assign w59659 = w59602 & w59626;
assign w59660 = ~w59612 & ~w59620;
assign w59661 = ~w59595 & ~w59660;
assign w59662 = ~w59648 & ~w59661;
assign w59663 = (w59642 & w64232) | (w59642 & w64233) | (w64232 & w64233);
assign w59664 = ~w59621 & ~w59659;
assign w59665 = (w59664 & w59642) | (w59664 & w63477) | (w59642 & w63477);
assign w59666 = ~w59658 & w59665;
assign w59667 = w59666 & w64234;
assign w59668 = (pi5098 & ~w59666) | (pi5098 & w64235) | (~w59666 & w64235);
assign w59669 = ~w59667 & ~w59668;
assign w59670 = w59252 & w59308;
assign w59671 = ~w59260 & w59274;
assign w59672 = w59251 & ~w59671;
assign w59673 = ~w59299 & ~w59671;
assign w59674 = ~w59672 & ~w59673;
assign w59675 = w59309 & ~w59674;
assign w59676 = (~w59295 & w59674) | (~w59295 & w64236) | (w59674 & w64236);
assign w59677 = ~w59287 & ~w59315;
assign w59678 = w59275 & ~w59677;
assign w59679 = ~w59253 & ~w59306;
assign w59680 = w59300 & w59672;
assign w59681 = ~w59252 & ~w59679;
assign w59682 = ~w59680 & w59681;
assign w59683 = ~w59670 & ~w59678;
assign w59684 = ~w59682 & w59683;
assign w59685 = w59676 & w59684;
assign w59686 = w59251 & w59283;
assign w59687 = ~w59280 & ~w59307;
assign w59688 = w59267 & ~w59687;
assign w59689 = w59275 & ~w59298;
assign w59690 = w59677 & w59689;
assign w59691 = w59295 & ~w59313;
assign w59692 = ~w59690 & w59691;
assign w59693 = ~w59688 & w59692;
assign w59694 = ~w59686 & w59693;
assign w59695 = ~w59685 & ~w59694;
assign w59696 = ~pi5183 & w59695;
assign w59697 = pi5183 & ~w59695;
assign w59698 = ~w59696 & ~w59697;
assign w59699 = ~w59045 & ~w59051;
assign w59700 = w59012 & ~w59699;
assign w59701 = ~w59538 & ~w59700;
assign w59702 = w59540 & ~w59701;
assign w59703 = w59002 & ~w59010;
assign w59704 = w58982 & w58996;
assign w59705 = ~w59047 & ~w59704;
assign w59706 = w59703 & ~w59705;
assign w59707 = ~w58976 & w59010;
assign w59708 = ~w59003 & ~w59522;
assign w59709 = ~w59538 & ~w59707;
assign w59710 = ~w59708 & w59709;
assign w59711 = w59020 & w59531;
assign w59712 = ~w59044 & ~w59711;
assign w59713 = w59002 & ~w59712;
assign w59714 = w59040 & ~w59699;
assign w59715 = ~w59520 & ~w59714;
assign w59716 = ~w59713 & w59715;
assign w59717 = w59010 & ~w59716;
assign w59718 = ~w59706 & ~w59710;
assign w59719 = ~w59056 & w59718;
assign w59720 = ~w59702 & w59719;
assign w59721 = ~w59717 & w59720;
assign w59722 = pi5428 & ~w59721;
assign w59723 = ~pi5428 & w59721;
assign w59724 = ~w59722 & ~w59723;
assign w59725 = w58983 & ~w59028;
assign w59726 = ~w59019 & ~w59057;
assign w59727 = ~w59711 & w59726;
assign w59728 = ~w59725 & w59727;
assign w59729 = w59010 & ~w59728;
assign w59730 = w58996 & w59703;
assign w59731 = ~w59048 & ~w59050;
assign w59732 = ~w59012 & w59022;
assign w59733 = w59731 & w59732;
assign w59734 = ~w59530 & ~w59730;
assign w59735 = (~w58982 & ~w59734) | (~w58982 & w64237) | (~w59734 & w64237);
assign w59736 = w58982 & ~w59731;
assign w59737 = ~w59541 & ~w59700;
assign w59738 = ~w59736 & w59737;
assign w59739 = ~w59010 & ~w59738;
assign w59740 = w58976 & ~w59052;
assign w59741 = ~w59525 & w59740;
assign w59742 = ~w59729 & ~w59735;
assign w59743 = ~w59739 & ~w59741;
assign w59744 = w59742 & w59743;
assign w59745 = pi5426 & w59744;
assign w59746 = ~pi5426 & ~w59744;
assign w59747 = ~w59745 & ~w59746;
assign w59748 = w59439 & w59568;
assign w59749 = ~w59466 & ~w59495;
assign w59750 = ~w59439 & w59446;
assign w59751 = ~w59749 & w59750;
assign w59752 = ~w59465 & ~w59748;
assign w59753 = w59752 & w64238;
assign w59754 = ~w59475 & ~w59753;
assign w59755 = w59452 & w59459;
assign w59756 = w59490 & w59755;
assign w59757 = ~w59468 & ~w59496;
assign w59758 = ~w59756 & w59757;
assign w59759 = w59497 & ~w59758;
assign w59760 = (w59439 & w59495) | (w59439 & w64239) | (w59495 & w64239);
assign w59761 = ~w59561 & ~w59760;
assign w59762 = w59475 & ~w59761;
assign w59763 = (~w59439 & ~w59490) | (~w59439 & w64240) | (~w59490 & w64240);
assign w59764 = ~w59461 & w59763;
assign w59765 = ~w59475 & ~w59764;
assign w59766 = w59478 & w59490;
assign w59767 = ~w59765 & w59766;
assign w59768 = ~w59759 & ~w59762;
assign w59769 = ~w59767 & w59768;
assign w59770 = ~w59754 & w59769;
assign w59771 = pi5427 & w59770;
assign w59772 = ~pi5427 & ~w59770;
assign w59773 = ~w59771 & ~w59772;
assign w59774 = w59375 & w59419;
assign w59775 = w59389 & w59403;
assign w59776 = w59359 & w59775;
assign w59777 = w59333 & ~w59389;
assign w59778 = w59339 & w59777;
assign w59779 = ~w59339 & ~w59366;
assign w59780 = ~w59403 & w59779;
assign w59781 = ~w59374 & ~w59776;
assign w59782 = ~w59778 & ~w59780;
assign w59783 = w59781 & w59782;
assign w59784 = w59381 & w59398;
assign w59785 = ~w59339 & ~w59359;
assign w59786 = w59382 & w59785;
assign w59787 = ~w59377 & ~w59388;
assign w59788 = w59359 & ~w59787;
assign w59789 = w59340 & ~w59362;
assign w59790 = ~w59786 & ~w59789;
assign w59791 = ~w59788 & w59790;
assign w59792 = w59339 & w59401;
assign w59793 = w59374 & ~w59784;
assign w59794 = w59791 & ~w59792;
assign w59795 = w59793 & w59794;
assign w59796 = ~w59783 & ~w59795;
assign w59797 = ~w59774 & ~w59796;
assign w59798 = ~pi5499 & w59797;
assign w59799 = pi5499 & ~w59797;
assign w59800 = ~w59798 & ~w59799;
assign w59801 = w59276 & w59312;
assign w59802 = ~w59310 & w59315;
assign w59803 = ~w59801 & ~w59802;
assign w59804 = w59310 & ~w59672;
assign w59805 = w59679 & w59804;
assign w59806 = (w59267 & ~w59804) | (w59267 & w64241) | (~w59804 & w64241);
assign w59807 = ~w59298 & ~w59299;
assign w59808 = ~w59254 & ~w59807;
assign w59809 = ~w59245 & w59315;
assign w59810 = ~w59267 & ~w59809;
assign w59811 = ~w59311 & ~w59808;
assign w59812 = w59810 & w59811;
assign w59813 = (w59803 & w59812) | (w59803 & w64242) | (w59812 & w64242);
assign w59814 = w59295 & ~w59813;
assign w59815 = ~w59274 & w59281;
assign w59816 = ~w59295 & ~w59802;
assign w59817 = ~w59804 & w59816;
assign w59818 = w59267 & ~w59815;
assign w59819 = ~w59817 & w59818;
assign w59820 = (~w59295 & w59805) | (~w59295 & w64243) | (w59805 & w64243);
assign w59821 = ~w59267 & w59803;
assign w59822 = ~w59820 & w59821;
assign w59823 = ~w59819 & ~w59822;
assign w59824 = ~w59814 & ~w59823;
assign w59825 = ~pi5349 & w59824;
assign w59826 = pi5349 & ~w59824;
assign w59827 = ~w59825 & ~w59826;
assign w59828 = w59439 & ~w59484;
assign w59829 = ~w59764 & ~w59828;
assign w59830 = ~w59480 & ~w59509;
assign w59831 = w59490 & ~w59830;
assign w59832 = w59440 & w59446;
assign w59833 = ~w59551 & w59832;
assign w59834 = w59439 & ~w59446;
assign w59835 = ~w59750 & ~w59834;
assign w59836 = w59551 & ~w59835;
assign w59837 = ~w59833 & ~w59836;
assign w59838 = w59476 & w59837;
assign w59839 = ~w59831 & w59838;
assign w59840 = ~w59758 & ~w59763;
assign w59841 = w59475 & ~w59557;
assign w59842 = ~w59840 & w59841;
assign w59843 = ~w59839 & ~w59842;
assign w59844 = ~w59498 & ~w59829;
assign w59845 = ~w59843 & w59844;
assign w59846 = pi5352 & ~w59845;
assign w59847 = ~pi5352 & w59845;
assign w59848 = ~w59846 & ~w59847;
assign w59849 = w59182 & w59201;
assign w59850 = w59160 & ~w59181;
assign w59851 = w59173 & w59850;
assign w59852 = ~w59849 & ~w59851;
assign w59853 = w59166 & ~w59852;
assign w59854 = ~w59181 & w59188;
assign w59855 = w59167 & w59854;
assign w59856 = w59209 & w64244;
assign w59857 = ~w59855 & ~w59856;
assign w59858 = w59166 & w59181;
assign w59859 = w59211 & w59858;
assign w59860 = ~w59198 & w59217;
assign w59861 = ~w59181 & w59860;
assign w59862 = ~w59175 & ~w59213;
assign w59863 = ~w59200 & w59862;
assign w59864 = ~w59196 & ~w59863;
assign w59865 = w59857 & ~w59859;
assign w59866 = ~w59861 & w59865;
assign w59867 = w59864 & w59866;
assign w59868 = ~w59173 & ~w59858;
assign w59869 = ~w59857 & w59868;
assign w59870 = w59213 & ~w59217;
assign w59871 = w59160 & w59166;
assign w59872 = ~w59182 & w59871;
assign w59873 = w59167 & w59197;
assign w59874 = ~w59166 & w59181;
assign w59875 = ~w59216 & w59874;
assign w59876 = ~w59199 & w59875;
assign w59877 = w59196 & ~w59872;
assign w59878 = ~w59873 & w59877;
assign w59879 = ~w59870 & ~w59876;
assign w59880 = w59878 & w59879;
assign w59881 = ~w59869 & w59880;
assign w59882 = ~w59867 & ~w59881;
assign w59883 = ~w59853 & ~w59882;
assign w59884 = ~pi5432 & w59883;
assign w59885 = pi5432 & ~w59883;
assign w59886 = ~w59884 & ~w59885;
assign w59887 = ~w59630 & ~w59650;
assign w59888 = (w59620 & w59887) | (w59620 & w63339) | (w59887 & w63339);
assign w59889 = ~w59636 & w59888;
assign w59890 = ~w59589 & ~w59622;
assign w59891 = w59888 & w63478;
assign w59892 = w59629 & w59891;
assign w59893 = (~w59648 & ~w59891) | (~w59648 & w64245) | (~w59891 & w64245);
assign w59894 = w59602 & ~w59608;
assign w59895 = ~w59620 & w59894;
assign w59896 = ~w59589 & ~w59608;
assign w59897 = w59630 & w59896;
assign w59898 = ~w59635 & ~w59897;
assign w59899 = w59620 & ~w59898;
assign w59900 = ~w59629 & ~w59895;
assign w59901 = ~w59899 & w59900;
assign w59902 = ~w59893 & ~w59901;
assign w59903 = (~w59642 & w64246) | (~w59642 & w64247) | (w64246 & w64247);
assign w59904 = ~w59620 & w59628;
assign w59905 = w59628 & w63479;
assign w59906 = ~w59633 & w63340;
assign w59907 = ~w59624 & ~w59636;
assign w59908 = w59614 & w59907;
assign w59909 = ~w59905 & w59908;
assign w59910 = ~w59906 & w59909;
assign w59911 = w59609 & w59611;
assign w59912 = w59648 & ~w59911;
assign w59913 = ~w59622 & ~w59896;
assign w59914 = w59660 & w59913;
assign w59915 = ~w59912 & w59914;
assign w59916 = (~w59915 & w59910) | (~w59915 & w63480) | (w59910 & w63480);
assign w59917 = ~w59902 & w59916;
assign w59918 = (pi5301 & ~w59917) | (pi5301 & w64248) | (~w59917 & w64248);
assign w59919 = w59917 & w64249;
assign w59920 = ~w59918 & ~w59919;
assign w59921 = w59279 & w59312;
assign w59922 = w59810 & ~w59921;
assign w59923 = ~w59278 & ~w59922;
assign w59924 = w59253 & w59308;
assign w59925 = ~w59317 & ~w59808;
assign w59926 = ~w59674 & ~w59925;
assign w59927 = (w59267 & w59925) | (w59267 & w63481) | (w59925 & w63481);
assign w59928 = ~w59296 & ~w59675;
assign w59929 = ~w59314 & w59928;
assign w59930 = w59295 & ~w59924;
assign w59931 = (w59930 & ~w59929) | (w59930 & w63482) | (~w59929 & w63482);
assign w59932 = w59300 & w59674;
assign w59933 = w59282 & ~w59686;
assign w59934 = ~w59926 & ~w59933;
assign w59935 = w59676 & ~w59932;
assign w59936 = ~w59934 & w59935;
assign w59937 = ~w59931 & ~w59936;
assign w59938 = ~w59937 & w64250;
assign w59939 = (pi5356 & w59937) | (pi5356 & w64251) | (w59937 & w64251);
assign w59940 = ~w59938 & ~w59939;
assign w59941 = w59374 & ~w59418;
assign w59942 = ~w59391 & w59941;
assign w59943 = ~w59379 & ~w59942;
assign w59944 = w59775 & w59785;
assign w59945 = ~w59374 & w59418;
assign w59946 = ~w59791 & w59945;
assign w59947 = ~w59390 & ~w59395;
assign w59948 = ~w59339 & ~w59947;
assign w59949 = ~w59389 & w59789;
assign w59950 = w59406 & ~w59949;
assign w59951 = ~w59948 & w59950;
assign w59952 = w59374 & ~w59951;
assign w59953 = ~w59364 & ~w59944;
assign w59954 = ~w59946 & w59953;
assign w59955 = ~w59943 & w59954;
assign w59956 = ~w59952 & w59955;
assign w59957 = pi5689 & ~w59956;
assign w59958 = ~pi5689 & w59956;
assign w59959 = ~w59957 & ~w59958;
assign w59960 = ~w59173 & ~w59854;
assign w59961 = w59217 & w59960;
assign w59962 = ~w59870 & ~w59961;
assign w59963 = ~w59196 & ~w59962;
assign w59964 = w59188 & w59851;
assign w59965 = ~w59229 & ~w59964;
assign w59966 = (~w59166 & w59963) | (~w59166 & w64252) | (w59963 & w64252);
assign w59967 = ~w59173 & w59854;
assign w59968 = ~w59863 & w64253;
assign w59969 = w59166 & ~w59209;
assign w59970 = w59230 & w59969;
assign w59971 = w59962 & w59970;
assign w59972 = ~w59202 & w59212;
assign w59973 = ~w59181 & w59201;
assign w59974 = w59181 & w59209;
assign w59975 = w59166 & ~w59973;
assign w59976 = ~w59974 & w59975;
assign w59977 = ~w59972 & ~w59976;
assign w59978 = w59160 & w59221;
assign w59979 = w59857 & ~w59978;
assign w59980 = w59965 & w59979;
assign w59981 = ~w59977 & w59980;
assign w59982 = w59196 & ~w59981;
assign w59983 = ~w59968 & ~w59971;
assign w59984 = ~w59966 & w59983;
assign w59985 = ~w59982 & w59984;
assign w59986 = pi5551 & ~w59985;
assign w59987 = ~pi5551 & w59985;
assign w59988 = ~w59986 & ~w59987;
assign w59989 = (~w59602 & ~w59628) | (~w59602 & w63483) | (~w59628 & w63483);
assign w59990 = (~w59608 & ~w59652) | (~w59608 & w63484) | (~w59652 & w63484);
assign w59991 = ~w59989 & w59990;
assign w59992 = w59609 & ~w59623;
assign w59993 = w59628 & w59992;
assign w59994 = ~w59991 & ~w59993;
assign w59995 = (w59648 & ~w59994) | (w59648 & w64254) | (~w59994 & w64254);
assign w59996 = ~w59660 & ~w59904;
assign w59997 = w59622 & w59896;
assign w59998 = ~w59613 & w59620;
assign w59999 = ~w59997 & w59998;
assign w60000 = w59996 & ~w59999;
assign w60001 = ~w59991 & w64255;
assign w60002 = ~w59996 & ~w60001;
assign w60003 = ~w59648 & ~w59889;
assign w60004 = ~w60002 & w60003;
assign w60005 = ~w59995 & ~w60000;
assign w60006 = ~w60004 & w60005;
assign w60007 = pi5300 & w60006;
assign w60008 = ~pi5300 & ~w60006;
assign w60009 = ~w60007 & ~w60008;
assign w60010 = ~w59390 & ~w59777;
assign w60011 = w59359 & ~w60010;
assign w60012 = w59393 & w59412;
assign w60013 = ~w59784 & ~w60012;
assign w60014 = ~w60011 & w60013;
assign w60015 = w59374 & ~w60014;
assign w60016 = w59339 & ~w59374;
assign w60017 = w59389 & w60016;
assign w60018 = ~w59784 & w60017;
assign w60019 = w59417 & ~w60018;
assign w60020 = w59374 & ~w59402;
assign w60021 = ~w59378 & w60020;
assign w60022 = ~w60019 & ~w60021;
assign w60023 = ~w60015 & ~w60022;
assign w60024 = pi5647 & w60023;
assign w60025 = ~pi5647 & ~w60023;
assign w60026 = ~w60024 & ~w60025;
assign w60027 = w59088 & w59095;
assign w60028 = w59103 & w59128;
assign w60029 = w59087 & w59141;
assign w60030 = ~w60028 & ~w60029;
assign w60031 = ~w59095 & w60030;
assign w60032 = w59072 & w59085;
assign w60033 = ~w59102 & w60032;
assign w60034 = w59095 & ~w60033;
assign w60035 = ~w59086 & w60034;
assign w60036 = ~w60031 & ~w60035;
assign w60037 = ~w59085 & w59095;
assign w60038 = w59102 & w59104;
assign w60039 = ~w60037 & w60038;
assign w60040 = ~w59089 & ~w59102;
assign w60041 = ~w59116 & ~w59118;
assign w60042 = ~w60039 & w60041;
assign w60043 = ~w60040 & w60042;
assign w60044 = ~w60036 & w60043;
assign w60045 = w59078 & w60032;
assign w60046 = ~w59072 & w59123;
assign w60047 = ~w59140 & ~w60045;
assign w60048 = ~w60046 & w60047;
assign w60049 = w59095 & ~w60048;
assign w60050 = ~w59123 & w59133;
assign w60051 = w59145 & w60050;
assign w60052 = ~w59087 & ~w60045;
assign w60053 = ~w59145 & ~w60052;
assign w60054 = w59116 & ~w60051;
assign w60055 = ~w60053 & w60054;
assign w60056 = ~w60049 & w60055;
assign w60057 = ~w60044 & ~w60056;
assign w60058 = w59104 & w59125;
assign w60059 = ~w60027 & ~w60058;
assign w60060 = ~w60057 & w60059;
assign w60061 = pi5467 & ~w60060;
assign w60062 = ~pi5467 & w60060;
assign w60063 = ~w60061 & ~w60062;
assign w60064 = w59127 & w60037;
assign w60065 = w59142 & w64256;
assign w60066 = w59133 & w59141;
assign w60067 = w60030 & ~w60066;
assign w60068 = ~w60065 & w60067;
assign w60069 = ~w59116 & ~w60068;
assign w60070 = ~w59119 & ~w59140;
assign w60071 = ~w59136 & w60070;
assign w60072 = ~w59088 & ~w60046;
assign w60073 = ~w60033 & w60072;
assign w60074 = ~w59095 & ~w60073;
assign w60075 = ~w59106 & ~w60032;
assign w60076 = w60034 & ~w60075;
assign w60077 = w60071 & ~w60076;
assign w60078 = ~w60074 & w60077;
assign w60079 = w59116 & ~w60078;
assign w60080 = ~w59095 & w59144;
assign w60081 = ~w59134 & ~w60064;
assign w60082 = ~w60080 & w60081;
assign w60083 = ~w60069 & w60082;
assign w60084 = ~w60079 & w60083;
assign w60085 = pi5497 & ~w60084;
assign w60086 = ~pi5497 & w60084;
assign w60087 = ~w60085 & ~w60086;
assign w60088 = ~pi7428 & pi9040;
assign w60089 = ~pi7401 & ~pi9040;
assign w60090 = ~w60088 & ~w60089;
assign w60091 = pi3930 & ~w60090;
assign w60092 = ~pi3930 & w60090;
assign w60093 = ~w60091 & ~w60092;
assign w60094 = ~pi7379 & pi9040;
assign w60095 = ~pi7428 & ~pi9040;
assign w60096 = ~w60094 & ~w60095;
assign w60097 = pi3852 & ~w60096;
assign w60098 = ~pi3852 & w60096;
assign w60099 = ~w60097 & ~w60098;
assign w60100 = ~w60093 & ~w60099;
assign w60101 = ~pi7430 & pi9040;
assign w60102 = ~pi7466 & ~pi9040;
assign w60103 = ~w60101 & ~w60102;
assign w60104 = pi3943 & ~w60103;
assign w60105 = ~pi3943 & w60103;
assign w60106 = ~w60104 & ~w60105;
assign w60107 = ~pi7528 & pi9040;
assign w60108 = ~pi7460 & ~pi9040;
assign w60109 = ~w60107 & ~w60108;
assign w60110 = pi3940 & ~w60109;
assign w60111 = ~pi3940 & w60109;
assign w60112 = ~w60110 & ~w60111;
assign w60113 = ~w60106 & w60112;
assign w60114 = w60100 & w60113;
assign w60115 = ~pi7366 & pi9040;
assign w60116 = ~pi7436 & ~pi9040;
assign w60117 = ~w60115 & ~w60116;
assign w60118 = pi3846 & ~w60117;
assign w60119 = ~pi3846 & w60117;
assign w60120 = ~w60118 & ~w60119;
assign w60121 = w60093 & w60120;
assign w60122 = ~w60099 & ~w60112;
assign w60123 = w60121 & w60122;
assign w60124 = ~w60114 & ~w60123;
assign w60125 = w60106 & ~w60112;
assign w60126 = w60093 & w60099;
assign w60127 = ~w60100 & ~w60126;
assign w60128 = ~w60120 & w60125;
assign w60129 = ~w60127 & w60128;
assign w60130 = w60124 & ~w60129;
assign w60131 = w60113 & w60126;
assign w60132 = ~w60113 & ~w60125;
assign w60133 = w60127 & w60132;
assign w60134 = ~w60131 & ~w60133;
assign w60135 = w60130 & w60134;
assign w60136 = ~pi7401 & pi9040;
assign w60137 = ~pi7396 & ~pi9040;
assign w60138 = ~w60136 & ~w60137;
assign w60139 = pi3840 & ~w60138;
assign w60140 = ~pi3840 & w60138;
assign w60141 = ~w60139 & ~w60140;
assign w60142 = ~w60135 & ~w60141;
assign w60143 = ~w60106 & ~w60112;
assign w60144 = ~w60093 & w60106;
assign w60145 = w60093 & ~w60106;
assign w60146 = w60099 & ~w60112;
assign w60147 = ~w60145 & ~w60146;
assign w60148 = ~w60144 & w60147;
assign w60149 = w60120 & w60148;
assign w60150 = w60126 & w60141;
assign w60151 = ~w60149 & ~w60150;
assign w60152 = w60143 & ~w60151;
assign w60153 = w60141 & ~w60143;
assign w60154 = w60099 & w60144;
assign w60155 = ~w60153 & ~w60154;
assign w60156 = ~w60120 & ~w60148;
assign w60157 = ~w60149 & ~w60155;
assign w60158 = ~w60156 & w60157;
assign w60159 = ~w60142 & ~w60152;
assign w60160 = ~w60158 & w60159;
assign w60161 = ~pi5433 & ~w60160;
assign w60162 = pi5433 & w60160;
assign w60163 = ~w60161 & ~w60162;
assign w60164 = w59198 & w59858;
assign w60165 = ~w59222 & ~w59231;
assign w60166 = ~w59219 & ~w60165;
assign w60167 = ~w59208 & ~w59871;
assign w60168 = w59198 & ~w60167;
assign w60169 = ~w59208 & ~w59850;
assign w60170 = w59868 & w60169;
assign w60171 = ~w59973 & ~w60168;
assign w60172 = ~w60170 & w60171;
assign w60173 = w59230 & w60172;
assign w60174 = w59166 & w59860;
assign w60175 = ~w59201 & ~w59854;
assign w60176 = w59174 & ~w60175;
assign w60177 = w59196 & ~w59849;
assign w60178 = ~w60176 & w60177;
assign w60179 = ~w60174 & w60178;
assign w60180 = ~w60173 & ~w60179;
assign w60181 = ~w60164 & ~w60166;
assign w60182 = ~w60180 & w60181;
assign w60183 = pi5603 & ~w60182;
assign w60184 = ~pi5603 & w60182;
assign w60185 = ~w60183 & ~w60184;
assign w60186 = w59108 & ~w60071;
assign w60187 = w59102 & w59108;
assign w60188 = ~w59108 & ~w59141;
assign w60189 = ~w59085 & ~w60187;
assign w60190 = ~w60188 & w60189;
assign w60191 = w59103 & w59117;
assign w60192 = ~w59078 & w60032;
assign w60193 = w59116 & ~w60191;
assign w60194 = ~w60192 & w60193;
assign w60195 = ~w60190 & w60194;
assign w60196 = (w59095 & ~w60075) | (w59095 & w64257) | (~w60075 & w64257);
assign w60197 = ~w59102 & w59104;
assign w60198 = (~w59085 & w60197) | (~w59085 & w64258) | (w60197 & w64258);
assign w60199 = ~w59116 & ~w60198;
assign w60200 = ~w60196 & w60199;
assign w60201 = ~w60195 & ~w60200;
assign w60202 = w59143 & ~w60072;
assign w60203 = ~w59086 & ~w60191;
assign w60204 = ~w60202 & w60203;
assign w60205 = ~w59095 & ~w60204;
assign w60206 = ~w60186 & ~w60201;
assign w60207 = ~w60205 & w60206;
assign w60208 = ~pi5691 & w60207;
assign w60209 = pi5691 & ~w60207;
assign w60210 = ~w60208 & ~w60209;
assign w60211 = ~w60093 & ~w60112;
assign w60212 = w60093 & w60112;
assign w60213 = w60106 & w60212;
assign w60214 = w60150 & ~w60213;
assign w60215 = w60099 & w60112;
assign w60216 = ~w60145 & ~w60215;
assign w60217 = ~w60120 & ~w60141;
assign w60218 = w60216 & w60217;
assign w60219 = ~w60214 & ~w60218;
assign w60220 = ~w60211 & ~w60219;
assign w60221 = w60099 & ~w60120;
assign w60222 = ~w60121 & w60143;
assign w60223 = ~w60099 & w60222;
assign w60224 = ~w60221 & ~w60223;
assign w60225 = ~w60216 & ~w60224;
assign w60226 = w60120 & ~w60213;
assign w60227 = w60099 & w60145;
assign w60228 = ~w60216 & ~w60227;
assign w60229 = w60226 & ~w60228;
assign w60230 = ~w60100 & w60132;
assign w60231 = ~w60132 & w60147;
assign w60232 = ~w60230 & ~w60231;
assign w60233 = w60229 & ~w60232;
assign w60234 = ~w60225 & ~w60233;
assign w60235 = w60141 & ~w60234;
assign w60236 = w60145 & w60221;
assign w60237 = w60141 & ~w60144;
assign w60238 = w60120 & ~w60237;
assign w60239 = w60228 & w60238;
assign w60240 = ~w60093 & ~w60141;
assign w60241 = w60232 & w60240;
assign w60242 = ~w60236 & ~w60239;
assign w60243 = ~w60220 & w60242;
assign w60244 = ~w60241 & w60243;
assign w60245 = ~w60235 & w60244;
assign w60246 = pi5646 & ~w60245;
assign w60247 = ~pi5646 & w60245;
assign w60248 = ~w60246 & ~w60247;
assign w60249 = w60124 & ~w60213;
assign w60250 = ~w60234 & ~w60249;
assign w60251 = (~w60120 & ~w60132) | (~w60120 & w64259) | (~w60132 & w64259);
assign w60252 = w60100 & ~w60125;
assign w60253 = ~w60093 & w60112;
assign w60254 = w60099 & ~w60143;
assign w60255 = ~w60253 & w60254;
assign w60256 = w60120 & ~w60252;
assign w60257 = ~w60255 & w60256;
assign w60258 = ~w60251 & ~w60257;
assign w60259 = (w60141 & w60130) | (w60141 & w64260) | (w60130 & w64260);
assign w60260 = ~w60258 & w60259;
assign w60261 = ~w60231 & w60251;
assign w60262 = ~w60212 & w60257;
assign w60263 = ~w60106 & ~w60212;
assign w60264 = w60215 & w60263;
assign w60265 = ~w60141 & ~w60264;
assign w60266 = ~w60261 & w60265;
assign w60267 = ~w60262 & w60266;
assign w60268 = ~w60260 & ~w60267;
assign w60269 = ~w60250 & ~w60268;
assign w60270 = ~pi5599 & w60269;
assign w60271 = pi5599 & ~w60269;
assign w60272 = ~w60270 & ~w60271;
assign w60273 = ~w59620 & ~w59654;
assign w60274 = ~w59612 & ~w59650;
assign w60275 = ~w59595 & ~w60274;
assign w60276 = ~w59648 & ~w60275;
assign w60277 = ~w59656 & w60276;
assign w60278 = ~w60273 & w60277;
assign w60279 = w59653 & w59888;
assign w60280 = ~w59659 & w59912;
assign w60281 = ~w59905 & w60280;
assign w60282 = ~w60279 & w60281;
assign w60283 = ~w60278 & ~w60282;
assign w60284 = (~w59997 & w59898) | (~w59997 & w64261) | (w59898 & w64261);
assign w60285 = ~w59620 & ~w60284;
assign w60286 = ~w59906 & ~w60285;
assign w60287 = ~w59892 & w60286;
assign w60288 = ~w60283 & w60287;
assign w60289 = pi5531 & w60288;
assign w60290 = ~pi5531 & ~w60288;
assign w60291 = ~w60289 & ~w60290;
assign w60292 = ~w60134 & w60229;
assign w60293 = ~w60211 & ~w60212;
assign w60294 = w60106 & ~w60293;
assign w60295 = ~w60293 & w64262;
assign w60296 = ~w60211 & ~w60263;
assign w60297 = w60226 & w60296;
assign w60298 = ~w60223 & ~w60295;
assign w60299 = ~w60297 & w60298;
assign w60300 = ~w60141 & ~w60299;
assign w60301 = w60125 & w60126;
assign w60302 = ~w60120 & ~w60254;
assign w60303 = ~w60301 & ~w60302;
assign w60304 = ~w60099 & ~w60113;
assign w60305 = ~w60303 & ~w60304;
assign w60306 = ~w60222 & w60263;
assign w60307 = ~w60294 & ~w60306;
assign w60308 = ~w60099 & ~w60307;
assign w60309 = ~w60305 & ~w60308;
assign w60310 = w60141 & ~w60309;
assign w60311 = w60221 & w60253;
assign w60312 = ~w60292 & ~w60311;
assign w60313 = ~w60300 & w60312;
assign w60314 = ~w60310 & w60313;
assign w60315 = pi5523 & ~w60314;
assign w60316 = ~pi5523 & w60314;
assign w60317 = ~w60315 & ~w60316;
assign w60318 = ~pi7745 & pi9040;
assign w60319 = ~pi7653 & ~pi9040;
assign w60320 = ~w60318 & ~w60319;
assign w60321 = pi5512 & ~w60320;
assign w60322 = ~pi5512 & w60320;
assign w60323 = ~w60321 & ~w60322;
assign w60324 = ~pi7648 & pi9040;
assign w60325 = ~pi7675 & ~pi9040;
assign w60326 = ~w60324 & ~w60325;
assign w60327 = pi5658 & ~w60326;
assign w60328 = ~pi5658 & w60326;
assign w60329 = ~w60327 & ~w60328;
assign w60330 = ~w60323 & w60329;
assign w60331 = ~pi7725 & pi9040;
assign w60332 = ~pi7662 & ~pi9040;
assign w60333 = ~w60331 & ~w60332;
assign w60334 = pi5856 & ~w60333;
assign w60335 = ~pi5856 & w60333;
assign w60336 = ~w60334 & ~w60335;
assign w60337 = ~pi7720 & pi9040;
assign w60338 = ~pi7739 & ~pi9040;
assign w60339 = ~w60337 & ~w60338;
assign w60340 = pi5431 & ~w60339;
assign w60341 = ~pi5431 & w60339;
assign w60342 = ~w60340 & ~w60341;
assign w60343 = ~w60336 & w60342;
assign w60344 = w60330 & w60343;
assign w60345 = ~pi7659 & pi9040;
assign w60346 = ~pi7666 & ~pi9040;
assign w60347 = ~w60345 & ~w60346;
assign w60348 = pi5607 & ~w60347;
assign w60349 = ~pi5607 & w60347;
assign w60350 = ~w60348 & ~w60349;
assign w60351 = ~w60336 & ~w60342;
assign w60352 = w60323 & w60351;
assign w60353 = w60336 & w60342;
assign w60354 = w60330 & w60353;
assign w60355 = ~w60351 & ~w60353;
assign w60356 = ~w60323 & ~w60329;
assign w60357 = w60355 & w60356;
assign w60358 = ~pi7739 & pi9040;
assign w60359 = ~pi7749 & ~pi9040;
assign w60360 = ~w60358 & ~w60359;
assign w60361 = pi5684 & ~w60360;
assign w60362 = ~pi5684 & w60360;
assign w60363 = ~w60361 & ~w60362;
assign w60364 = ~w60354 & w60363;
assign w60365 = ~w60357 & w60364;
assign w60366 = ~w60352 & w60365;
assign w60367 = w60329 & ~w60336;
assign w60368 = w60323 & w60367;
assign w60369 = w60323 & w60336;
assign w60370 = ~w60329 & ~w60336;
assign w60371 = w60329 & w60336;
assign w60372 = ~w60370 & ~w60371;
assign w60373 = (w60343 & w60372) | (w60343 & w63341) | (w60372 & w63341);
assign w60374 = ~w60369 & ~w60373;
assign w60375 = ~w60329 & w60342;
assign w60376 = (~w60368 & w60373) | (~w60368 & w64263) | (w60373 & w64263);
assign w60377 = w60366 & ~w60376;
assign w60378 = w60336 & ~w60363;
assign w60379 = w60323 & w60342;
assign w60380 = ~w60329 & w60379;
assign w60381 = ~w60330 & ~w60380;
assign w60382 = w60378 & ~w60381;
assign w60383 = w60351 & w60356;
assign w60384 = ~w60344 & w60350;
assign w60385 = ~w60383 & w60384;
assign w60386 = ~w60382 & w60385;
assign w60387 = ~w60377 & w60386;
assign w60388 = ~w60372 & w60379;
assign w60389 = ~w60329 & ~w60355;
assign w60390 = (w60363 & ~w60367) | (w60363 & w64264) | (~w60367 & w64264);
assign w60391 = w60336 & w60380;
assign w60392 = w60390 & ~w60391;
assign w60393 = w60355 & ~w60369;
assign w60394 = ~w60389 & ~w60393;
assign w60395 = w60392 & w60394;
assign w60396 = w60342 & w60363;
assign w60397 = w60336 & w60356;
assign w60398 = ~w60396 & w60397;
assign w60399 = w60370 & w60396;
assign w60400 = ~w60350 & ~w60399;
assign w60401 = ~w60388 & w60400;
assign w60402 = ~w60398 & w60401;
assign w60403 = ~w60395 & w60402;
assign w60404 = (w60363 & w60372) | (w60363 & w64264) | (w60372 & w64264);
assign w60405 = ~w60323 & ~w60342;
assign w60406 = ~w60367 & w60405;
assign w60407 = ~w60379 & ~w60405;
assign w60408 = w60367 & w60407;
assign w60409 = ~w60363 & ~w60406;
assign w60410 = ~w60408 & w60409;
assign w60411 = ~w60404 & ~w60410;
assign w60412 = (~w60411 & w60387) | (~w60411 & w64265) | (w60387 & w64265);
assign w60413 = ~pi8568 & w60412;
assign w60414 = pi8568 & ~w60412;
assign w60415 = ~w60413 & ~w60414;
assign w60416 = ~pi7650 & pi9040;
assign w60417 = ~pi7700 & ~pi9040;
assign w60418 = ~w60416 & ~w60417;
assign w60419 = pi5674 & ~w60418;
assign w60420 = ~pi5674 & w60418;
assign w60421 = ~w60419 & ~w60420;
assign w60422 = ~pi7742 & pi9040;
assign w60423 = ~pi7741 & ~pi9040;
assign w60424 = ~w60422 & ~w60423;
assign w60425 = pi5694 & ~w60424;
assign w60426 = ~pi5694 & w60424;
assign w60427 = ~w60425 & ~w60426;
assign w60428 = ~pi7752 & pi9040;
assign w60429 = ~pi7683 & ~pi9040;
assign w60430 = ~w60428 & ~w60429;
assign w60431 = pi5475 & ~w60430;
assign w60432 = ~pi5475 & w60430;
assign w60433 = ~w60431 & ~w60432;
assign w60434 = ~pi7689 & pi9040;
assign w60435 = ~pi7811 & ~pi9040;
assign w60436 = ~w60434 & ~w60435;
assign w60437 = pi5693 & ~w60436;
assign w60438 = ~pi5693 & w60436;
assign w60439 = ~w60437 & ~w60438;
assign w60440 = ~w60433 & ~w60439;
assign w60441 = ~pi7811 & pi9040;
assign w60442 = ~pi7742 & ~pi9040;
assign w60443 = ~w60441 & ~w60442;
assign w60444 = pi5703 & ~w60443;
assign w60445 = ~pi5703 & w60443;
assign w60446 = ~w60444 & ~w60445;
assign w60447 = ~w60427 & ~w60446;
assign w60448 = ~w60440 & w60447;
assign w60449 = ~w60433 & ~w60446;
assign w60450 = ~pi7661 & pi9040;
assign w60451 = ~pi7817 & ~pi9040;
assign w60452 = ~w60450 & ~w60451;
assign w60453 = pi5841 & ~w60452;
assign w60454 = ~pi5841 & w60452;
assign w60455 = ~w60453 & ~w60454;
assign w60456 = w60439 & w60455;
assign w60457 = w60449 & w60456;
assign w60458 = w60427 & w60446;
assign w60459 = ~w60455 & ~w60458;
assign w60460 = ~w60427 & w60433;
assign w60461 = w60455 & ~w60460;
assign w60462 = ~w60459 & ~w60461;
assign w60463 = ~w60448 & ~w60457;
assign w60464 = ~w60462 & w60463;
assign w60465 = w60440 & w60458;
assign w60466 = ~w60439 & ~w60446;
assign w60467 = ~w60455 & w60466;
assign w60468 = w60466 & w64266;
assign w60469 = ~w60465 & ~w60468;
assign w60470 = w60433 & w60446;
assign w60471 = ~w60449 & ~w60470;
assign w60472 = w60427 & ~w60455;
assign w60473 = ~w60439 & ~w60472;
assign w60474 = w60471 & w60473;
assign w60475 = w60469 & w60474;
assign w60476 = w60464 & ~w60475;
assign w60477 = w60421 & ~w60476;
assign w60478 = ~w60427 & w60457;
assign w60479 = ~w60427 & ~w60439;
assign w60480 = w60446 & w60455;
assign w60481 = w60479 & w60480;
assign w60482 = w60427 & ~w60433;
assign w60483 = ~w60460 & ~w60482;
assign w60484 = w60459 & w60483;
assign w60485 = ~w60427 & ~w60471;
assign w60486 = ~w60471 & w64267;
assign w60487 = ~w60484 & ~w60486;
assign w60488 = w60433 & w60439;
assign w60489 = ~w60440 & ~w60488;
assign w60490 = ~w60455 & ~w60489;
assign w60491 = w60487 & w60490;
assign w60492 = w60466 & w60482;
assign w60493 = w60439 & w60471;
assign w60494 = w60471 & w63486;
assign w60495 = w60471 & w64268;
assign w60496 = w60439 & w60446;
assign w60497 = w60484 & w60496;
assign w60498 = ~w60460 & w60467;
assign w60499 = w60470 & w60473;
assign w60500 = ~w60492 & ~w60498;
assign w60501 = ~w60499 & w60500;
assign w60502 = w60501 & w64269;
assign w60503 = ~w60421 & ~w60502;
assign w60504 = ~w60478 & ~w60481;
assign w60505 = ~w60491 & w60504;
assign w60506 = ~w60477 & w60505;
assign w60507 = ~w60503 & w60506;
assign w60508 = ~pi8556 & ~w60507;
assign w60509 = pi8556 & w60507;
assign w60510 = ~w60508 & ~w60509;
assign w60511 = ~w60355 & w64270;
assign w60512 = w60367 & w60405;
assign w60513 = ~w60511 & ~w60512;
assign w60514 = ~w60397 & w60513;
assign w60515 = ~w60342 & ~w60514;
assign w60516 = ~w60371 & w60407;
assign w60517 = w60363 & ~w60516;
assign w60518 = w60373 & ~w60390;
assign w60519 = ~w60350 & ~w60354;
assign w60520 = ~w60517 & w60519;
assign w60521 = ~w60518 & w60520;
assign w60522 = ~w60515 & w60521;
assign w60523 = w60344 & w60363;
assign w60524 = ~w60342 & w60371;
assign w60525 = w60376 & ~w60524;
assign w60526 = w60374 & ~w60525;
assign w60527 = ~w60369 & ~w60383;
assign w60528 = ~w60363 & ~w60527;
assign w60529 = w60350 & ~w60523;
assign w60530 = ~w60528 & w60529;
assign w60531 = ~w60526 & w60530;
assign w60532 = ~w60522 & ~w60531;
assign w60533 = ~pi8602 & w60532;
assign w60534 = pi8602 & ~w60532;
assign w60535 = ~w60533 & ~w60534;
assign w60536 = ~pi7679 & pi9040;
assign w60537 = ~pi7745 & ~pi9040;
assign w60538 = ~w60536 & ~w60537;
assign w60539 = pi5607 & ~w60538;
assign w60540 = ~pi5607 & w60538;
assign w60541 = ~w60539 & ~w60540;
assign w60542 = ~pi7675 & pi9040;
assign w60543 = ~pi7660 & ~pi9040;
assign w60544 = ~w60542 & ~w60543;
assign w60545 = pi5431 & ~w60544;
assign w60546 = ~pi5431 & w60544;
assign w60547 = ~w60545 & ~w60546;
assign w60548 = ~w60541 & ~w60547;
assign w60549 = ~pi7658 & pi9040;
assign w60550 = ~pi7821 & ~pi9040;
assign w60551 = ~w60549 & ~w60550;
assign w60552 = pi5694 & ~w60551;
assign w60553 = ~pi5694 & w60551;
assign w60554 = ~w60552 & ~w60553;
assign w60555 = w60548 & w60554;
assign w60556 = ~pi7813 & pi9040;
assign w60557 = ~pi7648 & ~pi9040;
assign w60558 = ~w60556 & ~w60557;
assign w60559 = pi5465 & ~w60558;
assign w60560 = ~pi5465 & w60558;
assign w60561 = ~w60559 & ~w60560;
assign w60562 = ~w60555 & w60561;
assign w60563 = ~pi7670 & pi9040;
assign w60564 = ~pi7720 & ~pi9040;
assign w60565 = ~w60563 & ~w60564;
assign w60566 = pi5895 & ~w60565;
assign w60567 = ~pi5895 & w60565;
assign w60568 = ~w60566 & ~w60567;
assign w60569 = ~w60554 & w60568;
assign w60570 = w60541 & ~w60547;
assign w60571 = w60569 & w60570;
assign w60572 = ~pi7744 & pi9040;
assign w60573 = ~pi7658 & ~pi9040;
assign w60574 = ~w60572 & ~w60573;
assign w60575 = pi5703 & ~w60574;
assign w60576 = ~pi5703 & w60574;
assign w60577 = ~w60575 & ~w60576;
assign w60578 = ~w60571 & ~w60577;
assign w60579 = w60562 & w60578;
assign w60580 = w60547 & w60554;
assign w60581 = ~w60561 & ~w60580;
assign w60582 = ~w60541 & ~w60554;
assign w60583 = w60568 & w60582;
assign w60584 = ~w60577 & w60581;
assign w60585 = ~w60583 & w60584;
assign w60586 = ~w60579 & ~w60585;
assign w60587 = w60568 & ~w60580;
assign w60588 = w60547 & ~w60554;
assign w60589 = w60541 & ~w60568;
assign w60590 = ~w60588 & ~w60589;
assign w60591 = ~w60568 & w60588;
assign w60592 = w60588 & w60589;
assign w60593 = w60561 & ~w60590;
assign w60594 = ~w60592 & w60593;
assign w60595 = w60541 & ~w60587;
assign w60596 = ~w60594 & w60595;
assign w60597 = ~w60586 & ~w60596;
assign w60598 = ~w60547 & ~w60568;
assign w60599 = ~w60541 & ~w60561;
assign w60600 = w60598 & w60599;
assign w60601 = ~w60541 & w60547;
assign w60602 = w60568 & w60601;
assign w60603 = w60554 & w60602;
assign w60604 = ~w60600 & ~w60603;
assign w60605 = ~w60547 & w60568;
assign w60606 = w60541 & ~w60561;
assign w60607 = w60605 & w60606;
assign w60608 = w60577 & ~w60607;
assign w60609 = ~w60594 & w60608;
assign w60610 = w60604 & w60609;
assign w60611 = ~w60597 & ~w60610;
assign w60612 = ~w60561 & ~w60592;
assign w60613 = w60554 & w60568;
assign w60614 = w60554 & w60598;
assign w60615 = ~w60602 & ~w60613;
assign w60616 = ~w60614 & w60615;
assign w60617 = (~w60590 & ~w60615) | (~w60590 & w64271) | (~w60615 & w64271);
assign w60618 = w60541 & w60561;
assign w60619 = ~w60601 & ~w60618;
assign w60620 = w60613 & w60619;
assign w60621 = ~w60554 & ~w60568;
assign w60622 = w60548 & w60621;
assign w60623 = w60561 & ~w60622;
assign w60624 = ~w60620 & w60623;
assign w60625 = ~w60617 & w60624;
assign w60626 = ~w60612 & ~w60625;
assign w60627 = ~w60611 & ~w60626;
assign w60628 = ~pi8557 & w60627;
assign w60629 = pi8557 & ~w60627;
assign w60630 = ~w60628 & ~w60629;
assign w60631 = ~pi7727 & pi9040;
assign w60632 = ~pi7736 & ~pi9040;
assign w60633 = ~w60631 & ~w60632;
assign w60634 = pi5550 & ~w60633;
assign w60635 = ~pi5550 & w60633;
assign w60636 = ~w60634 & ~w60635;
assign w60637 = ~pi7795 & pi9040;
assign w60638 = ~pi7664 & ~pi9040;
assign w60639 = ~w60637 & ~w60638;
assign w60640 = pi5585 & ~w60639;
assign w60641 = ~pi5585 & w60639;
assign w60642 = ~w60640 & ~w60641;
assign w60643 = ~pi7693 & pi9040;
assign w60644 = ~pi7727 & ~pi9040;
assign w60645 = ~w60643 & ~w60644;
assign w60646 = pi5512 & ~w60645;
assign w60647 = ~pi5512 & w60645;
assign w60648 = ~w60646 & ~w60647;
assign w60649 = w60642 & w60648;
assign w60650 = ~pi7663 & pi9040;
assign w60651 = ~pi7655 & ~pi9040;
assign w60652 = ~w60650 & ~w60651;
assign w60653 = pi5750 & ~w60652;
assign w60654 = ~pi5750 & w60652;
assign w60655 = ~w60653 & ~w60654;
assign w60656 = w60649 & ~w60655;
assign w60657 = (~w60636 & ~w60649) | (~w60636 & w60660) | (~w60649 & w60660);
assign w60658 = w60642 & ~w60655;
assign w60659 = w60657 & w60658;
assign w60660 = ~w60636 & w60655;
assign w60661 = ~pi7660 & pi9040;
assign w60662 = ~pi7693 & ~pi9040;
assign w60663 = ~w60661 & ~w60662;
assign w60664 = pi5813 & ~w60663;
assign w60665 = ~pi5813 & w60663;
assign w60666 = ~w60664 & ~w60665;
assign w60667 = w60648 & w60666;
assign w60668 = w60660 & w60667;
assign w60669 = ~w60636 & w60642;
assign w60670 = w60655 & ~w60669;
assign w60671 = ~w60649 & ~w60670;
assign w60672 = w60636 & w60649;
assign w60673 = w60636 & ~w60642;
assign w60674 = w60655 & w60673;
assign w60675 = (~w60666 & ~w60649) | (~w60666 & w60703) | (~w60649 & w60703);
assign w60676 = ~w60674 & w60675;
assign w60677 = ~w60671 & w60676;
assign w60678 = ~pi7664 & pi9040;
assign w60679 = ~pi7813 & ~pi9040;
assign w60680 = ~w60678 & ~w60679;
assign w60681 = pi5856 & ~w60680;
assign w60682 = ~pi5856 & w60680;
assign w60683 = ~w60681 & ~w60682;
assign w60684 = w60648 & ~w60655;
assign w60685 = w60673 & w60684;
assign w60686 = w60642 & ~w60648;
assign w60687 = w60655 & w60686;
assign w60688 = (w60666 & ~w60686) | (w60666 & w63487) | (~w60686 & w63487);
assign w60689 = ~w60642 & ~w60648;
assign w60690 = ~w60655 & w60689;
assign w60691 = w60636 & w60690;
assign w60692 = ~w60660 & w60689;
assign w60693 = ~w60672 & ~w60692;
assign w60694 = ~w60669 & w64272;
assign w60695 = w60693 & w60694;
assign w60696 = ~w60691 & ~w60695;
assign w60697 = ~w60684 & w60688;
assign w60698 = ~w60695 & w64273;
assign w60699 = ~w60683 & ~w60685;
assign w60700 = ~w60677 & w60699;
assign w60701 = ~w60698 & w60700;
assign w60702 = w60657 & w60684;
assign w60703 = ~w60636 & ~w60666;
assign w60704 = w60686 & w60703;
assign w60705 = w60649 & w64274;
assign w60706 = ~w60704 & ~w60705;
assign w60707 = ~w60702 & w60706;
assign w60708 = (w60683 & w60693) | (w60683 & w64275) | (w60693 & w64275);
assign w60709 = w60696 & w64276;
assign w60710 = ~w60701 & ~w60709;
assign w60711 = ~w60659 & ~w60668;
assign w60712 = ~w60710 & w60711;
assign w60713 = pi8605 & w60712;
assign w60714 = ~pi8605 & ~w60712;
assign w60715 = ~w60713 & ~w60714;
assign w60716 = ~w60642 & w60666;
assign w60717 = (~w60636 & w60687) | (~w60636 & w64277) | (w60687 & w64277);
assign w60718 = w60706 & ~w60717;
assign w60719 = ~w60683 & ~w60718;
assign w60720 = ~w60669 & ~w60673;
assign w60721 = ~w60666 & ~w60683;
assign w60722 = w60655 & w60721;
assign w60723 = ~w60720 & w60722;
assign w60724 = ~w60655 & ~w60669;
assign w60725 = w60689 & w60703;
assign w60726 = w60666 & ~w60683;
assign w60727 = ~w60689 & w60726;
assign w60728 = ~w60725 & ~w60727;
assign w60729 = w60724 & ~w60728;
assign w60730 = w60655 & w60689;
assign w60731 = w60689 & w60660;
assign w60732 = ~w60672 & ~w60731;
assign w60733 = w60666 & ~w60732;
assign w60734 = w60648 & w60655;
assign w60735 = ~w60642 & w60734;
assign w60736 = w60657 & ~w60735;
assign w60737 = w60676 & ~w60736;
assign w60738 = ~w60649 & ~w60658;
assign w60739 = ~w60684 & ~w60738;
assign w60740 = (~w60673 & w60738) | (~w60673 & w64278) | (w60738 & w64278);
assign w60741 = w60666 & ~w60724;
assign w60742 = ~w60740 & w60741;
assign w60743 = ~w60737 & ~w60742;
assign w60744 = w60683 & ~w60743;
assign w60745 = w60642 & ~w60660;
assign w60746 = ~w60690 & ~w60735;
assign w60747 = w60688 & w60746;
assign w60748 = (w60648 & ~w60746) | (w60648 & w63488) | (~w60746 & w63488);
assign w60749 = ~w60692 & ~w60745;
assign w60750 = ~w60748 & w60749;
assign w60751 = ~w60707 & w60750;
assign w60752 = ~w60723 & ~w60729;
assign w60753 = ~w60733 & w60752;
assign w60754 = ~w60719 & w60753;
assign w60755 = w60754 & w64279;
assign w60756 = pi8592 & ~w60755;
assign w60757 = ~pi8592 & w60755;
assign w60758 = ~w60756 & ~w60757;
assign w60759 = w60323 & w60355;
assign w60760 = w60355 & w64280;
assign w60761 = ~w60354 & ~w60760;
assign w60762 = ~w60363 & ~w60511;
assign w60763 = ~w60336 & w60356;
assign w60764 = ~w60524 & ~w60763;
assign w60765 = w60390 & w60764;
assign w60766 = ~w60759 & w60765;
assign w60767 = (w60761 & w60766) | (w60761 & w64281) | (w60766 & w64281);
assign w60768 = w60350 & ~w60767;
assign w60769 = ~w60350 & ~w60513;
assign w60770 = w60363 & w60761;
assign w60771 = ~w60769 & w60770;
assign w60772 = ~w60389 & ~w60760;
assign w60773 = w60519 & w60772;
assign w60774 = ~w60363 & ~w60512;
assign w60775 = ~w60773 & w60774;
assign w60776 = ~w60771 & ~w60775;
assign w60777 = ~w60768 & ~w60776;
assign w60778 = ~pi8550 & w60777;
assign w60779 = pi8550 & ~w60777;
assign w60780 = ~w60778 & ~w60779;
assign w60781 = ~pi7741 & pi9040;
assign w60782 = ~pi7846 & ~pi9040;
assign w60783 = ~w60781 & ~w60782;
assign w60784 = pi5795 & ~w60783;
assign w60785 = ~pi5795 & w60783;
assign w60786 = ~w60784 & ~w60785;
assign w60787 = ~pi7721 & pi9040;
assign w60788 = ~pi7674 & ~pi9040;
assign w60789 = ~w60787 & ~w60788;
assign w60790 = pi5805 & ~w60789;
assign w60791 = ~pi5805 & w60789;
assign w60792 = ~w60790 & ~w60791;
assign w60793 = w60786 & w60792;
assign w60794 = ~pi7817 & pi9040;
assign w60795 = ~pi7703 & ~pi9040;
assign w60796 = ~w60794 & ~w60795;
assign w60797 = pi5586 & ~w60796;
assign w60798 = ~pi5586 & w60796;
assign w60799 = ~w60797 & ~w60798;
assign w60800 = ~pi7651 & pi9040;
assign w60801 = ~pi7733 & ~pi9040;
assign w60802 = ~w60800 & ~w60801;
assign w60803 = pi5534 & ~w60802;
assign w60804 = ~pi5534 & w60802;
assign w60805 = ~w60803 & ~w60804;
assign w60806 = w60799 & ~w60805;
assign w60807 = ~pi7703 & pi9040;
assign w60808 = ~pi7752 & ~pi9040;
assign w60809 = ~w60807 & ~w60808;
assign w60810 = pi5748 & ~w60809;
assign w60811 = ~pi5748 & w60809;
assign w60812 = ~w60810 & ~w60811;
assign w60813 = w60805 & ~w60812;
assign w60814 = ~w60799 & w60813;
assign w60815 = ~w60806 & ~w60814;
assign w60816 = w60793 & ~w60815;
assign w60817 = w60792 & w60805;
assign w60818 = ~w60792 & ~w60805;
assign w60819 = ~w60817 & ~w60818;
assign w60820 = w60799 & w60812;
assign w60821 = ~w60819 & w60820;
assign w60822 = ~w60805 & ~w60812;
assign w60823 = ~w60799 & w60822;
assign w60824 = ~w60821 & ~w60823;
assign w60825 = ~w60786 & ~w60792;
assign w60826 = ~w60805 & w60812;
assign w60827 = ~w60799 & ~w60813;
assign w60828 = ~w60826 & ~w60827;
assign w60829 = ~w60827 & w64282;
assign w60830 = ~w60825 & ~w60829;
assign w60831 = ~w60824 & ~w60830;
assign w60832 = w60822 & w60825;
assign w60833 = ~pi7723 & pi9040;
assign w60834 = ~pi7651 & ~pi9040;
assign w60835 = ~w60833 & ~w60834;
assign w60836 = pi5749 & ~w60835;
assign w60837 = ~pi5749 & w60835;
assign w60838 = ~w60836 & ~w60837;
assign w60839 = ~w60832 & ~w60838;
assign w60840 = w60786 & ~w60792;
assign w60841 = w60805 & w60840;
assign w60842 = ~w60827 & w60841;
assign w60843 = w60792 & ~w60799;
assign w60844 = ~w60792 & w60799;
assign w60845 = w60822 & ~w60843;
assign w60846 = ~w60844 & w60845;
assign w60847 = w60805 & w60812;
assign w60848 = ~w60786 & w60847;
assign w60849 = w60786 & w60826;
assign w60850 = ~w60817 & ~w60848;
assign w60851 = ~w60849 & w60850;
assign w60852 = ~w60799 & ~w60851;
assign w60853 = w60839 & ~w60842;
assign w60854 = ~w60846 & w60853;
assign w60855 = ~w60852 & w60854;
assign w60856 = w60793 & w60822;
assign w60857 = w60786 & w60812;
assign w60858 = ~w60792 & ~w60799;
assign w60859 = w60805 & w60858;
assign w60860 = w60857 & w60859;
assign w60861 = w60813 & ~w60843;
assign w60862 = w60826 & w60843;
assign w60863 = ~w60861 & ~w60862;
assign w60864 = ~w60786 & ~w60863;
assign w60865 = w60838 & ~w60856;
assign w60866 = ~w60821 & w60865;
assign w60867 = ~w60860 & w60866;
assign w60868 = ~w60864 & w60867;
assign w60869 = ~w60855 & ~w60868;
assign w60870 = ~w60816 & ~w60831;
assign w60871 = ~w60869 & w60870;
assign w60872 = pi8554 & ~w60871;
assign w60873 = ~pi8554 & w60871;
assign w60874 = ~w60872 & ~w60873;
assign w60875 = w60793 & ~w60838;
assign w60876 = w60828 & w60875;
assign w60877 = ~w60840 & ~w60843;
assign w60878 = w60822 & ~w60877;
assign w60879 = w60792 & w60813;
assign w60880 = ~w60826 & ~w60879;
assign w60881 = w60799 & ~w60825;
assign w60882 = ~w60880 & w60881;
assign w60883 = ~w60793 & ~w60858;
assign w60884 = w60847 & ~w60883;
assign w60885 = ~w60806 & w60812;
assign w60886 = w60877 & w60885;
assign w60887 = ~w60884 & w60886;
assign w60888 = ~w60878 & ~w60882;
assign w60889 = ~w60887 & w60888;
assign w60890 = w60838 & ~w60889;
assign w60891 = ~w60814 & ~w60843;
assign w60892 = w60880 & ~w60891;
assign w60893 = ~w60792 & ~w60838;
assign w60894 = ~w60885 & w60893;
assign w60895 = ~w60892 & ~w60894;
assign w60896 = ~w60786 & ~w60895;
assign w60897 = w60838 & ~w60857;
assign w60898 = ~w60859 & ~w60862;
assign w60899 = ~w60897 & ~w60898;
assign w60900 = ~w60876 & ~w60899;
assign w60901 = ~w60896 & w60900;
assign w60902 = ~w60890 & w60901;
assign w60903 = ~pi8579 & ~w60902;
assign w60904 = pi8579 & w60902;
assign w60905 = ~w60903 & ~w60904;
assign w60906 = w60656 & w60703;
assign w60907 = w60636 & ~w60746;
assign w60908 = w60658 & ~w60666;
assign w60909 = w60683 & ~w60908;
assign w60910 = ~w60702 & w60909;
assign w60911 = ~w60907 & w60910;
assign w60912 = ~w60750 & w60911;
assign w60913 = w60636 & w60734;
assign w60914 = (~w60716 & ~w60746) | (~w60716 & w64283) | (~w60746 & w64283);
assign w60915 = ~w60730 & ~w60745;
assign w60916 = (~w60683 & w60915) | (~w60683 & w60721) | (w60915 & w60721);
assign w60917 = ~w60914 & w60916;
assign w60918 = ~w60751 & w60917;
assign w60919 = (~w60906 & w60918) | (~w60906 & w64284) | (w60918 & w64284);
assign w60920 = pi8633 & w60919;
assign w60921 = ~pi8633 & ~w60919;
assign w60922 = ~w60920 & ~w60921;
assign w60923 = ~pi7700 & pi9040;
assign w60924 = ~pi7721 & ~pi9040;
assign w60925 = ~w60923 & ~w60924;
assign w60926 = pi5446 & ~w60925;
assign w60927 = ~pi5446 & w60925;
assign w60928 = ~w60926 & ~w60927;
assign w60929 = ~pi7733 & pi9040;
assign w60930 = ~pi7677 & ~pi9040;
assign w60931 = ~w60929 & ~w60930;
assign w60932 = pi5798 & ~w60931;
assign w60933 = ~pi5798 & w60931;
assign w60934 = ~w60932 & ~w60933;
assign w60935 = ~pi7668 & pi9040;
assign w60936 = ~pi7803 & ~pi9040;
assign w60937 = ~w60935 & ~w60936;
assign w60938 = pi5650 & ~w60937;
assign w60939 = ~pi5650 & w60937;
assign w60940 = ~w60938 & ~w60939;
assign w60941 = w60934 & w60940;
assign w60942 = ~pi7683 & pi9040;
assign w60943 = ~pi7689 & ~pi9040;
assign w60944 = ~w60942 & ~w60943;
assign w60945 = pi5805 & ~w60944;
assign w60946 = ~pi5805 & w60944;
assign w60947 = ~w60945 & ~w60946;
assign w60948 = w60941 & ~w60947;
assign w60949 = ~w60928 & w60948;
assign w60950 = ~pi7686 & pi9040;
assign w60951 = ~pi7650 & ~pi9040;
assign w60952 = ~w60950 & ~w60951;
assign w60953 = pi5534 & ~w60952;
assign w60954 = ~pi5534 & w60952;
assign w60955 = ~w60953 & ~w60954;
assign w60956 = ~w60934 & ~w60940;
assign w60957 = ~pi7846 & pi9040;
assign w60958 = ~pi7686 & ~pi9040;
assign w60959 = ~w60957 & ~w60958;
assign w60960 = pi5587 & ~w60959;
assign w60961 = ~pi5587 & w60959;
assign w60962 = ~w60960 & ~w60961;
assign w60963 = w60947 & w60962;
assign w60964 = ~w60947 & ~w60962;
assign w60965 = ~w60963 & ~w60964;
assign w60966 = w60956 & ~w60965;
assign w60967 = ~w60934 & w60962;
assign w60968 = ~w60940 & ~w60962;
assign w60969 = ~w60967 & ~w60968;
assign w60970 = w60965 & w60969;
assign w60971 = ~w60966 & ~w60970;
assign w60972 = ~w60934 & ~w60971;
assign w60973 = w60934 & ~w60962;
assign w60974 = w60947 & w60973;
assign w60975 = (~w60928 & ~w60973) | (~w60928 & w64285) | (~w60973 & w64285);
assign w60976 = w60934 & ~w60947;
assign w60977 = ~w60940 & w60962;
assign w60978 = ~w60976 & w60977;
assign w60979 = w60975 & ~w60978;
assign w60980 = w60940 & w60962;
assign w60981 = ~w60976 & ~w60980;
assign w60982 = w60928 & w60981;
assign w60983 = ~w60948 & ~w60982;
assign w60984 = ~w60979 & w60983;
assign w60985 = ~w60972 & ~w60984;
assign w60986 = ~w60955 & ~w60985;
assign w60987 = w60940 & w60964;
assign w60988 = w60947 & w60968;
assign w60989 = ~w60987 & ~w60988;
assign w60990 = w60928 & ~w60989;
assign w60991 = ~w60947 & ~w60968;
assign w60992 = w60956 & w60991;
assign w60993 = w60928 & w60934;
assign w60994 = w60968 & w60993;
assign w60995 = ~w60992 & ~w60994;
assign w60996 = w60982 & ~w60995;
assign w60997 = ~w60990 & ~w60996;
assign w60998 = w60955 & ~w60997;
assign w60999 = ~w60934 & w60947;
assign w61000 = ~w60967 & ~w60973;
assign w61001 = ~w60981 & ~w61000;
assign w61002 = ~w60965 & w63489;
assign w61003 = w61001 & ~w61002;
assign w61004 = w60999 & w61003;
assign w61005 = ~w60928 & w60955;
assign w61006 = (w61005 & w61001) | (w61005 & w64286) | (w61001 & w64286);
assign w61007 = w60941 & w60955;
assign w61008 = ~w60963 & w61007;
assign w61009 = ~w60949 & ~w61008;
assign w61010 = ~w61006 & w61009;
assign w61011 = ~w61004 & w61010;
assign w61012 = ~w60986 & w61011;
assign w61013 = (pi8629 & ~w61012) | (pi8629 & w64287) | (~w61012 & w64287);
assign w61014 = w61012 & w64288;
assign w61015 = ~w61013 & ~w61014;
assign w61016 = ~w60336 & w60405;
assign w61017 = ~w60363 & ~w60380;
assign w61018 = ~w61016 & w61017;
assign w61019 = ~w60366 & ~w61018;
assign w61020 = ~w60404 & w60524;
assign w61021 = ~w60344 & ~w60363;
assign w61022 = ~w60392 & ~w61021;
assign w61023 = w60350 & ~w61020;
assign w61024 = ~w61022 & w61023;
assign w61025 = ~w61019 & w61024;
assign w61026 = w60369 & w60772;
assign w61027 = w60365 & ~w60407;
assign w61028 = w60378 & ~w60379;
assign w61029 = ~w60524 & w61028;
assign w61030 = ~w60350 & ~w60408;
assign w61031 = ~w61029 & w61030;
assign w61032 = ~w61027 & w61031;
assign w61033 = ~w61026 & w61032;
assign w61034 = ~w61025 & ~w61033;
assign w61035 = pi8561 & w61034;
assign w61036 = ~pi8561 & ~w61034;
assign w61037 = ~w61035 & ~w61036;
assign w61038 = w60688 & ~w60719;
assign w61039 = ~w60728 & ~w61038;
assign w61040 = ~w60685 & ~w60730;
assign w61041 = w60721 & ~w61040;
assign w61042 = ~w60667 & w60683;
assign w61043 = w60667 & ~w60683;
assign w61044 = ~w60636 & ~w60738;
assign w61045 = ~w61042 & ~w61043;
assign w61046 = w61044 & w61045;
assign w61047 = w60703 & w60738;
assign w61048 = ~w60731 & ~w60913;
assign w61049 = ~w61047 & w61048;
assign w61050 = w60683 & ~w61049;
assign w61051 = ~w60666 & ~w60739;
assign w61052 = w60636 & ~w60747;
assign w61053 = ~w61051 & w61052;
assign w61054 = ~w61041 & ~w61046;
assign w61055 = ~w61050 & w61054;
assign w61056 = ~w61053 & w61055;
assign w61057 = ~w61039 & w61056;
assign w61058 = pi8570 & ~w61057;
assign w61059 = ~pi8570 & w61057;
assign w61060 = ~w61058 & ~w61059;
assign w61061 = w60813 & w60844;
assign w61062 = ~w60823 & ~w61061;
assign w61063 = w60840 & ~w61062;
assign w61064 = w60817 & w60820;
assign w61065 = ~w60862 & ~w61064;
assign w61066 = w60799 & w60832;
assign w61067 = w61065 & ~w61066;
assign w61068 = w60838 & ~w61067;
assign w61069 = ~w60786 & ~w60799;
assign w61070 = w60819 & w61069;
assign w61071 = w60786 & ~w60819;
assign w61072 = ~w60880 & w61071;
assign w61073 = ~w61070 & ~w61072;
assign w61074 = ~w61068 & w61073;
assign w61075 = w60792 & w60814;
assign w61076 = ~w60838 & w61065;
assign w61077 = ~w61075 & w61076;
assign w61078 = ~w60786 & ~w60814;
assign w61079 = ~w60792 & w60812;
assign w61080 = ~w60861 & ~w61079;
assign w61081 = w61078 & ~w61080;
assign w61082 = w60786 & ~w61079;
assign w61083 = ~w60805 & ~w60843;
assign w61084 = w61082 & w61083;
assign w61085 = ~w60846 & ~w60884;
assign w61086 = ~w61084 & w61085;
assign w61087 = ~w61081 & w61086;
assign w61088 = ~w60838 & ~w61087;
assign w61089 = (~w61063 & w61074) | (~w61063 & w64289) | (w61074 & w64289);
assign w61090 = ~w61088 & w61089;
assign w61091 = ~pi8503 & w61090;
assign w61092 = pi8503 & ~w61090;
assign w61093 = ~w61091 & ~w61092;
assign w61094 = ~w60928 & ~w60980;
assign w61095 = w60991 & w61094;
assign w61096 = w60940 & w60974;
assign w61097 = w60962 & w60976;
assign w61098 = w60947 & ~w61000;
assign w61099 = ~w61097 & ~w61098;
assign w61100 = w60964 & ~w60993;
assign w61101 = ~w60940 & ~w61100;
assign w61102 = w61099 & w61101;
assign w61103 = w60955 & ~w61095;
assign w61104 = ~w61096 & w61103;
assign w61105 = ~w61102 & w61104;
assign w61106 = (w60928 & w61098) | (w60928 & w64290) | (w61098 & w64290);
assign w61107 = w60975 & ~w60991;
assign w61108 = ~w60967 & w61107;
assign w61109 = w60956 & w60964;
assign w61110 = ~w60955 & ~w61109;
assign w61111 = ~w61106 & w61110;
assign w61112 = ~w61108 & w61111;
assign w61113 = ~w61105 & ~w61112;
assign w61114 = ~w60928 & ~w60967;
assign w61115 = ~w60947 & w61000;
assign w61116 = w60928 & ~w61115;
assign w61117 = w60940 & ~w61114;
assign w61118 = ~w61116 & w61117;
assign w61119 = ~w61113 & ~w61118;
assign w61120 = ~pi8520 & w61119;
assign w61121 = pi8520 & ~w61119;
assign w61122 = ~w61120 & ~w61121;
assign w61123 = w60577 & ~w60605;
assign w61124 = ~w60591 & ~w61123;
assign w61125 = (w60561 & ~w60616) | (w60561 & w64291) | (~w60616 & w64291);
assign w61126 = w60541 & w60554;
assign w61127 = ~w60582 & ~w61126;
assign w61128 = w60547 & w60577;
assign w61129 = w61127 & w61128;
assign w61130 = w60612 & ~w61129;
assign w61131 = ~w60617 & w61130;
assign w61132 = ~w61125 & ~w61131;
assign w61133 = w60588 & w60599;
assign w61134 = ~w60620 & ~w61133;
assign w61135 = ~w60577 & ~w61134;
assign w61136 = w60601 & ~w60621;
assign w61137 = ~w60547 & ~w60555;
assign w61138 = w60561 & ~w61136;
assign w61139 = ~w61137 & w61138;
assign w61140 = ~w61127 & w61139;
assign w61141 = ~w60571 & ~w60614;
assign w61142 = w60604 & w61141;
assign w61143 = ~w61140 & w61142;
assign w61144 = w60577 & ~w61143;
assign w61145 = ~w61132 & ~w61135;
assign w61146 = ~w61144 & w61145;
assign w61147 = ~pi8685 & w61146;
assign w61148 = pi8685 & ~w61146;
assign w61149 = ~w61147 & ~w61148;
assign w61150 = ~pi7649 & pi9040;
assign w61151 = ~pi7708 & ~pi9040;
assign w61152 = ~w61150 & ~w61151;
assign w61153 = pi5674 & ~w61152;
assign w61154 = ~pi5674 & w61152;
assign w61155 = ~w61153 & ~w61154;
assign w61156 = ~pi7698 & pi9040;
assign w61157 = ~pi7649 & ~pi9040;
assign w61158 = ~w61156 & ~w61157;
assign w61159 = pi5475 & ~w61158;
assign w61160 = ~pi5475 & w61158;
assign w61161 = ~w61159 & ~w61160;
assign w61162 = w61155 & w61161;
assign w61163 = ~pi7803 & pi9040;
assign w61164 = ~pi7684 & ~pi9040;
assign w61165 = ~w61163 & ~w61164;
assign w61166 = pi5690 & ~w61165;
assign w61167 = ~pi5690 & w61165;
assign w61168 = ~w61166 & ~w61167;
assign w61169 = ~pi7674 & pi9040;
assign w61170 = ~pi7723 & ~pi9040;
assign w61171 = ~w61169 & ~w61170;
assign w61172 = pi5798 & ~w61171;
assign w61173 = ~pi5798 & w61171;
assign w61174 = ~w61172 & ~w61173;
assign w61175 = w61168 & ~w61174;
assign w61176 = w61162 & w61175;
assign w61177 = ~w61155 & ~w61161;
assign w61178 = w61168 & w61177;
assign w61179 = ~w61176 & ~w61178;
assign w61180 = ~pi7746 & pi9040;
assign w61181 = ~pi7661 & ~pi9040;
assign w61182 = ~w61180 & ~w61181;
assign w61183 = pi5587 & ~w61182;
assign w61184 = ~pi5587 & w61182;
assign w61185 = ~w61183 & ~w61184;
assign w61186 = w61174 & w61177;
assign w61187 = ~w61161 & ~w61168;
assign w61188 = ~w61174 & w61187;
assign w61189 = w61187 & w61203;
assign w61190 = ~w61162 & ~w61186;
assign w61191 = ~w61189 & w61190;
assign w61192 = ~w61185 & ~w61191;
assign w61193 = w61179 & ~w61192;
assign w61194 = ~pi7708 & pi9040;
assign w61195 = ~pi7705 & ~pi9040;
assign w61196 = ~w61194 & ~w61195;
assign w61197 = pi5598 & ~w61196;
assign w61198 = ~pi5598 & w61196;
assign w61199 = ~w61197 & ~w61198;
assign w61200 = ~w61193 & ~w61199;
assign w61201 = ~w61161 & w61168;
assign w61202 = ~w61155 & w61174;
assign w61203 = w61155 & ~w61174;
assign w61204 = ~w61202 & ~w61203;
assign w61205 = w61201 & w61204;
assign w61206 = ~w61155 & ~w61175;
assign w61207 = ~w61186 & w61206;
assign w61208 = w61199 & w61207;
assign w61209 = ~w61176 & ~w61185;
assign w61210 = ~w61205 & w61209;
assign w61211 = ~w61208 & w61210;
assign w61212 = w61177 & w64292;
assign w61213 = ~w61199 & w61207;
assign w61214 = w61161 & ~w61199;
assign w61215 = w61155 & w61174;
assign w61216 = ~w61214 & w61215;
assign w61217 = ~w61201 & w61216;
assign w61218 = w61155 & ~w61168;
assign w61219 = ~w61175 & ~w61218;
assign w61220 = w61179 & w61199;
assign w61221 = ~w61219 & w61220;
assign w61222 = w61185 & ~w61212;
assign w61223 = ~w61217 & w61222;
assign w61224 = ~w61213 & w61223;
assign w61225 = ~w61221 & w61224;
assign w61226 = ~w61211 & ~w61225;
assign w61227 = ~w61200 & ~w61226;
assign w61228 = ~pi8549 & w61227;
assign w61229 = pi8549 & ~w61227;
assign w61230 = ~w61228 & ~w61229;
assign w61231 = w60455 & w60492;
assign w61232 = ~w60464 & ~w60469;
assign w61233 = ~w60446 & ~w60483;
assign w61234 = ~w60484 & ~w61233;
assign w61235 = ~w60446 & ~w60479;
assign w61236 = w60470 & w60479;
assign w61237 = ~w61235 & ~w61236;
assign w61238 = w61234 & ~w61237;
assign w61239 = ~w60433 & w60495;
assign w61240 = ~w60483 & w64293;
assign w61241 = (w60421 & ~w60484) | (w60421 & w63490) | (~w60484 & w63490);
assign w61242 = ~w61240 & w61241;
assign w61243 = ~w61238 & w61242;
assign w61244 = ~w61239 & w61243;
assign w61245 = ~w60455 & w60496;
assign w61246 = ~w60483 & ~w61245;
assign w61247 = ~w60489 & ~w61246;
assign w61248 = ~w60482 & ~w60488;
assign w61249 = w60455 & ~w61237;
assign w61250 = ~w61248 & w61249;
assign w61251 = ~w60421 & ~w61247;
assign w61252 = ~w61250 & w61251;
assign w61253 = w60427 & w60488;
assign w61254 = w60421 & ~w61253;
assign w61255 = w60446 & w60472;
assign w61256 = ~w61254 & w61255;
assign w61257 = ~w60481 & ~w61231;
assign w61258 = ~w61256 & w61257;
assign w61259 = ~w61232 & w61258;
assign w61260 = (w61259 & w61244) | (w61259 & w64294) | (w61244 & w64294);
assign w61261 = ~pi8594 & w61260;
assign w61262 = pi8594 & ~w61260;
assign w61263 = ~w61261 & ~w61262;
assign w61264 = w60569 & ~w60601;
assign w61265 = ~w60605 & ~w60621;
assign w61266 = w60606 & ~w61265;
assign w61267 = (~w60571 & w61266) | (~w60571 & w64295) | (w61266 & w64295);
assign w61268 = w60555 & ~w60568;
assign w61269 = ~w60583 & ~w60589;
assign w61270 = w60547 & ~w61269;
assign w61271 = w60561 & w61265;
assign w61272 = ~w61270 & w61271;
assign w61273 = w60577 & ~w61268;
assign w61274 = ~w61267 & w61273;
assign w61275 = ~w61272 & w61274;
assign w61276 = ~w60580 & ~w60598;
assign w61277 = w60618 & w61276;
assign w61278 = w60599 & ~w61134;
assign w61279 = w60554 & ~w60561;
assign w61280 = ~w60580 & ~w61279;
assign w61281 = w60589 & ~w61280;
assign w61282 = ~w60602 & ~w60622;
assign w61283 = w60578 & w61282;
assign w61284 = ~w61277 & ~w61281;
assign w61285 = w61283 & w61284;
assign w61286 = ~w61278 & w61285;
assign w61287 = ~w61275 & ~w61286;
assign w61288 = ~w60568 & ~w60581;
assign w61289 = w60619 & w61288;
assign w61290 = ~w61287 & ~w61289;
assign w61291 = ~pi8559 & w61290;
assign w61292 = pi8559 & ~w61290;
assign w61293 = ~w61291 & ~w61292;
assign w61294 = w60480 & w60483;
assign w61295 = ~w60485 & ~w60492;
assign w61296 = ~w60455 & ~w61295;
assign w61297 = ~w60483 & w60493;
assign w61298 = ~w60421 & ~w61294;
assign w61299 = ~w61297 & w61298;
assign w61300 = ~w61296 & w61299;
assign w61301 = ~w61245 & w61254;
assign w61302 = w60469 & w61301;
assign w61303 = ~w61249 & w61302;
assign w61304 = ~w61300 & ~w61303;
assign w61305 = w60427 & w60455;
assign w61306 = ~w60476 & w61305;
assign w61307 = ~w61304 & ~w61306;
assign w61308 = ~pi8575 & w61307;
assign w61309 = pi8575 & ~w61307;
assign w61310 = ~w61308 & ~w61309;
assign w61311 = ~pi7726 & pi9040;
assign w61312 = ~pi7725 & ~pi9040;
assign w61313 = ~w61311 & ~w61312;
assign w61314 = pi5749 & ~w61313;
assign w61315 = ~pi5749 & w61313;
assign w61316 = ~w61314 & ~w61315;
assign w61317 = ~pi7711 & pi9040;
assign w61318 = ~pi7795 & ~pi9040;
assign w61319 = ~w61317 & ~w61318;
assign w61320 = pi5750 & ~w61319;
assign w61321 = ~pi5750 & w61319;
assign w61322 = ~w61320 & ~w61321;
assign w61323 = w61316 & w61322;
assign w61324 = ~pi7749 & pi9040;
assign w61325 = ~pi7659 & ~pi9040;
assign w61326 = ~w61324 & ~w61325;
assign w61327 = pi5888 & ~w61326;
assign w61328 = ~pi5888 & w61326;
assign w61329 = ~w61327 & ~w61328;
assign w61330 = ~pi7653 & pi9040;
assign w61331 = ~pi7711 & ~pi9040;
assign w61332 = ~w61330 & ~w61331;
assign w61333 = pi5748 & ~w61332;
assign w61334 = ~pi5748 & w61332;
assign w61335 = ~w61333 & ~w61334;
assign w61336 = ~w61329 & w61335;
assign w61337 = w61323 & w61336;
assign w61338 = w61329 & w61335;
assign w61339 = ~w61316 & ~w61335;
assign w61340 = ~w61338 & ~w61339;
assign w61341 = w61329 & ~w61335;
assign w61342 = w61316 & ~w61322;
assign w61343 = ~w61329 & ~w61335;
assign w61344 = w61342 & w61343;
assign w61345 = ~pi7666 & pi9040;
assign w61346 = ~pi7663 & ~pi9040;
assign w61347 = ~w61345 & ~w61346;
assign w61348 = pi5692 & ~w61347;
assign w61349 = ~pi5692 & w61347;
assign w61350 = ~w61348 & ~w61349;
assign w61351 = ~w61344 & w61350;
assign w61352 = w61323 & w61335;
assign w61353 = w61351 & ~w61352;
assign w61354 = w61323 & ~w61335;
assign w61355 = w61322 & ~w61329;
assign w61356 = ~w61342 & ~w61355;
assign w61357 = ~w61354 & ~w61356;
assign w61358 = (~w61341 & ~w61353) | (~w61341 & w63491) | (~w61353 & w63491);
assign w61359 = ~w61316 & w61322;
assign w61360 = w61341 & w61359;
assign w61361 = w61351 & ~w61360;
assign w61362 = w61335 & w61359;
assign w61363 = ~w61329 & ~w61350;
assign w61364 = ~w61362 & ~w61363;
assign w61365 = ~pi7662 & pi9040;
assign w61366 = ~pi7670 & ~pi9040;
assign w61367 = ~w61365 & ~w61366;
assign w61368 = pi5585 & ~w61367;
assign w61369 = ~pi5585 & w61367;
assign w61370 = ~w61368 & ~w61369;
assign w61371 = ~w61364 & ~w61370;
assign w61372 = (~w61371 & w61358) | (~w61371 & w64296) | (w61358 & w64296);
assign w61373 = ~w61340 & ~w61372;
assign w61374 = ~w61340 & ~w61362;
assign w61375 = ~w61342 & w61374;
assign w61376 = w61353 & ~w61375;
assign w61377 = ~w61316 & w61336;
assign w61378 = (~w61350 & ~w61323) | (~w61350 & w64297) | (~w61323 & w64297);
assign w61379 = ~w61377 & w61378;
assign w61380 = w61338 & w61342;
assign w61381 = w61335 & w61355;
assign w61382 = ~w61380 & ~w61381;
assign w61383 = (~w61376 & w64298) | (~w61376 & w64299) | (w64298 & w64299);
assign w61384 = w61316 & w61329;
assign w61385 = ~w61350 & w61384;
assign w61386 = ~w61335 & w61385;
assign w61387 = ~w61322 & w61350;
assign w61388 = w61336 & w61387;
assign w61389 = w61316 & w61335;
assign w61390 = ~w61338 & ~w61342;
assign w61391 = ~w61350 & ~w61389;
assign w61392 = ~w61390 & w61391;
assign w61393 = ~w61388 & ~w61392;
assign w61394 = ~w61370 & ~w61393;
assign w61395 = ~w61337 & ~w61386;
assign w61396 = ~w61394 & w61395;
assign w61397 = ~w61383 & w61396;
assign w61398 = ~w61373 & w61397;
assign w61399 = pi8547 & w61398;
assign w61400 = ~pi8547 & ~w61398;
assign w61401 = ~w61399 & ~w61400;
assign w61402 = w61254 & ~w61255;
assign w61403 = ~w60470 & w61234;
assign w61404 = ~w60459 & ~w61253;
assign w61405 = (w61404 & ~w61234) | (w61404 & w64300) | (~w61234 & w64300);
assign w61406 = w60487 & ~w61239;
assign w61407 = ~w61405 & w61406;
assign w61408 = ~w61402 & ~w61407;
assign w61409 = ~w60439 & ~w61403;
assign w61410 = w60421 & ~w60486;
assign w61411 = ~w60494 & w61410;
assign w61412 = ~w61409 & w61411;
assign w61413 = ~w61408 & ~w61412;
assign w61414 = ~pi8615 & w61413;
assign w61415 = pi8615 & ~w61413;
assign w61416 = ~w61414 & ~w61415;
assign w61417 = ~w60859 & w61082;
assign w61418 = w60830 & ~w61417;
assign w61419 = w60838 & ~w61418;
assign w61420 = w60786 & w61062;
assign w61421 = w60805 & w61079;
assign w61422 = w61078 & ~w61421;
assign w61423 = ~w61420 & ~w61422;
assign w61424 = w61077 & ~w61423;
assign w61425 = ~w61419 & ~w61424;
assign w61426 = ~w60819 & w60857;
assign w61427 = w60818 & ~w60839;
assign w61428 = ~w60875 & w60879;
assign w61429 = ~w60856 & ~w61426;
assign w61430 = ~w61428 & w61429;
assign w61431 = ~w61427 & w61430;
assign w61432 = w60799 & ~w61431;
assign w61433 = ~w61425 & ~w61432;
assign w61434 = pi8583 & w61433;
assign w61435 = ~pi8583 & ~w61433;
assign w61436 = ~w61434 & ~w61435;
assign w61437 = w61199 & ~w61202;
assign w61438 = ~w61187 & w61437;
assign w61439 = ~w61177 & ~w61218;
assign w61440 = w61438 & ~w61439;
assign w61441 = w61168 & ~w61199;
assign w61442 = ~w61162 & w61441;
assign w61443 = ~w61177 & ~w61442;
assign w61444 = ~w61161 & ~w61199;
assign w61445 = ~w61168 & w61174;
assign w61446 = w61444 & w61445;
assign w61447 = (~w61446 & ~w61207) | (~w61446 & w64301) | (~w61207 & w64301);
assign w61448 = ~w61443 & ~w61447;
assign w61449 = ~w61155 & ~w61444;
assign w61450 = w61188 & ~w61449;
assign w61451 = w61204 & w61442;
assign w61452 = w61162 & w61445;
assign w61453 = ~w61155 & w61168;
assign w61454 = w61161 & w61199;
assign w61455 = ~w61453 & w61454;
assign w61456 = w61185 & ~w61452;
assign w61457 = ~w61455 & w61456;
assign w61458 = ~w61450 & ~w61451;
assign w61459 = w61457 & w61458;
assign w61460 = ~w61448 & w61459;
assign w61461 = w61161 & ~w61174;
assign w61462 = ~w61186 & ~w61461;
assign w61463 = (~w61168 & w61186) | (~w61168 & w64302) | (w61186 & w64302);
assign w61464 = w61441 & ~w61451;
assign w61465 = w61219 & w61438;
assign w61466 = w61438 & w64303;
assign w61467 = ~w61185 & ~w61463;
assign w61468 = ~w61464 & w61467;
assign w61469 = w61447 & ~w61466;
assign w61470 = w61468 & w61469;
assign w61471 = ~w61460 & ~w61470;
assign w61472 = ~w61440 & ~w61471;
assign w61473 = pi8600 & ~w61472;
assign w61474 = ~pi8600 & w61472;
assign w61475 = ~w61473 & ~w61474;
assign w61476 = w60941 & w61107;
assign w61477 = w60941 & ~w60964;
assign w61478 = (~w60971 & w64304) | (~w60971 & w64305) | (w64304 & w64305);
assign w61479 = w60975 & w60988;
assign w61480 = ~w60992 & ~w61479;
assign w61481 = ~w61002 & w61480;
assign w61482 = ~w61478 & w61481;
assign w61483 = w60955 & ~w61482;
assign w61484 = ~w60928 & ~w60971;
assign w61485 = ~w60990 & ~w61003;
assign w61486 = ~w61484 & w61485;
assign w61487 = ~w60955 & ~w61486;
assign w61488 = ~w60996 & ~w61476;
assign w61489 = ~w61487 & w61488;
assign w61490 = w61489 & w64306;
assign w61491 = (~pi8528 & ~w61489) | (~pi8528 & w64307) | (~w61489 & w64307);
assign w61492 = ~w61490 & ~w61491;
assign w61493 = w60570 & ~w61123;
assign w61494 = ~w60613 & w61136;
assign w61495 = ~w60561 & ~w60622;
assign w61496 = ~w61493 & w61495;
assign w61497 = ~w61494 & w61496;
assign w61498 = w60561 & ~w60603;
assign w61499 = ~w61268 & w61498;
assign w61500 = ~w61497 & ~w61499;
assign w61501 = w60548 & w60562;
assign w61502 = ~w61126 & ~w61279;
assign w61503 = w60605 & ~w61502;
assign w61504 = w60577 & ~w61503;
assign w61505 = ~w61270 & w61504;
assign w61506 = ~w61501 & w61505;
assign w61507 = w60570 & w60621;
assign w61508 = ~w60577 & ~w61507;
assign w61509 = ~w61139 & w61508;
assign w61510 = ~w61506 & ~w61509;
assign w61511 = ~w61500 & ~w61510;
assign w61512 = ~pi8678 & w61511;
assign w61513 = pi8678 & ~w61511;
assign w61514 = ~w61512 & ~w61513;
assign w61515 = w61341 & w61342;
assign w61516 = ~w61350 & w61515;
assign w61517 = ~w61339 & ~w61384;
assign w61518 = ~w61342 & ~w61359;
assign w61519 = ~w61517 & w61518;
assign w61520 = w61374 & ~w61519;
assign w61521 = w61356 & w61520;
assign w61522 = (w61382 & ~w61520) | (w61382 & w64308) | (~w61520 & w64308);
assign w61523 = w61353 & ~w61522;
assign w61524 = ~w61316 & ~w61322;
assign w61525 = w61343 & w61524;
assign w61526 = ~w61354 & ~w61525;
assign w61527 = w61350 & ~w61526;
assign w61528 = w61316 & w61363;
assign w61529 = w61370 & ~w61528;
assign w61530 = ~w61527 & w61529;
assign w61531 = ~w61521 & w61530;
assign w61532 = w61341 & w61524;
assign w61533 = ~w61341 & w61359;
assign w61534 = w61378 & ~w61533;
assign w61535 = ~w61353 & ~w61534;
assign w61536 = ~w61370 & ~w61377;
assign w61537 = ~w61380 & ~w61532;
assign w61538 = w61536 & w61537;
assign w61539 = ~w61535 & w61538;
assign w61540 = ~w61531 & ~w61539;
assign w61541 = ~w61516 & ~w61523;
assign w61542 = ~w61540 & w61541;
assign w61543 = pi8548 & ~w61542;
assign w61544 = ~pi8548 & w61542;
assign w61545 = ~w61543 & ~w61544;
assign w61546 = ~w61176 & ~w61452;
assign w61547 = w61185 & w61546;
assign w61548 = w61199 & ~w61445;
assign w61549 = w61201 & ~w61202;
assign w61550 = ~w61548 & ~w61549;
assign w61551 = ~w61438 & ~w61550;
assign w61552 = ~w61155 & w61461;
assign w61553 = ~w61168 & w61552;
assign w61554 = w61547 & ~w61553;
assign w61555 = w61554 & w64309;
assign w61556 = ~w61189 & ~w61552;
assign w61557 = w61546 & w61556;
assign w61558 = w61437 & w61557;
assign w61559 = w61445 & w61449;
assign w61560 = ~w61185 & ~w61559;
assign w61561 = ~w61558 & w61560;
assign w61562 = ~w61555 & ~w61561;
assign w61563 = ~w61212 & w61557;
assign w61564 = ~w61199 & ~w61547;
assign w61565 = ~w61563 & w61564;
assign w61566 = ~w61562 & ~w61565;
assign w61567 = pi8585 & w61566;
assign w61568 = ~pi8585 & ~w61566;
assign w61569 = ~w61567 & ~w61568;
assign w61570 = w60964 & w61007;
assign w61571 = ~w60965 & w64310;
assign w61572 = ~w60928 & w61096;
assign w61573 = w60976 & w60980;
assign w61574 = ~w60994 & ~w61573;
assign w61575 = ~w61571 & w61574;
assign w61576 = ~w61572 & w61575;
assign w61577 = w61480 & w61576;
assign w61578 = ~w60955 & ~w61577;
assign w61579 = ~w60970 & ~w60999;
assign w61580 = (w60955 & w60970) | (w60955 & w64311) | (w60970 & w64311);
assign w61581 = w60940 & w60999;
assign w61582 = ~w61109 & ~w61581;
assign w61583 = ~w61580 & w61582;
assign w61584 = w60928 & ~w61583;
assign w61585 = ~w60964 & w61005;
assign w61586 = w61579 & w61585;
assign w61587 = ~w61570 & ~w61586;
assign w61588 = ~w61584 & w61587;
assign w61589 = ~w61578 & w61588;
assign w61590 = pi8582 & w61589;
assign w61591 = ~pi8582 & ~w61589;
assign w61592 = ~w61590 & ~w61591;
assign w61593 = (w61350 & ~w61336) | (w61350 & w64312) | (~w61336 & w64312);
assign w61594 = ~w61519 & w61593;
assign w61595 = w61340 & w61356;
assign w61596 = ~w61337 & ~w61350;
assign w61597 = ~w61344 & w61596;
assign w61598 = ~w61595 & w61597;
assign w61599 = (~w61594 & ~w61598) | (~w61594 & w63494) | (~w61598 & w63494);
assign w61600 = ~w61370 & ~w61599;
assign w61601 = ~w61322 & ~w61389;
assign w61602 = w61594 & ~w61601;
assign w61603 = w61323 & w61343;
assign w61604 = w61352 & w61385;
assign w61605 = w61336 & w61342;
assign w61606 = ~w61362 & ~w61525;
assign w61607 = w61363 & ~w61606;
assign w61608 = w61370 & ~w61515;
assign w61609 = ~w61603 & ~w61605;
assign w61610 = ~w61604 & w61608;
assign w61611 = w61609 & w61610;
assign w61612 = ~w61607 & w61611;
assign w61613 = ~w61602 & w61612;
assign w61614 = ~w61600 & ~w61613;
assign w61615 = ~w61532 & ~w61605;
assign w61616 = w61350 & ~w61615;
assign w61617 = ~w61350 & w61521;
assign w61618 = ~w61616 & ~w61617;
assign w61619 = ~w61614 & w64313;
assign w61620 = (pi8601 & w61614) | (pi8601 & w64314) | (w61614 & w64314);
assign w61621 = ~w61619 & ~w61620;
assign w61622 = w61202 & w61214;
assign w61623 = ~w61219 & ~w61461;
assign w61624 = ~w61220 & w61623;
assign w61625 = w61199 & ~w61462;
assign w61626 = w61185 & ~w61625;
assign w61627 = ~w61624 & w61626;
assign w61628 = ~w61201 & ~w61443;
assign w61629 = ~w61187 & w61216;
assign w61630 = ~w61188 & w61209;
assign w61631 = ~w61629 & w61630;
assign w61632 = ~w61628 & w61631;
assign w61633 = ~w61627 & ~w61632;
assign w61634 = ~w61465 & ~w61622;
assign w61635 = ~w61633 & w61634;
assign w61636 = ~pi8624 & ~w61635;
assign w61637 = pi8624 & w61635;
assign w61638 = ~w61636 & ~w61637;
assign w61639 = ~w61350 & w61362;
assign w61640 = w61350 & w61517;
assign w61641 = w61518 & w61640;
assign w61642 = ~w61337 & w61608;
assign w61643 = ~w61639 & w61642;
assign w61644 = ~w61641 & w61643;
assign w61645 = ~w61350 & ~w61357;
assign w61646 = ~w61358 & ~w61515;
assign w61647 = ~w61370 & ~w61645;
assign w61648 = ~w61646 & w61647;
assign w61649 = ~w61526 & ~w61603;
assign w61650 = ~w61350 & ~w61605;
assign w61651 = ~w61649 & w61650;
assign w61652 = ~w61361 & ~w61651;
assign w61653 = (~w61652 & w61648) | (~w61652 & w64315) | (w61648 & w64315);
assign w61654 = ~pi8622 & w61653;
assign w61655 = pi8622 & ~w61653;
assign w61656 = ~w61654 & ~w61655;
assign w61657 = ~pi7979 & pi9040;
assign w61658 = ~pi7999 & ~pi9040;
assign w61659 = ~w61657 & ~w61658;
assign w61660 = pi8803 & ~w61659;
assign w61661 = ~pi8803 & w61659;
assign w61662 = ~w61660 & ~w61661;
assign w61663 = ~pi7940 & pi9040;
assign w61664 = ~pi7997 & ~pi9040;
assign w61665 = ~w61663 & ~w61664;
assign w61666 = pi8727 & ~w61665;
assign w61667 = ~pi8727 & w61665;
assign w61668 = ~w61666 & ~w61667;
assign w61669 = w61662 & ~w61668;
assign w61670 = ~pi7978 & pi9040;
assign w61671 = ~pi7942 & ~pi9040;
assign w61672 = ~w61670 & ~w61671;
assign w61673 = pi8748 & ~w61672;
assign w61674 = ~pi8748 & w61672;
assign w61675 = ~w61673 & ~w61674;
assign w61676 = ~pi8033 & pi9040;
assign w61677 = ~pi7954 & ~pi9040;
assign w61678 = ~w61676 & ~w61677;
assign w61679 = pi8738 & ~w61678;
assign w61680 = ~pi8738 & w61678;
assign w61681 = ~w61679 & ~w61680;
assign w61682 = w61675 & w61681;
assign w61683 = w61669 & w61682;
assign w61684 = ~w61668 & ~w61675;
assign w61685 = ~pi8028 & pi9040;
assign w61686 = ~pi8004 & ~pi9040;
assign w61687 = ~w61685 & ~w61686;
assign w61688 = pi8742 & ~w61687;
assign w61689 = ~pi8742 & w61687;
assign w61690 = ~w61688 & ~w61689;
assign w61691 = ~w61681 & w61690;
assign w61692 = w61684 & w61691;
assign w61693 = w61675 & w61690;
assign w61694 = w61668 & w61693;
assign w61695 = w61693 & w63495;
assign w61696 = ~w61692 & ~w61695;
assign w61697 = w61668 & w61675;
assign w61698 = ~w61662 & ~w61690;
assign w61699 = ~w61684 & ~w61697;
assign w61700 = w61698 & w61699;
assign w61701 = w61696 & ~w61700;
assign w61702 = ~w61675 & ~w61690;
assign w61703 = ~w61669 & w61702;
assign w61704 = ~w61681 & ~w61703;
assign w61705 = ~w61694 & w61704;
assign w61706 = w61668 & ~w61690;
assign w61707 = w61662 & w61706;
assign w61708 = w61706 & w63496;
assign w61709 = ~w61668 & w61690;
assign w61710 = ~w61706 & ~w61709;
assign w61711 = w61662 & ~w61693;
assign w61712 = w61710 & w61711;
assign w61713 = w61681 & ~w61708;
assign w61714 = ~w61712 & w61713;
assign w61715 = ~w61705 & ~w61714;
assign w61716 = ~pi7991 & pi9040;
assign w61717 = ~pi7958 & ~pi9040;
assign w61718 = ~w61716 & ~w61717;
assign w61719 = pi8802 & ~w61718;
assign w61720 = ~pi8802 & w61718;
assign w61721 = ~w61719 & ~w61720;
assign w61722 = (w61721 & w61715) | (w61721 & w64316) | (w61715 & w64316);
assign w61723 = ~w61662 & w61675;
assign w61724 = w61662 & ~w61675;
assign w61725 = ~w61723 & ~w61724;
assign w61726 = w61690 & w61725;
assign w61727 = w61668 & ~w61693;
assign w61728 = (~w61707 & ~w61726) | (~w61707 & w63497) | (~w61726 & w63497);
assign w61729 = w61684 & ~w61728;
assign w61730 = w61697 & w61698;
assign w61731 = w61675 & w61709;
assign w61732 = (~w61681 & w61712) | (~w61681 & w63498) | (w61712 & w63498);
assign w61733 = ~w61703 & ~w61726;
assign w61734 = w61681 & ~w61700;
assign w61735 = ~w61733 & w61734;
assign w61736 = ~w61730 & ~w61732;
assign w61737 = ~w61735 & w61736;
assign w61738 = ~w61721 & ~w61737;
assign w61739 = ~w61683 & ~w61729;
assign w61740 = ~w61722 & w61739;
assign w61741 = ~w61738 & w61740;
assign w61742 = pi8696 & ~w61741;
assign w61743 = ~pi8696 & w61741;
assign w61744 = ~w61742 & ~w61743;
assign w61745 = (~w61681 & ~w61706) | (~w61681 & w64317) | (~w61706 & w64317);
assign w61746 = w61727 & w61745;
assign w61747 = ~w61681 & ~w61710;
assign w61748 = ~w61704 & ~w61747;
assign w61749 = ~w61728 & w61748;
assign w61750 = w61662 & w61668;
assign w61751 = w61710 & ~w61750;
assign w61752 = w61710 & w63499;
assign w61753 = ~w61723 & ~w61752;
assign w61754 = w61732 & ~w61753;
assign w61755 = w61682 & w61698;
assign w61756 = w61709 & w61724;
assign w61757 = ~w61755 & ~w61756;
assign w61758 = ~w61701 & ~w61757;
assign w61759 = w61721 & ~w61746;
assign w61760 = ~w61749 & w61759;
assign w61761 = ~w61754 & ~w61758;
assign w61762 = w61760 & w61761;
assign w61763 = w61662 & w61747;
assign w61764 = ~w61721 & w61757;
assign w61765 = w61696 & w61764;
assign w61766 = ~w61763 & w61765;
assign w61767 = ~w61762 & ~w61766;
assign w61768 = w61662 & w61702;
assign w61769 = ~w61668 & w61768;
assign w61770 = w61721 & ~w61769;
assign w61771 = w61751 & ~w61770;
assign w61772 = w61681 & ~w61694;
assign w61773 = ~w61771 & w61772;
assign w61774 = w61748 & ~w61773;
assign w61775 = (pi8716 & w61767) | (pi8716 & w64318) | (w61767 & w64318);
assign w61776 = ~w61767 & w64319;
assign w61777 = ~w61775 & ~w61776;
assign w61778 = ~pi7952 & pi9040;
assign w61779 = ~pi8005 & ~pi9040;
assign w61780 = ~w61778 & ~w61779;
assign w61781 = pi8796 & ~w61780;
assign w61782 = ~pi8796 & w61780;
assign w61783 = ~w61781 & ~w61782;
assign w61784 = ~pi7929 & pi9040;
assign w61785 = ~pi7935 & ~pi9040;
assign w61786 = ~w61784 & ~w61785;
assign w61787 = pi8798 & ~w61786;
assign w61788 = ~pi8798 & w61786;
assign w61789 = ~w61787 & ~w61788;
assign w61790 = w61783 & w61789;
assign w61791 = ~pi7975 & pi9040;
assign w61792 = ~pi8034 & ~pi9040;
assign w61793 = ~w61791 & ~w61792;
assign w61794 = pi8715 & ~w61793;
assign w61795 = ~pi8715 & w61793;
assign w61796 = ~w61794 & ~w61795;
assign w61797 = ~pi7972 & pi9040;
assign w61798 = ~pi7974 & ~pi9040;
assign w61799 = ~w61797 & ~w61798;
assign w61800 = pi8719 & ~w61799;
assign w61801 = ~pi8719 & w61799;
assign w61802 = ~w61800 & ~w61801;
assign w61803 = ~w61796 & ~w61802;
assign w61804 = w61790 & w61803;
assign w61805 = ~pi7931 & pi9040;
assign w61806 = ~pi8000 & ~pi9040;
assign w61807 = ~w61805 & ~w61806;
assign w61808 = pi8761 & ~w61807;
assign w61809 = ~pi8761 & w61807;
assign w61810 = ~w61808 & ~w61809;
assign w61811 = w61802 & ~w61810;
assign w61812 = ~w61789 & ~w61796;
assign w61813 = w61811 & w61812;
assign w61814 = ~w61804 & ~w61813;
assign w61815 = ~pi8016 & pi9040;
assign w61816 = ~pi7998 & ~pi9040;
assign w61817 = ~w61815 & ~w61816;
assign w61818 = pi8776 & ~w61817;
assign w61819 = ~pi8776 & w61817;
assign w61820 = ~w61818 & ~w61819;
assign w61821 = ~w61783 & ~w61810;
assign w61822 = w61789 & w61796;
assign w61823 = w61821 & w61822;
assign w61824 = w61783 & ~w61789;
assign w61825 = ~w61802 & w61810;
assign w61826 = ~w61824 & w61825;
assign w61827 = w61783 & w61810;
assign w61828 = ~w61821 & ~w61827;
assign w61829 = ~w61811 & w61828;
assign w61830 = ~w61783 & ~w61789;
assign w61831 = ~w61796 & ~w61830;
assign w61832 = w61829 & w61831;
assign w61833 = ~w61823 & ~w61826;
assign w61834 = ~w61832 & w61833;
assign w61835 = (w61820 & w61832) | (w61820 & w63500) | (w61832 & w63500);
assign w61836 = ~w61783 & w61802;
assign w61837 = ~w61790 & ~w61836;
assign w61838 = ~w61783 & ~w61803;
assign w61839 = ~w61802 & ~w61838;
assign w61840 = w61837 & ~w61839;
assign w61841 = ~w61811 & ~w61825;
assign w61842 = w61830 & ~w61841;
assign w61843 = w61796 & w61810;
assign w61844 = w61824 & w61843;
assign w61845 = ~w61820 & ~w61844;
assign w61846 = ~w61842 & w61845;
assign w61847 = (~w61846 & w61835) | (~w61846 & w64320) | (w61835 & w64320);
assign w61848 = ~w61802 & w61823;
assign w61849 = w61803 & w61827;
assign w61850 = ~w61783 & w61812;
assign w61851 = ~w61825 & w61850;
assign w61852 = w61796 & w61828;
assign w61853 = w61828 & w64321;
assign w61854 = w61802 & w61828;
assign w61855 = w61828 & w64322;
assign w61856 = ~w61853 & ~w61855;
assign w61857 = w61852 & ~w61856;
assign w61858 = ~w61796 & ~w61828;
assign w61859 = ~w61837 & w61858;
assign w61860 = ~w61849 & ~w61851;
assign w61861 = ~w61859 & w61860;
assign w61862 = ~w61857 & w61861;
assign w61863 = ~w61820 & ~w61862;
assign w61864 = w61814 & ~w61848;
assign w61865 = ~w61847 & w61864;
assign w61866 = ~w61863 & w61865;
assign w61867 = pi8754 & ~w61866;
assign w61868 = ~pi8754 & w61866;
assign w61869 = ~w61867 & ~w61868;
assign w61870 = ~pi8001 & pi9040;
assign w61871 = ~pi7965 & ~pi9040;
assign w61872 = ~w61870 & ~w61871;
assign w61873 = pi8705 & ~w61872;
assign w61874 = ~pi8705 & w61872;
assign w61875 = ~w61873 & ~w61874;
assign w61876 = ~pi8003 & pi9040;
assign w61877 = ~pi7991 & ~pi9040;
assign w61878 = ~w61876 & ~w61877;
assign w61879 = pi8719 & ~w61878;
assign w61880 = ~pi8719 & w61878;
assign w61881 = ~w61879 & ~w61880;
assign w61882 = w61875 & ~w61881;
assign w61883 = ~pi7946 & pi9040;
assign w61884 = ~pi7940 & ~pi9040;
assign w61885 = ~w61883 & ~w61884;
assign w61886 = pi8807 & ~w61885;
assign w61887 = ~pi8807 & w61885;
assign w61888 = ~w61886 & ~w61887;
assign w61889 = ~pi7954 & pi9040;
assign w61890 = ~pi7968 & ~pi9040;
assign w61891 = ~w61889 & ~w61890;
assign w61892 = pi8712 & ~w61891;
assign w61893 = ~pi8712 & w61891;
assign w61894 = ~w61892 & ~w61893;
assign w61895 = ~w61888 & w61894;
assign w61896 = ~w61882 & ~w61895;
assign w61897 = w61881 & w61888;
assign w61898 = ~w61875 & w61881;
assign w61899 = ~w61897 & ~w61898;
assign w61900 = w61875 & ~w61894;
assign w61901 = w61888 & w61900;
assign w61902 = w61899 & ~w61901;
assign w61903 = ~w61896 & ~w61902;
assign w61904 = ~w61881 & ~w61888;
assign w61905 = w61888 & w61898;
assign w61906 = ~w61904 & ~w61905;
assign w61907 = ~w61875 & ~w61894;
assign w61908 = ~w61906 & w61907;
assign w61909 = ~w61903 & ~w61908;
assign w61910 = ~pi8015 & pi9040;
assign w61911 = ~pi8013 & ~pi9040;
assign w61912 = ~w61910 & ~w61911;
assign w61913 = pi8766 & ~w61912;
assign w61914 = ~pi8766 & w61912;
assign w61915 = ~w61913 & ~w61914;
assign w61916 = ~w61909 & w61915;
assign w61917 = w61894 & ~w61915;
assign w61918 = ~w61906 & w61917;
assign w61919 = w61882 & w61918;
assign w61920 = ~w61894 & ~w61915;
assign w61921 = ~w61881 & w61888;
assign w61922 = w61920 & w61921;
assign w61923 = ~w61894 & w61915;
assign w61924 = w61898 & w61923;
assign w61925 = ~pi8039 & pi9040;
assign w61926 = ~pi8028 & ~pi9040;
assign w61927 = ~w61925 & ~w61926;
assign w61928 = pi8796 & ~w61927;
assign w61929 = ~pi8796 & w61927;
assign w61930 = ~w61928 & ~w61929;
assign w61931 = ~w61924 & ~w61930;
assign w61932 = w61875 & w61881;
assign w61933 = ~w61875 & w61915;
assign w61934 = ~w61881 & w61933;
assign w61935 = ~w61932 & ~w61934;
assign w61936 = w61888 & w61894;
assign w61937 = w61915 & ~w61936;
assign w61938 = ~w61935 & ~w61937;
assign w61939 = ~w61904 & w61915;
assign w61940 = w61895 & ~w61933;
assign w61941 = ~w61939 & w61940;
assign w61942 = ~w61922 & w61931;
assign w61943 = ~w61941 & w61942;
assign w61944 = ~w61938 & w61943;
assign w61945 = w61897 & w61900;
assign w61946 = ~w61888 & w61907;
assign w61947 = ~w61875 & w61894;
assign w61948 = w61888 & w61947;
assign w61949 = ~w61946 & ~w61948;
assign w61950 = ~w61915 & ~w61949;
assign w61951 = ~w61933 & ~w61939;
assign w61952 = ~w61923 & w61951;
assign w61953 = ~w61896 & ~w61952;
assign w61954 = w61930 & ~w61945;
assign w61955 = ~w61950 & w61954;
assign w61956 = ~w61953 & w61955;
assign w61957 = ~w61944 & ~w61956;
assign w61958 = ~w61916 & ~w61919;
assign w61959 = ~w61957 & w61958;
assign w61960 = ~pi8749 & ~w61959;
assign w61961 = pi8749 & w61959;
assign w61962 = ~w61960 & ~w61961;
assign w61963 = ~pi7968 & pi9040;
assign w61964 = ~pi7978 & ~pi9040;
assign w61965 = ~w61963 & ~w61964;
assign w61966 = pi8742 & ~w61965;
assign w61967 = ~pi8742 & w61965;
assign w61968 = ~w61966 & ~w61967;
assign w61969 = ~pi7999 & pi9040;
assign w61970 = ~pi8001 & ~pi9040;
assign w61971 = ~w61969 & ~w61970;
assign w61972 = pi8752 & ~w61971;
assign w61973 = ~pi8752 & w61971;
assign w61974 = ~w61972 & ~w61973;
assign w61975 = ~pi8004 & pi9040;
assign w61976 = ~pi8003 & ~pi9040;
assign w61977 = ~w61975 & ~w61976;
assign w61978 = pi8799 & ~w61977;
assign w61979 = ~pi8799 & w61977;
assign w61980 = ~w61978 & ~w61979;
assign w61981 = w61974 & w61980;
assign w61982 = ~pi7997 & pi9040;
assign w61983 = ~pi7966 & ~pi9040;
assign w61984 = ~w61982 & ~w61983;
assign w61985 = pi8781 & ~w61984;
assign w61986 = ~pi8781 & w61984;
assign w61987 = ~w61985 & ~w61986;
assign w61988 = ~w61980 & w61987;
assign w61989 = ~pi8013 & pi9040;
assign w61990 = ~pi7961 & ~pi9040;
assign w61991 = ~w61989 & ~w61990;
assign w61992 = pi8702 & ~w61991;
assign w61993 = ~pi8702 & w61991;
assign w61994 = ~w61992 & ~w61993;
assign w61995 = ~w61988 & w61994;
assign w61996 = ~pi7957 & pi9040;
assign w61997 = ~pi7943 & ~pi9040;
assign w61998 = ~w61996 & ~w61997;
assign w61999 = pi8803 & ~w61998;
assign w62000 = ~pi8803 & w61998;
assign w62001 = ~w61999 & ~w62000;
assign w62002 = ~w61974 & ~w61987;
assign w62003 = w61974 & w61987;
assign w62004 = ~w62002 & ~w62003;
assign w62005 = w62001 & w62004;
assign w62006 = ~w61981 & w61995;
assign w62007 = ~w62005 & w62006;
assign w62008 = ~w61974 & w61988;
assign w62009 = w61974 & ~w61987;
assign w62010 = w62001 & w62009;
assign w62011 = ~w62008 & ~w62010;
assign w62012 = ~w61994 & ~w62011;
assign w62013 = w61987 & w61994;
assign w62014 = w61974 & w62001;
assign w62015 = w62013 & w62014;
assign w62016 = ~w61974 & ~w62001;
assign w62017 = w61980 & w62001;
assign w62018 = ~w62016 & ~w62017;
assign w62019 = ~w61980 & ~w62001;
assign w62020 = w61987 & ~w62019;
assign w62021 = w62018 & w62020;
assign w62022 = ~w62015 & ~w62021;
assign w62023 = ~w62007 & ~w62012;
assign w62024 = w62022 & w62023;
assign w62025 = w61968 & ~w62024;
assign w62026 = w61980 & ~w61994;
assign w62027 = w62009 & w62026;
assign w62028 = w61980 & ~w62001;
assign w62029 = w62002 & w62028;
assign w62030 = ~w62014 & w62018;
assign w62031 = ~w62009 & ~w62017;
assign w62032 = w61994 & w62031;
assign w62033 = w62030 & w62032;
assign w62034 = ~w62029 & ~w62033;
assign w62035 = (w61995 & w62033) | (w61995 & w64323) | (w62033 & w64323);
assign w62036 = w61988 & w62014;
assign w62037 = ~w61994 & ~w62009;
assign w62038 = ~w61995 & ~w62001;
assign w62039 = ~w62037 & w62038;
assign w62040 = ~w61980 & ~w61994;
assign w62041 = w62002 & w62040;
assign w62042 = ~w61974 & w61987;
assign w62043 = w62013 & w62016;
assign w62044 = w61980 & w62042;
assign w62045 = ~w62043 & w62044;
assign w62046 = ~w62041 & ~w62045;
assign w62047 = ~w62039 & w62046;
assign w62048 = ~w61968 & ~w62047;
assign w62049 = ~w62027 & ~w62036;
assign w62050 = ~w62035 & w62049;
assign w62051 = ~w62048 & w62050;
assign w62052 = ~w62025 & w62051;
assign w62053 = pi8697 & ~w62052;
assign w62054 = ~pi8697 & w62052;
assign w62055 = ~w62053 & ~w62054;
assign w62056 = ~pi8017 & pi9040;
assign w62057 = ~pi7979 & ~pi9040;
assign w62058 = ~w62056 & ~w62057;
assign w62059 = pi8717 & ~w62058;
assign w62060 = ~pi8717 & w62058;
assign w62061 = ~w62059 & ~w62060;
assign w62062 = ~pi7966 & pi9040;
assign w62063 = ~pi8011 & ~pi9040;
assign w62064 = ~w62062 & ~w62063;
assign w62065 = pi8705 & ~w62064;
assign w62066 = ~pi8705 & w62064;
assign w62067 = ~w62065 & ~w62066;
assign w62068 = w62061 & w62067;
assign w62069 = ~pi8038 & pi9040;
assign w62070 = ~pi8033 & ~pi9040;
assign w62071 = ~w62069 & ~w62070;
assign w62072 = pi8802 & ~w62071;
assign w62073 = ~pi8802 & w62071;
assign w62074 = ~w62072 & ~w62073;
assign w62075 = ~pi7942 & pi9040;
assign w62076 = ~pi7946 & ~pi9040;
assign w62077 = ~w62075 & ~w62076;
assign w62078 = pi8748 & ~w62077;
assign w62079 = ~pi8748 & w62077;
assign w62080 = ~w62078 & ~w62079;
assign w62081 = ~w62074 & ~w62080;
assign w62082 = w62074 & w62080;
assign w62083 = ~w62081 & ~w62082;
assign w62084 = w62068 & w62083;
assign w62085 = ~w62067 & w62074;
assign w62086 = w62080 & w62085;
assign w62087 = w62085 & w63501;
assign w62088 = ~w62084 & ~w62087;
assign w62089 = ~pi7943 & pi9040;
assign w62090 = ~pi8039 & ~pi9040;
assign w62091 = ~w62089 & ~w62090;
assign w62092 = pi8710 & ~w62091;
assign w62093 = ~pi8710 & w62091;
assign w62094 = ~w62092 & ~w62093;
assign w62095 = (~w62094 & w62084) | (~w62094 & w64324) | (w62084 & w64324);
assign w62096 = w62067 & ~w62074;
assign w62097 = ~w62085 & ~w62096;
assign w62098 = w62061 & ~w62080;
assign w62099 = ~w62061 & ~w62081;
assign w62100 = ~w62061 & ~w62080;
assign w62101 = ~w62097 & w62100;
assign w62102 = w62067 & w62080;
assign w62103 = ~w62100 & ~w62102;
assign w62104 = ~w62067 & ~w62080;
assign w62105 = w62097 & ~w62104;
assign w62106 = w62103 & w62105;
assign w62107 = ~w62101 & ~w62106;
assign w62108 = w62099 & ~w62107;
assign w62109 = ~w62102 & ~w62104;
assign w62110 = ~w62094 & ~w62109;
assign w62111 = w62061 & ~w62074;
assign w62112 = w62080 & w62111;
assign w62113 = (~w62094 & ~w62111) | (~w62094 & w63502) | (~w62111 & w63502);
assign w62114 = ~w62099 & ~w62113;
assign w62115 = w62096 & w62114;
assign w62116 = ~pi7958 & pi9040;
assign w62117 = ~pi7937 & ~pi9040;
assign w62118 = ~w62116 & ~w62117;
assign w62119 = pi8712 & ~w62118;
assign w62120 = ~pi8712 & w62118;
assign w62121 = ~w62119 & ~w62120;
assign w62122 = (~w62121 & ~w62097) | (~w62121 & w64325) | (~w62097 & w64325);
assign w62123 = ~w62110 & w62122;
assign w62124 = ~w62095 & w62123;
assign w62125 = ~w62115 & w62124;
assign w62126 = ~w62108 & w62125;
assign w62127 = w62061 & ~w62067;
assign w62128 = w62083 & w62127;
assign w62129 = ~w62061 & w62067;
assign w62130 = w62083 & w62129;
assign w62131 = ~w62067 & w62100;
assign w62132 = ~w62074 & w62131;
assign w62133 = ~w62082 & ~w62132;
assign w62134 = w62094 & ~w62133;
assign w62135 = w62068 & w62081;
assign w62136 = w62121 & ~w62135;
assign w62137 = w62085 & ~w62100;
assign w62138 = ~w62074 & ~w62103;
assign w62139 = w62113 & ~w62137;
assign w62140 = ~w62138 & w62139;
assign w62141 = w62088 & w62140;
assign w62142 = w62121 & ~w62141;
assign w62143 = (~w62136 & w62141) | (~w62136 & w64326) | (w62141 & w64326);
assign w62144 = ~w62128 & ~w62130;
assign w62145 = ~w62134 & w62144;
assign w62146 = ~w62143 & w62145;
assign w62147 = ~w62126 & ~w62146;
assign w62148 = pi8788 & w62147;
assign w62149 = ~pi8788 & ~w62147;
assign w62150 = ~w62148 & ~w62149;
assign w62151 = w62074 & w62094;
assign w62152 = ~w62085 & ~w62151;
assign w62153 = w62100 & ~w62152;
assign w62154 = w62104 & w62111;
assign w62155 = ~w62086 & ~w62154;
assign w62156 = ~w62094 & ~w62155;
assign w62157 = w62068 & w62082;
assign w62158 = ~w62121 & ~w62157;
assign w62159 = ~w62061 & w62074;
assign w62160 = ~w62111 & ~w62159;
assign w62161 = w62067 & w62160;
assign w62162 = ~w62114 & w62161;
assign w62163 = ~w62153 & w62158;
assign w62164 = ~w62156 & w62163;
assign w62165 = ~w62162 & w62164;
assign w62166 = ~w62061 & w62102;
assign w62167 = ~w62098 & ~w62166;
assign w62168 = w62151 & ~w62167;
assign w62169 = (~w62094 & w62115) | (~w62094 & w64327) | (w62115 & w64327);
assign w62170 = ~w62132 & w62136;
assign w62171 = ~w62168 & w62170;
assign w62172 = ~w62169 & w62171;
assign w62173 = ~w62165 & ~w62172;
assign w62174 = w62080 & w62160;
assign w62175 = ~w62094 & ~w62174;
assign w62176 = w62094 & ~w62135;
assign w62177 = ~w62128 & ~w62131;
assign w62178 = w62176 & w62177;
assign w62179 = ~w62175 & ~w62178;
assign w62180 = ~w62173 & ~w62179;
assign w62181 = ~pi8709 & w62180;
assign w62182 = pi8709 & ~w62180;
assign w62183 = ~w62181 & ~w62182;
assign w62184 = ~pi7971 & pi9040;
assign w62185 = ~pi8025 & ~pi9040;
assign w62186 = ~w62184 & ~w62185;
assign w62187 = pi8773 & ~w62186;
assign w62188 = ~pi8773 & w62186;
assign w62189 = ~w62187 & ~w62188;
assign w62190 = ~pi7949 & pi9040;
assign w62191 = ~pi8036 & ~pi9040;
assign w62192 = ~w62190 & ~w62191;
assign w62193 = pi8772 & ~w62192;
assign w62194 = ~pi8772 & w62192;
assign w62195 = ~w62193 & ~w62194;
assign w62196 = ~pi7959 & pi9040;
assign w62197 = ~pi8023 & ~pi9040;
assign w62198 = ~w62196 & ~w62197;
assign w62199 = pi8778 & ~w62198;
assign w62200 = ~pi8778 & w62198;
assign w62201 = ~w62199 & ~w62200;
assign w62202 = ~pi8010 & pi9040;
assign w62203 = ~pi7972 & ~pi9040;
assign w62204 = ~w62202 & ~w62203;
assign w62205 = pi8775 & ~w62204;
assign w62206 = ~pi8775 & w62204;
assign w62207 = ~w62205 & ~w62206;
assign w62208 = ~w62201 & w62207;
assign w62209 = ~pi7998 & pi9040;
assign w62210 = ~pi8022 & ~pi9040;
assign w62211 = ~w62209 & ~w62210;
assign w62212 = pi8781 & ~w62211;
assign w62213 = ~pi8781 & w62211;
assign w62214 = ~w62212 & ~w62213;
assign w62215 = ~w62208 & ~w62214;
assign w62216 = w62201 & ~w62207;
assign w62217 = w62195 & ~w62216;
assign w62218 = w62215 & w62217;
assign w62219 = ~w62189 & w62218;
assign w62220 = ~w62207 & w62214;
assign w62221 = ~w62195 & ~w62201;
assign w62222 = w62189 & w62221;
assign w62223 = w62220 & w62222;
assign w62224 = w62207 & ~w62214;
assign w62225 = w62189 & w62195;
assign w62226 = w62224 & w62225;
assign w62227 = ~w62201 & w62226;
assign w62228 = w62216 & w62225;
assign w62229 = w62189 & ~w62207;
assign w62230 = ~w62189 & w62207;
assign w62231 = ~w62229 & ~w62230;
assign w62232 = w62195 & ~w62224;
assign w62233 = ~w62220 & w62232;
assign w62234 = w62231 & w62233;
assign w62235 = ~w62189 & ~w62195;
assign w62236 = ~w62189 & w62208;
assign w62237 = ~w62235 & ~w62236;
assign w62238 = w62214 & ~w62237;
assign w62239 = ~pi7963 & pi9040;
assign w62240 = ~pi7952 & ~pi9040;
assign w62241 = ~w62239 & ~w62240;
assign w62242 = pi8752 & ~w62241;
assign w62243 = ~pi8752 & w62241;
assign w62244 = ~w62242 & ~w62243;
assign w62245 = ~w62189 & ~w62214;
assign w62246 = ~w62207 & w62245;
assign w62247 = ~w62201 & w62246;
assign w62248 = w62201 & ~w62214;
assign w62249 = ~w62195 & w62207;
assign w62250 = ~w62229 & ~w62249;
assign w62251 = w62248 & ~w62250;
assign w62252 = ~w62228 & ~w62244;
assign w62253 = ~w62247 & w62252;
assign w62254 = ~w62251 & w62253;
assign w62255 = ~w62234 & ~w62238;
assign w62256 = w62254 & w62255;
assign w62257 = w62221 & ~w62231;
assign w62258 = w62244 & ~w62257;
assign w62259 = w62189 & w62214;
assign w62260 = ~w62208 & ~w62216;
assign w62261 = w62259 & w62260;
assign w62262 = w62195 & w62220;
assign w62263 = ~w62195 & w62248;
assign w62264 = w62231 & w62263;
assign w62265 = ~w62262 & ~w62264;
assign w62266 = ~w62189 & ~w62265;
assign w62267 = ~w62226 & ~w62261;
assign w62268 = w62258 & w62267;
assign w62269 = ~w62266 & w62268;
assign w62270 = ~w62256 & ~w62269;
assign w62271 = ~w62223 & ~w62227;
assign w62272 = ~w62219 & w62271;
assign w62273 = ~w62270 & w62272;
assign w62274 = pi8695 & ~w62273;
assign w62275 = ~pi8695 & w62273;
assign w62276 = ~w62274 & ~w62275;
assign w62277 = w61987 & w62028;
assign w62278 = ~w61974 & w62001;
assign w62279 = ~w61987 & w62278;
assign w62280 = ~w62277 & ~w62279;
assign w62281 = ~w62018 & ~w62280;
assign w62282 = ~w61994 & w62281;
assign w62283 = ~w62021 & w63503;
assign w62284 = (w61994 & ~w61988) | (w61994 & w64328) | (~w61988 & w64328);
assign w62285 = ~w62002 & ~w62017;
assign w62286 = ~w62278 & ~w62285;
assign w62287 = w62284 & ~w62286;
assign w62288 = ~w62001 & ~w62033;
assign w62289 = w62287 & ~w62288;
assign w62290 = ~w61994 & ~w62036;
assign w62291 = w62280 & w62290;
assign w62292 = w62040 & w62278;
assign w62293 = ~w62041 & ~w62292;
assign w62294 = w62291 & ~w62293;
assign w62295 = w62009 & ~w62017;
assign w62296 = ~w62019 & w62295;
assign w62297 = ~w62283 & ~w62296;
assign w62298 = ~w62294 & w62297;
assign w62299 = ~w62289 & w62298;
assign w62300 = w61968 & ~w62299;
assign w62301 = ~w62029 & ~w62283;
assign w62302 = w62284 & ~w62301;
assign w62303 = ~w61987 & w62017;
assign w62304 = ~w62019 & ~w62303;
assign w62305 = w62004 & ~w62304;
assign w62306 = w62291 & ~w62305;
assign w62307 = (~w61968 & w62286) | (~w61968 & w64329) | (w62286 & w64329);
assign w62308 = ~w62306 & w62307;
assign w62309 = ~w62282 & ~w62308;
assign w62310 = ~w62302 & w62309;
assign w62311 = ~w62300 & w62310;
assign w62312 = pi8793 & ~w62311;
assign w62313 = ~pi8793 & w62311;
assign w62314 = ~w62312 & ~w62313;
assign w62315 = w62295 & w64330;
assign w62316 = ~w62033 & ~w62315;
assign w62317 = ~w62284 & ~w62316;
assign w62318 = w62007 & w62009;
assign w62319 = ~w61994 & w62005;
assign w62320 = ~w62004 & w62028;
assign w62321 = (~w61968 & ~w61988) | (~w61968 & w64331) | (~w61988 & w64331);
assign w62322 = ~w62015 & ~w62292;
assign w62323 = w62321 & w62322;
assign w62324 = ~w62320 & w62323;
assign w62325 = ~w62319 & w62324;
assign w62326 = ~w62318 & w62325;
assign w62327 = ~w62004 & w62019;
assign w62328 = ~w62010 & ~w62327;
assign w62329 = w61995 & ~w62328;
assign w62330 = w61974 & w62040;
assign w62331 = w61968 & ~w62330;
assign w62332 = ~w62281 & w62331;
assign w62333 = ~w62329 & w62332;
assign w62334 = ~w62326 & ~w62333;
assign w62335 = w61980 & w61994;
assign w62336 = ~w62280 & w62335;
assign w62337 = ~w62317 & ~w62336;
assign w62338 = (~pi8744 & w62334) | (~pi8744 & w64332) | (w62334 & w64332);
assign w62339 = ~w62334 & w64333;
assign w62340 = ~w62338 & ~w62339;
assign w62341 = w62094 & w62154;
assign w62342 = ~w62084 & w63504;
assign w62343 = w62097 & w62099;
assign w62344 = ~w62061 & w62094;
assign w62345 = w62097 & w62344;
assign w62346 = (~w62345 & w62342) | (~w62345 & w64334) | (w62342 & w64334);
assign w62347 = ~w62154 & ~w62346;
assign w62348 = ~w62121 & ~w62347;
assign w62349 = w62342 & ~w62343;
assign w62350 = ~w62095 & ~w62341;
assign w62351 = (w62350 & ~w62142) | (w62350 & w64335) | (~w62142 & w64335);
assign w62352 = ~w62348 & w62351;
assign w62353 = pi8718 & w62352;
assign w62354 = ~pi8718 & ~w62352;
assign w62355 = ~w62353 & ~w62354;
assign w62356 = ~pi8000 & pi9040;
assign w62357 = ~pi7971 & ~pi9040;
assign w62358 = ~w62356 & ~w62357;
assign w62359 = pi8726 & ~w62358;
assign w62360 = ~pi8726 & w62358;
assign w62361 = ~w62359 & ~w62360;
assign w62362 = ~pi8023 & pi9040;
assign w62363 = ~pi8016 & ~pi9040;
assign w62364 = ~w62362 & ~w62363;
assign w62365 = pi8761 & ~w62364;
assign w62366 = ~pi8761 & w62364;
assign w62367 = ~w62365 & ~w62366;
assign w62368 = ~pi8005 & pi9040;
assign w62369 = ~pi8010 & ~pi9040;
assign w62370 = ~w62368 & ~w62369;
assign w62371 = pi8743 & ~w62370;
assign w62372 = ~pi8743 & w62370;
assign w62373 = ~w62371 & ~w62372;
assign w62374 = ~w62367 & w62373;
assign w62375 = ~pi8022 & pi9040;
assign w62376 = ~pi7986 & ~pi9040;
assign w62377 = ~w62375 & ~w62376;
assign w62378 = pi8776 & ~w62377;
assign w62379 = ~pi8776 & w62377;
assign w62380 = ~w62378 & ~w62379;
assign w62381 = ~w62374 & ~w62380;
assign w62382 = ~pi8030 & pi9040;
assign w62383 = ~pi7975 & ~pi9040;
assign w62384 = ~w62382 & ~w62383;
assign w62385 = pi8750 & ~w62384;
assign w62386 = ~pi8750 & w62384;
assign w62387 = ~w62385 & ~w62386;
assign w62388 = w62367 & ~w62387;
assign w62389 = w62367 & ~w62373;
assign w62390 = ~w62380 & ~w62387;
assign w62391 = ~w62389 & ~w62390;
assign w62392 = w62388 & w62391;
assign w62393 = ~w62380 & ~w62388;
assign w62394 = ~w62392 & ~w62393;
assign w62395 = ~w62381 & ~w62394;
assign w62396 = w62374 & ~w62387;
assign w62397 = w62380 & w62387;
assign w62398 = ~w62367 & w62397;
assign w62399 = (w62380 & ~w62397) | (w62380 & w64336) | (~w62397 & w64336);
assign w62400 = ~w62380 & w62387;
assign w62401 = ~w62367 & w62400;
assign w62402 = ~w62399 & ~w62401;
assign w62403 = ~pi8036 & pi9040;
assign w62404 = ~pi8007 & ~pi9040;
assign w62405 = ~w62403 & ~w62404;
assign w62406 = pi8713 & ~w62405;
assign w62407 = ~pi8713 & w62405;
assign w62408 = ~w62406 & ~w62407;
assign w62409 = ~w62396 & ~w62408;
assign w62410 = ~w62402 & w62409;
assign w62411 = ~w62395 & ~w62410;
assign w62412 = ~w62361 & ~w62411;
assign w62413 = ~w62373 & w62390;
assign w62414 = w62367 & w62400;
assign w62415 = ~w62413 & ~w62414;
assign w62416 = ~w62361 & ~w62415;
assign w62417 = w62361 & w62367;
assign w62418 = w62397 & w62417;
assign w62419 = w62373 & w62387;
assign w62420 = w62380 & w62419;
assign w62421 = w62389 & w62390;
assign w62422 = w62361 & ~w62420;
assign w62423 = ~w62421 & w62422;
assign w62424 = w62394 & w62423;
assign w62425 = w62374 & w62400;
assign w62426 = ~w62367 & ~w62373;
assign w62427 = w62397 & w62426;
assign w62428 = w62408 & ~w62418;
assign w62429 = ~w62425 & ~w62427;
assign w62430 = w62428 & w62429;
assign w62431 = ~w62416 & w62430;
assign w62432 = ~w62424 & w62431;
assign w62433 = w62374 & w62397;
assign w62434 = ~w62408 & ~w62433;
assign w62435 = ~w62392 & w62434;
assign w62436 = w62361 & ~w62415;
assign w62437 = ~w62380 & w62396;
assign w62438 = w62435 & ~w62437;
assign w62439 = ~w62436 & w62438;
assign w62440 = ~w62432 & ~w62439;
assign w62441 = ~w62412 & ~w62440;
assign w62442 = ~pi8771 & w62441;
assign w62443 = pi8771 & ~w62441;
assign w62444 = ~w62442 & ~w62443;
assign w62445 = w62195 & w62201;
assign w62446 = ~w62246 & ~w62262;
assign w62447 = ~w62445 & ~w62446;
assign w62448 = ~w62189 & w62195;
assign w62449 = w62208 & ~w62245;
assign w62450 = ~w62448 & w62449;
assign w62451 = ~w62201 & w62214;
assign w62452 = ~w62207 & ~w62248;
assign w62453 = ~w62451 & ~w62452;
assign w62454 = ~w62231 & ~w62249;
assign w62455 = w62453 & w62454;
assign w62456 = ~w62447 & ~w62450;
assign w62457 = (~w62244 & ~w62456) | (~w62244 & w64337) | (~w62456 & w64337);
assign w62458 = w62201 & w62231;
assign w62459 = w62231 & w64338;
assign w62460 = ~w62247 & ~w62459;
assign w62461 = ~w62195 & ~w62460;
assign w62462 = ~w62229 & ~w62236;
assign w62463 = w62233 & ~w62462;
assign w62464 = (~w62195 & ~w62221) | (~w62195 & w62235) | (~w62221 & w62235);
assign w62465 = w62224 & w62464;
assign w62466 = ~w62223 & ~w62459;
assign w62467 = ~w62463 & ~w62465;
assign w62468 = w62466 & w62467;
assign w62469 = w62244 & ~w62468;
assign w62470 = ~w62227 & ~w62228;
assign w62471 = ~w62461 & w62470;
assign w62472 = ~w62457 & w62471;
assign w62473 = ~w62469 & w62472;
assign w62474 = pi8722 & ~w62473;
assign w62475 = ~pi8722 & w62473;
assign w62476 = ~w62474 & ~w62475;
assign w62477 = w62189 & ~w62195;
assign w62478 = ~w62453 & w62477;
assign w62479 = ~w62220 & w62478;
assign w62480 = w62201 & w62220;
assign w62481 = ~w62246 & ~w62480;
assign w62482 = ~w62235 & ~w62481;
assign w62483 = w62214 & ~w62464;
assign w62484 = ~w62245 & w62260;
assign w62485 = ~w62483 & w62484;
assign w62486 = ~w62482 & ~w62485;
assign w62487 = w62244 & ~w62486;
assign w62488 = w62225 & ~w62244;
assign w62489 = w62453 & w62488;
assign w62490 = w62214 & ~w62216;
assign w62491 = w62235 & ~w62490;
assign w62492 = ~w62258 & w62491;
assign w62493 = ~w62232 & w62244;
assign w62494 = ~w62236 & ~w62451;
assign w62495 = ~w62462 & ~w62493;
assign w62496 = ~w62494 & w62495;
assign w62497 = ~w62479 & ~w62489;
assign w62498 = ~w62492 & ~w62496;
assign w62499 = w62497 & w62498;
assign w62500 = ~w62487 & w62499;
assign w62501 = pi8701 & ~w62500;
assign w62502 = ~pi8701 & w62500;
assign w62503 = ~w62501 & ~w62502;
assign w62504 = ~w61681 & w61710;
assign w62505 = w61690 & w61724;
assign w62506 = ~w61752 & ~w62505;
assign w62507 = w62504 & w62506;
assign w62508 = w61681 & w61727;
assign w62509 = (w62508 & w61715) | (w62508 & w64339) | (w61715 & w64339);
assign w62510 = w61681 & ~w61721;
assign w62511 = ~w61721 & ~w61731;
assign w62512 = ~w61730 & ~w61768;
assign w62513 = w62511 & w62512;
assign w62514 = ~w62510 & ~w62513;
assign w62515 = ~w61729 & ~w62514;
assign w62516 = w61681 & w61709;
assign w62517 = ~w61750 & ~w62516;
assign w62518 = w61675 & ~w62517;
assign w62519 = ~w61669 & w61690;
assign w62520 = ~w61692 & ~w62504;
assign w62521 = ~w62519 & ~w62520;
assign w62522 = w61770 & ~w62518;
assign w62523 = ~w62521 & w62522;
assign w62524 = ~w62515 & ~w62523;
assign w62525 = ~w62506 & w62510;
assign w62526 = ~w62507 & ~w62525;
assign w62527 = ~w62509 & w62526;
assign w62528 = ~w62524 & w62527;
assign w62529 = pi8790 & ~w62528;
assign w62530 = ~pi8790 & w62528;
assign w62531 = ~w62529 & ~w62530;
assign w62532 = w61903 & ~w61915;
assign w62533 = (~w61897 & w61948) | (~w61897 & w63342) | (w61948 & w63342);
assign w62534 = ~w61945 & ~w62533;
assign w62535 = w61882 & w61894;
assign w62536 = w61881 & w61900;
assign w62537 = ~w61946 & ~w62536;
assign w62538 = ~w62535 & w62537;
assign w62539 = ~w61894 & ~w61904;
assign w62540 = w61875 & w61915;
assign w62541 = ~w62539 & w62540;
assign w62542 = w62538 & w62541;
assign w62543 = ~w61915 & ~w62538;
assign w62544 = w62534 & ~w62542;
assign w62545 = (w61930 & ~w62544) | (w61930 & w64340) | (~w62544 & w64340);
assign w62546 = w61921 & w61933;
assign w62547 = w61930 & ~w62546;
assign w62548 = w61882 & w61920;
assign w62549 = w61902 & ~w61951;
assign w62550 = ~w61907 & ~w61917;
assign w62551 = w61897 & ~w62550;
assign w62552 = ~w62548 & ~w62551;
assign w62553 = ~w62549 & w62552;
assign w62554 = ~w62547 & ~w62553;
assign w62555 = ~w61919 & ~w62532;
assign w62556 = ~w62554 & w62555;
assign w62557 = ~w62545 & w62556;
assign w62558 = pi8755 & w62557;
assign w62559 = ~pi8755 & ~w62557;
assign w62560 = ~w62558 & ~w62559;
assign w62561 = ~pi8031 & pi9040;
assign w62562 = ~pi7949 & ~pi9040;
assign w62563 = ~w62561 & ~w62562;
assign w62564 = pi8750 & ~w62563;
assign w62565 = ~pi8750 & w62563;
assign w62566 = ~w62564 & ~w62565;
assign w62567 = ~pi8025 & pi9040;
assign w62568 = ~pi7939 & ~pi9040;
assign w62569 = ~w62567 & ~w62568;
assign w62570 = pi8773 & ~w62569;
assign w62571 = ~pi8773 & w62569;
assign w62572 = ~w62570 & ~w62571;
assign w62573 = ~w62566 & w62572;
assign w62574 = ~pi7986 & pi9040;
assign w62575 = ~pi7931 & ~pi9040;
assign w62576 = ~w62574 & ~w62575;
assign w62577 = pi8795 & ~w62576;
assign w62578 = ~pi8795 & w62576;
assign w62579 = ~w62577 & ~w62578;
assign w62580 = ~pi8034 & pi9040;
assign w62581 = ~pi7963 & ~pi9040;
assign w62582 = ~w62580 & ~w62581;
assign w62583 = pi8782 & ~w62582;
assign w62584 = ~pi8782 & w62582;
assign w62585 = ~w62583 & ~w62584;
assign w62586 = w62579 & w62585;
assign w62587 = w62573 & w62586;
assign w62588 = ~pi8020 & pi9040;
assign w62589 = ~pi7929 & ~pi9040;
assign w62590 = ~w62588 & ~w62589;
assign w62591 = pi8713 & ~w62590;
assign w62592 = ~pi8713 & w62590;
assign w62593 = ~w62591 & ~w62592;
assign w62594 = w62572 & w62593;
assign w62595 = ~w62585 & ~w62593;
assign w62596 = w62566 & w62593;
assign w62597 = ~w62572 & ~w62596;
assign w62598 = ~w62594 & ~w62595;
assign w62599 = ~w62597 & w62598;
assign w62600 = ~w62566 & ~w62585;
assign w62601 = ~w62572 & ~w62593;
assign w62602 = w62600 & w62601;
assign w62603 = ~w62599 & w64341;
assign w62604 = ~pi7977 & pi9040;
assign w62605 = ~pi7959 & ~pi9040;
assign w62606 = ~w62604 & ~w62605;
assign w62607 = pi8775 & ~w62606;
assign w62608 = ~pi8775 & w62606;
assign w62609 = ~w62607 & ~w62608;
assign w62610 = ~w62602 & ~w62609;
assign w62611 = w62579 & ~w62610;
assign w62612 = ~w62603 & w62611;
assign w62613 = w62566 & w62585;
assign w62614 = ~w62594 & w62613;
assign w62615 = ~w62594 & ~w62601;
assign w62616 = w62600 & ~w62615;
assign w62617 = ~w62599 & ~w62616;
assign w62618 = w62617 & w64342;
assign w62619 = w62614 & w62618;
assign w62620 = ~w62600 & ~w62613;
assign w62621 = w62579 & ~w62593;
assign w62622 = w62615 & ~w62621;
assign w62623 = ~w62599 & ~w62622;
assign w62624 = w62620 & ~w62623;
assign w62625 = ~w62620 & ~w62622;
assign w62626 = ~w62609 & ~w62625;
assign w62627 = ~w62624 & w62626;
assign w62628 = ~w62579 & w62609;
assign w62629 = ~w62601 & w62628;
assign w62630 = ~w62599 & w64343;
assign w62631 = ~w62587 & ~w62630;
assign w62632 = ~w62612 & w62631;
assign w62633 = ~w62627 & w62632;
assign w62634 = ~w62619 & w62633;
assign w62635 = pi8721 & ~w62634;
assign w62636 = ~pi8721 & w62634;
assign w62637 = ~w62635 & ~w62636;
assign w62638 = w61662 & w61694;
assign w62639 = ~w61768 & ~w62519;
assign w62640 = w61681 & ~w62639;
assign w62641 = ~w61681 & ~w61690;
assign w62642 = w61725 & w62641;
assign w62643 = ~w61721 & ~w62638;
assign w62644 = ~w62642 & w62643;
assign w62645 = ~w62640 & w62644;
assign w62646 = ~w61684 & ~w62516;
assign w62647 = w61662 & ~w62646;
assign w62648 = w61721 & ~w61755;
assign w62649 = ~w61700 & w62648;
assign w62650 = ~w61708 & w62649;
assign w62651 = ~w62647 & w62650;
assign w62652 = ~w62645 & ~w62651;
assign w62653 = ~w61662 & w61691;
assign w62654 = ~w62511 & w62653;
assign w62655 = ~w61758 & ~w62654;
assign w62656 = ~w62652 & w62655;
assign w62657 = pi8714 & ~w62656;
assign w62658 = ~pi8714 & w62656;
assign w62659 = ~w62657 & ~w62658;
assign w62660 = ~w62361 & ~w62367;
assign w62661 = w62373 & ~w62380;
assign w62662 = ~w62660 & ~w62661;
assign w62663 = w62387 & ~w62662;
assign w62664 = ~w62361 & w62373;
assign w62665 = w62367 & ~w62664;
assign w62666 = w62381 & ~w62665;
assign w62667 = w62663 & w62666;
assign w62668 = ~w62400 & w62664;
assign w62669 = ~w62399 & w62668;
assign w62670 = ~w62433 & ~w62668;
assign w62671 = ~w62669 & ~w62670;
assign w62672 = ~w62662 & w64344;
assign w62673 = ~w62408 & ~w62672;
assign w62674 = ~w62388 & ~w62401;
assign w62675 = w62373 & ~w62660;
assign w62676 = ~w62674 & ~w62675;
assign w62677 = ~w62671 & ~w62676;
assign w62678 = w62673 & w62677;
assign w62679 = ~w62387 & w62426;
assign w62680 = w62426 & w64345;
assign w62681 = w62390 & w62660;
assign w62682 = w62389 & w62397;
assign w62683 = w62417 & ~w62661;
assign w62684 = w62408 & ~w62681;
assign w62685 = ~w62682 & ~w62683;
assign w62686 = w62684 & w62685;
assign w62687 = ~w62680 & w62686;
assign w62688 = ~w62669 & w62687;
assign w62689 = ~w62678 & ~w62688;
assign w62690 = w62361 & ~w62381;
assign w62691 = ~w62391 & w62690;
assign w62692 = ~w62667 & ~w62691;
assign w62693 = ~w62689 & w62692;
assign w62694 = pi8765 & ~w62693;
assign w62695 = ~pi8765 & w62693;
assign w62696 = ~w62694 & ~w62695;
assign w62697 = (w62445 & ~w62467) | (w62445 & w64346) | (~w62467 & w64346);
assign w62698 = ~w62259 & w62458;
assign w62699 = ~w62215 & w62448;
assign w62700 = w62244 & ~w62699;
assign w62701 = ~w62478 & w62700;
assign w62702 = ~w62698 & w62701;
assign w62703 = w62218 & ~w62458;
assign w62704 = ~w62248 & w62249;
assign w62705 = ~w62259 & w62704;
assign w62706 = ~w62227 & ~w62244;
assign w62707 = ~w62261 & ~w62705;
assign w62708 = w62706 & w62707;
assign w62709 = ~w62703 & w62708;
assign w62710 = ~w62702 & ~w62709;
assign w62711 = ~w62264 & ~w62697;
assign w62712 = ~w62710 & w62711;
assign w62713 = pi8779 & ~w62712;
assign w62714 = ~pi8779 & w62712;
assign w62715 = ~w62713 & ~w62714;
assign w62716 = w62102 & w62159;
assign w62717 = w62113 & ~w62716;
assign w62718 = ~w62176 & ~w62717;
assign w62719 = (~w62067 & w62081) | (~w62067 & w62127) | (w62081 & w62127);
assign w62720 = ~w62112 & w62719;
assign w62721 = (w62094 & w62720) | (w62094 & w64347) | (w62720 & w64347);
assign w62722 = ~w62094 & ~w62107;
assign w62723 = ~w62087 & w62121;
assign w62724 = ~w62721 & w62723;
assign w62725 = ~w62722 & w62724;
assign w62726 = w62080 & ~w62160;
assign w62727 = ~w62127 & w62151;
assign w62728 = ~w62726 & ~w62727;
assign w62729 = ~w62102 & ~w62728;
assign w62730 = ~w62101 & w62110;
assign w62731 = ~w62135 & w62158;
assign w62732 = ~w62730 & w62731;
assign w62733 = ~w62729 & w62732;
assign w62734 = (~w62718 & w62725) | (~w62718 & w64348) | (w62725 & w64348);
assign w62735 = ~pi8787 & w62734;
assign w62736 = pi8787 & ~w62734;
assign w62737 = ~w62735 & ~w62736;
assign w62738 = ~w61834 & w61836;
assign w62739 = w61790 & w61841;
assign w62740 = ~w61802 & ~w61828;
assign w62741 = (~w61789 & w61859) | (~w61789 & w64349) | (w61859 & w64349);
assign w62742 = ~w61841 & w61852;
assign w62743 = ~w61820 & ~w62739;
assign w62744 = ~w62742 & w62743;
assign w62745 = ~w62741 & w62744;
assign w62746 = w61783 & ~w61796;
assign w62747 = w61811 & w62746;
assign w62748 = ~w61838 & ~w61849;
assign w62749 = w61789 & ~w62748;
assign w62750 = w61802 & w61843;
assign w62751 = w61820 & ~w62750;
assign w62752 = ~w61789 & ~w62746;
assign w62753 = ~w61838 & w62752;
assign w62754 = ~w62747 & w62751;
assign w62755 = ~w62753 & w62754;
assign w62756 = ~w62749 & w62755;
assign w62757 = ~w62745 & ~w62756;
assign w62758 = ~w62738 & ~w62757;
assign w62759 = ~pi8751 & w62758;
assign w62760 = pi8751 & ~w62758;
assign w62761 = ~w62759 & ~w62760;
assign w62762 = w62585 & w62593;
assign w62763 = ~w62579 & w62762;
assign w62764 = ~w62566 & w62763;
assign w62765 = ~w62566 & ~w62593;
assign w62766 = ~w62596 & ~w62765;
assign w62767 = w62572 & ~w62766;
assign w62768 = w62579 & ~w62597;
assign w62769 = ~w62767 & w62768;
assign w62770 = ~w62572 & w62595;
assign w62771 = ~w62767 & ~w62770;
assign w62772 = ~w62579 & ~w62771;
assign w62773 = w62610 & ~w62769;
assign w62774 = ~w62772 & w62773;
assign w62775 = w62566 & ~w62572;
assign w62776 = w62621 & w62775;
assign w62777 = (~w62585 & w62767) | (~w62585 & w64350) | (w62767 & w64350);
assign w62778 = ~w62572 & ~w62579;
assign w62779 = w62615 & w62766;
assign w62780 = ~w62778 & ~w62779;
assign w62781 = ~w62595 & ~w62762;
assign w62782 = ~w62780 & w62781;
assign w62783 = w62609 & ~w62777;
assign w62784 = ~w62782 & w62783;
assign w62785 = ~w62774 & ~w62784;
assign w62786 = ~w62572 & w62586;
assign w62787 = ~w62766 & w62786;
assign w62788 = ~w62764 & ~w62787;
assign w62789 = ~w62785 & w62788;
assign w62790 = pi8753 & ~w62789;
assign w62791 = ~pi8753 & w62789;
assign w62792 = ~w62790 & ~w62791;
assign w62793 = w61932 & w61941;
assign w62794 = w61900 & w61921;
assign w62795 = ~w61948 & ~w62794;
assign w62796 = ~w61936 & ~w62533;
assign w62797 = (~w62536 & w62796) | (~w62536 & w63505) | (w62796 & w63505);
assign w62798 = w61915 & ~w62797;
assign w62799 = w61921 & w62795;
assign w62800 = ~w61918 & ~w62799;
assign w62801 = (w61930 & w62798) | (w61930 & w64351) | (w62798 & w64351);
assign w62802 = w61881 & w61930;
assign w62803 = ~w61915 & ~w62802;
assign w62804 = w61946 & ~w62803;
assign w62805 = ~w61948 & ~w62535;
assign w62806 = w61915 & ~w62805;
assign w62807 = ~w61881 & ~w61949;
assign w62808 = w61888 & w61920;
assign w62809 = ~w61940 & ~w62808;
assign w62810 = w61881 & ~w62809;
assign w62811 = ~w61901 & ~w62548;
assign w62812 = ~w62806 & w62811;
assign w62813 = ~w62807 & ~w62810;
assign w62814 = w62812 & w62813;
assign w62815 = ~w62793 & ~w62804;
assign w62816 = (w62815 & w62814) | (w62815 & w64352) | (w62814 & w64352);
assign w62817 = ~w62801 & w62816;
assign w62818 = ~pi8725 & w62817;
assign w62819 = pi8725 & ~w62817;
assign w62820 = ~w62818 & ~w62819;
assign w62821 = w61923 & ~w62534;
assign w62822 = w61899 & ~w62537;
assign w62823 = w62795 & ~w62822;
assign w62824 = ~w61915 & ~w62823;
assign w62825 = ~w61895 & ~w61934;
assign w62826 = ~w61947 & ~w62825;
assign w62827 = w61905 & ~w61923;
assign w62828 = w61930 & ~w62794;
assign w62829 = ~w62827 & w62828;
assign w62830 = ~w62826 & w62829;
assign w62831 = ~w61939 & w61947;
assign w62832 = w61931 & ~w62541;
assign w62833 = ~w62831 & w62832;
assign w62834 = ~w62830 & ~w62833;
assign w62835 = ~w62821 & ~w62824;
assign w62836 = ~w62834 & w62835;
assign w62837 = pi8768 & w62836;
assign w62838 = ~pi8768 & ~w62836;
assign w62839 = ~w62837 & ~w62838;
assign w62840 = w61796 & ~w61854;
assign w62841 = ~w62740 & w62840;
assign w62842 = ~w62747 & ~w62841;
assign w62843 = w61820 & ~w62842;
assign w62844 = ~w61827 & w61841;
assign w62845 = ~w61796 & w61820;
assign w62846 = w62844 & w62845;
assign w62847 = ~w61820 & ~w61841;
assign w62848 = ~w62747 & w62847;
assign w62849 = ~w62846 & ~w62848;
assign w62850 = w61789 & ~w62849;
assign w62851 = ~w61789 & w62844;
assign w62852 = w61802 & ~w62746;
assign w62853 = ~w61803 & ~w61828;
assign w62854 = ~w62852 & w62853;
assign w62855 = ~w62851 & ~w62854;
assign w62856 = w61802 & w61824;
assign w62857 = w62751 & ~w62856;
assign w62858 = ~w62855 & ~w62857;
assign w62859 = ~w62850 & ~w62858;
assign w62860 = ~w62843 & w62859;
assign w62861 = pi8797 & w62860;
assign w62862 = ~pi8797 & ~w62860;
assign w62863 = ~w62861 & ~w62862;
assign w62864 = ~w62663 & ~w62679;
assign w62865 = w62361 & ~w62864;
assign w62866 = ~w62396 & ~w62398;
assign w62867 = ~w62361 & ~w62866;
assign w62868 = ~w62392 & ~w62682;
assign w62869 = ~w62421 & ~w62672;
assign w62870 = ~w62867 & w62868;
assign w62871 = w62869 & w62870;
assign w62872 = (w62408 & ~w62871) | (w62408 & w64353) | (~w62871 & w64353);
assign w62873 = w62367 & w62390;
assign w62874 = ~w62425 & ~w62873;
assign w62875 = (~w62408 & ~w62874) | (~w62408 & w64354) | (~w62874 & w64354);
assign w62876 = w62868 & ~w62875;
assign w62877 = ~w62361 & ~w62876;
assign w62878 = ~w62361 & ~w62414;
assign w62879 = w62673 & ~w62878;
assign w62880 = w62876 & w62879;
assign w62881 = ~w62877 & ~w62880;
assign w62882 = ~w62872 & w62881;
assign w62883 = ~pi8729 & w62882;
assign w62884 = pi8729 & ~w62882;
assign w62885 = ~w62883 & ~w62884;
assign w62886 = w61802 & ~w61822;
assign w62887 = w61820 & ~w62886;
assign w62888 = w61803 & ~w61810;
assign w62889 = (~w61811 & ~w61828) | (~w61811 & w64355) | (~w61828 & w64355);
assign w62890 = ~w61844 & ~w62888;
assign w62891 = (w62890 & ~w62749) | (w62890 & w64356) | (~w62749 & w64356);
assign w62892 = ~w62887 & ~w62891;
assign w62893 = ~w62750 & ~w62856;
assign w62894 = ~w61820 & ~w62893;
assign w62895 = w61814 & ~w61842;
assign w62896 = ~w61838 & ~w62895;
assign w62897 = ~w61856 & ~w62746;
assign w62898 = ~w61842 & ~w61849;
assign w62899 = ~w61848 & w62898;
assign w62900 = ~w62897 & w62899;
assign w62901 = w61820 & ~w62900;
assign w62902 = ~w62894 & ~w62896;
assign w62903 = ~w62892 & w62902;
assign w62904 = ~w62901 & w62903;
assign w62905 = pi8767 & ~w62904;
assign w62906 = ~pi8767 & w62904;
assign w62907 = ~w62905 & ~w62906;
assign w62908 = w62007 & ~w62031;
assign w62909 = ~w62036 & ~w62043;
assign w62910 = ~w62315 & w62909;
assign w62911 = w61968 & ~w62910;
assign w62912 = (~w62295 & w62327) | (~w62295 & w64357) | (w62327 & w64357);
assign w62913 = w61968 & w62001;
assign w62914 = w62042 & w62913;
assign w62915 = ~w62912 & ~w62914;
assign w62916 = ~w61994 & ~w62915;
assign w62917 = ~w62030 & w62290;
assign w62918 = ~w62303 & ~w62917;
assign w62919 = w62034 & w62918;
assign w62920 = ~w61968 & ~w62919;
assign w62921 = ~w62908 & ~w62911;
assign w62922 = ~w62916 & w62921;
assign w62923 = ~w62920 & w62922;
assign w62924 = pi8720 & ~w62923;
assign w62925 = ~pi8720 & w62923;
assign w62926 = ~w62924 & ~w62925;
assign w62927 = (w62586 & ~w62617) | (w62586 & w63343) | (~w62617 & w63343);
assign w62928 = (~w62600 & w62615) | (~w62600 & w64358) | (w62615 & w64358);
assign w62929 = (w62617 & w67187) | (w62617 & w67188) | (w67187 & w67188);
assign w62930 = ~w62927 & w63506;
assign w62931 = w62579 & ~w62617;
assign w62932 = w62617 & ~w62621;
assign w62933 = ~w62931 & ~w62932;
assign w62934 = ~w62930 & ~w62933;
assign w62935 = ~w62609 & ~w62934;
assign w62936 = w62763 & w62767;
assign w62937 = w62579 & ~w62585;
assign w62938 = w62779 & w62937;
assign w62939 = w62609 & ~w62933;
assign w62940 = ~w62936 & ~w62938;
assign w62941 = (w62940 & ~w62939) | (w62940 & w63507) | (~w62939 & w63507);
assign w62942 = ~w62935 & w62941;
assign w62943 = pi8747 & ~w62942;
assign w62944 = ~pi8747 & w62942;
assign w62945 = ~w62943 & ~w62944;
assign w62946 = ~w62423 & ~w62878;
assign w62947 = ~w62361 & w62380;
assign w62948 = ~w62388 & w62947;
assign w62949 = ~w62419 & w62948;
assign w62950 = w62361 & ~w62674;
assign w62951 = w62408 & ~w62437;
assign w62952 = ~w62949 & w62951;
assign w62953 = ~w62950 & w62952;
assign w62954 = ~w62418 & ~w62679;
assign w62955 = ~w62666 & w62954;
assign w62956 = w62435 & w62955;
assign w62957 = ~w62953 & ~w62956;
assign w62958 = ~w62946 & ~w62957;
assign w62959 = ~pi8693 & w62958;
assign w62960 = pi8693 & ~w62958;
assign w62961 = ~w62959 & ~w62960;
assign w62962 = ~w62762 & ~w62775;
assign w62963 = ~w62579 & ~w62765;
assign w62964 = w62962 & w62963;
assign w62965 = (~w62964 & w62617) | (~w62964 & w64359) | (w62617 & w64359);
assign w62966 = ~w62609 & ~w62965;
assign w62967 = ~w62593 & w62775;
assign w62968 = ~w62762 & ~w62967;
assign w62969 = w62628 & ~w62968;
assign w62970 = ~w62609 & ~w62778;
assign w62971 = w62614 & ~w62970;
assign w62972 = ~w62614 & ~w62962;
assign w62973 = ~w62573 & w62609;
assign w62974 = w62972 & w62973;
assign w62975 = ~w62618 & ~w62972;
assign w62976 = w62579 & ~w62974;
assign w62977 = ~w62975 & w62976;
assign w62978 = ~w62969 & ~w62971;
assign w62979 = ~w62966 & w62978;
assign w62980 = ~w62977 & w62979;
assign w62981 = ~pi8784 & w62980;
assign w62982 = pi8784 & ~w62980;
assign w62983 = ~w62981 & ~w62982;
assign w62984 = pi8895 & pi9040;
assign w62985 = pi9007 & ~pi9040;
assign w62986 = ~w62984 & ~w62985;
assign w62987 = pi9037 & pi9040;
assign w62988 = pi8925 & ~pi9040;
assign w62989 = ~w62987 & ~w62988;
assign w62990 = pi8881 & pi9040;
assign w62991 = pi8993 & ~pi9040;
assign w62992 = ~w62990 & ~w62991;
assign w62993 = pi9018 & pi9040;
assign w62994 = pi8906 & ~pi9040;
assign w62995 = ~w62993 & ~w62994;
assign w62996 = pi8912 & pi9040;
assign w62997 = pi9024 & ~pi9040;
assign w62998 = ~w62996 & ~w62997;
assign w62999 = pi8880 & pi9040;
assign w63000 = pi8992 & ~pi9040;
assign w63001 = ~w62999 & ~w63000;
assign w63002 = pi8897 & pi9040;
assign w63003 = pi9009 & ~pi9040;
assign w63004 = ~w63002 & ~w63003;
assign w63005 = pi8987 & pi9040;
assign w63006 = pi8875 & ~pi9040;
assign w63007 = ~w63005 & ~w63006;
assign w63008 = pi8917 & pi9040;
assign w63009 = pi9029 & ~pi9040;
assign w63010 = ~w63008 & ~w63009;
assign w63011 = pi9026 & pi9040;
assign w63012 = pi8914 & ~pi9040;
assign w63013 = ~w63011 & ~w63012;
assign w63014 = pi8882 & pi9040;
assign w63015 = pi8994 & ~pi9040;
assign w63016 = ~w63014 & ~w63015;
assign w63017 = pi8989 & pi9040;
assign w63018 = pi8877 & ~pi9040;
assign w63019 = ~w63017 & ~w63018;
assign w63020 = pi9028 & pi9040;
assign w63021 = pi8916 & ~pi9040;
assign w63022 = ~w63020 & ~w63021;
assign w63023 = pi8898 & pi9040;
assign w63024 = pi9010 & ~pi9040;
assign w63025 = ~w63023 & ~w63024;
assign w63026 = pi9014 & pi9040;
assign w63027 = pi8902 & ~pi9040;
assign w63028 = ~w63026 & ~w63027;
assign w63029 = pi9036 & pi9040;
assign w63030 = pi8924 & ~pi9040;
assign w63031 = ~w63029 & ~w63030;
assign w63032 = pi8927 & pi9040;
assign w63033 = pi9039 & ~pi9040;
assign w63034 = ~w63032 & ~w63033;
assign w63035 = pi8876 & pi9040;
assign w63036 = pi8988 & ~pi9040;
assign w63037 = ~w63035 & ~w63036;
assign w63038 = pi9021 & pi9040;
assign w63039 = pi8909 & ~pi9040;
assign w63040 = ~w63038 & ~w63039;
assign w63041 = pi8892 & pi9040;
assign w63042 = pi9004 & ~pi9040;
assign w63043 = ~w63041 & ~w63042;
assign w63044 = pi8890 & pi9040;
assign w63045 = pi9002 & ~pi9040;
assign w63046 = ~w63044 & ~w63045;
assign w63047 = pi9009 & pi9040;
assign w63048 = pi8897 & ~pi9040;
assign w63049 = ~w63047 & ~w63048;
assign w63050 = pi8906 & pi9040;
assign w63051 = pi9018 & ~pi9040;
assign w63052 = ~w63050 & ~w63051;
assign w63053 = pi8905 & pi9040;
assign w63054 = pi9017 & ~pi9040;
assign w63055 = ~w63053 & ~w63054;
assign w63056 = pi9024 & pi9040;
assign w63057 = pi8912 & ~pi9040;
assign w63058 = ~w63056 & ~w63057;
assign w63059 = pi8925 & pi9040;
assign w63060 = pi9037 & ~pi9040;
assign w63061 = ~w63059 & ~w63060;
assign w63062 = pi8993 & pi9040;
assign w63063 = pi8881 & ~pi9040;
assign w63064 = ~w63062 & ~w63063;
assign w63065 = pi8920 & pi9040;
assign w63066 = pi9032 & ~pi9040;
assign w63067 = ~w63065 & ~w63066;
assign w63068 = pi8923 & pi9040;
assign w63069 = pi9035 & ~pi9040;
assign w63070 = ~w63068 & ~w63069;
assign w63071 = pi9029 & pi9040;
assign w63072 = pi8917 & ~pi9040;
assign w63073 = ~w63071 & ~w63072;
assign w63074 = pi9019 & pi9040;
assign w63075 = pi8907 & ~pi9040;
assign w63076 = ~w63074 & ~w63075;
assign w63077 = pi9001 & pi9040;
assign w63078 = pi8889 & ~pi9040;
assign w63079 = ~w63077 & ~w63078;
assign w63080 = pi8873 & pi9040;
assign w63081 = pi8985 & ~pi9040;
assign w63082 = ~w63080 & ~w63081;
assign w63083 = pi8992 & pi9040;
assign w63084 = pi8880 & ~pi9040;
assign w63085 = ~w63083 & ~w63084;
assign w63086 = pi8914 & pi9040;
assign w63087 = pi9026 & ~pi9040;
assign w63088 = ~w63086 & ~w63087;
assign w63089 = pi9017 & pi9040;
assign w63090 = pi8905 & ~pi9040;
assign w63091 = ~w63089 & ~w63090;
assign w63092 = pi8879 & pi9040;
assign w63093 = pi8991 & ~pi9040;
assign w63094 = ~w63092 & ~w63093;
assign w63095 = pi9027 & pi9040;
assign w63096 = pi8915 & ~pi9040;
assign w63097 = ~w63095 & ~w63096;
assign w63098 = pi9015 & pi9040;
assign w63099 = pi8903 & ~pi9040;
assign w63100 = ~w63098 & ~w63099;
assign w63101 = pi8904 & pi9040;
assign w63102 = pi9016 & ~pi9040;
assign w63103 = ~w63101 & ~w63102;
assign w63104 = pi9000 & pi9040;
assign w63105 = pi8888 & ~pi9040;
assign w63106 = ~w63104 & ~w63105;
assign w63107 = pi8916 & pi9040;
assign w63108 = pi9028 & ~pi9040;
assign w63109 = ~w63107 & ~w63108;
assign w63110 = pi8887 & pi9040;
assign w63111 = pi8999 & ~pi9040;
assign w63112 = ~w63110 & ~w63111;
assign w63113 = pi9032 & pi9040;
assign w63114 = pi8920 & ~pi9040;
assign w63115 = ~w63113 & ~w63114;
assign w63116 = pi8988 & pi9040;
assign w63117 = pi8876 & ~pi9040;
assign w63118 = ~w63116 & ~w63117;
assign w63119 = pi8903 & pi9040;
assign w63120 = pi9015 & ~pi9040;
assign w63121 = ~w63119 & ~w63120;
assign w63122 = pi8995 & pi9040;
assign w63123 = pi8883 & ~pi9040;
assign w63124 = ~w63122 & ~w63123;
assign w63125 = pi9003 & pi9040;
assign w63126 = pi8891 & ~pi9040;
assign w63127 = ~w63125 & ~w63126;
assign w63128 = pi8907 & pi9040;
assign w63129 = pi9019 & ~pi9040;
assign w63130 = ~w63128 & ~w63129;
assign w63131 = pi8994 & pi9040;
assign w63132 = pi8882 & ~pi9040;
assign w63133 = ~w63131 & ~w63132;
assign w63134 = pi9007 & pi9040;
assign w63135 = pi8895 & ~pi9040;
assign w63136 = ~w63134 & ~w63135;
assign w63137 = pi9006 & pi9040;
assign w63138 = pi8894 & ~pi9040;
assign w63139 = ~w63137 & ~w63138;
assign w63140 = pi8926 & pi9040;
assign w63141 = pi9038 & ~pi9040;
assign w63142 = ~w63140 & ~w63141;
assign w63143 = pi8909 & pi9040;
assign w63144 = pi9021 & ~pi9040;
assign w63145 = ~w63143 & ~w63144;
assign w63146 = pi8875 & pi9040;
assign w63147 = pi8987 & ~pi9040;
assign w63148 = ~w63146 & ~w63147;
assign w63149 = pi8891 & pi9040;
assign w63150 = pi9003 & ~pi9040;
assign w63151 = ~w63149 & ~w63150;
assign w63152 = pi8884 & pi9040;
assign w63153 = pi8996 & ~pi9040;
assign w63154 = ~w63152 & ~w63153;
assign w63155 = pi8885 & pi9040;
assign w63156 = pi8997 & ~pi9040;
assign w63157 = ~w63155 & ~w63156;
assign w63158 = pi9011 & pi9040;
assign w63159 = pi8899 & ~pi9040;
assign w63160 = ~w63158 & ~w63159;
assign w63161 = pi8883 & pi9040;
assign w63162 = pi8995 & ~pi9040;
assign w63163 = ~w63161 & ~w63162;
assign w63164 = pi8901 & pi9040;
assign w63165 = pi9013 & ~pi9040;
assign w63166 = ~w63164 & ~w63165;
assign w63167 = pi8902 & pi9040;
assign w63168 = pi9014 & ~pi9040;
assign w63169 = ~w63167 & ~w63168;
assign w63170 = pi8913 & pi9040;
assign w63171 = pi9025 & ~pi9040;
assign w63172 = ~w63170 & ~w63171;
assign w63173 = pi9012 & pi9040;
assign w63174 = pi8900 & ~pi9040;
assign w63175 = ~w63173 & ~w63174;
assign w63176 = pi8893 & pi9040;
assign w63177 = pi9005 & ~pi9040;
assign w63178 = ~w63176 & ~w63177;
assign w63179 = pi8899 & pi9040;
assign w63180 = pi9011 & ~pi9040;
assign w63181 = ~w63179 & ~w63180;
assign w63182 = pi8900 & pi9040;
assign w63183 = pi9012 & ~pi9040;
assign w63184 = ~w63182 & ~w63183;
assign w63185 = pi8910 & pi9040;
assign w63186 = pi9022 & ~pi9040;
assign w63187 = ~w63185 & ~w63186;
assign w63188 = pi8894 & pi9040;
assign w63189 = pi9006 & ~pi9040;
assign w63190 = ~w63188 & ~w63189;
assign w63191 = pi9035 & pi9040;
assign w63192 = pi8923 & ~pi9040;
assign w63193 = ~w63191 & ~w63192;
assign w63194 = pi8997 & pi9040;
assign w63195 = pi8885 & ~pi9040;
assign w63196 = ~w63194 & ~w63195;
assign w63197 = pi9013 & pi9040;
assign w63198 = pi8901 & ~pi9040;
assign w63199 = ~w63197 & ~w63198;
assign w63200 = pi9025 & pi9040;
assign w63201 = pi8913 & ~pi9040;
assign w63202 = ~w63200 & ~w63201;
assign w63203 = pi9020 & pi9040;
assign w63204 = pi8908 & ~pi9040;
assign w63205 = ~w63203 & ~w63204;
assign w63206 = pi8878 & pi9040;
assign w63207 = pi8990 & ~pi9040;
assign w63208 = ~w63206 & ~w63207;
assign w63209 = pi9005 & pi9040;
assign w63210 = pi8893 & ~pi9040;
assign w63211 = ~w63209 & ~w63210;
assign w63212 = pi8998 & pi9040;
assign w63213 = pi8886 & ~pi9040;
assign w63214 = ~w63212 & ~w63213;
assign w63215 = pi9031 & pi9040;
assign w63216 = pi8919 & ~pi9040;
assign w63217 = ~w63215 & ~w63216;
assign w63218 = pi8908 & pi9040;
assign w63219 = pi9020 & ~pi9040;
assign w63220 = ~w63218 & ~w63219;
assign w63221 = pi9023 & pi9040;
assign w63222 = pi8911 & ~pi9040;
assign w63223 = ~w63221 & ~w63222;
assign w63224 = pi8896 & pi9040;
assign w63225 = pi9008 & ~pi9040;
assign w63226 = ~w63224 & ~w63225;
assign w63227 = pi8888 & pi9040;
assign w63228 = pi9000 & ~pi9040;
assign w63229 = ~w63227 & ~w63228;
assign w63230 = pi9038 & pi9040;
assign w63231 = pi8926 & ~pi9040;
assign w63232 = ~w63230 & ~w63231;
assign w63233 = pi9022 & pi9040;
assign w63234 = pi8910 & ~pi9040;
assign w63235 = ~w63233 & ~w63234;
assign w63236 = pi8877 & pi9040;
assign w63237 = pi8989 & ~pi9040;
assign w63238 = ~w63236 & ~w63237;
assign w63239 = pi8985 & pi9040;
assign w63240 = pi8873 & ~pi9040;
assign w63241 = ~w63239 & ~w63240;
assign w63242 = pi8886 & pi9040;
assign w63243 = pi8998 & ~pi9040;
assign w63244 = ~w63242 & ~w63243;
assign w63245 = pi9033 & pi9040;
assign w63246 = pi8921 & ~pi9040;
assign w63247 = ~w63245 & ~w63246;
assign w63248 = pi8990 & pi9040;
assign w63249 = pi8878 & ~pi9040;
assign w63250 = ~w63248 & ~w63249;
assign w63251 = pi8999 & pi9040;
assign w63252 = pi8887 & ~pi9040;
assign w63253 = ~w63251 & ~w63252;
assign w63254 = pi8918 & pi9040;
assign w63255 = pi9030 & ~pi9040;
assign w63256 = ~w63254 & ~w63255;
assign w63257 = pi8922 & pi9040;
assign w63258 = pi9034 & ~pi9040;
assign w63259 = ~w63257 & ~w63258;
assign w63260 = pi9030 & pi9040;
assign w63261 = pi8918 & ~pi9040;
assign w63262 = ~w63260 & ~w63261;
assign w63263 = pi8911 & pi9040;
assign w63264 = pi9023 & ~pi9040;
assign w63265 = ~w63263 & ~w63264;
assign w63266 = pi9004 & pi9040;
assign w63267 = pi8892 & ~pi9040;
assign w63268 = ~w63266 & ~w63267;
assign w63269 = pi9008 & pi9040;
assign w63270 = pi8896 & ~pi9040;
assign w63271 = ~w63269 & ~w63270;
assign w63272 = pi8921 & pi9040;
assign w63273 = pi9033 & ~pi9040;
assign w63274 = ~w63272 & ~w63273;
assign w63275 = pi9039 & pi9040;
assign w63276 = pi8927 & ~pi9040;
assign w63277 = ~w63275 & ~w63276;
assign w63278 = pi8874 & pi9040;
assign w63279 = pi8986 & ~pi9040;
assign w63280 = ~w63278 & ~w63279;
assign w63281 = pi8919 & pi9040;
assign w63282 = pi9031 & ~pi9040;
assign w63283 = ~w63281 & ~w63282;
assign w63284 = pi8991 & pi9040;
assign w63285 = pi8879 & ~pi9040;
assign w63286 = ~w63284 & ~w63285;
assign w63287 = pi8924 & pi9040;
assign w63288 = pi9036 & ~pi9040;
assign w63289 = ~w63287 & ~w63288;
assign w63290 = pi8996 & pi9040;
assign w63291 = pi8884 & ~pi9040;
assign w63292 = ~w63290 & ~w63291;
assign w63293 = pi9002 & pi9040;
assign w63294 = pi8890 & ~pi9040;
assign w63295 = ~w63293 & ~w63294;
assign w63296 = pi8889 & pi9040;
assign w63297 = pi9001 & ~pi9040;
assign w63298 = ~w63296 & ~w63297;
assign w63299 = pi8986 & pi9040;
assign w63300 = pi8874 & ~pi9040;
assign w63301 = ~w63299 & ~w63300;
assign w63302 = pi9010 & pi9040;
assign w63303 = pi8898 & ~pi9040;
assign w63304 = ~w63302 & ~w63303;
assign w63305 = pi8915 & pi9040;
assign w63306 = pi9027 & ~pi9040;
assign w63307 = ~w63305 & ~w63306;
assign w63308 = pi9016 & pi9040;
assign w63309 = pi8904 & ~pi9040;
assign w63310 = ~w63308 & ~w63309;
assign w63311 = pi8872 & pi9040;
assign w63312 = pi8984 & ~pi9040;
assign w63313 = ~w63311 & ~w63312;
assign w63314 = pi9034 & pi9040;
assign w63315 = pi8922 & ~pi9040;
assign w63316 = ~w63314 & ~w63315;
assign w63317 = pi8984 & pi9040;
assign w63318 = pi8872 & ~pi9040;
assign w63319 = ~w63317 & ~w63318;
assign w63320 = (w5625 & ~w5561) | (w5625 & w63344) | (~w5561 & w63344);
assign w63321 = ~w10704 & ~w10579;
assign w63322 = w13560 & w13571;
assign w63323 = w13576 & ~w13572;
assign w63324 = ~w14558 & ~w14567;
assign w63325 = w19726 & ~w19742;
assign w63326 = (~w19774 & w19777) | (~w19774 & w63345) | (w19777 & w63345);
assign w63327 = ~w23992 & w23941;
assign w63328 = ~w26591 & w26607;
assign w63329 = w30682 & w30675;
assign w63330 = w44157 & w63346;
assign w63331 = w50482 & ~w50502;
assign w63332 = w52762 & w52775;
assign w63333 = w55588 & w63347;
assign w63334 = w58034 & w58052;
assign w63335 = ~w63334 & ~w58049;
assign w63336 = w58072 & ~w58083;
assign w63337 = ~w58331 & w58358;
assign w63338 = ~w58331 & ~w58344;
assign w63339 = w59651 & w59620;
assign w63340 = w59620 & w59894;
assign w63341 = ~w60323 & w60343;
assign w63342 = w61898 & ~w61897;
assign w63343 = w62596 & w62586;
assign w63344 = ~w5567 & w5625;
assign w63345 = ~w19720 & ~w19774;
assign w63346 = w44143 & w44128;
assign w63347 = ~w55571 & w55585;
assign w63348 = ~w1392 & ~w1403;
assign w63349 = w2146 & ~w2151;
assign w63350 = w2607 & ~w2599;
assign w63351 = w2857 & ~w2844;
assign w63352 = w4599 & ~w4448;
assign w63353 = ~w63320 & ~w5652;
assign w63354 = w5691 & w5678;
assign w63355 = w6041 & w6058;
assign w63356 = w6188 & ~w6187;
assign w63357 = ~w6464 & w63508;
assign w63358 = ~w6553 & w6565;
assign w63359 = w6537 & ~w6577;
assign w63360 = w6652 & w6660;
assign w63361 = ~w6993 & w6982;
assign w63362 = w6555 & ~w7256;
assign w63363 = ~w6582 & w6551;
assign w63364 = ~w7180 & ~w7138;
assign w63365 = w8653 & w8628;
assign w63366 = ~w8269 & ~w8282;
assign w63367 = w9341 & ~w9348;
assign w63368 = ~w9407 & ~w9363;
assign w63369 = ~w10404 & ~w10411;
assign w63370 = w10575 & ~w10573;
assign w63371 = ~w10534 & w10579;
assign w63372 = ~w10534 & ~w63321;
assign w63373 = ~w10714 & ~w10571;
assign w63374 = (w13953 & ~w13689) | (w13953 & w63509) | (~w13689 & w63509);
assign w63375 = w14106 & ~w14104;
assign w63376 = w14546 & ~w14581;
assign w63377 = ~w15914 & w15892;
assign w63378 = w15958 & ~w15975;
assign w63379 = w16006 & w15988;
assign w63380 = w15975 & w15968;
assign w63381 = ~w16723 & ~w16722;
assign w63382 = w17808 & ~w17654;
assign w63383 = (~w18031 & ~w18072) | (~w18031 & w63510) | (~w18072 & w63510);
assign w63384 = ~w18756 & ~w18768;
assign w63385 = ~w63326 & w19772;
assign w63386 = ~w19948 & ~w19933;
assign w63387 = ~w19940 & w19926;
assign w63388 = w24152 & w63511;
assign w63389 = w24403 & w24465;
assign w63390 = ~w23971 & ~w24645;
assign w63391 = ~w23971 & ~w24001;
assign w63392 = w25333 & w25324;
assign w63393 = w25360 & ~w25938;
assign w63394 = w26569 & w26582;
assign w63395 = ~w26726 & w63512;
assign w63396 = ~w27817 & ~w27798;
assign w63397 = w27798 & w27804;
assign w63398 = ~w28195 & ~w28247;
assign w63399 = w29136 & w63513;
assign w63400 = w29134 & w29148;
assign w63401 = ~w29327 & ~w29325;
assign w63402 = w63329 & w30656;
assign w63403 = ~w30693 & w30656;
assign w63404 = ~w30704 & w63514;
assign w63405 = ~w31057 & w31061;
assign w63406 = (~w31839 & ~w31879) | (~w31839 & w31846) | (~w31879 & w31846);
assign w63407 = w32713 & ~w32732;
assign w63408 = ~w33320 & w33288;
assign w63409 = w32788 & ~w32815;
assign w63410 = ~w33338 & ~w33487;
assign w63411 = ~w33845 & ~w33867;
assign w63412 = ~w36918 & ~w36888;
assign w63413 = ~w37859 & ~w37842;
assign w63414 = ~w38114 & ~w38090;
assign w63415 = w38135 & ~w38129;
assign w63416 = w39434 & ~w39419;
assign w63417 = w39443 & ~w39441;
assign w63418 = ~w40148 & w63515;
assign w63419 = ~w42601 & ~w42593;
assign w63420 = w42578 & w42612;
assign w63421 = ~w42992 & ~w43133;
assign w63422 = ~w43136 & ~w42944;
assign w63423 = w43134 & ~w43129;
assign w63424 = ~w43767 & w43704;
assign w63425 = w44036 & ~w44034;
assign w63426 = w43589 & w43564;
assign w63427 = w43538 & ~w44057;
assign w63428 = ~w44156 & w44163;
assign w63429 = ~w45342 & w45325;
assign w63430 = w46606 & w63516;
assign w63431 = w49465 & ~w49448;
assign w63432 = w49465 & ~w49491;
assign w63433 = ~w49360 & ~w49362;
assign w63434 = (~w49373 & ~w49379) | (~w49373 & w63517) | (~w49379 & w63517);
assign w63435 = w49628 & w49373;
assign w63436 = w49978 & ~w49983;
assign w63437 = w50492 & ~w50505;
assign w63438 = w52791 & w63518;
assign w63439 = (w52798 & w63519) | (w52798 & w63520) | (w63519 & w63520);
assign w63440 = w52788 & w52813;
assign w63441 = ~w53036 & ~w53053;
assign w63442 = ~w53614 & ~w53615;
assign w63443 = w55377 & w55422;
assign w63444 = ~w55586 & ~w55585;
assign w63445 = ~w55586 & ~w63333;
assign w63446 = w55564 & w55570;
assign w63447 = ~w56531 & w56525;
assign w63448 = w57023 & ~w57016;
assign w63449 = w57423 & w57469;
assign w63450 = w57815 & w57775;
assign w63451 = ~w57811 & w57807;
assign w63452 = w57822 & ~w57781;
assign w63453 = ~w57866 & ~w57871;
assign w63454 = ~w57869 & ~pi3783;
assign w63455 = w57869 & pi3783;
assign w63456 = w57915 & w57893;
assign w63457 = w58035 & w58050;
assign w63458 = ~w58051 & ~w58096;
assign w63459 = ~w58108 & ~pi3759;
assign w63460 = w58108 & pi3759;
assign w63461 = ~w58243 & w58221;
assign w63462 = w58214 & w58221;
assign w63463 = w58289 & w58300;
assign w63464 = ~w57703 & w57717;
assign w63465 = w58374 & ~w58338;
assign w63466 = w58375 & w58408;
assign w63467 = ~w63334 & ~w58055;
assign w63468 = ~w58415 & w58408;
assign w63469 = ~w57944 & w57902;
assign w63470 = w58761 & ~w58765;
assign w63471 = ~w58568 & ~w58392;
assign w63472 = ~w59280 & ~w59274;
assign w63473 = w59280 & ~w59267;
assign w63474 = w59313 & w59309;
assign w63475 = w59362 & ~w59346;
assign w63476 = w59660 & w59631;
assign w63477 = ~w59648 & w59664;
assign w63478 = ~w59636 & ~w59890;
assign w63479 = ~w59620 & w59651;
assign w63480 = w59648 & ~w59915;
assign w63481 = w59674 & w59267;
assign w63482 = w59927 & w59930;
assign w63483 = w59620 & ~w59602;
assign w63484 = w59596 & ~w59608;
assign w63485 = ~w60369 & w60375;
assign w63486 = w60439 & w60427;
assign w63487 = ~w60655 & w60666;
assign w63488 = ~w60688 & w60648;
assign w63489 = ~w60956 & ~w60928;
assign w63490 = ~w60496 & w60421;
assign w63491 = ~w61357 & ~w61341;
assign w63492 = w61379 & w61382;
assign w63493 = w60934 & ~w61477;
assign w63494 = w61520 & ~w61594;
assign w63495 = w61668 & ~w61662;
assign w63496 = w61662 & w61675;
assign w63497 = w61727 & ~w61707;
assign w63498 = w61731 & ~w61681;
assign w63499 = ~w61750 & w61675;
assign w63500 = ~w61833 & w61820;
assign w63501 = w62080 & w62061;
assign w63502 = ~w62080 & ~w62094;
assign w63503 = ~w62015 & w62003;
assign w63504 = ~w62087 & w62094;
assign w63505 = ~w62795 & ~w62536;
assign w63506 = w62928 & ~w62566;
assign w63507 = w62929 & w62940;
assign w63508 = w6423 & w6386;
assign w63509 = ~w13690 & w13953;
assign w63510 = ~w18043 & ~w18031;
assign w63511 = w24119 & ~w24125;
assign w63512 = ~w26563 & w26604;
assign w63513 = ~w29134 & w29142;
assign w63514 = ~w31051 & w30669;
assign w63515 = ~w40142 & ~w40140;
assign w63516 = ~w46611 & ~w46602;
assign w63517 = w49350 & ~w49373;
assign w63518 = ~w52768 & ~w52776;
assign w63519 = w52769 & ~w52776;
assign w63520 = w52769 & w63438;
assign w63521 = w1459 & w1452;
assign w63522 = w1647 & w1662;
assign w63523 = w1669 & ~w1679;
assign w63524 = w1716 & ~w1420;
assign w63525 = w1420 & w1715;
assign w63526 = w1883 & ~w1876;
assign w63527 = ~w2129 & ~w2136;
assign w63528 = (~w2162 & ~w2149) | (~w2162 & w64360) | (~w2149 & w64360);
assign w63529 = ~w2381 & ~w2361;
assign w63530 = ~w2346 & ~w2347;
assign w63531 = ~w63350 & ~w2624;
assign w63532 = ~w2628 & ~w2623;
assign w63533 = ~w2599 & w2622;
assign w63534 = w2873 & w2844;
assign w63535 = ~w2856 & w2844;
assign w63536 = w2856 & ~w2899;
assign w63537 = w3057 & w64361;
assign w63538 = ~w3049 & w3056;
assign w63539 = ~w3074 & ~w3056;
assign w63540 = ~w3213 & ~w3205;
assign w63541 = w3194 & w3160;
assign w63542 = ~w2968 & w2955;
assign w63543 = ~w3257 & w3279;
assign w63544 = ~w2992 & ~w3005;
assign w63545 = ~w3337 & ~w3070;
assign w63546 = ~w3403 & w3400;
assign w63547 = ~w2775 & ~w3475;
assign w63548 = ~w2881 & w2856;
assign w63549 = ~w3543 & ~w2856;
assign w63550 = ~w3477 & w64362;
assign w63551 = w3696 & w3693;
assign w63552 = w3651 & ~w3688;
assign w63553 = ~w3667 & ~w3651;
assign w63554 = w4448 & ~w4438;
assign w63555 = (w4465 & w4616) | (w4465 & w64363) | (w4616 & w64363);
assign w63556 = ~w4815 & ~w4770;
assign w63557 = ~w4899 & ~w4898;
assign w63558 = ~w5646 & ~w5581;
assign w63559 = ~w5552 & w64364;
assign w63560 = w5551 & w5560;
assign w63561 = w5615 & w64365;
assign w63562 = ~w5698 & ~w5672;
assign w63563 = w5716 & ~w5706;
assign w63564 = w5706 & w5712;
assign w63565 = w5851 & w5848;
assign w63566 = w5528 & w5480;
assign w63567 = ~w5911 & w6007;
assign w63568 = w5648 & w64366;
assign w63569 = ~w6041 & w6058;
assign w63570 = w5724 & ~w5736;
assign w63571 = w5780 & w64367;
assign w63572 = ~w6154 & ~w5748;
assign w63573 = (w6049 & ~w6208) | (w6049 & w64368) | (~w6208 & w64368);
assign w63574 = w6459 & ~w6423;
assign w63575 = ~w6474 & w64369;
assign w63576 = (pi0371 & w6474) | (pi0371 & w64370) | (w6474 & w64370);
assign w63577 = w6666 & w6663;
assign w63578 = w6670 & ~w6682;
assign w63579 = w6828 & ~w6793;
assign w63580 = w6969 & w6993;
assign w63581 = ~w7021 & w64371;
assign w63582 = w7058 & w7017;
assign w63583 = ~w7138 & w7157;
assign w63584 = w7144 & w7163;
assign w63585 = ~w7235 & ~w7193;
assign w63586 = w7253 & w6588;
assign w63587 = w7036 & ~w7055;
assign w63588 = w7151 & w7181;
assign w63589 = w7151 & ~w63364;
assign w63590 = w7479 & w7503;
assign w63591 = ~w7518 & w7512;
assign w63592 = w7572 & ~w7466;
assign w63593 = ~w7951 & w7931;
assign w63594 = ~w7937 & ~w7931;
assign w63595 = w8122 & w8158;
assign w63596 = ~w8034 & ~w8018;
assign w63597 = w7951 & w7918;
assign w63598 = w7924 & ~w7918;
assign w63599 = w8311 & w8314;
assign w63600 = w8685 & w8651;
assign w63601 = ~w8628 & w8663;
assign w63602 = w7985 & w8859;
assign w63603 = ~w8675 & w8627;
assign w63604 = w8946 & ~w8640;
assign w63605 = ~w8985 & w8972;
assign w63606 = ~w8218 & ~w9109;
assign w63607 = ~w9039 & w64372;
assign w63608 = w9163 & ~w9162;
assign w63609 = w9148 & w9164;
assign w63610 = (~w9180 & w9203) | (~w9180 & w64373) | (w9203 & w64373);
assign w63611 = w9355 & ~w9335;
assign w63612 = w9393 & ~w9384;
assign w63613 = ~w9411 & ~w9335;
assign w63614 = ~w9355 & w9341;
assign w63615 = w9367 & w64374;
assign w63616 = w9390 & w9517;
assign w63617 = w9409 & w9406;
assign w63618 = w9727 & w9708;
assign w63619 = ~w9987 & ~w9964;
assign w63620 = w9727 & ~w9708;
assign w63621 = ~w9841 & ~w10142;
assign w63622 = w10075 & w10188;
assign w63623 = w9993 & w9995;
assign w63624 = ~w10403 & w64375;
assign w63625 = ~w10416 & ~w9964;
assign w63626 = ~w10446 & w10453;
assign w63627 = ~w10528 & w10541;
assign w63628 = ~w10563 & ~w10549;
assign w63629 = ~w10558 & w10528;
assign w63630 = ~w10572 & ~w10581;
assign w63631 = w10735 & w64376;
assign w63632 = w10776 & ~w10752;
assign w63633 = w10776 & ~w10760;
assign w63634 = w10982 & ~w10961;
assign w63635 = w11108 & w10499;
assign w63636 = (~w10493 & w11105) | (~w10493 & w64377) | (w11105 & w64377);
assign w63637 = ~w11143 & w11146;
assign w63638 = w11441 & w11400;
assign w63639 = w11360 & w11379;
assign w63640 = w10919 & ~w10808;
assign w63641 = w11746 & w11768;
assign w63642 = w11949 & ~w11972;
assign w63643 = w12059 & w12050;
assign w63644 = w11886 & w11875;
assign w63645 = ~w12118 & ~w12107;
assign w63646 = w11939 & ~w11932;
assign w63647 = ~w12139 & ~w11932;
assign w63648 = w12218 & w12202;
assign w63649 = (w12181 & w12196) | (w12181 & w64378) | (w12196 & w64378);
assign w63650 = ~w12000 & ~w11950;
assign w63651 = w12483 & w12440;
assign w63652 = (w11758 & ~w11778) | (w11758 & w64379) | (~w11778 & w64379);
assign w63653 = ~w12578 & w64380;
assign w63654 = ~w12337 & w12325;
assign w63655 = (~w12667 & w12261) | (~w12667 & w64381) | (w12261 & w64381);
assign w63656 = w12850 & ~w12862;
assign w63657 = ~w12904 & ~w12923;
assign w63658 = w12361 & w64382;
assign w63659 = ~w12378 & w64383;
assign w63660 = w13085 & ~w13091;
assign w63661 = ~w13238 & w64384;
assign w63662 = w13199 & w13152;
assign w63663 = ~w13158 & ~w13178;
assign w63664 = w13371 & w13358;
assign w63665 = w13372 & w13435;
assign w63666 = w13299 & ~w13284;
assign w63667 = (~w13565 & w13589) | (~w13565 & w64385) | (w13589 & w64385);
assign w63668 = w13606 & w13600;
assign w63669 = ~w13684 & ~w13687;
assign w63670 = ~w13695 & ~w13674;
assign w63671 = (w13561 & ~w13612) | (w13561 & w64386) | (~w13612 & w64386);
assign w63672 = ~w13632 & w13663;
assign w63673 = ~w13632 & ~w13645;
assign w63674 = ~w13645 & w13653;
assign w63675 = ~w63374 & ~w13656;
assign w63676 = w13645 & ~w13700;
assign w63677 = w13491 & w13314;
assign w63678 = w13076 & ~w13061;
assign w63679 = ~w14113 & w13780;
assign w63680 = (~w13780 & w14105) | (~w13780 & w64387) | (w14105 & w64387);
assign w63681 = ~w13067 & ~w13091;
assign w63682 = (~w14053 & w14057) | (~w14053 & w64388) | (w14057 & w64388);
assign w63683 = w13911 & ~w13883;
assign w63684 = w14567 & w14545;
assign w63685 = w14580 & ~w14578;
assign w63686 = ~w14584 & ~w14576;
assign w63687 = w14580 & w14612;
assign w63688 = ~w14655 & w14660;
assign w63689 = w14692 & ~w14707;
assign w63690 = w14748 & w14751;
assign w63691 = w14903 & w14896;
assign w63692 = w14908 & w14896;
assign w63693 = ~w15487 & w14746;
assign w63694 = ~w15565 & w15549;
assign w63695 = w15563 & w64389;
assign w63696 = w15549 & ~w15560;
assign w63697 = ~w15660 & w15667;
assign w63698 = ~w15822 & ~w15820;
assign w63699 = w15893 & ~w15878;
assign w63700 = ~w15884 & w15902;
assign w63701 = w15884 & w15890;
assign w63702 = ~w63377 & w15912;
assign w63703 = ~w15981 & w64390;
assign w63704 = w16021 & w15987;
assign w63705 = (w16013 & w16018) | (w16013 & w64391) | (w16018 & w64391);
assign w63706 = w16015 & w64392;
assign w63707 = ~w15905 & w15906;
assign w63708 = w16514 & w16516;
assign w63709 = (~w16493 & ~w16513) | (~w16493 & w64393) | (~w16513 & w64393);
assign w63710 = ~w16006 & w16608;
assign w63711 = (~w16702 & w16723) | (~w16702 & w64394) | (w16723 & w64394);
assign w63712 = w16702 & ~w16748;
assign w63713 = (w16821 & w16817) | (w16821 & w64395) | (w16817 & w64395);
assign w63714 = w16835 & w16812;
assign w63715 = w16134 & ~w16170;
assign w63716 = ~w16723 & w16702;
assign w63717 = (~w16832 & w16834) | (~w16832 & w64396) | (w16834 & w64396);
assign w63718 = ~w17415 & w17402;
assign w63719 = ~w17689 & ~w17920;
assign w63720 = ~w18073 & ~w18067;
assign w63721 = w18150 & ~w18066;
assign w63722 = w18073 & ~w18204;
assign w63723 = ~w18205 & w18206;
assign w63724 = (~w18398 & ~w18463) | (~w18398 & w64397) | (~w18463 & w64397);
assign w63725 = ~w18505 & ~w18552;
assign w63726 = w18560 & ~w18581;
assign w63727 = ~w18770 & w18774;
assign w63728 = ~w18751 & w18768;
assign w63729 = ~w18778 & w18782;
assign w63730 = w18441 & ~w18410;
assign w63731 = w18914 & w18908;
assign w63732 = w19583 & w64398;
assign w63733 = ~w19799 & ~w19811;
assign w63734 = w19977 & ~w19932;
assign w63735 = w19948 & w19962;
assign w63736 = ~w19967 & ~w19939;
assign w63737 = w20374 & w20188;
assign w63738 = ~w20383 & ~w20375;
assign w63739 = w20302 & w20289;
assign w63740 = ~w19720 & ~w19742;
assign w63741 = ~w20544 & w20537;
assign w63742 = w20561 & ~w20569;
assign w63743 = ~w20587 & ~w20676;
assign w63744 = ~w20692 & ~w20472;
assign w63745 = w20789 & ~w20853;
assign w63746 = (~w20799 & ~w20790) | (~w20799 & w64399) | (~w20790 & w64399);
assign w63747 = ~w21017 & w21002;
assign w63748 = ~w21133 & w21139;
assign w63749 = w20944 & w20956;
assign w63750 = w21301 & w21281;
assign w63751 = w21471 & w21454;
assign w63752 = ~w21766 & ~w21758;
assign w63753 = w21789 & w64400;
assign w63754 = w22210 & w22238;
assign w63755 = ~w22210 & w22216;
assign w63756 = ~w22242 & ~w22216;
assign w63757 = w22267 & w22233;
assign w63758 = ~w22463 & w22455;
assign w63759 = w22833 & w22829;
assign w63760 = w22653 & w64401;
assign w63761 = w23073 & ~w23063;
assign w63762 = ~w23027 & ~w23088;
assign w63763 = w23108 & w23115;
assign w63764 = w23137 & w23040;
assign w63765 = w23077 & ~w23039;
assign w63766 = (w23027 & w23144) | (w23027 & w64402) | (w23144 & w64402);
assign w63767 = w22925 & w22931;
assign w63768 = w22965 & ~w23187;
assign w63769 = ~w23542 & ~w23549;
assign w63770 = ~w23718 & ~w23714;
assign w63771 = w23947 & ~w23954;
assign w63772 = ~w23992 & ~w23997;
assign w63773 = w23715 & ~w23698;
assign w63774 = w24030 & ~w23706;
assign w63775 = w24031 & ~w23712;
assign w63776 = ~w24144 & ~w24170;
assign w63777 = w24148 & w24187;
assign w63778 = (w24125 & ~w24159) | (w24125 & w64403) | (~w24159 & w64403);
assign w63779 = ~w24230 & ~w63388;
assign w63780 = w24378 & w24403;
assign w63781 = w24411 & w24371;
assign w63782 = ~w24411 & w24414;
assign w63783 = w24469 & ~w24471;
assign w63784 = w24365 & ~w24494;
assign w63785 = (w24510 & ~w24598) | (w24510 & w64404) | (~w24598 & w64404);
assign w63786 = w24565 & ~w24543;
assign w63787 = (w24645 & w24646) | (w24645 & w64405) | (w24646 & w64405);
assign w63788 = ~w24647 & ~w63390;
assign w63789 = w24125 & w24159;
assign w63790 = (w24184 & w24671) | (w24184 & w64406) | (w24671 & w64406);
assign w63791 = w24170 & w24119;
assign w63792 = w24601 & ~w24539;
assign w63793 = w23987 & ~w24001;
assign w63794 = w23987 & w63391;
assign w63795 = ~w24841 & w24828;
assign w63796 = w25156 & w25143;
assign w63797 = w25166 & w25137;
assign w63798 = (w25360 & w25352) | (w25360 & w64407) | (w25352 & w64407);
assign w63799 = w24841 & w24834;
assign w63800 = (~w25536 & ~w25572) | (~w25536 & w64408) | (~w25572 & w64408);
assign w63801 = ~w25542 & ~w25549;
assign w63802 = w25868 & w25857;
assign w63803 = w25870 & w25820;
assign w63804 = ~w25886 & ~w25880;
assign w63805 = ~w25943 & ~w25935;
assign w63806 = ~w25886 & ~w25896;
assign w63807 = w25849 & w64409;
assign w63808 = ~w26386 & w26369;
assign w63809 = ~w26480 & ~w26486;
assign w63810 = ~w26488 & w26445;
assign w63811 = ~w26454 & w26471;
assign w63812 = w26501 & ~w26460;
assign w63813 = w26480 & w26504;
assign w63814 = ~w26476 & ~w26471;
assign w63815 = w26476 & ~w26445;
assign w63816 = ~w26582 & ~w26589;
assign w63817 = (w26603 & w26593) | (w26603 & w64410) | (w26593 & w64410);
assign w63818 = w26766 & ~w26604;
assign w63819 = w26766 & ~w63395;
assign w63820 = w26762 & w26773;
assign w63821 = w26659 & ~w26681;
assign w63822 = w27054 & w27047;
assign w63823 = ~w27054 & w27056;
assign w63824 = w27169 & w27158;
assign w63825 = ~w26366 & ~w27240;
assign w63826 = w26589 & ~w27255;
assign w63827 = w26835 & w26653;
assign w63828 = ~w27649 & ~w27643;
assign w63829 = w27696 & w27702;
assign w63830 = w27836 & ~w27777;
assign w63831 = ~w27854 & w27856;
assign w63832 = ~w27898 & ~w27906;
assign w63833 = w27466 & w64411;
assign w63834 = ~w27741 & ~w27702;
assign w63835 = ~w27690 & w27749;
assign w63836 = ~w27742 & w64412;
assign w63837 = ~w27619 & w27625;
assign w63838 = w27854 & w28167;
assign w63839 = ~w27783 & ~w27798;
assign w63840 = ~w28188 & ~w28214;
assign w63841 = w27750 & w27719;
assign w63842 = (w28208 & w28222) | (w28208 & w64413) | (w28222 & w64413);
assign w63843 = (w28357 & ~w28354) | (w28357 & w64414) | (~w28354 & w64414);
assign w63844 = ~w28172 & w64415;
assign w63845 = w27619 & ~w27584;
assign w63846 = w27740 & ~w27718;
assign w63847 = w28864 & ~w28871;
assign w63848 = w29064 & ~w29089;
assign w63849 = w29334 & w29148;
assign w63850 = ~w29647 & w29643;
assign w63851 = ~w29640 & ~w29574;
assign w63852 = w29588 & w29608;
assign w63853 = w30149 & w30126;
assign w63854 = (w30246 & w30251) | (w30246 & w64416) | (w30251 & w64416);
assign w63855 = ~w30247 & ~w30252;
assign w63856 = w30272 & ~w30251;
assign w63857 = w30376 & w64417;
assign w63858 = w30682 & w30719;
assign w63859 = ~w30693 & w30806;
assign w63860 = ~w30963 & w64418;
assign w63861 = ~w31060 & ~w31059;
assign w63862 = (pi1648 & w31065) | (pi1648 & w64419) | (w31065 & w64419);
assign w63863 = ~w31065 & w64420;
assign w63864 = ~w30225 & ~w30243;
assign w63865 = ~w31073 & w64421;
assign w63866 = (~pi1651 & w31073) | (~pi1651 & w64422) | (w31073 & w64422);
assign w63867 = ~w31142 & w31161;
assign w63868 = (~w31122 & ~w31165) | (~w31122 & w64423) | (~w31165 & w64423);
assign w63869 = ~w30807 & ~w30800;
assign w63870 = w31486 & ~w31501;
assign w63871 = w31862 & ~w63406;
assign w63872 = w31862 & w31880;
assign w63873 = w31887 & w31833;
assign w63874 = w31893 & w64424;
assign w63875 = w31852 & ~w31845;
assign w63876 = w31933 & ~w31939;
assign w63877 = w31783 & ~w31757;
assign w63878 = w32076 & ~w31982;
assign w63879 = ~w32089 & ~w32086;
assign w63880 = (w32178 & w32190) | (w32178 & w64425) | (w32190 & w64425);
assign w63881 = w32155 & w32184;
assign w63882 = w32210 & ~w32149;
assign w63883 = w32212 & w32215;
assign w63884 = ~w31652 & w31665;
assign w63885 = (w31706 & ~w32248) | (w31706 & w64426) | (~w32248 & w64426);
assign w63886 = w32342 & ~w32354;
assign w63887 = ~w32913 & ~w32920;
assign w63888 = ~w33279 & ~w33288;
assign w63889 = ~w33454 & ~w32788;
assign w63890 = w33325 & w33479;
assign w63891 = ~w33496 & w64427;
assign w63892 = w33696 & w32699;
assign w63893 = w33863 & w33826;
assign w63894 = ~w34179 & ~w34140;
assign w63895 = ~w34293 & w34292;
assign w63896 = ~w34277 & w34270;
assign w63897 = ~w34649 & w34613;
assign w63898 = w34650 & ~w34672;
assign w63899 = ~w34779 & ~w34772;
assign w63900 = ~w34916 & ~w34912;
assign w63901 = (~w34517 & w35096) | (~w34517 & w64428) | (w35096 & w64428);
assign w63902 = w35159 & w64429;
assign w63903 = w35387 & ~w35378;
assign w63904 = ~w35465 & w35472;
assign w63905 = w35665 & w35696;
assign w63906 = ~w35711 & ~w35702;
assign w63907 = ~w35737 & w64430;
assign w63908 = ~w35790 & w64431;
assign w63909 = ~w36046 & ~w36029;
assign w63910 = w35732 & w35701;
assign w63911 = ~w36401 & ~w36395;
assign w63912 = w36404 & w36224;
assign w63913 = w35472 & w35446;
assign w63914 = ~w36797 & w36785;
assign w63915 = ~w36902 & w36875;
assign w63916 = w36888 & w36937;
assign w63917 = ~w36951 & w64432;
assign w63918 = ~w36974 & ~w36981;
assign w63919 = w36974 & w36998;
assign w63920 = w37029 & ~w37006;
assign w63921 = w37113 & w37112;
assign w63922 = ~w37133 & w64433;
assign w63923 = ~w37190 & ~w37198;
assign w63924 = w37177 & ~w37222;
assign w63925 = w36797 & w36805;
assign w63926 = (~w36778 & ~w36846) | (~w36778 & w64434) | (~w36846 & w64434);
assign w63927 = w37022 & w36974;
assign w63928 = ~w37472 & w64435;
assign w63929 = w36917 & w36881;
assign w63930 = w36948 & w64436;
assign w63931 = w37395 & w37357;
assign w63932 = ~w37344 & ~w37401;
assign w63933 = w37522 & ~w37532;
assign w63934 = w37089 & w37076;
assign w63935 = w37121 & ~w37063;
assign w63936 = w37119 & w37101;
assign w63937 = ~w37472 & w64437;
assign w63938 = w37262 & w37222;
assign w63939 = w37644 & w37208;
assign w63940 = w36734 & w36687;
assign w63941 = ~w37720 & ~w37709;
assign w63942 = w36712 & ~w36699;
assign w63943 = (~w36752 & w37736) | (~w36752 & w64438) | (w37736 & w64438);
assign w63944 = w37723 & ~w36693;
assign w63945 = (w37738 & w64439) | (w37738 & w64440) | (w64439 & w64440);
assign w63946 = ~w37745 & w36752;
assign w63947 = w37320 & ~w36805;
assign w63948 = ~w36845 & w37785;
assign w63949 = ~w37821 & w37842;
assign w63950 = (w37828 & w37919) | (w37828 & w64441) | (w37919 & w64441);
assign w63951 = w38149 & w64442;
assign w63952 = ~w38191 & w38197;
assign w63953 = w38479 & w38485;
assign w63954 = w38559 & w38555;
assign w63955 = w38746 & w64443;
assign w63956 = ~w38954 & w38973;
assign w63957 = w38986 & ~w38947;
assign w63958 = w38559 & w38586;
assign w63959 = ~w39201 & w39206;
assign w63960 = w39443 & ~w39432;
assign w63961 = w39453 & ~w39441;
assign w63962 = w39453 & w39445;
assign w63963 = ~w39475 & ~w39452;
assign w63964 = ~w39857 & ~w39862;
assign w63965 = (~w39770 & ~w39806) | (~w39770 & w64444) | (~w39806 & w64444);
assign w63966 = ~w63418 & ~w40138;
assign w63967 = (w40160 & w40148) | (w40160 & w64445) | (w40148 & w64445);
assign w63968 = w39820 & ~w40044;
assign w63969 = w40025 & w39750;
assign w63970 = ~w40310 & ~w40329;
assign w63971 = ~w39464 & ~w40464;
assign w63972 = w40475 & w39472;
assign w63973 = ~w40470 & w64446;
assign w63974 = (~pi2200 & w40470) | (~pi2200 & w64447) | (w40470 & w64447);
assign w63975 = ~w40725 & w40712;
assign w63976 = w40829 & ~w40887;
assign w63977 = w40972 & w40958;
assign w63978 = ~w40860 & ~w40848;
assign w63979 = ~w41372 & ~w41354;
assign w63980 = w41427 & ~w40759;
assign w63981 = ~w41361 & ~w41340;
assign w63982 = w41670 & w64448;
assign w63983 = w41953 & w41986;
assign w63984 = w41960 & ~w41986;
assign w63985 = ~w42004 & w42012;
assign w63986 = w42625 & w42616;
assign w63987 = w42629 & w42633;
assign w63988 = w42944 & w43133;
assign w63989 = (~w42992 & ~w43125) | (~w42992 & w64449) | (~w43125 & w64449);
assign w63990 = ~w43137 & w43171;
assign w63991 = ~w43266 & ~w43251;
assign w63992 = w43250 & w43266;
assign w63993 = w43282 & w64450;
assign w63994 = w43529 & w43563;
assign w63995 = w43745 & w64451;
assign w63996 = ~w43736 & ~w43773;
assign w63997 = ~w43822 & w43795;
assign w63998 = ~w43723 & w43732;
assign w63999 = w44022 & w43744;
assign w64000 = ~w44039 & ~w44032;
assign w64001 = ~w43559 & ~w43564;
assign w64002 = ~w43559 & ~w63426;
assign w64003 = w43574 & w43573;
assign w64004 = w44065 & w44071;
assign w64005 = ~w44128 & ~w44161;
assign w64006 = (~w44149 & w44137) | (~w44149 & w64452) | (w44137 & w64452);
assign w64007 = w44359 & ~w44281;
assign w64008 = w44450 & w44135;
assign w64009 = (w44182 & w44513) | (w44182 & w64453) | (w44513 & w64453);
assign w64010 = ~w44650 & w44641;
assign w64011 = w44675 & ~w44627;
assign w64012 = w44643 & ~w44614;
assign w64013 = w44824 & ~w44804;
assign w64014 = ~w44842 & ~w44845;
assign w64015 = ~w44871 & ~w44878;
assign w64016 = ~w44547 & ~w44574;
assign w64017 = w44564 & w64454;
assign w64018 = ~w45034 & w64455;
assign w64019 = w45183 & ~w45229;
assign w64020 = w45233 & w45190;
assign w64021 = ~w45325 & ~w45306;
assign w64022 = w45397 & ~w45372;
assign w64023 = w45342 & w45333;
assign w64024 = (~w45879 & w45881) | (~w45879 & w64456) | (w45881 & w64456);
assign w64025 = ~w45881 & w64457;
assign w64026 = ~w45854 & ~w45876;
assign w64027 = ~w45942 & w64458;
assign w64028 = (~pi2474 & w45942) | (~pi2474 & w64459) | (w45942 & w64459);
assign w64029 = w46385 & w46322;
assign w64030 = w46427 & w46209;
assign w64031 = ~w46603 & w46602;
assign w64032 = ~w46603 & ~w63430;
assign w64033 = w46777 & w46763;
assign w64034 = ~w47296 & w47324;
assign w64035 = w47324 & w47315;
assign w64036 = w47437 & ~w47458;
assign w64037 = ~w47570 & w47586;
assign w64038 = ~w47596 & ~w47569;
assign w64039 = w47597 & ~w47623;
assign w64040 = w47920 & ~w47925;
assign w64041 = w48439 & ~w48436;
assign w64042 = w48531 & ~w48553;
assign w64043 = ~w48816 & w48797;
assign w64044 = w48898 & ~w48911;
assign w64045 = w48841 & w48861;
assign w64046 = ~w49204 & ~w48985;
assign w64047 = w49258 & w49295;
assign w64048 = (w48937 & w48966) | (w48937 & w64460) | (w48966 & w64460);
assign w64049 = w49493 & ~w49442;
assign w64050 = w49475 & ~w49485;
assign w64051 = w49448 & ~w49491;
assign w64052 = w49534 & ~w49541;
assign w64053 = ~w49343 & w49360;
assign w64054 = w49343 & w49362;
assign w64055 = w49343 & ~w63433;
assign w64056 = w49624 & w49634;
assign w64057 = w49636 & ~w49625;
assign w64058 = ~w49373 & ~w49777;
assign w64059 = w49942 & w49936;
assign w64060 = ~w49958 & w64461;
assign w64061 = w50199 & ~w50190;
assign w64062 = w50212 & ~w50171;
assign w64063 = ~w50225 & w50224;
assign w64064 = ~w50165 & w50177;
assign w64065 = w50242 & ~w50208;
assign w64066 = ~w50285 & ~w50300;
assign w64067 = w50521 & ~w50514;
assign w64068 = w50827 & ~w50824;
assign w64069 = w50500 & w50505;
assign w64070 = w50500 & ~w63437;
assign w64071 = ~w50492 & ~w50472;
assign w64072 = w51129 & ~w51160;
assign w64073 = w51129 & ~w51148;
assign w64074 = w51129 & w51142;
assign w64075 = w51282 & ~w51308;
assign w64076 = w51129 & ~w51123;
assign w64077 = ~w51671 & w51677;
assign w64078 = w51465 & w51533;
assign w64079 = ~w51845 & w51852;
assign w64080 = w51604 & ~w52113;
assign w64081 = w51364 & w51395;
assign w64082 = w52141 & w64462;
assign w64083 = ~w52216 & ~w52210;
assign w64084 = ~w52544 & w52531;
assign w64085 = ~w52442 & ~w52436;
assign w64086 = w52448 & ~w52460;
assign w64087 = w52606 & w52613;
assign w64088 = w52604 & ~w52622;
assign w64089 = w52782 & ~w52788;
assign w64090 = (~w52756 & ~w52824) | (~w52756 & w64463) | (~w52824 & w64463);
assign w64091 = ~w52838 & w52840;
assign w64092 = ~w53052 & ~w53050;
assign w64093 = ~w53163 & ~w53160;
assign w64094 = w53182 & ~w53188;
assign w64095 = ~w53216 & ~w53090;
assign w64096 = ~w53017 & ~w53208;
assign w64097 = ~w53045 & w64464;
assign w64098 = w52782 & w52768;
assign w64099 = ~w53242 & ~w52756;
assign w64100 = w52788 & w52762;
assign w64101 = ~w52794 & w52820;
assign w64102 = ~w53156 & ~w53122;
assign w64103 = w53030 & ~w53017;
assign w64104 = ~w52954 & ~w52917;
assign w64105 = w53438 & w64465;
assign w64106 = ~w53305 & w64466;
assign w64107 = ~w53513 & w53510;
assign w64108 = w53562 & ~w53561;
assign w64109 = ~w53479 & ~w53509;
assign w64110 = (w53531 & w64467) | (w53531 & w64468) | (w64467 & w64468);
assign w64111 = w53731 & w53751;
assign w64112 = (w54020 & w54014) | (w54020 & w64469) | (w54014 & w64469);
assign w64113 = w54138 & w54142;
assign w64114 = w54113 & w64470;
assign w64115 = ~w53996 & ~w54291;
assign w64116 = w54089 & ~w54124;
assign w64117 = w54942 & w54944;
assign w64118 = ~w55079 & w55078;
assign w64119 = ~w55579 & w55558;
assign w64120 = ~w55628 & w64471;
assign w64121 = w55390 & w55377;
assign w64122 = w55845 & w55410;
assign w64123 = ~w55848 & ~w55399;
assign w64124 = ~w55858 & w67189;
assign w64125 = ~w55438 & w55383;
assign w64126 = ~w55603 & w55831;
assign w64127 = ~w55596 & w64472;
assign w64128 = ~w56254 & w56258;
assign w64129 = w56271 & ~w56040;
assign w64130 = ~w56541 & ~w56524;
assign w64131 = w56524 & w56541;
assign w64132 = ~w56576 & w64473;
assign w64133 = (w56558 & ~w56551) | (w56558 & w64474) | (~w56551 & w64474);
assign w64134 = ~w56653 & w56641;
assign w64135 = ~w56594 & w56562;
assign w64136 = w57023 & w57016;
assign w64137 = ~w57278 & ~w57046;
assign w64138 = ~w56461 & w56448;
assign w64139 = ~w57424 & w57416;
assign w64140 = w57471 & ~w57463;
assign w64141 = w57478 & ~w57428;
assign w64142 = ~w57577 & w64475;
assign w64143 = ~w57687 & ~w57702;
assign w64144 = ~w57663 & w57710;
assign w64145 = ~w57731 & ~w57727;
assign w64146 = ~w57737 & w57725;
assign w64147 = w57813 & w57840;
assign w64148 = w57844 & ~w57840;
assign w64149 = w57848 & w57840;
assign w64150 = w57848 & ~w64148;
assign w64151 = w57849 & ~pi3763;
assign w64152 = ~w57849 & pi3763;
assign w64153 = ~w57857 & ~w57798;
assign w64154 = w57864 & w57840;
assign w64155 = w57908 & w57893;
assign w64156 = ~w57934 & ~w57999;
assign w64157 = ~w58105 & w58106;
assign w64158 = w58123 & ~w57807;
assign w64159 = ~w57833 & w58132;
assign w64160 = ~w58133 & pi3778;
assign w64161 = w58133 & ~pi3778;
assign w64162 = ~w58160 & ~w58146;
assign w64163 = w57725 & ~w57710;
assign w64164 = w58172 & w57717;
assign w64165 = w57744 & ~w57717;
assign w64166 = w57754 & pi3849;
assign w64167 = ~w57754 & ~pi3849;
assign w64168 = w58201 & ~w58233;
assign w64169 = ~w58233 & ~w58247;
assign w64170 = w58215 & w58257;
assign w64171 = w58243 & w58233;
assign w64172 = ~w58240 & ~w58300;
assign w64173 = ~w58240 & ~w63463;
assign w64174 = ~w58301 & ~pi3843;
assign w64175 = w58301 & pi3843;
assign w64176 = w58358 & w58350;
assign w64177 = w58358 & w58364;
assign w64178 = ~w58417 & pi3764;
assign w64179 = w58417 & ~pi3764;
assign w64180 = ~w58425 & w58092;
assign w64181 = w58430 & ~w58092;
assign w64182 = ~w57928 & ~w57893;
assign w64183 = w58449 & w58455;
assign w64184 = w58514 & w58520;
assign w64185 = w58527 & ~w58548;
assign w64186 = w58380 & ~w58358;
assign w64187 = w58605 & ~w57717;
assign w64188 = ~w58291 & ~w58240;
assign w64189 = w58291 & ~w58632;
assign w64190 = w58633 & w58240;
assign w64191 = w58640 & pi3864;
assign w64192 = ~w58640 & ~pi3864;
assign w64193 = w58358 & w58331;
assign w64194 = w58650 & w58408;
assign w64195 = ~w58686 & ~w58715;
assign w64196 = w57934 & ~w57935;
assign w64197 = ~w57923 & ~w58770;
assign w64198 = ~w58794 & ~w58492;
assign w64199 = w58797 & ~w58537;
assign w64200 = w58819 & w58706;
assign w64201 = w58686 & w58840;
assign w64202 = w58847 & ~w58706;
assign w64203 = w58679 & w58686;
assign w64204 = w58868 & ~w58706;
assign w64205 = w58891 & ~w58408;
assign w64206 = w58886 & pi3841;
assign w64207 = ~w58886 & ~pi3841;
assign w64208 = w58221 & w58233;
assign w64209 = w58931 & w58240;
assign w64210 = w58641 & ~w58233;
assign w64211 = ~w59023 & ~w59022;
assign w64212 = w58976 & ~w59002;
assign w64213 = w59053 & ~w59010;
assign w64214 = w59078 & w59095;
assign w64215 = ~w59085 & ~w59102;
assign w64216 = w59140 & ~w59105;
assign w64217 = w59132 & ~w59134;
assign w64218 = w59160 & ~w59166;
assign w64219 = w59181 & w59173;
assign w64220 = w59378 & w59333;
assign w64221 = ~w59333 & w59381;
assign w64222 = w59466 & ~w59439;
assign w64223 = w59433 & w59459;
assign w64224 = ~w59433 & ~w59484;
assign w64225 = w59515 & ~w59465;
assign w64226 = w59522 & w58982;
assign w64227 = w59527 & pi5191;
assign w64228 = ~w59527 & ~pi5191;
assign w64229 = w59479 & w59560;
assign w64230 = w59651 & ~w59650;
assign w64231 = w59596 & w59620;
assign w64232 = w59662 & ~w59631;
assign w64233 = w59662 & ~w63476;
assign w64234 = ~w59663 & ~pi5098;
assign w64235 = w59663 & pi5098;
assign w64236 = ~w59309 & ~w59295;
assign w64237 = w59733 & ~w58982;
assign w64238 = ~w59751 & w59485;
assign w64239 = w59466 & w59439;
assign w64240 = ~w59755 & ~w59439;
assign w64241 = ~w59679 & w59267;
assign w64242 = w59806 & w59803;
assign w64243 = w59815 & ~w59295;
assign w64244 = w59160 & w59181;
assign w64245 = ~w59629 & ~w59648;
assign w64246 = w59655 & w59631;
assign w64247 = w59655 & w63476;
assign w64248 = w59903 & pi5301;
assign w64249 = ~w59903 & ~pi5301;
assign w64250 = ~w59923 & ~pi5356;
assign w64251 = w59923 & pi5356;
assign w64252 = ~w59965 & ~w59166;
assign w64253 = ~w59196 & w59967;
assign w64254 = w59891 & w59648;
assign w64255 = ~w59993 & ~w59612;
assign w64256 = ~w59140 & w59107;
assign w64257 = w59135 & w59095;
assign w64258 = w59133 & ~w59085;
assign w64259 = w60100 & ~w60120;
assign w64260 = w60093 & w60141;
assign w64261 = w59894 & ~w59997;
assign w64262 = w60106 & ~w60120;
assign w64263 = ~w63485 & ~w60368;
assign w64264 = ~w60323 & w60363;
assign w64265 = w60403 & ~w60411;
assign w64266 = ~w60455 & ~w60427;
assign w64267 = ~w60427 & w60439;
assign w64268 = w63486 & w60455;
assign w64269 = ~w60497 & ~w60495;
assign w64270 = ~w60329 & ~w60405;
assign w64271 = w60614 & ~w60590;
assign w64272 = w60655 & w60666;
assign w64273 = ~w60691 & w60697;
assign w64274 = w60636 & ~w60655;
assign w64275 = w60666 & w60683;
assign w64276 = w60708 & w60707;
assign w64277 = w60716 & ~w60636;
assign w64278 = w60684 & ~w60673;
assign w64279 = ~w60744 & ~w60751;
assign w64280 = w60323 & w60329;
assign w64281 = w60762 & w60761;
assign w64282 = ~w60826 & ~w60786;
assign w64283 = w60913 & ~w60716;
assign w64284 = w60912 & ~w60906;
assign w64285 = ~w60947 & ~w60928;
assign w64286 = w60980 & w61005;
assign w64287 = w60998 & pi8629;
assign w64288 = ~w60998 & ~pi8629;
assign w64289 = w61077 & ~w61063;
assign w64290 = w61097 & w60928;
assign w64291 = ~w61124 & w60561;
assign w64292 = w61168 & w61174;
assign w64293 = ~w60446 & ~w60455;
assign w64294 = w61252 & w61259;
assign w64295 = w61264 & ~w60571;
assign w64296 = ~w61361 & ~w61371;
assign w64297 = w61335 & ~w61350;
assign w64298 = w61370 & ~w61382;
assign w64299 = w61370 & ~w63492;
assign w64300 = w60470 & w61404;
assign w64301 = ~w61168 & ~w61446;
assign w64302 = w61461 & ~w61168;
assign w64303 = w61219 & w61201;
assign w64304 = w60928 & w61477;
assign w64305 = w60928 & ~w63493;
assign w64306 = ~w61483 & pi8528;
assign w64307 = w61483 & ~pi8528;
assign w64308 = ~w61356 & w61382;
assign w64309 = ~w61551 & w61447;
assign w64310 = ~w60956 & ~w60941;
assign w64311 = w60999 & w60955;
assign w64312 = w61316 & w61350;
assign w64313 = w61618 & ~pi8601;
assign w64314 = ~w61618 & pi8601;
assign w64315 = w61644 & ~w61652;
assign w64316 = ~w61701 & w61721;
assign w64317 = ~w61662 & ~w61681;
assign w64318 = w61774 & pi8716;
assign w64319 = ~w61774 & ~pi8716;
assign w64320 = w61840 & ~w61846;
assign w64321 = ~w61811 & w61824;
assign w64322 = w61802 & w61789;
assign w64323 = w62029 & w61995;
assign w64324 = w62087 & ~w62094;
assign w64325 = ~w62098 & ~w62121;
assign w64326 = ~w62121 & ~w62136;
assign w64327 = w62130 & ~w62094;
assign w64328 = w61974 & w61994;
assign w64329 = ~w62284 & ~w61968;
assign w64330 = ~w62019 & ~w62040;
assign w64331 = w61974 & ~w61968;
assign w64332 = ~w62337 & ~pi8744;
assign w64333 = w62337 & pi8744;
assign w64334 = w62343 & ~w62345;
assign w64335 = w62349 & w62350;
assign w64336 = w62367 & w62380;
assign w64337 = w62455 & ~w62244;
assign w64338 = w62201 & w62214;
assign w64339 = ~w61701 & w62508;
assign w64340 = w62543 & w61930;
assign w64341 = ~w62573 & ~w62602;
assign w64342 = ~w62596 & w62609;
assign w64343 = ~w62573 & w62629;
assign w64344 = w62387 & ~w62374;
assign w64345 = ~w62387 & w62380;
assign w64346 = ~w62466 & w62445;
assign w64347 = w62166 & w62094;
assign w64348 = w62733 & ~w62718;
assign w64349 = w62740 & ~w61789;
assign w64350 = w62776 & ~w62585;
assign w64351 = ~w62800 & w61930;
assign w64352 = w61930 & w62815;
assign w64353 = w62865 & w62408;
assign w64354 = w62680 & ~w62408;
assign w64355 = ~w61796 & ~w61811;
assign w64356 = w62889 & w62890;
assign w64357 = w62010 & ~w62295;
assign w64358 = w62579 & ~w62600;
assign w64359 = w62566 & ~w62964;
assign w64360 = w2145 & ~w2162;
assign w64361 = ~w3082 & ~w3065;
assign w64362 = ~w2758 & w2792;
assign w64363 = ~w4617 & w4465;
assign w64364 = ~w5560 & w5581;
assign w64365 = w5629 & w5581;
assign w64366 = ~w5609 & w5573;
assign w64367 = w5707 & ~w5678;
assign w64368 = w6202 & w6049;
assign w64369 = ~w6412 & ~pi0371;
assign w64370 = w6412 & pi0371;
assign w64371 = ~w7020 & ~w6976;
assign w64372 = w8225 & ~w8245;
assign w64373 = w9197 & ~w9180;
assign w64374 = w63614 & w9335;
assign w64375 = ~w10235 & w9964;
assign w64376 = ~w10734 & w10522;
assign w64377 = w10486 & ~w10493;
assign w64378 = ~w12202 & w12181;
assign w64379 = w11746 & w11758;
assign w64380 = w11761 & w11787;
assign w64381 = w12257 & ~w12667;
assign w64382 = ~w12331 & ~w12370;
assign w64383 = ~w13009 & w12370;
assign w64384 = ~w13185 & ~w13199;
assign w64385 = w13561 & ~w13565;
assign w64386 = w13724 & w13561;
assign w64387 = ~w13742 & ~w13780;
assign w64388 = w14058 & ~w14053;
assign w64389 = w15560 & ~w15549;
assign w64390 = ~w15987 & ~w16013;
assign w64391 = w16016 & w16013;
assign w64392 = w15957 & ~w15975;
assign w64393 = ~w16465 & ~w16493;
assign w64394 = w16722 & ~w16702;
assign w64395 = w16702 & w16821;
assign w64396 = ~w16702 & ~w16832;
assign w64397 = ~w18423 & ~w18398;
assign w64398 = w19421 & ~w19262;
assign w64399 = w20789 & ~w20799;
assign w64400 = ~w21766 & w21783;
assign w64401 = ~w22634 & w22641;
assign w64402 = w23072 & w23027;
assign w64403 = w24119 & w24125;
assign w64404 = ~w24522 & w24510;
assign w64405 = ~w23971 & w24645;
assign w64406 = w24679 & w24184;
assign w64407 = w25353 & w25360;
assign w64408 = w25555 & ~w25536;
assign w64409 = ~w25858 & ~w25820;
assign w64410 = ~w26583 & w26603;
assign w64411 = ~w27474 & w27493;
assign w64412 = w27709 & w27715;
assign w64413 = ~w28195 & w28208;
assign w64414 = w28343 & w28357;
assign w64415 = w27783 & w27777;
assign w64416 = w30255 & w30246;
assign w64417 = w30310 & ~w30379;
assign w64418 = ~w30745 & ~w30558;
assign w64419 = ~w31069 & pi1648;
assign w64420 = w31069 & ~pi1648;
assign w64421 = ~w31091 & pi1651;
assign w64422 = w31091 & ~pi1651;
assign w64423 = ~w31135 & ~w31122;
assign w64424 = w31894 & ~w31827;
assign w64425 = w32192 & w32178;
assign w64426 = ~w32251 & w31706;
assign w64427 = ~w33288 & w33296;
assign w64428 = w34503 & ~w34517;
assign w64429 = ~w35127 & ~w35156;
assign w64430 = ~w35708 & w35719;
assign w64431 = ~w35787 & ~w35758;
assign w64432 = w36958 & w36869;
assign w64433 = w37144 & ~w37103;
assign w64434 = ~w36805 & ~w36778;
assign w64435 = w36998 & w37006;
assign w64436 = w36919 & w36869;
assign w64437 = w36998 & w37024;
assign w64438 = w36763 & ~w36752;
assign w64439 = w37747 & ~w36752;
assign w64440 = w37747 & w63943;
assign w64441 = w37920 & w37828;
assign w64442 = w38148 & ~w38126;
assign w64443 = w38450 & ~w38459;
assign w64444 = ~w39783 & ~w39770;
assign w64445 = w40142 & w40160;
assign w64446 = ~w39472 & pi2200;
assign w64447 = w39472 & ~pi2200;
assign w64448 = ~w41669 & w41646;
assign w64449 = w43123 & ~w42992;
assign w64450 = w63992 & ~w43244;
assign w64451 = ~w43704 & w43717;
assign w64452 = ~w44150 & ~w44149;
assign w64453 = w44511 & w44182;
assign w64454 = w44554 & w44547;
assign w64455 = ~w45029 & ~w45012;
assign w64456 = ~w45882 & ~w45879;
assign w64457 = w45882 & w45876;
assign w64458 = ~w45894 & pi2474;
assign w64459 = w45894 & ~pi2474;
assign w64460 = w49420 & w48937;
assign w64461 = ~w49930 & ~w49917;
assign w64462 = w51424 & w51422;
assign w64463 = w52819 & ~w52756;
assign w64464 = w53030 & w53017;
assign w64465 = ~w53363 & w53447;
assign w64466 = ~w53156 & w53129;
assign w64467 = w53613 & w53509;
assign w64468 = w53613 & ~w64109;
assign w64469 = w54011 & w54020;
assign w64470 = w54082 & ~w54069;
assign w64471 = ~w55585 & w55558;
assign w64472 = ~w55579 & w55621;
assign w64473 = ~w56535 & ~w56531;
assign w64474 = w56550 & w56558;
assign w64475 = w57464 & ~w57413;
assign w64476 = ~w18 & ~w46;
assign w64477 = ~w168 & w194;
assign w64478 = w475 & ~w456;
assign w64479 = ~w475 & ~w468;
assign w64480 = ~w826 & ~w504;
assign w64481 = ~w838 & w841;
assign w64482 = ~w231 & w237;
assign w64483 = ~w786 & w779;
assign w64484 = ~w1116 & ~w1128;
assign w64485 = ~w1307 & ~w1296;
assign w64486 = w1306 & ~w1317;
assign w64487 = ~w1324 & w1315;
assign w64488 = ~w1268 & ~w1274;
assign w64489 = ~w1379 & ~w1389;
assign w64490 = ~w1401 & ~w1425;
assign w64491 = ~w1459 & ~w1473;
assign w64492 = w1523 & ~w1446;
assign w64493 = ~w1474 & w1490;
assign w64494 = ~w1607 & ~w1347;
assign w64495 = w1685 & ~w1640;
assign w64496 = ~w1687 & w1679;
assign w64497 = w1722 & ~w1387;
assign w64498 = ~w1392 & w1399;
assign w64499 = ~w1387 & w1741;
assign w64500 = w1452 & ~w1459;
assign w64501 = w1543 & w1490;
assign w64502 = ~w1667 & ~w1662;
assign w64503 = ~w1640 & ~w1679;
assign w64504 = w1669 & ~w1816;
assign w64505 = ~w1836 & ~w1830;
assign w64506 = w1836 & w1830;
assign w64507 = ~w1836 & w1849;
assign w64508 = w1901 & w1902;
assign w64509 = ~w1392 & w1408;
assign w64510 = w1366 & ~w1399;
assign w64511 = ~w1387 & ~w1956;
assign w64512 = w1973 & w1974;
assign w64513 = ~w2010 & w1984;
assign w64514 = ~w2041 & ~w2048;
assign w64515 = ~w2075 & ~w1871;
assign w64516 = ~w2087 & ~w1868;
assign w64517 = w1860 & w1868;
assign w64518 = w2078 & ~w2097;
assign w64519 = ~w63528 & w2116;
assign w64520 = w2144 & w2136;
assign w64521 = w2150 & w2171;
assign w64522 = ~w1984 & w2048;
assign w64523 = ~w1655 & ~w1816;
assign w64524 = ~w2245 & ~w2244;
assign w64525 = w1647 & w1640;
assign w64526 = w2251 & w1679;
assign w64527 = ~w1849 & w2195;
assign w64528 = ~w1830 & w1868;
assign w64529 = w2280 & ~pi0175;
assign w64530 = ~w2280 & pi0175;
assign w64531 = ~w2293 & w2145;
assign w64532 = ~w2299 & ~w2297;
assign w64533 = ~w2149 & ~w2285;
assign w64534 = w2301 & pi0170;
assign w64535 = ~w2301 & ~pi0170;
assign w64536 = w2347 & w2356;
assign w64537 = ~w2348 & ~w2356;
assign w64538 = w2346 & ~w2388;
assign w64539 = ~w2064 & w1991;
assign w64540 = w1984 & w2010;
assign w64541 = w2295 & ~w2171;
assign w64542 = w2293 & w2298;
assign w64543 = w2442 & pi0178;
assign w64544 = ~w2442 & ~pi0178;
assign w64545 = w2222 & ~w2058;
assign w64546 = ~w2346 & w2468;
assign w64547 = ~w2346 & ~w2380;
assign w64548 = w2373 & ~w2484;
assign w64549 = w2337 & ~w2468;
assign w64550 = w2381 & w2373;
assign w64551 = w2607 & ~w2638;
assign w64552 = ~w2599 & ~w2607;
assign w64553 = w2656 & ~w2628;
assign w64554 = w2607 & w2599;
assign w64555 = w2657 & pi0233;
assign w64556 = ~w2657 & ~pi0233;
assign w64557 = ~w2651 & w2587;
assign w64558 = w2656 & ~w2587;
assign w64559 = ~w2587 & ~w2718;
assign w64560 = w2880 & w2879;
assign w64561 = w2883 & ~w2872;
assign w64562 = w2863 & w2869;
assign w64563 = w2801 & w2744;
assign w64564 = ~w3059 & w3057;
assign w64565 = w3072 & ~w3037;
assign w64566 = w3037 & w3059;
assign w64567 = ~w3125 & pi0228;
assign w64568 = w3125 & ~pi0228;
assign w64569 = w3103 & ~w3037;
assign w64570 = w3210 & w3173;
assign w64571 = ~w3227 & ~w3154;
assign w64572 = w3213 & w3154;
assign w64573 = w3228 & pi0226;
assign w64574 = ~w3228 & ~pi0226;
assign w64575 = ~w2962 & ~w2982;
assign w64576 = ~w3281 & ~w3014;
assign w64577 = w3275 & ~w2974;
assign w64578 = ~w3297 & pi0235;
assign w64579 = w3297 & ~pi0235;
assign w64580 = w3302 & ~w3154;
assign w64581 = w3304 & w3154;
assign w64582 = w3082 & w3097;
assign w64583 = w3355 & ~pi0238;
assign w64584 = ~w3355 & pi0238;
assign w64585 = ~w3364 & w3377;
assign w64586 = ~w3385 & ~w3377;
assign w64587 = w3402 & ~w3389;
assign w64588 = ~w3469 & pi0239;
assign w64589 = w3469 & ~pi0239;
assign w64590 = ~w2775 & w2751;
assign w64591 = ~w2729 & ~w2762;
assign w64592 = w2735 & ~w2751;
assign w64593 = w3488 & w2792;
assign w64594 = w3235 & ~w3154;
assign w64595 = ~w2850 & w2863;
assign w64596 = w3542 & ~w3514;
assign w64597 = w2880 & w3550;
assign w64598 = w3546 & ~w3541;
assign w64599 = ~w2885 & w3563;
assign w64600 = ~w3619 & ~w2929;
assign w64601 = ~w3634 & ~w2792;
assign w64602 = ~w3634 & ~w63550;
assign w64603 = w3669 & w3680;
assign w64604 = ~w3658 & w3667;
assign w64605 = w3672 & w3651;
assign w64606 = ~w3688 & w3659;
assign w64607 = ~w3645 & ~w3732;
assign w64608 = ~w3740 & w3680;
assign w64609 = w3747 & ~w3680;
assign w64610 = ~w3652 & w3692;
assign w64611 = ~w3789 & ~w3795;
assign w64612 = ~w3797 & pi0260;
assign w64613 = w3797 & ~pi0260;
assign w64614 = ~w3688 & w3807;
assign w64615 = w3412 & ~w3392;
assign w64616 = w3832 & w3421;
assign w64617 = ~w3951 & w3907;
assign w64618 = w3953 & w3926;
assign w64619 = w4137 & w4113;
assign w64620 = w3890 & ~w3884;
assign w64621 = ~w4223 & pi0290;
assign w64622 = w4223 & ~pi0290;
assign w64623 = w4228 & w4045;
assign w64624 = w4332 & w4344;
assign w64625 = w4378 & ~w4300;
assign w64626 = w4204 & ~w3926;
assign w64627 = w4392 & w3907;
assign w64628 = ~w4451 & w4425;
assign w64629 = w4424 & w4473;
assign w64630 = ~w4562 & ~w4539;
assign w64631 = ~w4594 & pi0299;
assign w64632 = w4594 & ~pi0299;
assign w64633 = w4437 & ~w4431;
assign w64634 = w4619 & pi0289;
assign w64635 = ~w4619 & ~pi0289;
assign w64636 = ~w4370 & w4325;
assign w64637 = ~w4343 & ~w4656;
assign w64638 = w4651 & pi0297;
assign w64639 = ~w4651 & ~pi0297;
assign w64640 = ~w4356 & w4343;
assign w64641 = ~w4672 & w4306;
assign w64642 = ~w4670 & ~pi0307;
assign w64643 = w4670 & pi0307;
assign w64644 = w4731 & ~w4706;
assign w64645 = ~w4809 & ~w4751;
assign w64646 = w4797 & w4706;
assign w64647 = w4807 & ~w4825;
assign w64648 = ~w4831 & w4560;
assign w64649 = w4897 & ~w4912;
assign w64650 = w4883 & ~w4902;
assign w64651 = w4914 & w4883;
assign w64652 = w4928 & ~w4931;
assign w64653 = w4913 & pi0298;
assign w64654 = ~w4913 & ~pi0298;
assign w64655 = ~w4950 & ~w4912;
assign w64656 = w4971 & ~pi0320;
assign w64657 = ~w4971 & pi0320;
assign w64658 = w4125 & w4113;
assign w64659 = ~w4437 & ~w4424;
assign w64660 = ~w4456 & ~w4424;
assign w64661 = ~w4873 & ~w4859;
assign w64662 = w4873 & w4859;
assign w64663 = ~w4454 & w4424;
assign w64664 = w4602 & w5213;
assign w64665 = w5237 & w5244;
assign w64666 = ~w5448 & ~w5483;
assign w64667 = w5455 & w5494;
assign w64668 = w5489 & ~w5480;
assign w64669 = w5493 & w5509;
assign w64670 = ~w5590 & w5586;
assign w64671 = w5551 & w5608;
assign w64672 = ~w5614 & ~w5581;
assign w64673 = ~w5618 & ~w5575;
assign w64674 = ~w5600 & ~w63559;
assign w64675 = ~w5600 & ~w5582;
assign w64676 = ~w5661 & pi0367;
assign w64677 = w5661 & ~pi0367;
assign w64678 = ~w5736 & ~w5751;
assign w64679 = w5758 & pi0360;
assign w64680 = ~w5758 & ~pi0360;
assign w64681 = w5775 & w5736;
assign w64682 = ~w5822 & ~w5845;
assign w64683 = ~w5854 & ~w5847;
assign w64684 = ~w5882 & pi0364;
assign w64685 = w5882 & ~pi0364;
assign w64686 = w5906 & pi0381;
assign w64687 = ~w5906 & ~pi0381;
assign w64688 = w5995 & ~w5993;
assign w64689 = w5996 & w5999;
assign w64690 = w5551 & ~w5583;
assign w64691 = w5560 & w5574;
assign w64692 = ~w6004 & ~w6007;
assign w64693 = ~w6004 & ~w63567;
assign w64694 = ~w6011 & ~w5573;
assign w64695 = ~w6011 & ~w63568;
assign w64696 = w6061 & ~w6049;
assign w64697 = ~w6035 & w6022;
assign w64698 = ~w6078 & ~w6084;
assign w64699 = w6113 & ~w5267;
assign w64700 = w5775 & w5715;
assign w64701 = w5679 & w5692;
assign w64702 = w6149 & pi0362;
assign w64703 = ~w6149 & ~pi0362;
assign w64704 = w6169 & ~w5855;
assign w64705 = ~w6035 & ~w6022;
assign w64706 = w6028 & ~w6058;
assign w64707 = w6049 & w6212;
assign w64708 = w6213 & ~pi0365;
assign w64709 = ~w6213 & pi0365;
assign w64710 = ~w5323 & w5353;
assign w64711 = w5329 & w5336;
assign w64712 = w5382 & ~w6243;
assign w64713 = w6220 & w6241;
assign w64714 = w6255 & ~w6251;
assign w64715 = w6270 & ~w6262;
assign w64716 = w6035 & w6058;
assign w64717 = ~w6041 & ~w6058;
assign w64718 = w6041 & ~w6049;
assign w64719 = ~w5336 & w5353;
assign w64720 = ~w6316 & ~w5361;
assign w64721 = w6424 & w6412;
assign w64722 = w6434 & w6433;
assign w64723 = ~w6434 & w6400;
assign w64724 = w6449 & ~pi0369;
assign w64725 = ~w6449 & pi0369;
assign w64726 = w6508 & w6423;
assign w64727 = w6582 & ~w6588;
assign w64728 = w6670 & w6676;
assign w64729 = ~w6700 & pi0422;
assign w64730 = w6700 & ~pi0422;
assign w64731 = w6664 & ~w6660;
assign w64732 = ~w6651 & w6629;
assign w64733 = ~w6649 & ~w6660;
assign w64734 = ~w6724 & w6623;
assign w64735 = ~w6718 & pi0420;
assign w64736 = w6718 & ~pi0420;
assign w64737 = w6833 & w6786;
assign w64738 = w6812 & w6799;
assign w64739 = w6836 & ~w6776;
assign w64740 = w6931 & w6919;
assign w64741 = w6908 & w6939;
assign w64742 = w6919 & w6956;
assign w64743 = ~w6993 & ~w7001;
assign w64744 = w7028 & ~w7022;
assign w64745 = w7028 & ~w63581;
assign w64746 = w7035 & w7034;
assign w64747 = w7040 & w7039;
assign w64748 = ~w7029 & ~pi0429;
assign w64749 = w7029 & pi0429;
assign w64750 = w7061 & ~w7028;
assign w64751 = ~w6982 & ~w7008;
assign w64752 = w7152 & w7163;
assign w64753 = w7173 & ~w7176;
assign w64754 = ~w7199 & w7145;
assign w64755 = ~w6606 & w6557;
assign w64756 = w6573 & ~w6588;
assign w64757 = ~w7281 & pi0445;
assign w64758 = w7281 & ~pi0445;
assign w64759 = ~w6590 & w6588;
assign w64760 = w7057 & w6993;
assign w64761 = ~w7311 & w7028;
assign w64762 = ~w6993 & ~w6983;
assign w64763 = ~w7355 & ~w7369;
assign w64764 = w7430 & pi0431;
assign w64765 = ~w7430 & ~pi0431;
assign w64766 = ~w6893 & ~w6886;
assign w64767 = ~w7438 & ~pi0426;
assign w64768 = w7438 & pi0426;
assign w64769 = ~w7479 & w7507;
assign w64770 = w7508 & w7466;
assign w64771 = w7518 & w7520;
assign w64772 = w7530 & ~w7503;
assign w64773 = w6994 & w7028;
assign w64774 = ~w6982 & ~w7007;
assign w64775 = w6994 & ~w7305;
assign w64776 = w7353 & w7333;
assign w64777 = w7648 & w7333;
assign w64778 = w7649 & ~w7346;
assign w64779 = ~w7673 & w6588;
assign w64780 = w6565 & w6550;
assign w64781 = w7678 & ~w6588;
assign w64782 = w7486 & ~w7694;
assign w64783 = ~w7503 & ~w7524;
assign w64784 = w7495 & ~w7503;
assign w64785 = ~w6919 & ~w7101;
assign w64786 = w6795 & w6783;
assign w64787 = ~w7878 & w7836;
assign w64788 = w7856 & w7904;
assign w64789 = ~w7918 & ~w7955;
assign w64790 = ~w7981 & ~w7945;
assign w64791 = w7985 & w7945;
assign w64792 = ~w8034 & ~w8033;
assign w64793 = ~w8036 & w7999;
assign w64794 = ~w8117 & w8110;
assign w64795 = w8103 & w8110;
assign w64796 = w8153 & ~w8129;
assign w64797 = ~w63596 & ~w8040;
assign w64798 = w8185 & ~w8077;
assign w64799 = w8031 & w7999;
assign w64800 = w8193 & ~w8055;
assign w64801 = w8183 & ~pi0490;
assign w64802 = ~w8183 & pi0490;
assign w64803 = w8258 & ~w8212;
assign w64804 = ~w7951 & w7918;
assign w64805 = w8301 & ~w7945;
assign w64806 = ~w8311 & w7945;
assign w64807 = ~w8363 & ~w8336;
assign w64808 = ~w8103 & ~w8117;
assign w64809 = ~w8117 & w8090;
assign w64810 = ~w8141 & ~w8140;
assign w64811 = w8430 & w8429;
assign w64812 = ~w8386 & ~w8348;
assign w64813 = ~w8457 & ~pi0492;
assign w64814 = w8457 & pi0492;
assign w64815 = ~w8416 & w8140;
assign w64816 = w8117 & ~w8103;
assign w64817 = w8026 & ~w8012;
assign w64818 = w8517 & w8055;
assign w64819 = ~w8190 & ~w8055;
assign w64820 = w8564 & ~w8309;
assign w64821 = w8565 & ~w7945;
assign w64822 = w7904 & w7870;
assign w64823 = ~w8677 & w8675;
assign w64824 = w8678 & w8685;
assign w64825 = ~w8678 & ~w8621;
assign w64826 = w8700 & w8704;
assign w64827 = w8706 & pi0501;
assign w64828 = ~w8706 & ~pi0501;
assign w64829 = w8723 & ~w8735;
assign w64830 = w8806 & ~w8808;
assign w64831 = w8759 & w8820;
assign w64832 = w8810 & ~w8795;
assign w64833 = w8830 & w8831;
assign w64834 = w8826 & pi0484;
assign w64835 = ~w8826 & ~pi0484;
assign w64836 = ~w8313 & ~w8572;
assign w64837 = w8858 & w7918;
assign w64838 = w8562 & ~w7945;
assign w64839 = w8869 & w7945;
assign w64840 = w8416 & w8423;
assign w64841 = w8910 & ~w7878;
assign w64842 = w7829 & w7844;
assign w64843 = ~w8189 & w8024;
assign w64844 = w8055 & ~w8523;
assign w64845 = w8930 & ~w8055;
assign w64846 = ~w8964 & w8661;
assign w64847 = w8971 & ~w8372;
assign w64848 = w8391 & w8336;
assign w64849 = ~w8363 & ~w8348;
assign w64850 = w8984 & w8372;
assign w64851 = ~w9021 & w8795;
assign w64852 = w8765 & ~w9025;
assign w64853 = ~w9030 & ~w8795;
assign w64854 = ~w9022 & ~pi0488;
assign w64855 = w9022 & pi0488;
assign w64856 = ~w8231 & w9109;
assign w64857 = ~w8231 & ~w63606;
assign w64858 = ~w9119 & ~w9115;
assign w64859 = ~w9120 & ~w8212;
assign w64860 = w9149 & w9180;
assign w64861 = ~w9585 & ~w9186;
assign w64862 = ~w9141 & w9155;
assign w64863 = ~w9220 & pi0553;
assign w64864 = w9220 & ~pi0553;
assign w64865 = w9256 & w9262;
assign w64866 = w9276 & ~w9269;
assign w64867 = w9269 & ~w9250;
assign w64868 = ~w9299 & ~pi0551;
assign w64869 = w9299 & pi0551;
assign w64870 = ~w9348 & w9355;
assign w64871 = ~w9383 & w9384;
assign w64872 = ~w9383 & ~w63612;
assign w64873 = w9531 & w9382;
assign w64874 = (w9382 & w9531) | (w9382 & w9407) | (w9531 & w9407);
assign w64875 = w9405 & pi0549;
assign w64876 = ~w9405 & ~pi0549;
assign w64877 = w9447 & w9457;
assign w64878 = w9457 & ~w9475;
assign w64879 = w9485 & w9457;
assign w64880 = ~w9464 & w9457;
assign w64881 = ~w9348 & ~w9335;
assign w64882 = w9520 & ~w9382;
assign w64883 = w9394 & w9335;
assign w64884 = w9527 & w9382;
assign w64885 = ~w9283 & ~w9262;
assign w64886 = w9561 & ~w9543;
assign w64887 = ~w9204 & w9180;
assign w64888 = ~w9585 & w9600;
assign w64889 = w9655 & ~w9647;
assign w64890 = w9727 & ~w9734;
assign w64891 = ~w9749 & ~w9748;
assign w64892 = ~w9752 & ~w9740;
assign w64893 = w9792 & ~w9788;
assign w64894 = w9791 & w9382;
assign w64895 = ~w9813 & ~w9702;
assign w64896 = ~w9720 & ~w9708;
assign w64897 = ~w9773 & ~w9807;
assign w64898 = ~w9856 & ~w9863;
assign w64899 = ~w9871 & ~w9904;
assign w64900 = w9882 & w9863;
assign w64901 = ~w9939 & w9926;
assign w64902 = w9995 & w9964;
assign w64903 = ~w9997 & ~w9989;
assign w64904 = ~w9977 & ~pi0548;
assign w64905 = w9977 & pi0548;
assign w64906 = w10020 & w9639;
assign w64907 = ~w10039 & pi0554;
assign w64908 = w10039 & ~pi0554;
assign w64909 = w9527 & w10092;
assign w64910 = ~w9364 & w9342;
assign w64911 = w9373 & w9335;
assign w64912 = ~w9364 & ~w9382;
assign w64913 = w9292 & w10112;
assign w64914 = ~w9276 & w9250;
assign w64915 = w10122 & w9292;
assign w64916 = ~w9878 & ~w9863;
assign w64917 = ~w10146 & ~w10141;
assign w64918 = ~w10147 & ~w9870;
assign w64919 = w9870 & ~w10169;
assign w64920 = ~w10191 & w9702;
assign w64921 = ~w10075 & ~w9776;
assign w64922 = ~w9939 & ~w9957;
assign w64923 = w9932 & w9926;
assign w64924 = ~w9992 & w10231;
assign w64925 = ~w10228 & w9926;
assign w64926 = ~w10252 & pi0546;
assign w64927 = w10252 & ~pi0546;
assign w64928 = ~w9850 & w9870;
assign w64929 = w9458 & w9440;
assign w64930 = w9498 & w9457;
assign w64931 = w9485 & w9428;
assign w64932 = w10371 & ~w9428;
assign w64933 = ~w10389 & ~w9964;
assign w64934 = ~w10226 & w9964;
assign w64935 = ~w10410 & ~w9964;
assign w64936 = ~w10410 & ~w63624;
assign w64937 = w10418 & ~pi0567;
assign w64938 = ~w10418 & pi0567;
assign w64939 = w10453 & w10427;
assign w64940 = w10578 & ~w10522;
assign w64941 = ~w10591 & w10595;
assign w64942 = ~w10606 & w10522;
assign w64943 = ~w10644 & ~w10638;
assign w64944 = ~w10662 & w10677;
assign w64945 = ~w10632 & w10670;
assign w64946 = ~w10606 & w10704;
assign w64947 = ~w10563 & ~w10547;
assign w64948 = w10729 & w10522;
assign w64949 = ~w10732 & ~pi0629;
assign w64950 = w10732 & pi0629;
assign w64951 = w10753 & w10768;
assign w64952 = w10759 & ~w10776;
assign w64953 = w10779 & w10776;
assign w64954 = w10830 & pi0621;
assign w64955 = ~w10830 & ~pi0621;
assign w64956 = w10846 & ~w10840;
assign w64957 = ~w10840 & w10881;
assign w64958 = w10810 & ~w10752;
assign w64959 = ~w10746 & ~w10752;
assign w64960 = w10961 & w10955;
assign w64961 = ~w10968 & w11010;
assign w64962 = w10840 & w10846;
assign w64963 = ~w10859 & w10853;
assign w64964 = w11072 & ~w11075;
assign w64965 = ~w10439 & ~w10433;
assign w64966 = w11107 & w10493;
assign w64967 = w63636 | ~w10493;
assign w64968 = (~w10493 & w63636) | (~w10493 & w11129) | (w63636 & w11129);
assign w64969 = w11143 & ~w10522;
assign w64970 = w11145 & w10522;
assign w64971 = ~w11148 & ~pi0623;
assign w64972 = w11148 & pi0623;
assign w64973 = ~w10968 & ~w10955;
assign w64974 = ~w11161 & w10968;
assign w64975 = ~w11233 & ~w11239;
assign w64976 = w11259 & ~w11249;
assign w64977 = ~w11290 & ~w11286;
assign w64978 = w11226 & w11239;
assign w64979 = ~w11307 & ~w11272;
assign w64980 = w11321 & ~w11248;
assign w64981 = w11373 & w11397;
assign w64982 = w11410 & w11415;
assign w64983 = w11440 & ~w11397;
assign w64984 = w11452 & pi0630;
assign w64985 = ~w11452 & ~pi0630;
assign w64986 = ~w11064 & ~w10861;
assign w64987 = ~w10875 & ~w11046;
assign w64988 = ~w11478 & w10867;
assign w64989 = w10776 & w10759;
assign w64990 = w11503 & ~w10788;
assign w64991 = w11527 & ~w11519;
assign w64992 = ~w10937 & ~w10752;
assign w64993 = w11542 & w10788;
assign w64994 = ~w10629 & ~w10683;
assign w64995 = w11559 & w11083;
assign w64996 = ~w11372 & ~w11420;
assign w64997 = ~w11622 & ~w11620;
assign w64998 = w11638 & w11009;
assign w64999 = ~w11239 & ~w11246;
assign w65000 = w11667 & ~w11666;
assign w65001 = ~w11672 & ~w11673;
assign w65002 = w11698 & ~w10638;
assign w65003 = w11709 & ~w11689;
assign w65004 = w11769 & w11740;
assign w65005 = ~w11746 & w11758;
assign w65006 = ~w11746 & ~w11758;
assign w65007 = w11746 & ~w11758;
assign w65008 = ~w11758 & w11768;
assign w65009 = w11825 & ~w11787;
assign w65010 = w11837 & w11857;
assign w65011 = ~w11863 & w11857;
assign w65012 = w11862 & w11875;
assign w65013 = w11906 & w11881;
assign w65014 = w11949 & ~w11940;
assign w65015 = w11932 & w11962;
assign w65016 = ~w11962 & ~w11991;
assign w65017 = ~w12032 & ~w12025;
assign w65018 = w12066 & ~w12059;
assign w65019 = w12026 & w12032;
assign w65020 = ~w12039 & ~w12059;
assign w65021 = w12125 & ~w11881;
assign w65022 = w12118 & w11881;
assign w65023 = w12126 & pi0682;
assign w65024 = ~w12126 & ~pi0682;
assign w65025 = w11984 & ~w12151;
assign w65026 = ~w12157 & w11980;
assign w65027 = ~w12244 & ~w12175;
assign w65028 = ~w12245 & pi0675;
assign w65029 = w12245 & ~pi0675;
assign w65030 = w12299 & ~w12234;
assign w65031 = w12181 & w12193;
assign w65032 = ~w12344 & ~w12325;
assign w65033 = w12344 & ~w12325;
assign w65034 = w12381 & ~w12370;
assign w65035 = w12408 & ~w12412;
assign w65036 = ~w12482 & ~w12489;
assign w65037 = ~w12514 & w12515;
assign w65038 = ~w12498 & ~w12470;
assign w65039 = w12083 & ~w12066;
assign w65040 = ~w11746 & ~w11768;
assign w65041 = w12569 & ~w11787;
assign w65042 = ~w12581 & w11787;
assign w65043 = ~w12576 & ~w11787;
assign w65044 = ~w12576 & ~w63653;
assign w65045 = ~w12389 & ~w12352;
assign w65046 = w12257 & w12222;
assign w65047 = w12674 & ~w12175;
assign w65048 = ~w12568 & ~w11787;
assign w65049 = ~w12715 & pi0693;
assign w65050 = w12715 & ~pi0693;
assign w65051 = w12492 & ~w12498;
assign w65052 = ~w12723 & ~w12728;
assign w65053 = w12731 & w12498;
assign w65054 = w12806 & ~w12059;
assign w65055 = ~w12059 & w12083;
assign w65056 = w12038 & w12032;
assign w65057 = ~w12072 & ~w12083;
assign w65058 = ~w12837 & w12859;
assign w65059 = w12851 & ~w12836;
assign w65060 = w12919 & w12889;
assign w65061 = ~w12929 & ~w12904;
assign w65062 = w12934 & ~w12878;
assign w65063 = ~w12935 & pi0702;
assign w65064 = w12935 & ~pi0702;
assign w65065 = ~w12490 & ~w12498;
assign w65066 = w12751 & w12476;
assign w65067 = w12731 & w12991;
assign w65068 = w13014 & pi0687;
assign w65069 = ~w13014 & ~pi0687;
assign w65070 = w13022 & ~w12858;
assign w65071 = w12895 & ~w12836;
assign w65072 = w13049 & ~pi0707;
assign w65073 = ~w13049 & pi0707;
assign w65074 = w13067 & ~w13076;
assign w65075 = ~w13076 & w13091;
assign w65076 = w13099 & ~w13104;
assign w65077 = ~w13083 & w13091;
assign w65078 = w13061 & ~w13076;
assign w65079 = ~w13200 & w13152;
assign w65080 = ~w13184 & w13193;
assign w65081 = w13152 & ~w13181;
assign w65082 = w13202 & ~w13183;
assign w65083 = w13200 & ~w13178;
assign w65084 = ~w13182 & w13199;
assign w65085 = ~w13182 & ~w63661;
assign w65086 = w13185 & w13152;
assign w65087 = w13185 & w63662;
assign w65088 = ~w13258 & w13259;
assign w65089 = w13260 & w13261;
assign w65090 = ~w13349 & ~pi0740;
assign w65091 = w13349 & pi0740;
assign w65092 = ~w13414 & ~w13435;
assign w65093 = ~w13414 & ~w63665;
assign w65094 = ~w13447 & pi0742;
assign w65095 = w13447 & ~pi0742;
assign w65096 = w13519 & w13193;
assign w65097 = ~w13603 & ~w13608;
assign w65098 = ~w13547 & ~w13571;
assign w65099 = w13614 & ~w13600;
assign w65100 = ~w13594 & ~pi0756;
assign w65101 = w13594 & pi0756;
assign w65102 = ~w13688 & w13690;
assign w65103 = ~w13692 & ~w13691;
assign w65104 = w13671 & w13674;
assign w65105 = w13671 & w13694;
assign w65106 = ~w13561 & ~w13714;
assign w65107 = w13713 & w13600;
assign w65108 = ~w13729 & ~w13600;
assign w65109 = w13769 & ~w13755;
assign w65110 = ~w13748 & ~w13798;
assign w65111 = w13939 & w13647;
assign w65112 = w13671 & ~w13970;
assign w65113 = ~w13967 & pi0743;
assign w65114 = w13967 & ~pi0743;
assign w65115 = w13211 & w13152;
assign w65116 = w13997 & ~pi0741;
assign w65117 = ~w13997 & pi0741;
assign w65118 = ~w13284 & w13271;
assign w65119 = w14005 & w14009;
assign w65120 = w14011 & ~pi0765;
assign w65121 = ~w14011 & pi0765;
assign w65122 = w13645 & w13653;
assign w65123 = w13687 & w13939;
assign w65124 = w14034 & ~w13671;
assign w65125 = w13126 & w13091;
assign w65126 = ~w13102 & w13111;
assign w65127 = ~w13076 & ~w13083;
assign w65128 = ~w13380 & ~w13364;
assign w65129 = w13402 & ~w13358;
assign w65130 = w14094 & pi0755;
assign w65131 = ~w14094 & ~pi0755;
assign w65132 = ~w13583 & ~w13600;
assign w65133 = ~w14157 & ~w14147;
assign w65134 = w14159 & pi0754;
assign w65135 = ~w14159 & ~pi0754;
assign w65136 = w13866 & ~w13859;
assign w65137 = w14232 & ~w14233;
assign w65138 = ~w14236 & ~w14223;
assign w65139 = w14272 & w14053;
assign w65140 = w14272 & ~w63682;
assign w65141 = ~w14279 & ~w13671;
assign w65142 = w13688 & w14281;
assign w65143 = ~w14302 & ~pi0770;
assign w65144 = w14302 & pi0770;
assign w65145 = w14228 & w13905;
assign w65146 = w14327 & ~w13905;
assign w65147 = w14243 & w13859;
assign w65148 = w14347 & w14352;
assign w65149 = w14364 & w14379;
assign w65150 = w14390 & w14406;
assign w65151 = w14611 & w14610;
assign w65152 = w14539 & w14608;
assign w65153 = w14618 & ~pi0811;
assign w65154 = ~w14618 & pi0811;
assign w65155 = ~w14667 & ~w14459;
assign w65156 = ~w14673 & w14459;
assign w65157 = ~w14707 & ~w14714;
assign w65158 = w14763 & ~pi0805;
assign w65159 = ~w14763 & pi0805;
assign w65160 = ~w14778 & ~w14798;
assign w65161 = ~w14798 & w14772;
assign w65162 = w14827 & w14809;
assign w65163 = w14791 & ~w14798;
assign w65164 = w14879 & ~w14886;
assign w65165 = ~w14902 & w14879;
assign w65166 = w14935 & w14867;
assign w65167 = w14957 & ~w14867;
assign w65168 = w14993 & ~w15022;
assign w65169 = ~w14993 & w15022;
assign w65170 = w14791 & w15072;
assign w65171 = ~w14459 & ~w15113;
assign w65172 = w15142 & ~pi0830;
assign w65173 = ~w15142 & pi0830;
assign w65174 = ~w15012 & ~w14993;
assign w65175 = ~w15022 & ~w15039;
assign w65176 = w15232 & w15237;
assign w65177 = w15247 & w15250;
assign w65178 = ~w15243 & ~w14867;
assign w65179 = w15291 & ~w15295;
assign w65180 = ~w15297 & ~w15308;
assign w65181 = w14398 & w15356;
assign w65182 = ~w15390 & w15391;
assign w65183 = ~w14429 & ~w14406;
assign w65184 = w15435 & w15436;
assign w65185 = w14839 & w14772;
assign w65186 = w14747 & ~w14726;
assign w65187 = w15495 & ~w14686;
assign w65188 = w15514 & w14686;
assign w65189 = w15564 & ~w15530;
assign w65190 = w15572 & w15581;
assign w65191 = w15563 & ~w15605;
assign w65192 = w15621 & ~w15551;
assign w65193 = w15635 & w15549;
assign w65194 = w15536 & w15581;
assign w65195 = w15660 & ~w15581;
assign w65196 = w15669 & pi0832;
assign w65197 = ~w15669 & ~pi0832;
assign w65198 = w15728 & ~w15729;
assign w65199 = w15800 & w15836;
assign w65200 = w15840 & ~w15817;
assign w65201 = ~w15890 & ~w15914;
assign w65202 = ~w15884 & ~w15890;
assign w65203 = ~w15914 & ~w15902;
assign w65204 = w15942 & pi0869;
assign w65205 = ~w15942 & ~pi0869;
assign w65206 = w16032 & ~w15975;
assign w65207 = w16032 & w63706;
assign w65208 = ~w16029 & w16037;
assign w65209 = w16038 & pi0867;
assign w65210 = ~w16038 & ~pi0867;
assign w65211 = w16079 & w15737;
assign w65212 = ~w15728 & ~w15696;
assign w65213 = ~w16152 & ~pi0864;
assign w65214 = w16152 & pi0864;
assign w65215 = w16194 & w15865;
assign w65216 = w16199 & w15902;
assign w65217 = w16209 & ~w15902;
assign w65218 = ~w15871 & w15902;
assign w65219 = w16211 & ~w15865;
assign w65220 = w16234 & w16244;
assign w65221 = ~w16019 & w15991;
assign w65222 = w16302 & ~w16295;
assign w65223 = w16307 & ~w16305;
assign w65224 = ~w16337 & ~pi0868;
assign w65225 = w16337 & pi0868;
assign w65226 = w15719 & w15696;
assign w65227 = w16437 & ~w15865;
assign w65228 = ~w16437 & ~w16201;
assign w65229 = ~w16222 & ~w16450;
assign w65230 = w16495 & ~w16480;
assign w65231 = ~w16518 & ~w16471;
assign w65232 = w16521 & w16509;
assign w65233 = ~w16532 & w16493;
assign w65234 = ~w16532 & w16494;
assign w65235 = w16471 & ~w16493;
assign w65236 = w16549 & ~pi0875;
assign w65237 = ~w16549 & pi0875;
assign w65238 = ~w16471 & w16493;
assign w65239 = w16580 & ~w16585;
assign w65240 = ~w16589 & w16509;
assign w65241 = ~w16619 & pi0882;
assign w65242 = w16619 & ~pi0882;
assign w65243 = ~w16629 & w16509;
assign w65244 = ~w16544 & ~w16537;
assign w65245 = w16509 & ~w16502;
assign w65246 = ~w15690 & ~w16689;
assign w65247 = w16715 & w16741;
assign w65248 = w16725 & w16750;
assign w65249 = ~w16725 & ~w16750;
assign w65250 = w15785 & w15793;
assign w65251 = ~w15785 & ~w15818;
assign w65252 = ~w16797 & pi0877;
assign w65253 = w16797 & ~pi0877;
assign w65254 = ~w16809 & ~w16702;
assign w65255 = ~w16809 & w63711;
assign w65256 = ~w16748 & ~w16751;
assign w65257 = ~w16741 & ~w63713;
assign w65258 = ~w16741 & w16818;
assign w65259 = ~w16830 & pi0887;
assign w65260 = w16830 & ~pi0887;
assign w65261 = ~w16846 & ~w16146;
assign w65262 = ~w16660 & ~w16326;
assign w65263 = w16288 & w16275;
assign w65264 = w16877 & ~w16346;
assign w65265 = w16868 & w16648;
assign w65266 = ~w63381 & w16731;
assign w65267 = w16931 & w16937;
assign w65268 = w63716 & ~w16716;
assign w65269 = w16741 & w16832;
assign w65270 = w16741 & ~w63717;
assign w65271 = w16981 & w16984;
assign w65272 = w16985 & ~w16971;
assign w65273 = w17025 & w17012;
assign w65274 = ~w17025 & ~w17006;
assign w65275 = ~w17033 & w17053;
assign w65276 = w17078 & pi0928;
assign w65277 = ~w17078 & ~pi0928;
assign w65278 = ~w17101 & w17127;
assign w65279 = w17128 & ~w17130;
assign w65280 = w17146 & ~w17127;
assign w65281 = w17164 & ~w17159;
assign w65282 = ~w17180 & pi0947;
assign w65283 = w17180 & ~pi0947;
assign w65284 = w17152 & w17186;
assign w65285 = w17127 & w17089;
assign w65286 = w17101 & w17108;
assign w65287 = w17194 & w17201;
assign w65288 = w17202 & w17203;
assign w65289 = w17237 & w17252;
assign w65290 = ~w17213 & w17226;
assign w65291 = ~w17277 & ~w17274;
assign w65292 = w17309 & w17327;
assign w65293 = w17368 & w17373;
assign w65294 = w17381 & ~w17128;
assign w65295 = w17392 & ~w17379;
assign w65296 = w17436 & ~w17421;
assign w65297 = w17421 & w17436;
assign w65298 = w17449 & w17456;
assign w65299 = ~w17466 & w17429;
assign w65300 = w17470 & ~w17468;
assign w65301 = ~w17533 & w17520;
assign w65302 = ~w17553 & ~w17495;
assign w65303 = ~w17523 & ~w17508;
assign w65304 = w17572 & w17495;
assign w65305 = ~w17514 & w17501;
assign w65306 = w17213 & ~w17251;
assign w65307 = w17657 & ~w17621;
assign w65308 = w17733 & ~w17703;
assign w65309 = ~w17143 & ~w17738;
assign w65310 = w17742 & pi0938;
assign w65311 = ~w17742 & ~pi0938;
assign w65312 = w17621 & w17627;
assign w65313 = w17767 & w17614;
assign w65314 = w17634 & w17628;
assign w65315 = w17780 & w17668;
assign w65316 = w17806 & ~w17653;
assign w65317 = ~w17822 & ~w17829;
assign w65318 = ~w17370 & w17866;
assign w65319 = ~w17436 & w17446;
assign w65320 = w17450 & ~w17895;
assign w65321 = w17893 & w17429;
assign w65322 = ~w17784 & w17660;
assign w65323 = ~w17621 & ~w17654;
assign w65324 = w17803 & ~w17917;
assign w65325 = w17922 & pi0948;
assign w65326 = ~w17922 & ~pi0948;
assign w65327 = ~w17957 & w17962;
assign w65328 = w17953 & ~w17941;
assign w65329 = ~w17938 & ~w17068;
assign w65330 = w17252 & ~w18004;
assign w65331 = w18031 & ~w18076;
assign w65332 = w18099 & w18031;
assign w65333 = w18096 & pi0966;
assign w65334 = ~w18096 & ~pi0966;
assign w65335 = w18140 & ~w17577;
assign w65336 = ~w18173 & ~w18058;
assign w65337 = ~w18208 & w18058;
assign w65338 = w18205 & ~w18058;
assign w65339 = w18133 & w17850;
assign w65340 = w17236 & ~w17251;
assign w65341 = w18284 & ~w18291;
assign w65342 = w18292 & w17251;
assign w65343 = w18322 & ~w18329;
assign w65344 = ~w18448 & ~pi1061;
assign w65345 = w18448 & pi1061;
assign w65346 = ~w18511 & w18517;
assign w65347 = w18490 & w18505;
assign w65348 = ~w18505 & ~w18517;
assign w65349 = w18584 & pi1071;
assign w65350 = ~w18584 & ~pi1071;
assign w65351 = w18599 & ~w18606;
assign w65352 = ~w18641 & ~w18636;
assign w65353 = w18633 & w18655;
assign w65354 = ~w18738 & w18768;
assign w65355 = ~w18808 & ~w18777;
assign w65356 = w18816 & pi1062;
assign w65357 = ~w18816 & ~pi1062;
assign w65358 = ~w18847 & w18885;
assign w65359 = ~w18906 & w18439;
assign w65360 = w18468 & ~w18919;
assign w65361 = w18917 & pi1072;
assign w65362 = ~w18917 & ~pi1072;
assign w65363 = w18631 & w18634;
assign w65364 = w18965 & ~w18825;
assign w65365 = w18620 & ~w19012;
assign w65366 = w18751 & ~w18768;
assign w65367 = w18807 & ~w19033;
assign w65368 = w18807 & ~w19037;
assign w65369 = w18732 & w18786;
assign w65370 = ~w19035 & ~w19024;
assign w65371 = ~w19048 & pi1077;
assign w65372 = w19048 & ~pi1077;
assign w65373 = w18860 & ~w18857;
assign w65374 = ~w18808 & ~w18804;
assign w65375 = ~w18533 & w18552;
assign w65376 = w19130 & w19143;
assign w65377 = w19165 & w19153;
assign w65378 = w19130 & w19193;
assign w65379 = w19266 & w19262;
assign w65380 = w19264 & w19289;
assign w65381 = ~w18464 & w18426;
assign w65382 = w18906 & w19305;
assign w65383 = w19176 & ~w19325;
assign w65384 = w19165 & w19150;
assign w65385 = ~w19143 & w19164;
assign w65386 = w19185 & w19143;
assign w65387 = w19352 & ~w19176;
assign w65388 = ~w19358 & ~w19360;
assign w65389 = ~w19371 & w19376;
assign w65390 = w19217 & w19262;
assign w65391 = ~w18309 & w18329;
assign w65392 = w18347 & w18316;
assign w65393 = w18346 & ~w18365;
assign w65394 = ~w19493 & ~w18346;
assign w65395 = ~w19224 & ~w19238;
assign w65396 = w19584 & w19262;
assign w65397 = w19238 & ~w19239;
assign w65398 = ~w19595 & ~w19262;
assign w65399 = w19610 & ~w19238;
assign w65400 = ~w19612 & ~w19609;
assign w65401 = ~w19615 & pi1068;
assign w65402 = w19615 & ~pi1068;
assign w65403 = ~w19647 & w19654;
assign w65404 = ~w19754 & w19789;
assign w65405 = ~w19766 & ~pi0993;
assign w65406 = w19766 & pi0993;
assign w65407 = ~w19948 & ~w19955;
assign w65408 = w19939 & ~w20003;
assign w65409 = ~w20006 & pi1027;
assign w65410 = w20006 & ~pi1027;
assign w65411 = ~w19939 & w20016;
assign w65412 = w19962 & ~w63736;
assign w65413 = w19962 & w20018;
assign w65414 = ~w20032 & ~w19962;
assign w65415 = w20052 & ~w20051;
assign w65416 = w19684 & w19641;
assign w65417 = w20154 & w19673;
assign w65418 = ~w20222 & w20202;
assign w65419 = w19681 & w19673;
assign w65420 = w20302 & ~w20308;
assign w65421 = w20372 & ~w20221;
assign w65422 = ~w20374 & w20387;
assign w65423 = w20383 & w20221;
assign w65424 = ~w20379 & ~w20373;
assign w65425 = w20289 & ~w20326;
assign w65426 = ~w20465 & w20466;
assign w65427 = w20413 & w20188;
assign w65428 = w20244 & ~w20188;
assign w65429 = w19778 & w19789;
assign w65430 = w20562 & ~w20554;
assign w65431 = ~w20585 & ~w20566;
assign w65432 = ~w20544 & w20531;
assign w65433 = w20663 & ~w20552;
assign w65434 = ~w20684 & w20685;
assign w65435 = ~w20667 & ~pi1019;
assign w65436 = w20667 & pi1019;
assign w65437 = w20347 & ~w20308;
assign w65438 = ~w20701 & ~w20699;
assign w65439 = w20718 & ~w19742;
assign w65440 = w19727 & ~w19790;
assign w65441 = w20721 & w19789;
assign w65442 = w20728 & ~w19792;
assign w65443 = ~w19726 & ~w19742;
assign w65444 = w20773 & w20781;
assign w65445 = w20805 & w20809;
assign w65446 = ~w20805 & w20783;
assign w65447 = w20799 & w20809;
assign w65448 = w20870 & w20804;
assign w65449 = w20891 & pi1036;
assign w65450 = ~w20891 & ~pi1036;
assign w65451 = ~w20791 & ~w20780;
assign w65452 = ~w21146 & ~w21152;
assign w65453 = w21139 & w21152;
assign w65454 = ~w21146 & w21127;
assign w65455 = w21001 & ~w20962;
assign w65456 = ~w21250 & ~pi1227;
assign w65457 = w21250 & pi1227;
assign w65458 = ~w21288 & ~w21281;
assign w65459 = w21318 & ~w21313;
assign w65460 = w21164 & ~w21127;
assign w65461 = ~w21164 & w21166;
assign w65462 = ~w21418 & ~w21192;
assign w65463 = w21424 & ~pi1232;
assign w65464 = ~w21424 & pi1232;
assign w65465 = w21471 & ~w21504;
assign w65466 = w21791 & w21777;
assign w65467 = w21911 & ~w21783;
assign w65468 = ~w21916 & ~w21803;
assign w65469 = ~w22042 & w21462;
assign w65470 = ~w22043 & ~w21520;
assign w65471 = w22081 & ~w21977;
assign w65472 = w22237 & w22244;
assign w65473 = ~w22235 & w22216;
assign w65474 = ~w22254 & w22255;
assign w65475 = w22216 & w22233;
assign w65476 = w22310 & ~w22305;
assign w65477 = w22308 & w22324;
assign w65478 = w22397 & w22398;
assign w65479 = w22417 & w22233;
assign w65480 = ~w22448 & w22455;
assign w65481 = ~w22567 & w22539;
assign w65482 = w22656 & ~w22662;
assign w65483 = w22681 & ~w22676;
assign w65484 = ~w22746 & w22731;
assign w65485 = w22267 & ~w22808;
assign w65486 = w22828 & w22492;
assign w65487 = ~w22833 & ~w22492;
assign w65488 = w22835 & pi1252;
assign w65489 = ~w22835 & ~pi1252;
assign w65490 = w22989 & ~w22963;
assign w65491 = ~w22311 & w22331;
assign w65492 = w22996 & ~w22324;
assign w65493 = ~w22282 & w22324;
assign w65494 = ~w22331 & w23015;
assign w65495 = ~w23081 & ~w23027;
assign w65496 = ~w23090 & w23088;
assign w65497 = ~w23090 & ~w63762;
assign w65498 = ~w22641 & ~w22635;
assign w65499 = w22676 & ~w22641;
assign w65500 = w22676 & ~w63760;
assign w65501 = ~w22852 & w22662;
assign w65502 = w23121 & ~w23106;
assign w65503 = ~w23073 & w23050;
assign w65504 = ~w23138 & w23151;
assign w65505 = w23153 & w23155;
assign w65506 = w22975 & ~w22919;
assign w65507 = w23186 & ~w22958;
assign w65508 = w23193 & ~w23168;
assign w65509 = ~w23141 & ~w23279;
assign w65510 = w23285 & pi1274;
assign w65511 = ~w23285 & ~pi1274;
assign w65512 = w22356 & ~w22331;
assign w65513 = w23316 & w22324;
assign w65514 = w22887 & w23340;
assign w65515 = ~w22749 & ~w23349;
assign w65516 = w22475 & ~w23364;
assign w65517 = w23365 & w22492;
assign w65518 = w22482 & w23376;
assign w65519 = w22857 & ~w22662;
assign w65520 = w22634 & w22662;
assign w65521 = ~w23408 & ~w22676;
assign w65522 = w22964 & ~w22958;
assign w65523 = ~w22938 & ~w22931;
assign w65524 = ~w22958 & ~w23442;
assign w65525 = w23468 & w23475;
assign w65526 = w22513 & ~w23483;
assign w65527 = ~w23566 & w23557;
assign w65528 = w23568 & ~w23530;
assign w65529 = ~w23563 & ~w23542;
assign w65530 = w23603 & w23536;
assign w65531 = w23549 & w23569;
assign w65532 = w23734 & ~w23735;
assign w65533 = w23737 & w23679;
assign w65534 = w23743 & ~w23679;
assign w65535 = ~w23774 & w23767;
assign w65536 = w23794 & ~w23782;
assign w65537 = w23812 & w23755;
assign w65538 = w23873 & ~w23879;
assign w65539 = ~w23961 & ~w23948;
assign w65540 = w23960 & ~w23947;
assign w65541 = ~w23992 & ~w24002;
assign w65542 = w24021 & pi1314;
assign w65543 = ~w24021 & ~pi1314;
assign w65544 = ~w23679 & ~w23735;
assign w65545 = w23699 & ~w24054;
assign w65546 = ~w24058 & ~pi1322;
assign w65547 = w24058 & pi1322;
assign w65548 = w24068 & w23706;
assign w65549 = ~w23699 & ~w23706;
assign w65550 = w23799 & w24093;
assign w65551 = ~w24165 & w24156;
assign w65552 = w24176 & ~w24125;
assign w65553 = w24186 & pi1313;
assign w65554 = ~w24186 & ~pi1313;
assign w65555 = w23827 & w23794;
assign w65556 = ~w23780 & ~w23794;
assign w65557 = w24204 & w23755;
assign w65558 = w23761 & w23819;
assign w65559 = w24157 & ~w24229;
assign w65560 = w23881 & w23879;
assign w65561 = ~w24278 & ~pi1337;
assign w65562 = w24278 & pi1337;
assign w65563 = w24103 & w23794;
assign w65564 = ~w23861 & w24250;
assign w65565 = ~w23861 & ~w23920;
assign w65566 = ~w24378 & w24407;
assign w65567 = w24408 & w24365;
assign w65568 = ~w24435 & ~w24394;
assign w65569 = ~w24371 & ~w24385;
assign w65570 = w24463 & ~w24365;
assign w65571 = ~w24469 & w24365;
assign w65572 = ~w24473 & pi1332;
assign w65573 = w24473 & ~pi1332;
assign w65574 = w24423 & w24411;
assign w65575 = ~w24498 & w24365;
assign w65576 = w24499 & ~pi1342;
assign w65577 = ~w24499 & pi1342;
assign w65578 = ~w24565 & ~w24559;
assign w65579 = w24574 & w24565;
assign w65580 = ~w24590 & ~w24578;
assign w65581 = ~w24601 & w24565;
assign w65582 = w24530 & w24536;
assign w65583 = w24597 & pi1328;
assign w65584 = ~w24597 & ~pi1328;
assign w65585 = w23907 & w24256;
assign w65586 = ~w24641 & pi1344;
assign w65587 = w24641 & ~pi1344;
assign w65588 = w24649 & ~w23997;
assign w65589 = ~w24650 & w23978;
assign w65590 = ~w24692 & pi1331;
assign w65591 = w24692 & ~pi1331;
assign w65592 = w24522 & ~w24510;
assign w65593 = ~w24699 & ~w24704;
assign w65594 = w24720 & pi1325;
assign w65595 = ~w24720 & ~pi1325;
assign w65596 = w24729 & ~w24001;
assign w65597 = w24729 & w63391;
assign w65598 = ~w23960 & w23947;
assign w65599 = w23992 & ~w24003;
assign w65600 = ~w24743 & ~pi1349;
assign w65601 = w24743 & pi1349;
assign w65602 = w24776 & ~w24119;
assign w65603 = w24794 & pi1324;
assign w65604 = ~w24794 & ~pi1324;
assign w65605 = w24812 & ~w24813;
assign w65606 = w24880 & w24849;
assign w65607 = w24895 & w24849;
assign w65608 = ~w24974 & w24973;
assign w65609 = w25056 & ~w25042;
assign w65610 = w25076 & w25036;
assign w65611 = ~w25105 & w25085;
assign w65612 = ~w25093 & ~w25094;
assign w65613 = ~w25156 & w25130;
assign w65614 = ~w25156 & w25143;
assign w65615 = w25212 & w25211;
assign w65616 = w25184 & pi1376;
assign w65617 = ~w25184 & ~pi1376;
assign w65618 = w25234 & w25254;
assign w65619 = ~w25287 & ~w25272;
assign w65620 = w25366 & ~w25342;
assign w65621 = ~w25360 & ~w25318;
assign w65622 = w25360 & ~w25378;
assign w65623 = w25333 & w25360;
assign w65624 = ~w25400 & w25401;
assign w65625 = w25227 & ~w25258;
assign w65626 = ~w25156 & w25149;
assign w65627 = w25480 & ~w24869;
assign w65628 = w24841 & w24849;
assign w65629 = w24828 & ~w24890;
assign w65630 = w24878 & ~w25506;
assign w65631 = ~w24841 & w24867;
assign w65632 = w25556 & ~w25543;
assign w65633 = ~w25585 & w25562;
assign w65634 = w25536 & w25568;
assign w65635 = ~w25610 & pi1394;
assign w65636 = w25610 & ~pi1394;
assign w65637 = ~w25334 & ~w25360;
assign w65638 = w24899 & w24867;
assign w65639 = ~w24939 & ~w24958;
assign w65640 = w25661 & w25660;
assign w65641 = ~w25692 & ~w25562;
assign w65642 = ~w25693 & ~w25584;
assign w65643 = w25710 & ~w25687;
assign w65644 = w25717 & ~w25164;
assign w65645 = ~w25166 & w25149;
assign w65646 = ~w25287 & w25744;
assign w65647 = ~w25409 & ~w25263;
assign w65648 = w25741 & w25283;
assign w65649 = w25793 & ~w24958;
assign w65650 = w25810 & ~w25791;
assign w65651 = w25841 & ~w25855;
assign w65652 = w25891 & ~w25820;
assign w65653 = w25892 & pi1398;
assign w65654 = ~w25892 & ~pi1398;
assign w65655 = ~w25196 & ~w25728;
assign w65656 = w25912 & w25164;
assign w65657 = w25931 & w25360;
assign w65658 = w25373 & ~w25950;
assign w65659 = w25951 & ~pi1391;
assign w65660 = ~w25951 & pi1391;
assign w65661 = w25962 & ~w25049;
assign w65662 = ~w25967 & ~w25085;
assign w65663 = w25969 & w25085;
assign w65664 = ~w25975 & pi1396;
assign w65665 = w25975 & ~pi1396;
assign w65666 = w25820 & w25896;
assign w65667 = w25820 & ~w63806;
assign w65668 = w25988 & w25820;
assign w65669 = w25986 & pi1408;
assign w65670 = ~w25986 & ~pi1408;
assign w65671 = w26004 & ~w25820;
assign w65672 = ~w26042 & ~w25536;
assign w65673 = ~w25354 & w26067;
assign w65674 = ~w26112 & w25820;
assign w65675 = w26118 & ~w25820;
assign w65676 = w25692 & w25536;
assign w65677 = w26194 & w26188;
assign w65678 = w26274 & w26251;
assign w65679 = w26298 & w26283;
assign w65680 = w26304 & w26323;
assign w65681 = w26320 & pi1441;
assign w65682 = ~w26320 & ~pi1441;
assign w65683 = ~w26345 & ~w26358;
assign w65684 = w26380 & w26386;
assign w65685 = w26391 & w26389;
assign w65686 = w26405 & ~w26386;
assign w65687 = ~w26366 & ~w26409;
assign w65688 = ~w63809 & ~w26473;
assign w65689 = w26492 & ~w26507;
assign w65690 = ~w26499 & ~pi1452;
assign w65691 = w26499 & pi1452;
assign w65692 = w26500 & ~w26486;
assign w65693 = w26510 & ~w26488;
assign w65694 = ~w26552 & ~pi1449;
assign w65695 = w26552 & pi1449;
assign w65696 = ~w26589 & w26583;
assign w65697 = ~w26736 & ~w26594;
assign w65698 = ~w26731 & ~pi1446;
assign w65699 = w26731 & pi1446;
assign w65700 = w26756 & w26621;
assign w65701 = ~w26769 & ~w26772;
assign w65702 = pi1450 & ~w26773;
assign w65703 = pi1450 & ~w63820;
assign w65704 = ~pi1450 & w26773;
assign w65705 = ~pi1450 & w63820;
assign w65706 = w26681 & w26666;
assign w65707 = w26685 & w26830;
assign w65708 = ~w26831 & ~w26836;
assign w65709 = ~w26659 & ~w26666;
assign w65710 = ~w26842 & ~w26694;
assign w65711 = w26848 & ~w26829;
assign w65712 = ~w26866 & ~w26868;
assign w65713 = ~w26880 & ~w26876;
assign w65714 = w26934 & ~w26936;
assign w65715 = w26910 & ~w26934;
assign w65716 = ~w26938 & ~w26943;
assign w65717 = ~w27070 & w27077;
assign w65718 = ~w26267 & w26283;
assign w65719 = w26158 & w26178;
assign w65720 = ~w26178 & ~w26165;
assign w65721 = ~w26158 & ~w26152;
assign w65722 = w27130 & w27127;
assign w65723 = w27152 & ~w27037;
assign w65724 = w27157 & w27174;
assign w65725 = w27161 & pi1454;
assign w65726 = ~w27161 & ~pi1454;
assign w65727 = w27182 & w26283;
assign w65728 = w26934 & ~w26959;
assign w65729 = ~w27200 & ~w27199;
assign w65730 = w27198 & ~w26891;
assign w65731 = w26421 & w26386;
assign w65732 = w26371 & ~w26403;
assign w65733 = w26378 & w26386;
assign w65734 = w27254 & w27258;
assign w65735 = w26583 & w26589;
assign w65736 = w26603 & w26563;
assign w65737 = ~w26755 & ~w26733;
assign w65738 = ~w27278 & ~pi1465;
assign w65739 = w27278 & pi1465;
assign w65740 = w26836 & w26666;
assign w65741 = ~w26667 & ~w27303;
assign w65742 = ~w27316 & pi1472;
assign w65743 = w27316 & ~pi1472;
assign w65744 = w26368 & w27321;
assign w65745 = w26193 & ~w26777;
assign w65746 = ~w27343 & w26184;
assign w65747 = w27371 & ~w27368;
assign w65748 = w27391 & ~w27038;
assign w65749 = ~w26910 & ~w26949;
assign w65750 = w27520 & ~w27493;
assign w65751 = ~w27528 & ~w27641;
assign w65752 = ~w27653 & ~w27535;
assign w65753 = w27649 & w27535;
assign w65754 = w27732 & ~w27690;
assign w65755 = ~w27696 & w27709;
assign w65756 = ~w63831 & w27777;
assign w65757 = ~w27857 & ~pi1508;
assign w65758 = w27857 & pi1508;
assign w65759 = ~w27909 & w27908;
assign w65760 = ~w27898 & ~w27882;
assign w65761 = ~w27889 & w27908;
assign w65762 = ~w27917 & pi1514;
assign w65763 = w27917 & ~pi1514;
assign w65764 = w27963 & ~w27967;
assign w65765 = ~w27465 & w27493;
assign w65766 = w28038 & w27989;
assign w65767 = w27909 & w28077;
assign w65768 = ~w27882 & ~w27889;
assign w65769 = w27882 & w27889;
assign w65770 = w27753 & w27690;
assign w65771 = ~w27728 & ~w27735;
assign w65772 = w28124 & pi1513;
assign w65773 = ~w28124 & ~pi1513;
assign w65774 = ~w27577 & ~w27584;
assign w65775 = ~w27568 & ~w27619;
assign w65776 = w28142 & w28135;
assign w65777 = ~w27812 & ~w27806;
assign w65778 = w28171 & ~w27798;
assign w65779 = w28171 & w63839;
assign w65780 = ~w28178 & ~pi1510;
assign w65781 = w28178 & pi1510;
assign w65782 = w28214 & ~w28194;
assign w65783 = ~w28188 & ~w28194;
assign w65784 = w27728 & w28306;
assign w65785 = ~w27690 & ~w28310;
assign w65786 = w27898 & w27876;
assign w65787 = w28355 & ~w28232;
assign w65788 = w28366 & ~pi1517;
assign w65789 = ~w28366 & pi1517;
assign w65790 = ~w28394 & ~w27798;
assign w65791 = ~w28394 & w63839;
assign w65792 = ~w28399 & ~w27777;
assign w65793 = ~w28399 & ~w63844;
assign w65794 = w28416 & ~w28444;
assign w65795 = ~w28448 & w28444;
assign w65796 = ~w28416 & ~w28455;
assign w65797 = ~w28463 & ~w28456;
assign w65798 = ~w28422 & w28472;
assign w65799 = w28437 & ~w28416;
assign w65800 = w28194 & w28214;
assign w65801 = w28529 & w28232;
assign w65802 = w28585 & ~w27936;
assign w65803 = ~w28021 & ~w27989;
assign w65804 = w28602 & w28049;
assign w65805 = w28622 & pi1527;
assign w65806 = ~w28622 & ~pi1527;
assign w65807 = w27568 & w27584;
assign w65808 = w28632 & ~w28633;
assign w65809 = w27600 & ~w28640;
assign w65810 = w28654 & ~w27690;
assign w65811 = w28661 & pi1540;
assign w65812 = ~w28661 & ~pi1540;
assign w65813 = w28443 & w28416;
assign w65814 = w28699 & ~w28437;
assign w65815 = ~w28410 & ~w28464;
assign w65816 = w28830 & w28839;
assign w65817 = ~w28924 & ~w28898;
assign w65818 = w28951 & ~w28938;
assign w65819 = ~w28973 & w28967;
assign w65820 = ~w28962 & w28991;
assign w65821 = ~w29062 & ~w29037;
assign w65822 = ~w29095 & w29089;
assign w65823 = ~w29095 & ~w63848;
assign w65824 = ~w29050 & w29062;
assign w65825 = w29100 & w29099;
assign w65826 = ~w29096 & pi1570;
assign w65827 = w29096 & ~pi1570;
assign w65828 = w29271 & w29261;
assign w65829 = ~w29267 & w29287;
assign w65830 = ~w29297 & w29291;
assign w65831 = w29307 & ~w29282;
assign w65832 = w29338 & ~w29154;
assign w65833 = ~w29134 & ~w29148;
assign w65834 = ~w29134 & ~w29142;
assign w65835 = ~w29353 & ~w29350;
assign w65836 = w29184 & w29148;
assign w65837 = w29378 & w29384;
assign w65838 = w29507 & w29236;
assign w65839 = w29504 & w29282;
assign w65840 = ~w29051 & w29036;
assign w65841 = ~w29044 & ~w29062;
assign w65842 = ~w29044 & w29062;
assign w65843 = ~w29546 & ~w29554;
assign w65844 = w29602 & ~w29608;
assign w65845 = w29646 & ~w29594;
assign w65846 = w29664 & pi1581;
assign w65847 = ~w29664 & ~pi1581;
assign w65848 = w29598 & ~w29627;
assign w65849 = w29044 & w29036;
assign w65850 = ~w29051 & ~w29053;
assign w65851 = w29099 & ~w29069;
assign w65852 = ~w29450 & ~w29464;
assign w65853 = ~w29483 & ~w29427;
assign w65854 = ~w29761 & w29760;
assign w65855 = ~w28918 & w28883;
assign w65856 = w28792 & w29828;
assign w65857 = w29829 & w29832;
assign w65858 = ~w29003 & ~w28991;
assign w65859 = ~w28972 & w28984;
assign w65860 = w29009 & w28992;
assign w65861 = ~w28973 & w28991;
assign w65862 = w29857 & ~w29873;
assign w65863 = w29880 & w29282;
assign w65864 = w29269 & w29261;
assign w65865 = w29965 & ~w29948;
assign w65866 = w29984 & ~w29973;
assign w65867 = w30026 & w29095;
assign w65868 = w29865 & w28991;
assign w65869 = ~w30094 & w30151;
assign w65870 = w30143 & w30164;
assign w65871 = ~w30088 & w30094;
assign w65872 = ~w30233 & ~w30236;
assign w65873 = ~w30247 & w30211;
assign w65874 = ~w30263 & ~w30256;
assign w65875 = ~w30289 & w30291;
assign w65876 = ~w30293 & ~w30282;
assign w65877 = ~w30294 & ~pi1635;
assign w65878 = w30294 & pi1635;
assign w65879 = ~w30330 & w30323;
assign w65880 = w30359 & w30336;
assign w65881 = w30338 & w30366;
assign w65882 = w30378 & ~w30352;
assign w65883 = w30477 & w30480;
assign w65884 = w30337 & ~w30310;
assign w65885 = w30514 & pi1660;
assign w65886 = ~w30514 & ~pi1660;
assign w65887 = w30624 & w30379;
assign w65888 = w30624 & ~w63857;
assign w65889 = w30716 & w30650;
assign w65890 = w30733 & w30741;
assign w65891 = ~w30558 & ~w30541;
assign w65892 = w30565 & ~w30595;
assign w65893 = w30753 & w30555;
assign w65894 = ~w30797 & ~w30650;
assign w65895 = ~w30803 & w30650;
assign w65896 = ~w30095 & w30082;
assign w65897 = ~w30920 & pi1658;
assign w65898 = w30920 & ~pi1658;
assign w65899 = w30412 & w30399;
assign w65900 = w30961 & w30555;
assign w65901 = ~w63860 & ~w30752;
assign w65902 = ~w30966 & pi1636;
assign w65903 = w30966 & ~pi1636;
assign w65904 = ~w30998 & ~w30821;
assign w65905 = ~w31005 & ~pi1638;
assign w65906 = w31005 & pi1638;
assign w65907 = w30445 & w30429;
assign w65908 = w31009 & w30938;
assign w65909 = w30445 & ~w30423;
assign w65910 = w31027 & ~w30821;
assign w65911 = w31038 & w31031;
assign w65912 = ~w31042 & w31043;
assign w65913 = ~w30231 & ~w30278;
assign w65914 = ~w63854 & ~w31095;
assign w65915 = ~w31112 & pi1671;
assign w65916 = w31112 & ~pi1671;
assign w65917 = w31129 & w31142;
assign w65918 = ~w31129 & w31192;
assign w65919 = ~w31142 & w31122;
assign w65920 = ~w31226 & pi1673;
assign w65921 = w31226 & ~pi1673;
assign w65922 = w31182 & ~w31169;
assign w65923 = w30692 & w30723;
assign w65924 = w31263 & pi1650;
assign w65925 = ~w31263 & ~pi1650;
assign w65926 = w31287 & w30461;
assign w65927 = ~w30429 & ~w30471;
assign w65928 = w31299 & ~w30461;
assign w65929 = w31320 & ~w31182;
assign w65930 = w31333 & ~w30243;
assign w65931 = w31083 & w30278;
assign w65932 = w31402 & ~w31399;
assign w65933 = w31444 & w31435;
assign w65934 = w31440 & ~w31446;
assign w65935 = ~w31473 & w31493;
assign w65936 = ~w31525 & w31479;
assign w65937 = w31531 & w31524;
assign w65938 = ~w31584 & ~w31571;
assign w65939 = ~w31711 & w31652;
assign w65940 = ~w31778 & w31757;
assign w65941 = w31787 & w31772;
assign w65942 = w31772 & w31790;
assign w65943 = w31788 & w31745;
assign w65944 = w31880 & ~w31839;
assign w65945 = w31911 & ~pi1708;
assign w65946 = ~w31911 & pi1708;
assign w65947 = ~w31933 & w31939;
assign w65948 = w31959 & ~w31939;
assign w65949 = ~w31940 & w31958;
assign w65950 = ~w31972 & ~w31927;
assign w65951 = w31988 & pi1710;
assign w65952 = ~w31988 & ~pi1710;
assign w65953 = ~w31764 & w31778;
assign w65954 = ~w31778 & ~w31757;
assign w65955 = ~w31772 & w31757;
assign w65956 = w32041 & w31779;
assign w65957 = ~w32037 & ~pi1716;
assign w65958 = w32037 & pi1716;
assign w65959 = ~w32073 & ~w32081;
assign w65960 = ~w32082 & w31958;
assign w65961 = w31958 & w32091;
assign w65962 = ~w32035 & ~w31772;
assign w65963 = w31486 & w31493;
assign w65964 = ~w32122 & ~w32124;
assign w65965 = w32156 & ~w32178;
assign w65966 = ~w32149 & ~w32184;
assign w65967 = w32184 & ~w32178;
assign w65968 = ~w32228 & pi1727;
assign w65969 = w32228 & ~pi1727;
assign w65970 = w32252 & ~w31704;
assign w65971 = w31682 & ~w32258;
assign w65972 = ~w32261 & w31704;
assign w65973 = w31652 & ~w32258;
assign w65974 = ~w32262 & pi1711;
assign w65975 = w32262 & ~pi1711;
assign w65976 = ~w31665 & ~w31708;
assign w65977 = ~w32303 & ~pi1721;
assign w65978 = w32303 & pi1721;
assign w65979 = w31577 & ~w31595;
assign w65980 = ~w32342 & ~w31524;
assign w65981 = ~w32356 & w31524;
assign w65982 = w32191 & w32223;
assign w65983 = w32187 & w32178;
assign w65984 = w32379 & pi1726;
assign w65985 = ~w32379 & ~pi1726;
assign w65986 = w32407 & ~w31839;
assign w65987 = w32446 & ~w32442;
assign w65988 = ~w31392 & ~w31379;
assign w65989 = w32457 & ~w31423;
assign w65990 = w32479 & pi1717;
assign w65991 = ~w32479 & ~pi1717;
assign w65992 = ~w32503 & ~w31958;
assign w65993 = w32506 & w31958;
assign w65994 = w31425 & ~w31416;
assign w65995 = ~w31583 & ~w31571;
assign w65996 = w31634 & w31583;
assign w65997 = w32566 & ~w32567;
assign w65998 = ~w32184 & w32590;
assign w65999 = ~w31608 & ~w31595;
assign w66000 = w32612 & w31603;
assign w66001 = w32543 & ~w31427;
assign w66002 = w32705 & w32712;
assign w66003 = w32800 & w32788;
assign w66004 = w32825 & w32844;
assign w66005 = w32849 & w32833;
assign w66006 = ~w32782 & w32861;
assign w66007 = ~w32849 & ~w32782;
assign w66008 = w32938 & ~w32905;
assign w66009 = ~w32946 & ~w32953;
assign w66010 = w32960 & ~w32933;
assign w66011 = ~w33013 & ~w33022;
assign w66012 = ~w33022 & ~w33006;
assign w66013 = w33031 & ~w33022;
assign w66014 = ~w33000 & w33022;
assign w66015 = w33087 & w32994;
assign w66016 = ~w33080 & ~w32994;
assign w66017 = w33102 & ~w33098;
assign w66018 = w33022 & ~w33045;
assign w66019 = w33058 & w32994;
assign w66020 = w32955 & ~w32936;
assign w66021 = w33223 & w33233;
assign w66022 = w33315 & ~w33288;
assign w66023 = w33324 & w33344;
assign w66024 = ~w33423 & ~w33418;
assign w66025 = w33425 & w33442;
assign w66026 = ~w33484 & ~w33296;
assign w66027 = ~w33180 & ~w33174;
assign w66028 = w32953 & w33584;
assign w66029 = w33399 & w33634;
assign w66030 = w33297 & ~w33288;
assign w66031 = w33668 & pi1767;
assign w66032 = ~w33668 & ~pi1767;
assign w66033 = w33518 & ~w33679;
assign w66034 = w32722 & w32734;
assign w66035 = ~w33704 & w32758;
assign w66036 = w33721 & w32692;
assign w66037 = w33081 & ~w33022;
assign w66038 = ~w33167 & ~w33198;
assign w66039 = w33167 & w33180;
assign w66040 = w33770 & w33778;
assign w66041 = w33872 & ~w33826;
assign w66042 = ~w33874 & w33820;
assign w66043 = w33845 & w33857;
assign w66044 = ~w33889 & ~w33887;
assign w66045 = w33696 & ~w32723;
assign w66046 = w33929 & w33930;
assign w66047 = ~w33966 & pi1782;
assign w66048 = w33966 & ~pi1782;
assign w66049 = w33847 & w33820;
assign w66050 = w33977 & ~w33820;
assign w66051 = w33864 & ~w33848;
assign w66052 = w34049 & w34033;
assign w66053 = ~w34026 & w34039;
assign w66054 = ~w34065 & ~w34074;
assign w66055 = w34072 & ~w34078;
assign w66056 = ~w34091 & w34057;
assign w66057 = w34168 & w34148;
assign w66058 = w34113 & w34140;
assign w66059 = ~w34132 & ~w34140;
assign w66060 = ~w34132 & ~w34120;
assign w66061 = ~w34091 & ~w34234;
assign w66062 = w34237 & w34026;
assign w66063 = w34239 & w34057;
assign w66064 = w34245 & ~w34057;
assign w66065 = ~w34303 & w34322;
assign w66066 = w34306 & ~w34283;
assign w66067 = ~w34264 & w34270;
assign w66068 = w34098 & ~w34026;
assign w66069 = w34372 & ~pi1863;
assign w66070 = ~w34372 & pi1863;
assign w66071 = w34495 & ~w34501;
assign w66072 = w34534 & ~w34495;
assign w66073 = w34533 & w34476;
assign w66074 = w34555 & ~w34554;
assign w66075 = w34176 & w34132;
assign w66076 = w34588 & ~w34587;
assign w66077 = ~w34626 & ~w34648;
assign w66078 = w34632 & w34670;
assign w66079 = w34723 & ~w34725;
assign w66080 = ~w34765 & w34772;
assign w66081 = w34153 & ~w34847;
assign w66082 = ~w34853 & ~w34164;
assign w66083 = w34203 & ~w34856;
assign w66084 = ~w34909 & w34935;
assign w66085 = ~w34936 & pi1827;
assign w66086 = w34936 & ~pi1827;
assign w66087 = ~w34963 & pi1840;
assign w66088 = w34963 & ~pi1840;
assign w66089 = ~w34632 & ~w34642;
assign w66090 = ~w34659 & ~w34969;
assign w66091 = w35050 & w34642;
assign w66092 = w35063 & ~w35058;
assign w66093 = w35097 & w35100;
assign w66094 = w35102 & w34517;
assign w66095 = w35102 & ~w63901;
assign w66096 = ~w35158 & w35136;
assign w66097 = w35135 & ~w35156;
assign w66098 = w35135 & w63902;
assign w66099 = w35208 & w35121;
assign w66100 = ~w35204 & w35218;
assign w66101 = w35235 & ~w35121;
assign w66102 = ~w35255 & ~w35261;
assign w66103 = ~w35305 & w35121;
assign w66104 = w34442 & ~w34943;
assign w66105 = w34445 & ~w35313;
assign w66106 = ~w35325 & w34416;
assign w66107 = w34502 & ~w34521;
assign w66108 = ~w35372 & w35378;
assign w66109 = w35365 & w35359;
assign w66110 = w35365 & ~w35378;
assign w66111 = w35408 & w35416;
assign w66112 = w35378 & w35414;
assign w66113 = w35432 & w35431;
assign w66114 = ~w35465 & w35446;
assign w66115 = w35518 & ~w35508;
assign w66116 = ~w35414 & ~w35545;
assign w66117 = w35700 & ~w35698;
assign w66118 = ~w35705 & ~w35722;
assign w66119 = ~w35695 & ~w35746;
assign w66120 = w35720 & ~pi1897;
assign w66121 = ~w35720 & pi1897;
assign w66122 = ~w35803 & ~w35758;
assign w66123 = ~w35803 & w63908;
assign w66124 = w35785 & w35765;
assign w66125 = w35427 & w35378;
assign w66126 = w35535 & ~w35852;
assign w66127 = w35406 & w35378;
assign w66128 = w35856 & w35378;
assign w66129 = ~w35365 & ~w35378;
assign w66130 = w35547 & w35414;
assign w66131 = ~w36070 & w36060;
assign w66132 = ~w36046 & w36038;
assign w66133 = w36117 & w36132;
assign w66134 = w36177 & w36184;
assign w66135 = w36198 & w35596;
assign w66136 = w35613 & ~w36193;
assign w66137 = w36267 & w36224;
assign w66138 = w36272 & ~w36251;
assign w66139 = ~w36093 & ~w36065;
assign w66140 = w36093 & w36081;
assign w66141 = ~w35596 & w35589;
assign w66142 = ~w36365 & ~w36362;
assign w66143 = ~w35709 & ~w36372;
assign w66144 = ~w35692 & ~w35689;
assign w66145 = ~w36378 & pi1913;
assign w66146 = w36378 & ~pi1913;
assign w66147 = w36254 & w36395;
assign w66148 = w36254 & ~w63911;
assign w66149 = w36415 & ~w36264;
assign w66150 = w36445 & w36448;
assign w66151 = w36449 & w36264;
assign w66152 = w35823 & ~w35758;
assign w66153 = ~w35771 & ~w35788;
assign w66154 = w36511 & w36509;
assign w66155 = w36265 & w36286;
assign w66156 = ~w35518 & w35489;
assign w66157 = w36562 & pi1902;
assign w66158 = ~w36562 & ~pi1902;
assign w66159 = ~w35573 & w35596;
assign w66160 = ~w36642 & ~w36066;
assign w66161 = ~w36693 & w36687;
assign w66162 = ~w36734 & ~w36755;
assign w66163 = ~w36687 & ~w36760;
assign w66164 = pi1960 & w63917;
assign w66165 = pi1960 & w36959;
assign w66166 = ~pi1960 & ~w63917;
assign w66167 = ~pi1960 & ~w36959;
assign w66168 = w37022 & w36998;
assign w66169 = ~w36981 & w36998;
assign w66170 = w37052 & pi1953;
assign w66171 = ~w37052 & ~pi1953;
assign w66172 = pi1952 & ~w37103;
assign w66173 = pi1952 & w63922;
assign w66174 = ~pi1952 & w37103;
assign w66175 = ~pi1952 & ~w63922;
assign w66176 = w37208 & ~w37210;
assign w66177 = ~w37177 & w37190;
assign w66178 = ~w37241 & ~w37231;
assign w66179 = ~w36797 & ~w36785;
assign w66180 = w36845 & w36848;
assign w66181 = ~w37329 & pi1955;
assign w66182 = w37329 & ~pi1955;
assign w66183 = ~w37344 & w37373;
assign w66184 = ~w37461 & w37463;
assign w66185 = ~w37488 & pi1957;
assign w66186 = w37488 & ~pi1957;
assign w66187 = w63916 & w36919;
assign w66188 = ~w37511 & w37351;
assign w66189 = w37374 & ~w37378;
assign w66190 = w37536 & w37532;
assign w66191 = w37536 & ~w63933;
assign w66192 = ~w36888 & w36869;
assign w66193 = w37542 & pi1963;
assign w66194 = ~w37542 & ~pi1963;
assign w66195 = w37557 & w37100;
assign w66196 = ~w37551 & ~w37562;
assign w66197 = w37564 & ~pi1964;
assign w66198 = ~w37564 & pi1964;
assign w66199 = ~w37338 & w37568;
assign w66200 = ~w37580 & ~w37577;
assign w66201 = w37583 & w37401;
assign w66202 = w36981 & ~w36998;
assign w66203 = ~w37613 & ~w37006;
assign w66204 = ~w36981 & w37614;
assign w66205 = ~w37630 & pi1958;
assign w66206 = w37630 & ~pi1958;
assign w66207 = ~w37634 & ~w37222;
assign w66208 = w37651 & pi1986;
assign w66209 = ~w37651 & ~pi1986;
assign w66210 = ~w37659 & w37006;
assign w66211 = w37307 & w37318;
assign w66212 = ~w36845 & ~w36832;
assign w66213 = w37344 & w37401;
assign w66214 = ~w37701 & w37702;
assign w66215 = ~w37727 & ~w36752;
assign w66216 = w37737 & ~w37723;
assign w66217 = w37748 & pi1984;
assign w66218 = ~w37748 & ~pi1984;
assign w66219 = w36693 & w37729;
assign w66220 = ~w36738 & ~w37729;
assign w66221 = ~w37764 & ~pi1996;
assign w66222 = w37764 & pi1996;
assign w66223 = w37780 & w37781;
assign w66224 = w37298 & w36791;
assign w66225 = w37782 & ~w37774;
assign w66226 = w37833 & ~w37808;
assign w66227 = w37821 & ~w37831;
assign w66228 = w63950 & w37828;
assign w66229 = (w37828 & w63950) | (w37828 & w37932) | (w63950 & w37932);
assign w66230 = ~w37938 & ~w37828;
assign w66231 = w38019 & w38000;
assign w66232 = ~w38006 & w38012;
assign w66233 = ~w38037 & w38031;
assign w66234 = ~w38000 & ~w38023;
assign w66235 = w38045 & w38063;
assign w66236 = ~w38084 & ~w38090;
assign w66237 = w38167 & w38168;
assign w66238 = ~w38191 & ~w38219;
assign w66239 = ~w38178 & w38229;
assign w66240 = w38242 & w38208;
assign w66241 = w38253 & w38245;
assign w66242 = w38254 & ~w38208;
assign w66243 = ~w38208 & w38191;
assign w66244 = ~w38210 & w38229;
assign w66245 = w38099 & w38090;
assign w66246 = ~w38336 & w38370;
assign w66247 = w38447 & w38441;
assign w66248 = ~w38441 & ~w38447;
assign w66249 = ~w38474 & w38479;
assign w66250 = ~w38488 & w38459;
assign w66251 = w38441 & w38421;
assign w66252 = w38467 & w38421;
assign w66253 = w38459 & ~w38453;
assign w66254 = w38528 & w38597;
assign w66255 = ~w38450 & w38427;
assign w66256 = ~w38441 & w38421;
assign w66257 = ~w38622 & ~w38505;
assign w66258 = ~w38178 & ~w38230;
assign w66259 = w38669 & ~w38682;
assign w66260 = w38006 & w37994;
assign w66261 = w38792 & ~w38764;
assign w66262 = ~w38028 & ~w38066;
assign w66263 = w38043 & ~w37994;
assign w66264 = w38806 & w38818;
assign w66265 = w38135 & w38321;
assign w66266 = ~w38544 & ~w38528;
assign w66267 = w38858 & ~w38838;
assign w66268 = ~w38253 & ~w38229;
assign w66269 = ~w38972 & ~w39007;
assign w66270 = w38982 & ~w38976;
assign w66271 = ~w39013 & pi2034;
assign w66272 = w39013 & ~pi2034;
assign w66273 = w38954 & ~w38960;
assign w66274 = w39021 & ~w38982;
assign w66275 = w39033 & w38972;
assign w66276 = w38689 & w38663;
assign w66277 = ~w38663 & w38669;
assign w66278 = ~w39051 & ~w39061;
assign w66279 = w39067 & ~w39048;
assign w66280 = w39085 & ~w38363;
assign w66281 = w39087 & ~w39091;
assign w66282 = w39090 & ~w39103;
assign w66283 = ~w39137 & ~w38572;
assign w66284 = ~w39150 & ~w38543;
assign w66285 = w39155 & pi2050;
assign w66286 = ~w39155 & ~pi2050;
assign w66287 = w38051 & w37994;
assign w66288 = w39032 & w38982;
assign w66289 = ~w38560 & ~w38528;
assign w66290 = w39200 & w38572;
assign w66291 = w39209 & ~w39210;
assign w66292 = ~w39222 & w38982;
assign w66293 = w38987 & ~w38972;
assign w66294 = ~w38693 & w38691;
assign w66295 = ~w39068 & ~w38699;
assign w66296 = w38370 & ~w38891;
assign w66297 = ~w39310 & ~w39317;
assign w66298 = w39421 & ~w39429;
assign w66299 = w39441 & w39419;
assign w66300 = w39441 & w39430;
assign w66301 = w39443 & w39445;
assign w66302 = w39455 & w39472;
assign w66303 = w39429 & w39450;
assign w66304 = w39487 & pi2152;
assign w66305 = ~w39487 & ~pi2152;
assign w66306 = w39496 & ~w39509;
assign w66307 = ~w39594 & pi2169;
assign w66308 = w39594 & ~pi2169;
assign w66309 = w39615 & w39365;
assign w66310 = w39619 & ~w39375;
assign w66311 = ~w39696 & w39661;
assign w66312 = ~w39727 & w39531;
assign w66313 = w39509 & w39503;
assign w66314 = ~w39742 & w39743;
assign w66315 = w39729 & w39509;
assign w66316 = w39783 & ~w39764;
assign w66317 = ~w39791 & w39770;
assign w66318 = w39828 & w39813;
assign w66319 = w39813 & w39849;
assign w66320 = w39317 & ~w39338;
assign w66321 = ~w39304 & w39862;
assign w66322 = ~w39304 & ~w63964;
assign w66323 = w39863 & ~w39872;
assign w66324 = w39680 & w39678;
assign w66325 = ~w39927 & ~w39936;
assign w66326 = w39927 & w39942;
assign w66327 = ~w39978 & ~w39983;
assign w66328 = w39522 & ~w39509;
assign w66329 = w39496 & w39516;
assign w66330 = w40025 & w39531;
assign w66331 = ~w39954 & w39943;
assign w66332 = ~w39942 & w39914;
assign w66333 = ~w40062 & ~w39942;
assign w66334 = w39920 & ~w39976;
assign w66335 = ~w40081 & ~w39963;
assign w66336 = ~w40143 & w40104;
assign w66337 = w40152 & ~w40137;
assign w66338 = ~w40160 & w40138;
assign w66339 = ~w40160 & ~w40154;
assign w66340 = w40178 & w40197;
assign w66341 = ~w40211 & ~pi2148;
assign w66342 = w40211 & pi2148;
assign w66343 = w40196 & w40223;
assign w66344 = ~w40162 & w40160;
assign w66345 = w40224 & w40237;
assign w66346 = ~w40244 & ~w39813;
assign w66347 = ~w39826 & ~w39835;
assign w66348 = ~w40255 & w39813;
assign w66349 = w40256 & pi2151;
assign w66350 = ~w40256 & ~pi2151;
assign w66351 = w40271 & w39531;
assign w66352 = ~w40269 & ~pi2161;
assign w66353 = w40269 & pi2161;
assign w66354 = ~w40304 & w40310;
assign w66355 = w39648 & w39642;
assign w66356 = ~w39642 & ~w39712;
assign w66357 = w40365 & w40362;
assign w66358 = w40311 & w40314;
assign w66359 = w40389 & w40325;
assign w66360 = w40318 & ~w40395;
assign w66361 = ~w40284 & ~w40291;
assign w66362 = w39479 & w40477;
assign w66363 = w39481 & w39441;
assign w66364 = ~w40503 & ~w39951;
assign w66365 = ~w40507 & pi2157;
assign w66366 = w40507 & ~pi2157;
assign w66367 = ~w40332 & w40524;
assign w66368 = w40528 & ~w40297;
assign w66369 = w40552 & ~w40562;
assign w66370 = ~w40624 & ~w40653;
assign w66371 = w40753 & ~w40759;
assign w66372 = ~w40725 & w40731;
assign w66373 = ~w40706 & ~w40765;
assign w66374 = w40777 & w40706;
assign w66375 = w40676 & w40610;
assign w66376 = ~w40643 & w40633;
assign w66377 = ~w40810 & ~w40804;
assign w66378 = w40829 & ~w40842;
assign w66379 = w40855 & ~w40860;
assign w66380 = w41000 & w40982;
assign w66381 = w40688 & ~w40674;
assign w66382 = w40829 & w40823;
assign w66383 = ~w63978 & w40864;
assign w66384 = ~w41108 & pi2085;
assign w66385 = w41108 & ~pi2085;
assign w66386 = w41218 & ~w41216;
assign w66387 = ~w41063 & w40952;
assign w66388 = ~w41030 & w40989;
assign w66389 = w40999 & ~w40982;
assign w66390 = w41255 & ~w41242;
assign w66391 = ~w41333 & w41347;
assign w66392 = ~w41334 & ~w41375;
assign w66393 = w41411 & w40706;
assign w66394 = w40761 & w40759;
assign w66395 = w41420 & pi2101;
assign w66396 = ~w41420 & ~pi2101;
assign w66397 = w41466 & w40706;
assign w66398 = w41472 & ~w41464;
assign w66399 = ~w40706 & ~w40725;
assign w66400 = w40777 & ~w40718;
assign w66401 = w41479 & ~w40759;
assign w66402 = w41528 & ~w41496;
assign w66403 = w41508 & w41544;
assign w66404 = w41548 & ~w41543;
assign w66405 = w41543 & ~w41557;
assign w66406 = ~w41562 & ~w41534;
assign w66407 = ~w41588 & ~w41168;
assign w66408 = ~w41588 & w41593;
assign w66409 = w41649 & w41612;
assign w66410 = w41675 & ~w41646;
assign w66411 = w41624 & ~w41637;
assign w66412 = ~w41705 & w41646;
assign w66413 = w41702 & w41612;
assign w66414 = ~w41698 & ~w41700;
assign w66415 = ~w41367 & ~w41361;
assign w66416 = w41357 & ~w41386;
assign w66417 = w41646 & w41660;
assign w66418 = w41825 & ~w41612;
assign w66419 = ~w41652 & w41631;
assign w66420 = w41831 & ~w41646;
assign w66421 = w41827 & pi2127;
assign w66422 = ~w41827 & ~pi2127;
assign w66423 = w41842 & ~w41646;
assign w66424 = w41669 & w41652;
assign w66425 = ~w41612 & ~w41668;
assign w66426 = ~w41849 & w41646;
assign w66427 = ~w41528 & ~w41548;
assign w66428 = ~w41523 & ~w41546;
assign w66429 = w41527 & w41543;
assign w66430 = w41543 & ~w41564;
assign w66431 = ~w41333 & ~w41354;
assign w66432 = w41888 & w41890;
assign w66433 = w41354 & ~w41897;
assign w66434 = ~w41333 & ~w41347;
assign w66435 = w41910 & w41386;
assign w66436 = ~w41918 & w41355;
assign w66437 = w41989 & w41986;
assign w66438 = w41989 & w63983;
assign w66439 = ~w41993 & w41988;
assign w66440 = w42000 & ~w42018;
assign w66441 = w42021 & ~w41986;
assign w66442 = w42000 & w42051;
assign w66443 = w42578 & ~w42616;
assign w66444 = w42578 & ~w63986;
assign w66445 = w42637 & w42641;
assign w66446 = ~w42468 & ~w42516;
assign w66447 = ~w42822 & ~w42406;
assign w66448 = w42872 & w42886;
assign w66449 = w42425 & ~w42359;
assign w66450 = w43014 & w43017;
assign w66451 = w43063 & ~w42640;
assign w66452 = w42981 & w43152;
assign w66453 = ~w43153 & pi2297;
assign w66454 = w43153 & ~pi2297;
assign w66455 = w43158 & w63989;
assign w66456 = w43158 & ~w43126;
assign w66457 = w42981 & ~w43133;
assign w66458 = w42981 & ~w63988;
assign w66459 = w42944 & ~w42981;
assign w66460 = w43164 & pi2289;
assign w66461 = ~w43164 & ~pi2289;
assign w66462 = w42578 & w42649;
assign w66463 = w43220 & ~pi2311;
assign w66464 = ~w43220 & pi2311;
assign w66465 = w43244 & ~w43274;
assign w66466 = w43244 & w43299;
assign w66467 = w43273 & ~w43244;
assign w66468 = w43260 & ~w43266;
assign w66469 = w43317 & ~w43305;
assign w66470 = w43294 & ~w43285;
assign w66471 = ~w43373 & ~w43307;
assign w66472 = w43360 & pi2368;
assign w66473 = ~w43360 & ~pi2368;
assign w66474 = w43416 & ~w43403;
assign w66475 = w43501 & ~w43437;
assign w66476 = w43507 & ~w43447;
assign w66477 = ~w43538 & w43523;
assign w66478 = w43558 & w43544;
assign w66479 = w43529 & ~w43554;
assign w66480 = ~w43554 & ~w43529;
assign w66481 = ~w43532 & ~w43557;
assign w66482 = ~w43589 & w43596;
assign w66483 = w43597 & ~w43603;
assign w66484 = w43644 & w43626;
assign w66485 = ~w43638 & w43619;
assign w66486 = ~w43717 & ~w43732;
assign w66487 = w43766 & w43785;
assign w66488 = ~w43855 & w43858;
assign w66489 = ~w43801 & ~w43841;
assign w66490 = w43857 & w43866;
assign w66491 = ~w43801 & ~w43828;
assign w66492 = w43822 & ~w43841;
assign w66493 = w43918 & ~w43841;
assign w66494 = w43941 & ~w43841;
assign w66495 = ~w43842 & w43841;
assign w66496 = w43945 & w43957;
assign w66497 = w43767 & w43732;
assign w66498 = ~w43767 & w43723;
assign w66499 = w43737 & w43732;
assign w66500 = w43976 & ~w43967;
assign w66501 = ~w43717 & w43732;
assign w66502 = w43992 & ~w43995;
assign w66503 = w44002 & ~w43744;
assign w66504 = w43746 & ~w43744;
assign w66505 = w44016 & ~w43771;
assign w66506 = w44017 & ~w44027;
assign w66507 = ~w43573 & w44032;
assign w66508 = ~w43573 & ~w64000;
assign w66509 = w44052 & pi2345;
assign w66510 = ~w44052 & ~pi2345;
assign w66511 = w44063 & w43573;
assign w66512 = ~pi2350 & ~w44071;
assign w66513 = ~pi2350 & ~w64004;
assign w66514 = pi2350 & w44071;
assign w66515 = pi2350 & w64004;
assign w66516 = w43587 & w44077;
assign w66517 = w44075 & pi2362;
assign w66518 = ~w44075 & ~pi2362;
assign w66519 = w43816 & w43831;
assign w66520 = w44166 & ~w44163;
assign w66521 = ~w44169 & w44135;
assign w66522 = ~w43639 & w43625;
assign w66523 = ~w43639 & ~w43643;
assign w66524 = ~w44248 & ~w44251;
assign w66525 = w44253 & ~w44223;
assign w66526 = ~w44244 & w43625;
assign w66527 = w44244 & ~w43656;
assign w66528 = w44271 & ~w44260;
assign w66529 = ~w44314 & w44308;
assign w66530 = ~w44361 & ~w44333;
assign w66531 = w44313 & w44301;
assign w66532 = ~w44281 & ~w44308;
assign w66533 = w44406 & pi2356;
assign w66534 = ~w44406 & ~pi2356;
assign w66535 = w44308 & ~w44412;
assign w66536 = w44157 & ~w44143;
assign w66537 = ~w44135 & ~w44448;
assign w66538 = w44482 & ~w44481;
assign w66539 = ~w44156 & ~w44182;
assign w66540 = w44182 & ~w44518;
assign w66541 = w44519 & ~pi2354;
assign w66542 = ~w44519 & pi2354;
assign w66543 = w44567 & ~w44528;
assign w66544 = ~w44547 & ~w44585;
assign w66545 = w44561 & w44554;
assign w66546 = ~w44594 & ~w44547;
assign w66547 = w44650 & w44652;
assign w66548 = w44672 & ~w44655;
assign w66549 = ~w44699 & ~pi2425;
assign w66550 = w44699 & pi2425;
assign w66551 = ~w44675 & ~w44680;
assign w66552 = w44733 & ~w44528;
assign w66553 = w44808 & w44779;
assign w66554 = ~w44801 & ~w44816;
assign w66555 = ~w44773 & w44779;
assign w66556 = w44816 & ~w44819;
assign w66557 = w44823 & w44854;
assign w66558 = ~w44878 & ~w44908;
assign w66559 = w44878 & w44894;
assign w66560 = ~w44931 & w44903;
assign w66561 = w44564 & ~w44547;
assign w66562 = w44564 & ~w64017;
assign w66563 = ~w44953 & w44954;
assign w66564 = ~w45059 & ~pi2407;
assign w66565 = w45059 & pi2407;
assign w66566 = w45070 & ~w44547;
assign w66567 = w45071 & w44528;
assign w66568 = w45085 & w44627;
assign w66569 = w44627 & ~w44662;
assign w66570 = w45090 & w45084;
assign w66571 = w44915 & ~w44878;
assign w66572 = w45120 & ~w44919;
assign w66573 = w44894 & w44884;
assign w66574 = w45207 & ~w45190;
assign w66575 = ~w45247 & ~w45190;
assign w66576 = w45280 & ~w45214;
assign w66577 = ~w45259 & w45215;
assign w66578 = w45287 & w45214;
assign w66579 = ~w45352 & ~w45370;
assign w66580 = ~w45333 & w45379;
assign w66581 = w45346 & w45358;
assign w66582 = w45418 & ~w45396;
assign w66583 = ~w45012 & ~w45025;
assign w66584 = w45033 & w44975;
assign w66585 = w45442 & w45012;
assign w66586 = ~w45035 & w45451;
assign w66587 = w45467 & pi2416;
assign w66588 = ~w45467 & ~pi2416;
assign w66589 = w45475 & pi2446;
assign w66590 = ~w45475 & ~pi2446;
assign w66591 = ~w45562 & w45130;
assign w66592 = w45115 & ~w44903;
assign w66593 = w45637 & ~w45670;
assign w66594 = w45644 & w45694;
assign w66595 = w45716 & ~w45706;
assign w66596 = ~w45395 & ~w45333;
assign w66597 = ~w45759 & w45651;
assign w66598 = w45650 & ~w45637;
assign w66599 = ~w45637 & ~w45623;
assign w66600 = w45899 & w45904;
assign w66601 = w45919 & ~w45870;
assign w66602 = w45921 & w45894;
assign w66603 = w64024 & ~w45934;
assign w66604 = w45957 & ~w45951;
assign w66605 = w45935 & w45894;
assign w66606 = ~w45990 & ~w45876;
assign w66607 = ~w45945 & w45867;
assign w66608 = ~w46004 & ~pi2495;
assign w66609 = w46004 & pi2495;
assign w66610 = w46027 & w46020;
assign w66611 = ~w46033 & w46044;
assign w66612 = w46057 & ~w46037;
assign w66613 = w46196 & ~w46209;
assign w66614 = ~w46107 & ~w46131;
assign w66615 = w46350 & ~w46358;
assign w66616 = ~w46362 & ~w46331;
assign w66617 = ~w46402 & pi2489;
assign w66618 = w46402 & ~pi2489;
assign w66619 = w46406 & w46413;
assign w66620 = ~w46337 & ~w46375;
assign w66621 = w46481 & ~w46329;
assign w66622 = ~w46354 & ~w46471;
assign w66623 = w46381 & ~w46337;
assign w66624 = w46044 & w46514;
assign w66625 = ~w46067 & ~w46064;
assign w66626 = ~w46517 & ~pi2471;
assign w66627 = w46517 & pi2471;
assign w66628 = ~w46600 & pi2470;
assign w66629 = w46600 & ~pi2470;
assign w66630 = w46675 & ~w46658;
assign w66631 = ~w46639 & ~w46674;
assign w66632 = ~w46658 & w46696;
assign w66633 = ~w46757 & ~w46785;
assign w66634 = w46785 & ~w46763;
assign w66635 = w46637 & w46674;
assign w66636 = w46900 & ~w46898;
assign w66637 = ~w46936 & w46938;
assign w66638 = w46939 & ~w46190;
assign w66639 = ~w64033 & ~w46816;
assign w66640 = ~w46771 & ~w46998;
assign w66641 = w46988 & pi2483;
assign w66642 = ~w46988 & ~pi2483;
assign w66643 = w46994 & w46809;
assign w66644 = ~w46660 & ~w46650;
assign w66645 = w47042 & pi2485;
assign w66646 = ~w47042 & ~pi2485;
assign w66647 = ~w46869 & ~w46883;
assign w66648 = ~w47050 & ~pi2503;
assign w66649 = w47050 & pi2503;
assign w66650 = w46784 & ~w47012;
assign w66651 = w47100 & ~w46809;
assign w66652 = w47124 & ~w47137;
assign w66653 = ~w47174 & ~w47187;
assign w66654 = ~w47208 & ~w47181;
assign w66655 = w47324 & w47303;
assign w66656 = ~w64034 & ~w47315;
assign w66657 = ~w64035 & ~w47351;
assign w66658 = w47277 & w47201;
assign w66659 = w47352 & ~w47302;
assign w66660 = w47403 & ~w47337;
assign w66661 = ~w47485 & ~w47458;
assign w66662 = ~w47437 & ~w47478;
assign w66663 = ~w47495 & ~w47437;
assign w66664 = ~w47520 & ~w47501;
assign w66665 = w47532 & ~w47437;
assign w66666 = w47480 & ~w47517;
assign w66667 = w47592 & ~w47586;
assign w66668 = ~w47555 & ~w47568;
assign w66669 = w47614 & ~w47549;
assign w66670 = ~w47635 & pi2544;
assign w66671 = w47635 & ~pi2544;
assign w66672 = w47685 & w47680;
assign w66673 = w47690 & ~w47644;
assign w66674 = ~w47735 & ~w47195;
assign w66675 = w47705 & w47657;
assign w66676 = w47753 & w47644;
assign w66677 = ~w47691 & w47671;
assign w66678 = ~w47707 & ~w47773;
assign w66679 = ~w47774 & ~w47644;
assign w66680 = ~w47324 & ~w47415;
assign w66681 = ~w47826 & w47843;
assign w66682 = w47889 & pi2535;
assign w66683 = ~w47889 & ~pi2535;
assign w66684 = ~w47561 & w47568;
assign w66685 = ~w47596 & w47908;
assign w66686 = w47910 & w47911;
assign w66687 = ~w47920 & ~w47644;
assign w66688 = w47928 & w47644;
assign w66689 = ~w47561 & ~w47586;
assign w66690 = ~w47607 & ~w48010;
assign w66691 = ~w47561 & w47586;
assign w66692 = ~w48027 & ~w47549;
assign w66693 = w48041 & w47478;
assign w66694 = w47502 & ~w47437;
assign w66695 = ~w48052 & ~w48036;
assign w66696 = w48117 & ~w48124;
assign w66697 = w48140 & ~w48124;
assign w66698 = ~w48099 & ~w48107;
assign w66699 = w48204 & w48211;
assign w66700 = w47826 & w47843;
assign w66701 = ~w47807 & ~w47843;
assign w66702 = w48247 & w48250;
assign w66703 = ~w48269 & w47867;
assign w66704 = ~w48323 & w48297;
assign w66705 = w48345 & ~w48342;
assign w66706 = w48305 & ~w48330;
assign w66707 = w48373 & w48339;
assign w66708 = w48383 & ~pi2555;
assign w66709 = ~w48383 & pi2555;
assign w66710 = w48398 & w48124;
assign w66711 = w48399 & pi2543;
assign w66712 = ~w48399 & ~pi2543;
assign w66713 = ~w48424 & pi2550;
assign w66714 = w48424 & ~pi2550;
assign w66715 = ~w48359 & w48445;
assign w66716 = ~w48446 & pi2551;
assign w66717 = w48446 & ~pi2551;
assign w66718 = w48346 & w48450;
assign w66719 = ~w48373 & ~w48359;
assign w66720 = ~w48477 & ~w47843;
assign w66721 = ~w48509 & ~w48516;
assign w66722 = ~w48531 & w48490;
assign w66723 = ~w48526 & w48516;
assign w66724 = w48552 & ~w48490;
assign w66725 = w48559 & w48516;
assign w66726 = ~w48595 & ~w48601;
assign w66727 = w48627 & ~w48576;
assign w66728 = w48595 & w48588;
assign w66729 = ~w48588 & ~w48638;
assign w66730 = w48665 & w48662;
assign w66731 = w48711 & w48490;
assign w66732 = w48722 & ~w48744;
assign w66733 = w48776 & ~w48601;
assign w66734 = ~w48601 & w48778;
assign w66735 = w48843 & ~w48845;
assign w66736 = ~w48904 & ~w48898;
assign w66737 = ~w48947 & ~w48911;
assign w66738 = w48927 & w48904;
assign w66739 = w49083 & w49041;
assign w66740 = ~w48918 & w48937;
assign w66741 = ~w48929 & w49112;
assign w66742 = w48503 & w48557;
assign w66743 = ~w48831 & w48797;
assign w66744 = ~w48831 & w64043;
assign w66745 = w48857 & w48868;
assign w66746 = w49164 & ~w49160;
assign w66747 = ~w48852 & w49176;
assign w66748 = w49187 & ~w49198;
assign w66749 = ~w49004 & ~w48991;
assign w66750 = w48985 & ~w48997;
assign w66751 = w49252 & w49291;
assign w66752 = ~w49305 & ~w49291;
assign w66753 = w49363 & ~w49373;
assign w66754 = w49375 & w49365;
assign w66755 = ~w49383 & ~w49374;
assign w66756 = w49389 & w49331;
assign w66757 = ~w48948 & ~w48954;
assign w66758 = ~w49428 & pi2615;
assign w66759 = w49428 & ~pi2615;
assign w66760 = ~w49476 & w49442;
assign w66761 = w49499 & w49501;
assign w66762 = ~w49521 & w49522;
assign w66763 = w49502 & pi2618;
assign w66764 = ~w49502 & ~pi2618;
assign w66765 = w49442 & w49541;
assign w66766 = w49442 & ~w64052;
assign w66767 = w49542 & pi2620;
assign w66768 = ~w49542 & ~pi2620;
assign w66769 = ~w48852 & ~w49171;
assign w66770 = w49559 & w48852;
assign w66771 = ~w49565 & ~w48852;
assign w66772 = w49251 & w49309;
assign w66773 = ~w49600 & pi2611;
assign w66774 = w49600 & ~pi2611;
assign w66775 = ~w49624 & w49621;
assign w66776 = w49626 & w49331;
assign w66777 = ~w49645 & pi2606;
assign w66778 = w49645 & ~pi2606;
assign w66779 = w49405 & ~w49331;
assign w66780 = ~w49398 & w49656;
assign w66781 = ~w49373 & w49402;
assign w66782 = w49653 & w49663;
assign w66783 = w49205 & w49059;
assign w66784 = w48991 & ~w49015;
assign w66785 = ~w48991 & ~w49021;
assign w66786 = w49206 & ~w49049;
assign w66787 = w49679 & w49049;
assign w66788 = w49580 & ~w49258;
assign w66789 = w49406 & w49337;
assign w66790 = w49773 & ~w49397;
assign w66791 = w49776 & ~w49624;
assign w66792 = ~w49818 & ~w49853;
assign w66793 = w49811 & ~w49802;
assign w66794 = ~w49832 & ~pi2669;
assign w66795 = w49832 & pi2669;
assign w66796 = ~w49830 & ~w49833;
assign w66797 = w50014 & w50021;
assign w66798 = w50031 & ~w49853;
assign w66799 = ~w50081 & w50075;
assign w66800 = ~w50062 & ~w50093;
assign w66801 = ~w50082 & ~w50132;
assign w66802 = w50082 & ~w50130;
assign w66803 = ~w50158 & ~w50152;
assign w66804 = ~w50203 & ~w50180;
assign w66805 = w50159 & ~w50165;
assign w66806 = ~w50214 & ~w50218;
assign w66807 = w50152 & w50165;
assign w66808 = ~w50152 & ~w50165;
assign w66809 = ~w50206 & ~pi2663;
assign w66810 = w50206 & pi2663;
assign w66811 = w50282 & w50307;
assign w66812 = w50283 & ~w50294;
assign w66813 = w50317 & w50294;
assign w66814 = ~w50277 & w50294;
assign w66815 = w50354 & ~w50353;
assign w66816 = w50177 & w50165;
assign w66817 = w50075 & w50093;
assign w66818 = w50388 & ~w50378;
assign w66819 = ~w50402 & ~w50400;
assign w66820 = w50357 & w50224;
assign w66821 = ~w50075 & ~w50069;
assign w66822 = w50492 & w50459;
assign w66823 = w50482 & w50508;
assign w66824 = ~w50496 & ~w50479;
assign w66825 = ~w50515 & ~w50520;
assign w66826 = ~w50541 & ~w50224;
assign w66827 = ~w50224 & ~w50213;
assign w66828 = ~w49971 & ~w50551;
assign w66829 = w50479 & ~w50520;
assign w66830 = w50522 & ~w50479;
assign w66831 = ~w50576 & w50517;
assign w66832 = w50580 & ~w50452;
assign w66833 = w50104 & ~w50084;
assign w66834 = ~w50651 & w50665;
assign w66835 = ~w50718 & ~pi2685;
assign w66836 = w50718 & pi2685;
assign w66837 = ~w50769 & w50743;
assign w66838 = w50835 & w49979;
assign w66839 = ~w50835 & w49949;
assign w66840 = ~w50850 & pi2681;
assign w66841 = w50850 & ~pi2681;
assign w66842 = w50871 & ~w50872;
assign w66843 = w50880 & w50665;
assign w66844 = ~w50693 & ~w50697;
assign w66845 = w50934 & ~w50937;
assign w66846 = ~w50755 & ~w50761;
assign w66847 = ~w50911 & w50974;
assign w66848 = w50975 & w50961;
assign w66849 = ~w50258 & w50294;
assign w66850 = w50990 & ~w50987;
assign w66851 = w51041 & ~w51042;
assign w66852 = ~w51049 & ~w51045;
assign w66853 = ~w50996 & w50252;
assign w66854 = w51063 & ~w50314;
assign w66855 = ~w50297 & ~w51080;
assign w66856 = ~w51142 & w51129;
assign w66857 = w51161 & w51182;
assign w66858 = w51181 & ~w51123;
assign w66859 = w51172 & ~w51155;
assign w66860 = w51180 & ~w51202;
assign w66861 = w51282 & ~w51291;
assign w66862 = ~w51289 & ~w51312;
assign w66863 = ~w51289 & ~w51346;
assign w66864 = ~w51325 & ~w51343;
assign w66865 = w51352 & pi2726;
assign w66866 = ~w51352 & ~pi2726;
assign w66867 = ~w51383 & ~w51395;
assign w66868 = ~w51377 & w51395;
assign w66869 = w51384 & w51442;
assign w66870 = w51497 & w51472;
assign w66871 = w51516 & ~w51497;
assign w66872 = ~w51517 & ~w51486;
assign w66873 = w51180 & ~w51149;
assign w66874 = w51200 & ~w51123;
assign w66875 = w51200 & ~w51158;
assign w66876 = w51549 & pi2750;
assign w66877 = ~w51549 & ~pi2750;
assign w66878 = w51604 & w51581;
assign w66879 = ~w51604 & ~w51613;
assign w66880 = w51650 & w51642;
assign w66881 = w51650 & ~w51629;
assign w66882 = w51671 & w51319;
assign w66883 = w51669 & ~w51289;
assign w66884 = ~w51679 & ~w51319;
assign w66885 = ~w51532 & w51706;
assign w66886 = ~w51763 & ~w51740;
assign w66887 = w51747 & w51740;
assign w66888 = ~w51782 & ~w51748;
assign w66889 = w51819 & ~w51342;
assign w66890 = ~w51839 & ~w51852;
assign w66891 = ~w51852 & ~w51845;
assign w66892 = ~w51881 & ~w51845;
assign w66893 = ~w51852 & ~w51869;
assign w66894 = ~w51876 & ~w51900;
assign w66895 = ~w51905 & ~w51914;
assign w66896 = w51816 & ~w51326;
assign w66897 = w51334 & ~w51929;
assign w66898 = w51951 & ~w51962;
assign w66899 = w51747 & ~w51726;
assign w66900 = ~w51860 & w51869;
assign w66901 = w52004 & ~w51900;
assign w66902 = ~w51999 & ~w52011;
assign w66903 = w52029 & w51626;
assign w66904 = ~w52048 & w51486;
assign w66905 = w51690 & w51696;
assign w66906 = ~w52060 & pi2743;
assign w66907 = w52060 & ~pi2743;
assign w66908 = ~w51739 & ~w51779;
assign w66909 = w52065 & w52071;
assign w66910 = w51869 & ~w52086;
assign w66911 = ~w51876 & ~w51880;
assign w66912 = w51660 & w51626;
assign w66913 = ~w51370 & w51395;
assign w66914 = ~w51425 & ~w51400;
assign w66915 = ~w52130 & ~w51422;
assign w66916 = ~w52130 & ~w64082;
assign w66917 = w52209 & ~w52205;
assign w66918 = ~w51761 & ~w51726;
assign w66919 = w52244 & w51759;
assign w66920 = ~w51981 & w52251;
assign w66921 = w51597 & ~w52028;
assign w66922 = ~w52277 & ~pi2751;
assign w66923 = w52277 & pi2751;
assign w66924 = ~w52209 & ~w52201;
assign w66925 = ~w52209 & ~w52183;
assign w66926 = w52337 & ~w52177;
assign w66927 = ~w52337 & w52348;
assign w66928 = w52342 & pi2746;
assign w66929 = ~w52342 & ~pi2746;
assign w66930 = w52128 & ~w51395;
assign w66931 = w52361 & w51422;
assign w66932 = w52429 & ~w52460;
assign w66933 = w52518 & ~w52537;
assign w66934 = w52524 & w52544;
assign w66935 = w52577 & w52544;
assign w66936 = ~w52436 & w52460;
assign w66937 = w52622 & w52476;
assign w66938 = ~w52647 & w52684;
assign w66939 = ~w52681 & ~w52680;
assign w66940 = w52688 & ~w52694;
assign w66941 = ~w52694 & w52678;
assign w66942 = ~w52604 & ~w52460;
assign w66943 = w52469 & ~w52611;
assign w66944 = w52740 & w52742;
assign w66945 = ~w52746 & pi2806;
assign w66946 = w52746 & ~pi2806;
assign w66947 = w52830 & ~w52829;
assign w66948 = ~w52842 & w52756;
assign w66949 = ~w52850 & ~pi2795;
assign w66950 = w52850 & pi2795;
assign w66951 = w52862 & w52678;
assign w66952 = w52694 & w52870;
assign w66953 = ~w52923 & ~w52917;
assign w66954 = w53196 & w53188;
assign w66955 = w53198 & pi2784;
assign w66956 = ~w53198 & ~pi2784;
assign w66957 = ~w53017 & ~w53215;
assign w66958 = w53065 & w53228;
assign w66959 = w52799 & w52756;
assign w66960 = w53235 & pi2799;
assign w66961 = ~w53235 & ~pi2799;
assign w66962 = w53274 & ~w52544;
assign w66963 = w52566 & w52544;
assign w66964 = w53293 & w53300;
assign w66965 = w53179 & w53129;
assign w66966 = w53195 & ~w53188;
assign w66967 = ~w53036 & ~w53051;
assign w66968 = ~w53336 & ~w53335;
assign w66969 = w53344 & ~w53065;
assign w66970 = ~w53371 & w53372;
assign w66971 = w53376 & ~w52954;
assign w66972 = ~w52670 & ~w52659;
assign w66973 = ~w52862 & w52864;
assign w66974 = ~w52581 & ~w53412;
assign w66975 = w52537 & ~w52553;
assign w66976 = ~w53434 & ~w53447;
assign w66977 = ~w53434 & ~w64105;
assign w66978 = ~w53163 & ~w53462;
assign w66979 = w53509 & ~w53493;
assign w66980 = w53545 & ~w53524;
assign w66981 = ~w53559 & w53065;
assign w66982 = ~w64097 & ~w53072;
assign w66983 = ~w53560 & ~pi2800;
assign w66984 = w53560 & pi2800;
assign w66985 = ~w53585 & ~pi2843;
assign w66986 = w53585 & pi2843;
assign w66987 = w53524 & ~w53629;
assign w66988 = w53630 & pi2805;
assign w66989 = ~w53630 & ~pi2805;
assign w66990 = w53529 & ~w53486;
assign w66991 = ~w53479 & ~w53643;
assign w66992 = w53648 & ~w53529;
assign w66993 = ~w53614 & ~w53666;
assign w66994 = w53667 & ~w53524;
assign w66995 = ~w53503 & ~w53675;
assign w66996 = w53136 & ~w53129;
assign w66997 = w53686 & ~w53685;
assign w66998 = w53310 & ~w53130;
assign w66999 = w53731 & ~w53712;
assign w67000 = w53764 & ~w53746;
assign w67001 = w53783 & w53785;
assign w67002 = w53797 & w53734;
assign w67003 = w53804 & w53772;
assign w67004 = w53810 & w53745;
assign w67005 = ~w53811 & w53817;
assign w67006 = ~w53864 & ~w53856;
assign w67007 = w53883 & w53837;
assign w67008 = w53849 & w53837;
assign w67009 = ~w53896 & w53882;
assign w67010 = ~w53901 & ~w53904;
assign w67011 = w53810 & w53718;
assign w67012 = ~w53954 & w53772;
assign w67013 = ~w53950 & ~w53772;
assign w67014 = w53731 & w53800;
assign w67015 = w53955 & pi2869;
assign w67016 = ~w53955 & ~pi2869;
assign w67017 = w53990 & w53996;
assign w67018 = ~w54020 & w54042;
assign w67019 = w54048 & w54022;
assign w67020 = w54111 & ~w54107;
assign w67021 = w54152 & w54069;
assign w67022 = w54160 & pi2848;
assign w67023 = ~w54160 & ~pi2848;
assign w67024 = ~w54116 & w54126;
assign w67025 = w54164 & w54069;
assign w67026 = w54089 & ~w54099;
assign w67027 = w53977 & w54020;
assign w67028 = w53977 & w64112;
assign w67029 = w54274 & ~w54004;
assign w67030 = w54048 & w53996;
assign w67031 = ~w54004 & ~w54283;
assign w67032 = ~w54279 & pi2855;
assign w67033 = w54279 & ~pi2855;
assign w67034 = ~w54363 & ~w54362;
assign w67035 = ~w54344 & ~w54375;
assign w67036 = ~w54304 & w54378;
assign w67037 = ~w54383 & ~w54385;
assign w67038 = ~w53837 & ~w54408;
assign w67039 = w54583 & ~w54591;
assign w67040 = w54435 & w54459;
assign w67041 = ~w54482 & w54487;
assign w67042 = ~w54663 & w54655;
assign w67043 = w54699 & ~w54069;
assign w67044 = w54178 & ~w54106;
assign w67045 = ~w54712 & ~pi2856;
assign w67046 = w54712 & pi2856;
assign w67047 = ~w54486 & ~w54450;
assign w67048 = ~w54435 & w54459;
assign w67049 = ~w54717 & ~w54722;
assign w67050 = ~w54476 & w54766;
assign w67051 = w54657 & ~w54449;
assign w67052 = ~w54048 & ~w54004;
assign w67053 = w53996 & ~w54020;
assign w67054 = w54048 & ~w54828;
assign w67055 = ~w54020 & w54022;
assign w67056 = w54570 & w54563;
assign w67057 = w54840 & ~w54557;
assign w67058 = ~w54617 & ~w54557;
assign w67059 = ~w54363 & ~w54788;
assign w67060 = w54362 & ~w54340;
assign w67061 = ~w54915 & ~pi2883;
assign w67062 = w54915 & pi2883;
assign w67063 = w54048 & ~w54927;
assign w67064 = w54038 & ~w54814;
assign w67065 = ~w54069 & ~w54944;
assign w67066 = ~w54069 & ~w64117;
assign w67067 = ~w54081 & ~w54948;
assign w67068 = ~w54945 & pi2859;
assign w67069 = w54945 & ~pi2859;
assign w67070 = w54600 & w54981;
assign w67071 = ~w54576 & ~w54557;
assign w67072 = ~w54990 & w54600;
assign w67073 = ~w55003 & ~w53902;
assign w67074 = ~w55077 & ~w55074;
assign w67075 = w55098 & ~w55110;
assign w67076 = w55118 & w55110;
assign w67077 = ~w55090 & ~w55091;
assign w67078 = ~w55198 & ~w55194;
assign w67079 = ~w55170 & ~w55164;
assign w67080 = w55177 & ~w55170;
assign w67081 = ~w55170 & ~w55194;
assign w67082 = w55243 & ~w55195;
assign w67083 = w55304 & w55302;
assign w67084 = w55259 & w55266;
assign w67085 = ~w55283 & ~w55268;
assign w67086 = w55340 & ~w55290;
assign w67087 = w55283 & ~w55260;
assign w67088 = w55353 & w55290;
assign w67089 = w55438 & w55410;
assign w67090 = w55393 & ~w55458;
assign w67091 = ~w55500 & w55533;
assign w67092 = w55540 & w55548;
assign w67093 = w55638 & w55621;
assign w67094 = w55671 & w55677;
assign w67095 = ~w55722 & ~w55726;
assign w67096 = ~w55699 & ~w55693;
assign w67097 = ~w55207 & ~w55164;
assign w67098 = ~w55781 & ~w55206;
assign w67099 = w55835 & ~w55823;
assign w67100 = ~w55845 & w55429;
assign w67101 = w55845 & ~w55410;
assign w67102 = w55297 & w55283;
assign w67103 = w55626 & w55621;
assign w67104 = ~w55602 & w55621;
assign w67105 = w55305 & w55290;
assign w67106 = w55895 & ~w55283;
assign w67107 = w55852 & w55439;
assign w67108 = w55844 & w55410;
assign w67109 = w55972 & ~w55419;
assign w67110 = w56000 & pi2932;
assign w67111 = ~w56000 & ~pi2932;
assign w67112 = ~w55090 & ~w55064;
assign w67113 = ~w55477 & ~w55491;
assign w67114 = w55490 & w55477;
assign w67115 = w56107 & w56117;
assign w67116 = ~w56076 & ~w56068;
assign w67117 = w55700 & w55665;
assign w67118 = w55715 & ~w55700;
assign w67119 = w55709 & ~w55707;
assign w67120 = ~w56224 & ~w56061;
assign w67121 = w56181 & w55665;
assign w67122 = ~w56260 & w55699;
assign w67123 = w55699 & ~w56263;
assign w67124 = ~w56283 & pi2927;
assign w67125 = w56283 & ~pi2927;
assign w67126 = ~w56298 & ~pi2931;
assign w67127 = w56298 & pi2931;
assign w67128 = ~w56387 & w56393;
assign w67129 = ~w56473 & w56479;
assign w67130 = ~w56442 & w56448;
assign w67131 = w56489 & ~w56501;
assign w67132 = ~w56567 & w56570;
assign w67133 = w56574 & w56598;
assign w67134 = ~w56368 & ~w56344;
assign w67135 = ~w56614 & ~w56400;
assign w67136 = ~w56616 & ~w56393;
assign w67137 = ~w56619 & w56411;
assign w67138 = ~w56614 & w56401;
assign w67139 = w56671 & w56689;
assign w67140 = w56641 & ~w56647;
assign w67141 = w56698 & ~w56635;
assign w67142 = ~w56681 & w56676;
assign w67143 = w56795 & ~w56750;
assign w67144 = w56805 & ~w56793;
assign w67145 = ~w56855 & pi3190;
assign w67146 = w56855 & ~pi3190;
assign w67147 = ~w56877 & w56884;
assign w67148 = w56957 & ~w56635;
assign w67149 = ~w56532 & w56558;
assign w67150 = w57001 & pi3193;
assign w67151 = ~w57001 & ~pi3193;
assign w67152 = ~w57023 & w57010;
assign w67153 = ~w57052 & ~w57056;
assign w67154 = ~w57047 & ~w57029;
assign w67155 = ~w57016 & w57029;
assign w67156 = ~w56641 & ~w56701;
assign w67157 = w56703 & ~w56674;
assign w67158 = ~w56359 & ~w56396;
assign w67159 = w57120 & w56393;
assign w67160 = ~w56368 & ~w56350;
assign w67161 = w57140 & ~pi3249;
assign w67162 = ~w57140 & pi3249;
assign w67163 = w57197 & w56793;
assign w67164 = w56712 & ~w56676;
assign w67165 = w57236 & w56635;
assign w67166 = ~w57255 & ~w56535;
assign w67167 = w57283 & w57046;
assign w67168 = w57286 & ~w57290;
assign w67169 = ~w56594 & w56532;
assign w67170 = ~w56994 & w57306;
assign w67171 = ~w57307 & ~pi3231;
assign w67172 = w57307 & pi3231;
assign w67173 = w57326 & ~w57323;
assign w67174 = w57376 & w57377;
assign w67175 = w57460 & ~w57413;
assign w67176 = w57474 & pi3331;
assign w67177 = ~w57474 & ~pi3331;
assign w67178 = w57313 & ~w56923;
assign w67179 = w57558 & ~w57569;
assign w67180 = w57394 & ~w57576;
assign w67181 = ~w57585 & w57413;
assign w67182 = ~w57585 & ~w64142;
assign w67183 = w57400 & ~w57620;
assign w67184 = ~w57690 & w57689;
assign w67185 = ~w57711 & pi3762;
assign w67186 = w57711 & ~pi3762;
assign w67187 = w62928 & ~w62586;
assign w67188 = w62928 & ~w63343;
assign w67189 = w55863 & w55866;
assign w67190 = pi2913 & ~w55866;
assign w67191 = pi2913 & ~w64124;
assign w67192 = ~pi2913 & w55866;
assign w67193 = ~pi2913 & w64124;
assign one = 1;
assign po0000 = pi0012;// level 0
assign po0001 = pi0046;// level 0
assign po0002 = pi0001;// level 0
assign po0003 = pi0042;// level 0
assign po0004 = pi0003;// level 0
assign po0005 = pi0057;// level 0
assign po0006 = pi0014;// level 0
assign po0007 = pi0041;// level 0
assign po0008 = pi0020;// level 0
assign po0009 = pi0040;// level 0
assign po0010 = pi0023;// level 0
assign po0011 = pi0082;// level 0
assign po0012 = pi0018;// level 0
assign po0013 = pi0054;// level 0
assign po0014 = pi0013;// level 0
assign po0015 = pi0039;// level 0
assign po0016 = pi0026;// level 0
assign po0017 = pi0047;// level 0
assign po0018 = pi0011;// level 0
assign po0019 = pi0072;// level 0
assign po0020 = pi0015;// level 0
assign po0021 = pi0062;// level 0
assign po0022 = pi0022;// level 0
assign po0023 = pi0073;// level 0
assign po0024 = pi0005;// level 0
assign po0025 = pi0037;// level 0
assign po0026 = pi0008;// level 0
assign po0027 = pi0033;// level 0
assign po0028 = pi0016;// level 0
assign po0029 = pi0034;// level 0
assign po0030 = pi0007;// level 0
assign po0031 = pi0045;// level 0
assign po0032 = pi0010;// level 0
assign po0033 = pi0043;// level 0
assign po0034 = pi0024;// level 0
assign po0035 = pi0038;// level 0
assign po0036 = pi0002;// level 0
assign po0037 = pi0056;// level 0
assign po0038 = pi0019;// level 0
assign po0039 = pi0032;// level 0
assign po0040 = pi0030;// level 0
assign po0041 = pi0081;// level 0
assign po0042 = pi0004;// level 0
assign po0043 = pi0044;// level 0
assign po0044 = pi0009;// level 0
assign po0045 = pi0079;// level 0
assign po0046 = pi0029;// level 0
assign po0047 = pi0078;// level 0
assign po0048 = pi0000;// level 0
assign po0049 = pi0053;// level 0
assign po0050 = pi0006;// level 0
assign po0051 = pi0080;// level 0
assign po0052 = pi0028;// level 0
assign po0053 = pi0048;// level 0
assign po0054 = pi0025;// level 0
assign po0055 = pi0055;// level 0
assign po0056 = pi0021;// level 0
assign po0057 = pi0035;// level 0
assign po0058 = pi0027;// level 0
assign po0059 = pi0052;// level 0
assign po0060 = pi0031;// level 0
assign po0061 = pi0063;// level 0
assign po0062 = pi0017;// level 0
assign po0063 = pi0051;// level 0
assign po0064 = one;// level 0
assign po0065 = pi9041;// level 0
assign po0066 = ~w100;// level 14
assign po0067 = pi0113;// level 0
assign po0068 = w100;// level 14
assign po0069 = pi0105;// level 0
assign po0070 = w117;// level 13
assign po0071 = ~pi0105;// level 0
assign po0072 = pi0110;// level 0
assign po0073 = ~w207;// level 13
assign po0074 = ~pi0110;// level 0
assign po0075 = pi0108;// level 0
assign po0076 = w225;// level 12
assign po0077 = ~pi0108;// level 0
assign po0078 = pi0104;// level 0
assign po0079 = w315;// level 13
assign po0080 = ~pi0104;// level 0
assign po0081 = pi0103;// level 0
assign po0082 = ~w343;// level 13
assign po0083 = ~pi0103;// level 0
assign po0084 = pi0125;// level 0
assign po0085 = ~w360;// level 14
assign po0086 = ~pi0125;// level 0
assign po0087 = pi0100;// level 0
assign po0088 = w444;// level 14
assign po0089 = ~pi0100;// level 0
assign po0090 = pi0099;// level 0
assign po0091 = w538;// level 14
assign po0092 = ~pi0099;// level 0
assign po0093 = pi0139;// level 0
assign po0094 = w624;// level 13
assign po0095 = ~pi0139;// level 0
assign po0096 = pi0096;// level 0
assign po0097 = ~w655;// level 13
assign po0098 = ~pi0096;// level 0
assign po0099 = pi0102;// level 0
assign po0100 = ~w676;// level 14
assign po0101 = ~pi0102;// level 0
assign po0102 = pi0111;// level 0
assign po0103 = ~w707;// level 14
assign po0104 = ~pi0111;// level 0
assign po0105 = pi0115;// level 0
assign po0106 = ~w729;// level 14
assign po0107 = ~pi0115;// level 0
assign po0108 = pi0117;// level 0
assign po0109 = ~w752;// level 13
assign po0110 = ~pi0117;// level 0
assign po0111 = pi0098;// level 0
assign po0112 = ~w774;// level 14
assign po0113 = ~pi0098;// level 0
assign po0114 = pi0097;// level 0
assign po0115 = ~w798;// level 13
assign po0116 = ~pi0097;// level 0
assign po0117 = pi0121;// level 0
assign po0118 = ~w824;// level 14
assign po0119 = ~pi0121;// level 0
assign po0120 = pi0116;// level 0
assign po0121 = ~w849;// level 14
assign po0122 = ~pi0116;// level 0
assign po0123 = pi0101;// level 0
assign po0124 = ~w939;// level 14
assign po0125 = ~pi0101;// level 0
assign po0126 = pi0126;// level 0
assign po0127 = w957;// level 13
assign po0128 = ~pi0126;// level 0
assign po0129 = pi0123;// level 0
assign po0130 = ~w985;// level 13
assign po0131 = ~pi0123;// level 0
assign po0132 = pi0158;// level 0
assign po0133 = ~w1005;// level 14
assign po0134 = ~pi0158;// level 0
assign po0135 = pi0137;// level 0
assign po0136 = ~w1021;// level 13
assign po0137 = ~pi0137;// level 0
assign po0138 = w1050;// level 13
assign po0139 = pi0118;// level 0
assign po0140 = ~w1050;// level 13
assign po0141 = pi0128;// level 0
assign po0142 = ~w1067;// level 14
assign po0143 = ~pi0128;// level 0
assign po0144 = pi0135;// level 0
assign po0145 = ~w1090;// level 14
assign po0146 = ~pi0135;// level 0
assign po0147 = pi0124;// level 0
assign po0148 = ~w1177;// level 13
assign po0149 = ~pi0124;// level 0
assign po0150 = pi0130;// level 0
assign po0151 = ~w1192;// level 13
assign po0152 = ~pi0130;// level 0
assign po0153 = pi0136;// level 0
assign po0154 = ~w1221;// level 14
assign po0155 = ~pi0136;// level 0
assign po0156 = pi0138;// level 0
assign po0157 = ~w1238;// level 12
assign po0158 = ~pi0138;// level 0
assign po0159 = pi0109;// level 0
assign po0160 = ~w1262;// level 13
assign po0161 = ~pi0109;// level 0
assign po0162 = pi0036;// level 0
assign po0163 = pi0058;// level 0
assign po0164 = pi0049;// level 0
assign po0165 = pi0070;// level 0
assign po0166 = w1354;// level 14
assign po0167 = pi0061;// level 0
assign po0168 = pi0060;// level 0
assign po0169 = pi0067;// level 0
assign po0170 = pi0050;// level 0
assign po0171 = pi0066;// level 0
assign po0172 = pi0083;// level 0
assign po0173 = pi0068;// level 0
assign po0174 = pi0064;// level 0
assign po0175 = pi0077;// level 0
assign po0176 = pi0076;// level 0
assign po0177 = ~pi0069;// level 0
assign po0178 = pi0059;// level 0
assign po0179 = w1440;// level 14
assign po0180 = w1534;// level 14
assign po0181 = pi0086;// level 0
assign po0182 = pi0087;// level 0
assign po0183 = pi0074;// level 0
assign po0184 = pi0065;// level 0
assign po0185 = pi0071;// level 0
assign po0186 = pi0084;// level 0
assign po0187 = pi0088;// level 0
assign po0188 = ~w1571;// level 14
assign po0189 = w1600;// level 14
assign po0190 = w1628;// level 14
assign po0191 = ~w1713;// level 14
assign po0192 = pi0075;// level 0
assign po0193 = pi0092;// level 0
assign po0194 = w1747;// level 14
assign po0195 = w1770;// level 14
assign po0196 = ~w1791;// level 14
assign po0197 = w1824;// level 14
assign po0198 = ~w1909;// level 14
assign po0199 = ~w1934;// level 14
assign po0200 = ~w1961;// level 14
assign po0201 = w1978;// level 14
assign po0202 = pi0085;// level 0
assign po0203 = pi0095;// level 0
assign po0204 = ~w2074;// level 14
assign po0205 = ~w2110;// level 14
assign po0206 = ~w2190;// level 14
assign po0207 = w2218;// level 14
assign po0208 = pi0091;// level 0
assign po0209 = pi0089;// level 0
assign po0210 = pi0090;// level 0
assign po0211 = pi0093;// level 0
assign po0212 = pi0094;// level 0
assign po0213 = ~w2242;// level 14
assign po0214 = w2263;// level 14
assign po0215 = w2283;// level 14
assign po0216 = w2317;// level 14
assign po0217 = ~w2402;// level 14
assign po0218 = ~w2424;// level 14
assign po0219 = ~w2446;// level 14
assign po0220 = ~w2466;// level 14
assign po0221 = w2494;// level 14
assign po0222 = w2518;// level 14
assign po0223 = ~w2539;// level 14
assign po0224 = w2560;// level 13
assign po0225 = ~w2581;// level 14
assign po0226 = pi0107;// level 0
assign po0227 = pi0122;// level 0
assign po0228 = pi0106;// level 0
assign po0229 = pi0132;// level 0
assign po0230 = pi0119;// level 0
assign po0231 = pi0120;// level 0
assign po0232 = pi0112;// level 0
assign po0233 = pi0127;// level 0
assign po0234 = pi0114;// level 0
assign po0235 = pi0131;// level 0
assign po0236 = w2678;// level 14
assign po0237 = ~w2706;// level 14
assign po0238 = pi0152;// level 0
assign po0239 = pi0153;// level 0
assign po0240 = pi0140;// level 0
assign po0241 = pi0142;// level 0
assign po0242 = w2723;// level 14
assign po0243 = pi0129;// level 0
assign po0244 = w2814;// level 14
assign po0245 = pi0133;// level 0
assign po0246 = pi0134;// level 0
assign po0247 = pi0146;// level 0
assign po0248 = pi0147;// level 0
assign po0249 = ~w2838;// level 14
assign po0250 = ~w2922;// level 14
assign po0251 = pi0148;// level 0
assign po0252 = ~w2949;// level 14
assign po0253 = pi0150;// level 0
assign po0254 = pi0155;// level 0
assign po0255 = pi0141;// level 0
assign po0256 = pi0143;// level 0
assign po0257 = w3031;// level 14
assign po0258 = pi0144;// level 0
assign po0259 = w3128;// level 14
assign po0260 = pi0145;// level 0
assign po0261 = ~w3148;// level 14
assign po0262 = w3253;// level 14
assign po0263 = ~w3300;// level 14
assign po0264 = ~w3318;// level 14
assign po0265 = pi0149;// level 0
assign po0266 = pi0151;// level 0
assign po0267 = pi0154;// level 0
assign po0268 = pi0156;// level 0
assign po0269 = pi0157;// level 0
assign po0270 = ~w3336;// level 14
assign po0271 = ~w3358;// level 14
assign po0272 = w3448;// level 14
assign po0273 = ~w3474;// level 14
assign po0274 = ~w3497;// level 14
assign po0275 = w3523;// level 14
assign po0276 = ~w3539;// level 14
assign po0277 = w3569;// level 14
assign po0278 = w3594;// level 14
assign po0279 = w3618;// level 14
assign po0280 = w3639;// level 14
assign po0281 = w3719;// level 14
assign po0282 = ~w3731;// level 14
assign po0283 = w3757;// level 14
assign po0284 = ~w3779;// level 13
assign po0285 = ~w3801;// level 14
assign po0286 = ~w3823;// level 14
assign po0287 = ~w3854;// level 14
assign po0288 = pi0159;// level 0
assign po0289 = w3878;// level 14
assign po0290 = pi0177;// level 0
assign po0291 = pi0176;// level 0
assign po0292 = pi0180;// level 0
assign po0293 = pi0181;// level 0
assign po0294 = pi0182;// level 0
assign po0295 = pi0198;// level 0
assign po0296 = pi0203;// level 0
assign po0297 = pi0193;// level 0
assign po0298 = pi0184;// level 0
assign po0299 = pi0196;// level 0
assign po0300 = pi0205;// level 0
assign po0301 = pi0201;// level 0
assign po0302 = pi0202;// level 0
assign po0303 = pi0204;// level 0
assign po0304 = pi0207;// level 0
assign po0305 = pi0185;// level 0
assign po0306 = w3980;// level 14
assign po0307 = ~w4081;// level 14
assign po0308 = pi0206;// level 0
assign po0309 = pi0208;// level 0
assign po0310 = ~w4168;// level 14
assign po0311 = ~w4198;// level 14
assign po0312 = ~w4226;// level 14
assign po0313 = pi0221;// level 0
assign po0314 = ~w4249;// level 14
assign po0315 = w4272;// level 14
assign po0316 = pi0211;// level 0
assign po0317 = pi0212;// level 0
assign po0318 = pi0213;// level 0
assign po0319 = pi0214;// level 0
assign po0320 = pi0215;// level 0
assign po0321 = pi0216;// level 0
assign po0322 = pi0217;// level 0
assign po0323 = w4294;// level 14
assign po0324 = pi0209;// level 0
assign po0325 = pi0218;// level 0
assign po0326 = w4389;// level 14
assign po0327 = pi0223;// level 0
assign po0328 = w4412;// level 14
assign po0329 = pi0219;// level 0
assign po0330 = pi0220;// level 0
assign po0331 = w4499;// level 14
assign po0332 = w4597;// level 14
assign po0333 = ~w4622;// level 14
assign po0334 = ~w4642;// level 14
assign po0335 = w4669;// level 14
assign po0336 = ~w4700;// level 14
assign po0337 = w4789;// level 14
assign po0338 = w4829;// level 14
assign po0339 = w4847;// level 14
assign po0340 = pi0222;// level 0
assign po0341 = ~w4938;// level 14
assign po0342 = ~w4966;// level 14
assign po0343 = ~w4988;// level 14
assign po0344 = ~w5008;// level 14
assign po0345 = w5041;// level 14
assign po0346 = w5075;// level 14
assign po0347 = w5094;// level 14
assign po0348 = w5119;// level 14
assign po0349 = ~w5135;// level 14
assign po0350 = ~w5159;// level 14
assign po0351 = w5184;// level 14
assign po0352 = w5203;// level 14
assign po0353 = ~w5225;// level 14
assign po0354 = pi0251;// level 0
assign po0355 = pi0245;// level 0
assign po0356 = pi0256;// level 0
assign po0357 = pi0250;// level 0
assign po0358 = pi0254;// level 0
assign po0359 = pi0255;// level 0
assign po0360 = pi0257;// level 0
assign po0361 = pi0266;// level 0
assign po0362 = pi0274;// level 0
assign po0363 = pi0261;// level 0
assign po0364 = pi0262;// level 0
assign po0365 = pi0263;// level 0
assign po0366 = pi0275;// level 0
assign po0367 = pi0271;// level 0
assign po0368 = pi0264;// level 0
assign po0369 = pi0265;// level 0
assign po0370 = pi0269;// level 0
assign po0371 = pi0270;// level 0
assign po0372 = pi0272;// level 0
assign po0373 = pi0280;// level 0
assign po0374 = pi0273;// level 0
assign po0375 = w5311;// level 14
assign po0376 = pi0277;// level 0
assign po0377 = pi0278;// level 0
assign po0378 = pi0276;// level 0
assign po0379 = pi0279;// level 0
assign po0380 = w5392;// level 14
assign po0381 = w5423;// level 14
assign po0382 = pi0281;// level 0
assign po0383 = pi0286;// level 0
assign po0384 = w5513;// level 14
assign po0385 = ~w5539;// level 14
assign po0386 = ~w5624;// level 14
assign po0387 = w5666;// level 14
assign po0388 = pi0283;// level 0
assign po0389 = pi0284;// level 0
assign po0390 = pi0285;// level 0
assign po0391 = w5763;// level 14
assign po0392 = ~w5789;// level 14
assign po0393 = w5885;// level 14
assign po0394 = ~w5909;// level 14
assign po0395 = w5930;// level 14
assign po0396 = w5958;// level 14
assign po0397 = pi0282;// level 0
assign po0398 = pi0287;// level 0
assign po0399 = w5980;// level 14
assign po0400 = w6003;// level 14
assign po0401 = ~w6016;// level 14
assign po0402 = w6106;// level 14
assign po0403 = w6131;// level 14
assign po0404 = ~w6146;// level 14
assign po0405 = w6165;// level 14
assign po0406 = ~w6183;// level 14
assign po0407 = ~w6216;// level 14
assign po0408 = w6249;// level 14
assign po0409 = w6278;// level 14
assign po0410 = w6302;// level 14
assign po0411 = ~w6327;// level 14
assign po0412 = w6348;// level 14
assign po0413 = w6367;// level 14
assign po0414 = ~w6457;// level 14
assign po0415 = w6484;// level 15
assign po0416 = w6506;// level 14
assign po0417 = ~w6523;// level 14
assign po0418 = pi0302;// level 0
assign po0419 = pi0323;// level 0
assign po0420 = pi0312;// level 0
assign po0421 = pi0315;// level 0
assign po0422 = pi0322;// level 0
assign po0423 = pi0326;// level 0
assign po0424 = pi0335;// level 0
assign po0425 = pi0329;// level 0
assign po0426 = pi0324;// level 0
assign po0427 = pi0330;// level 0
assign po0428 = pi0341;// level 0
assign po0429 = pi0325;// level 0
assign po0430 = pi0327;// level 0
assign po0431 = pi0328;// level 0
assign po0432 = ~w6617;// level 14
assign po0433 = pi0344;// level 0
assign po0434 = pi0346;// level 0
assign po0435 = pi0332;// level 0
assign po0436 = pi0342;// level 0
assign po0437 = pi0331;// level 0
assign po0438 = pi0333;// level 0
assign po0439 = pi0336;// level 0
assign po0440 = pi0334;// level 0
assign po0441 = pi0337;// level 0
assign po0442 = ~w6703;// level 14
assign po0443 = pi0338;// level 0
assign po0444 = pi0339;// level 0
assign po0445 = ~w6741;// level 14
assign po0446 = pi0343;// level 0
assign po0447 = pi0345;// level 0
assign po0448 = pi0350;// level 0
assign po0449 = pi0347;// level 0
assign po0450 = pi0348;// level 0
assign po0451 = pi0349;// level 0
assign po0452 = w6826;// level 14
assign po0453 = w6852;// level 14
assign po0454 = w6874;// level 14
assign po0455 = w6963;// level 14
assign po0456 = w7054;// level 14
assign po0457 = ~w7081;// level 14
assign po0458 = ~w7113;// level 14
assign po0459 = w7132;// level 14
assign po0460 = w7222;// level 14
assign po0461 = ~w7252;// level 15
assign po0462 = w7284;// level 14
assign po0463 = w7304;// level 14
assign po0464 = w7327;// level 14
assign po0465 = w7415;// level 14
assign po0466 = w7436;// level 14
assign po0467 = ~w7460;// level 14
assign po0468 = ~w7546;// level 14
assign po0469 = w7566;// level 14
assign po0470 = pi0351;// level 0
assign po0471 = ~w7592;// level 15
assign po0472 = w7613;// level 14
assign po0473 = w7647;// level 14
assign po0474 = w7670;// level 14
assign po0475 = w7689;// level 14
assign po0476 = w7712;// level 14
assign po0477 = ~w7732;// level 14
assign po0478 = w7757;// level 14
assign po0479 = ~w7775;// level 14
assign po0480 = w7801;// level 14
assign po0481 = ~w7823;// level 14
assign po0482 = pi0376;// level 0
assign po0483 = pi0386;// level 0
assign po0484 = pi0382;// level 0
assign po0485 = pi0395;// level 0
assign po0486 = pi0383;// level 0
assign po0487 = pi0384;// level 0
assign po0488 = pi0389;// level 0
assign po0489 = pi0387;// level 0
assign po0490 = pi0388;// level 0
assign po0491 = pi0391;// level 0
assign po0492 = pi0404;// level 0
assign po0493 = pi0408;// level 0
assign po0494 = pi0392;// level 0
assign po0495 = pi0394;// level 0
assign po0496 = pi0396;// level 0
assign po0497 = pi0393;// level 0
assign po0498 = pi0397;// level 0
assign po0499 = pi0399;// level 0
assign po0500 = pi0413;// level 0
assign po0501 = pi0400;// level 0
assign po0502 = pi0401;// level 0
assign po0503 = pi0402;// level 0
assign po0504 = pi0403;// level 0
assign po0505 = pi0405;// level 0
assign po0506 = w7912;// level 14
assign po0507 = pi0406;// level 0
assign po0508 = pi0407;// level 0
assign po0509 = pi0410;// level 0
assign po0510 = pi0409;// level 0
assign po0511 = pi0411;// level 0
assign po0512 = ~w7993;// level 14
assign po0513 = ~w8084;// level 14
assign po0514 = ~w8170;// level 14
assign po0515 = pi0412;// level 0
assign po0516 = ~w8206;// level 14
assign po0517 = w8297;// level 14
assign po0518 = w8330;// level 14
assign po0519 = ~w8414;// level 14
assign po0520 = pi0415;// level 0
assign po0521 = w8453;// level 14
assign po0522 = w8490;// level 14
assign po0523 = ~w8512;// level 14
assign po0524 = ~w8534;// level 14
assign po0525 = w8561;// level 13
assign po0526 = w8583;// level 14
assign po0527 = w8615;// level 14
assign po0528 = pi0414;// level 0
assign po0529 = w8698;// level 14
assign po0530 = ~w8722;// level 14
assign po0531 = w8740;// level 14
assign po0532 = w8838;// level 14
assign po0533 = ~w8856;// level 14
assign po0534 = w8879;// level 14
assign po0535 = w8899;// level 14
assign po0536 = w8924;// level 14
assign po0537 = w8945;// level 14
assign po0538 = w8970;// level 14
assign po0539 = ~w8994;// level 14
assign po0540 = ~w9018;// level 14
assign po0541 = ~w9038;// level 14
assign po0542 = ~w9065;// level 14
assign po0543 = ~w9084;// level 14
assign po0544 = w9106;// level 14
assign po0545 = w9129;// level 14
assign po0546 = pi0443;// level 0
assign po0547 = pi0455;// level 0
assign po0548 = pi0440;// level 0
assign po0549 = pi0442;// level 0
assign po0550 = pi0446;// level 0
assign po0551 = pi0448;// level 0
assign po0552 = pi0450;// level 0
assign po0553 = pi0451;// level 0
assign po0554 = pi0466;// level 0
assign po0555 = pi0467;// level 0
assign po0556 = pi0453;// level 0
assign po0557 = pi0460;// level 0
assign po0558 = pi0468;// level 0
assign po0559 = pi0463;// level 0
assign po0560 = pi0472;// level 0
assign po0561 = pi0457;// level 0
assign po0562 = pi0456;// level 0
assign po0563 = pi0459;// level 0
assign po0564 = pi0461;// level 0
assign po0565 = pi0462;// level 0
assign po0566 = pi0464;// level 0
assign po0567 = pi0465;// level 0
assign po0568 = pi0469;// level 0
assign po0569 = pi0470;// level 0
assign po0570 = w9224;// level 14
assign po0571 = pi0473;// level 0
assign po0572 = ~w9244;// level 14
assign po0573 = w9329;// level 14
assign po0574 = pi0474;// level 0
assign po0575 = pi0475;// level 0
assign po0576 = w9422;// level 14
assign po0577 = pi0476;// level 0
assign po0578 = ~w9513;// level 14
assign po0579 = pi0477;// level 0
assign po0580 = w9539;// level 14
assign po0581 = ~w9574;// level 14
assign po0582 = pi0478;// level 0
assign po0583 = w9599;// level 14
assign po0584 = pi0471;// level 0
assign po0585 = w9614;// level 14
assign po0586 = ~w9696;// level 14
assign po0587 = w9786;// level 14
assign po0588 = pi0479;// level 0
assign po0589 = w9805;// level 14
assign po0590 = ~w9835;// level 14
assign po0591 = ~w9920;// level 14
assign po0592 = w10004;// level 14
assign po0593 = w10042;// level 14
assign po0594 = ~w10067;// level 14
assign po0595 = ~w10091;// level 14
assign po0596 = ~w10110;// level 14
assign po0597 = ~w10133;// level 14
assign po0598 = ~w10165;// level 14
assign po0599 = ~w10185;// level 14
assign po0600 = ~w10206;// level 14
assign po0601 = w10225;// level 14
assign po0602 = ~w10255;// level 14
assign po0603 = w10278;// level 14
assign po0604 = w10300;// level 14
assign po0605 = ~w10330;// level 14
assign po0606 = w10359;// level 14
assign po0607 = ~w10382;// level 14
assign po0608 = w10400;// level 14
assign po0609 = w10421;// level 14
assign po0610 = pi0494;// level 0
assign po0611 = pi0520;// level 0
assign po0612 = pi0515;// level 0
assign po0613 = pi0524;// level 0
assign po0614 = pi0509;// level 0
assign po0615 = pi0510;// level 0
assign po0616 = pi0512;// level 0
assign po0617 = pi0517;// level 0
assign po0618 = pi0513;// level 0
assign po0619 = pi0514;// level 0
assign po0620 = pi0528;// level 0
assign po0621 = pi0518;// level 0
assign po0622 = pi0519;// level 0
assign po0623 = pi0521;// level 0
assign po0624 = w10516;// level 14
assign po0625 = pi0537;// level 0
assign po0626 = pi0525;// level 0
assign po0627 = pi0526;// level 0
assign po0628 = pi0527;// level 0
assign po0629 = pi0529;// level 0
assign po0630 = pi0530;// level 0
assign po0631 = pi0531;// level 0
assign po0632 = pi0540;// level 0
assign po0633 = pi0534;// level 0
assign po0634 = pi0533;// level 0
assign po0635 = pi0535;// level 0
assign po0636 = pi0532;// level 0
assign po0637 = pi0536;// level 0
assign po0638 = pi0539;// level 0
assign po0639 = w10617;// level 14
assign po0640 = w10703;// level 14
assign po0641 = pi0541;// level 0
assign po0642 = w10725;// level 14
assign po0643 = ~w10740;// level 14
assign po0644 = w10834;// level 14
assign po0645 = w10918;// level 14
assign po0646 = pi0542;// level 0
assign po0647 = w10949;// level 14
assign po0648 = w11036;// level 14
assign po0649 = w11079;// level 14
assign po0650 = ~w11103;// level 14
assign po0651 = w11141;// level 14
assign po0652 = pi0543;// level 0
assign po0653 = pi0538;// level 0
assign po0654 = w11153;// level 14
assign po0655 = w11194;// level 14
assign po0656 = w11214;// level 14
assign po0657 = w11301;// level 14
assign po0658 = w11332;// level 14
assign po0659 = w11354;// level 14
assign po0660 = w11431;// level 14
assign po0661 = ~w11467;// level 14
assign po0662 = ~w11491;// level 14
assign po0663 = ~w11517;// level 14
assign po0664 = w11540;// level 14
assign po0665 = w11557;// level 14
assign po0666 = ~w11580;// level 14
assign po0667 = ~w11601;// level 14
assign po0668 = ~w11617;// level 14
assign po0669 = ~w11637;// level 14
assign po0670 = ~w11663;// level 14
assign po0671 = ~w11686;// level 14
assign po0672 = w11713;// level 14
assign po0673 = w11734;// level 14
assign po0674 = pi0558;// level 0
assign po0675 = pi0575;// level 0
assign po0676 = pi0582;// level 0
assign po0677 = pi0572;// level 0
assign po0678 = pi0576;// level 0
assign po0679 = pi0577;// level 0
assign po0680 = pi0579;// level 0
assign po0681 = pi0584;// level 0
assign po0682 = pi0592;// level 0
assign po0683 = pi0581;// level 0
assign po0684 = pi0596;// level 0
assign po0685 = pi0583;// level 0
assign po0686 = pi0585;// level 0
assign po0687 = pi0586;// level 0
assign po0688 = w11831;// level 14
assign po0689 = pi0587;// level 0
assign po0690 = pi0588;// level 0
assign po0691 = pi0602;// level 0
assign po0692 = pi0590;// level 0
assign po0693 = pi0591;// level 0
assign po0694 = pi0605;// level 0
assign po0695 = pi0593;// level 0
assign po0696 = pi0594;// level 0
assign po0697 = pi0599;// level 0
assign po0698 = pi0606;// level 0
assign po0699 = pi0595;// level 0
assign po0700 = pi0597;// level 0
assign po0701 = pi0598;// level 0
assign po0702 = ~w11920;// level 14
assign po0703 = pi0600;// level 0
assign po0704 = pi0601;// level 0
assign po0705 = w12013;// level 14
assign po0706 = w12105;// level 14
assign po0707 = w12138;// level 14
assign po0708 = pi0604;// level 0
assign po0709 = ~w12169;// level 14
assign po0710 = pi0607;// level 0
assign po0711 = ~w12268;// level 14
assign po0712 = w12296;// level 14
assign po0713 = ~w12319;// level 14
assign po0714 = w12407;// level 14
assign po0715 = w12434;// level 14
assign po0716 = ~w12523;// level 14
assign po0717 = ~w12545;// level 14
assign po0718 = ~w12565;// level 14
assign po0719 = pi0603;// level 0
assign po0720 = w12597;// level 14
assign po0721 = ~w12632;// level 14
assign po0722 = w12661;// level 14
assign po0723 = ~w12683;// level 15
assign po0724 = w12696;// level 14
assign po0725 = w12718;// level 14
assign po0726 = w12746;// level 14
assign po0727 = ~w12774;// level 14
assign po0728 = w12801;// level 14
assign po0729 = w12824;// level 14
assign po0730 = w12915;// level 14
assign po0731 = w12947;// level 14
assign po0732 = ~w12963;// level 14
assign po0733 = w12982;// level 14
assign po0734 = w13002;// level 14
assign po0735 = ~w13018;// level 14
assign po0736 = ~w13039;// level 14
assign po0737 = w13055;// level 14
assign po0738 = pi0634;// level 0
assign po0739 = pi0646;// level 0
assign po0740 = pi0639;// level 0
assign po0741 = pi0651;// level 0
assign po0742 = pi0636;// level 0
assign po0743 = pi0638;// level 0
assign po0744 = pi0654;// level 0
assign po0745 = pi0648;// level 0
assign po0746 = pi0642;// level 0
assign po0747 = pi0643;// level 0
assign po0748 = pi0653;// level 0
assign po0749 = pi0644;// level 0
assign po0750 = pi0645;// level 0
assign po0751 = pi0647;// level 0
assign po0752 = pi0650;// level 0
assign po0753 = pi0664;// level 0
assign po0754 = pi0652;// level 0
assign po0755 = pi0656;// level 0
assign po0756 = pi0666;// level 0
assign po0757 = pi0655;// level 0
assign po0758 = pi0657;// level 0
assign po0759 = pi0658;// level 0
assign po0760 = pi0660;// level 0
assign po0761 = pi0661;// level 0
assign po0762 = pi0662;// level 0
assign po0763 = pi0668;// level 0
assign po0764 = ~w13146;// level 14
assign po0765 = pi0663;// level 0
assign po0766 = ~w13234;// level 14
assign po0767 = pi0667;// level 0
assign po0768 = w13265;// level 14
assign po0769 = w13352;// level 14
assign po0770 = pi0669;// level 0
assign po0771 = pi0670;// level 0
assign po0772 = w13450;// level 14
assign po0773 = ~w13476;// level 14
assign po0774 = w13513;// level 14
assign po0775 = ~w13535;// level 14
assign po0776 = w13626;// level 14
assign po0777 = w13710;// level 14
assign po0778 = ~w13736;// level 14
assign po0779 = pi0665;// level 0
assign po0780 = w13810;// level 14
assign po0781 = w13847;// level 14
assign po0782 = ~w13936;// level 14
assign po0783 = ~w13975;// level 14
assign po0784 = w14000;// level 14
assign po0785 = w14024;// level 14
assign po0786 = ~w14042;// level 14
assign po0787 = w14079;// level 14
assign po0788 = ~w14098;// level 14
assign po0789 = pi0671;// level 0
assign po0790 = w14125;// level 15
assign po0791 = ~w14146;// level 14
assign po0792 = ~w14164;// level 14
assign po0793 = w14184;// level 14
assign po0794 = ~w14202;// level 14
assign po0795 = w14218;// level 14
assign po0796 = w14258;// level 14
assign po0797 = w14278;// level 14
assign po0798 = w14295;// level 14
assign po0799 = w14316;// level 14
assign po0800 = ~w14336;// level 14
assign po0801 = w14358;// level 14
assign po0802 = pi0691;// level 0
assign po0803 = pi0703;// level 0
assign po0804 = pi0717;// level 0
assign po0805 = pi0704;// level 0
assign po0806 = pi0710;// level 0
assign po0807 = pi0718;// level 0
assign po0808 = pi0705;// level 0
assign po0809 = pi0706;// level 0
assign po0810 = pi0723;// level 0
assign po0811 = pi0708;// level 0
assign po0812 = pi0709;// level 0
assign po0813 = pi0711;// level 0
assign po0814 = pi0712;// level 0
assign po0815 = pi0713;// level 0
assign po0816 = pi0728;// level 0
assign po0817 = pi0715;// level 0
assign po0818 = pi0716;// level 0
assign po0819 = pi0719;// level 0
assign po0820 = pi0720;// level 0
assign po0821 = ~w14447;// level 14
assign po0822 = pi0721;// level 0
assign po0823 = pi0722;// level 0
assign po0824 = pi0724;// level 0
assign po0825 = pi0725;// level 0
assign po0826 = pi0726;// level 0
assign po0827 = pi0727;// level 0
assign po0828 = pi0729;// level 0
assign po0829 = pi0731;// level 0
assign po0830 = pi0730;// level 0
assign po0831 = pi0734;// level 0
assign po0832 = pi0735;// level 0
assign po0833 = w14533;// level 14
assign po0834 = w14621;// level 14
assign po0835 = w14645;// level 14
assign po0836 = w14680;// level 14
assign po0837 = pi0732;// level 0
assign po0838 = w14766;// level 14
assign po0839 = w14861;// level 14
assign po0840 = w14955;// level 14
assign po0841 = ~w14981;// level 14
assign po0842 = w15065;// level 14
assign po0843 = ~w15098;// level 14
assign po0844 = pi0733;// level 0
assign po0845 = ~w15122;// level 14
assign po0846 = ~w15145;// level 14
assign po0847 = ~w15181;// level 14
assign po0848 = w15219;// level 14
assign po0849 = ~w15241;// level 14
assign po0850 = ~w15265;// level 14
assign po0851 = w15290;// level 14
assign po0852 = w15313;// level 14
assign po0853 = w15328;// level 14
assign po0854 = w15348;// level 14
assign po0855 = w15387;// level 14
assign po0856 = ~w15409;// level 14
assign po0857 = w15440;// level 14
assign po0858 = w15467;// level 14
assign po0859 = w15486;// level 14
assign po0860 = ~w15503;// level 14
assign po0861 = w15524;// level 14
assign po0862 = ~w15603;// level 14
assign po0863 = w15628;// level 14
assign po0864 = ~w15659;// level 14
assign po0865 = ~w15677;// level 14
assign po0866 = pi0745;// level 0
assign po0867 = pi0772;// level 0
assign po0868 = pi0762;// level 0
assign po0869 = pi0766;// level 0
assign po0870 = pi0774;// level 0
assign po0871 = pi0781;// level 0
assign po0872 = pi0771;// level 0
assign po0873 = pi0778;// level 0
assign po0874 = pi0773;// level 0
assign po0875 = ~w15772;// level 14
assign po0876 = pi0775;// level 0
assign po0877 = pi0791;// level 0
assign po0878 = pi0776;// level 0
assign po0879 = pi0777;// level 0
assign po0880 = pi0779;// level 0
assign po0881 = pi0780;// level 0
assign po0882 = pi0782;// level 0
assign po0883 = pi0797;// level 0
assign po0884 = pi0784;// level 0
assign po0885 = pi0785;// level 0
assign po0886 = pi0786;// level 0
assign po0887 = pi0787;// level 0
assign po0888 = pi0788;// level 0
assign po0889 = pi0789;// level 0
assign po0890 = pi0790;// level 0
assign po0891 = pi0792;// level 0
assign po0892 = ~w15859;// level 14
assign po0893 = pi0794;// level 0
assign po0894 = pi0795;// level 0
assign po0895 = pi0793;// level 0
assign po0896 = w15945;// level 14
assign po0897 = pi0796;// level 0
assign po0898 = pi0783;// level 0
assign po0899 = pi0798;// level 0
assign po0900 = pi0799;// level 0
assign po0901 = ~w16041;// level 14
assign po0902 = ~w16067;// level 14
assign po0903 = w16100;// level 14
assign po0904 = w16190;// level 14
assign po0905 = w16221;// level 14
assign po0906 = ~w16248;// level 14
assign po0907 = w16269;// level 14
assign po0908 = w16376;// level 14
assign po0909 = w16410;// level 14
assign po0910 = w16436;// level 14
assign po0911 = ~w16459;// level 14
assign po0912 = ~w16554;// level 14
assign po0913 = w16574;// level 14
assign po0914 = ~w16602;// level 14
assign po0915 = ~w16622;// level 14
assign po0916 = w16645;// level 14
assign po0917 = w16675;// level 14
assign po0918 = ~w16696;// level 14
assign po0919 = w16767;// level 14
assign po0920 = w16792;// level 14
assign po0921 = ~w16805;// level 14
assign po0922 = w16842;// level 14
assign po0923 = w16864;// level 14
assign po0924 = w16888;// level 14
assign po0925 = w16902;// level 14
assign po0926 = w16927;// level 14
assign po0927 = w16954;// level 14
assign po0928 = w16970;// level 14
assign po0929 = w16994;// level 14
assign po0930 = pi0819;// level 0
assign po0931 = pi0826;// level 0
assign po0932 = pi0828;// level 0
assign po0933 = pi0842;// level 0
assign po0934 = pi0835;// level 0
assign po0935 = pi0834;// level 0
assign po0936 = pi0840;// level 0
assign po0937 = pi0848;// level 0
assign po0938 = pi0836;// level 0
assign po0939 = pi0837;// level 0
assign po0940 = pi0845;// level 0
assign po0941 = pi0838;// level 0
assign po0942 = pi0839;// level 0
assign po0943 = pi0841;// level 0
assign po0944 = pi0843;// level 0
assign po0945 = pi0844;// level 0
assign po0946 = pi0858;// level 0
assign po0947 = pi0861;// level 0
assign po0948 = pi0847;// level 0
assign po0949 = ~w17083;// level 14
assign po0950 = pi0849;// level 0
assign po0951 = pi0850;// level 0
assign po0952 = pi0851;// level 0
assign po0953 = pi0852;// level 0
assign po0954 = pi0853;// level 0
assign po0955 = pi0854;// level 0
assign po0956 = w17183;// level 14
assign po0957 = pi0855;// level 0
assign po0958 = ~w17207;// level 14
assign po0959 = pi0863;// level 0
assign po0960 = pi0856;// level 0
assign po0961 = pi0857;// level 0
assign po0962 = pi0859;// level 0
assign po0963 = pi0860;// level 0
assign po0964 = w17291;// level 14
assign po0965 = w17377;// level 14
assign po0966 = w17396;// level 14
assign po0967 = w17489;// level 14
assign po0968 = w17584;// level 14
assign po0969 = ~w17602;// level 14
assign po0970 = ~w17701;// level 14
assign po0971 = w17737;// level 14
assign po0972 = w17762;// level 14
assign po0973 = ~w17793;// level 14
assign po0974 = w17818;// level 14
assign po0975 = ~w17840;// level 14
assign po0976 = pi0862;// level 0
assign po0977 = ~w17863;// level 14
assign po0978 = ~w17887;// level 14
assign po0979 = ~w17914;// level 14
assign po0980 = w17927;// level 14
assign po0981 = w17971;// level 14
assign po0982 = w17993;// level 14
assign po0983 = w18025;// level 14
assign po0984 = ~w18107;// level 14
assign po0985 = w18127;// level 14
assign po0986 = w18146;// level 14
assign po0987 = ~w18179;// level 14
assign po0988 = w18202;// level 14
assign po0989 = w18218;// level 14
assign po0990 = w18240;// level 14
assign po0991 = w18259;// level 14
assign po0992 = w18278;// level 14
assign po0993 = ~w18303;// level 14
assign po0994 = pi0891;// level 0
assign po0995 = pi0905;// level 0
assign po0996 = pi0890;// level 0
assign po0997 = pi0893;// level 0
assign po0998 = pi0904;// level 0
assign po0999 = pi0895;// level 0
assign po1000 = pi0897;// level 0
assign po1001 = pi0896;// level 0
assign po1002 = pi0899;// level 0
assign po1003 = pi0901;// level 0
assign po1004 = pi0898;// level 0
assign po1005 = pi0909;// level 0
assign po1006 = pi0916;// level 0
assign po1007 = pi0918;// level 0
assign po1008 = pi0903;// level 0
assign po1009 = pi0920;// level 0
assign po1010 = pi0906;// level 0
assign po1011 = pi0907;// level 0
assign po1012 = pi0910;// level 0
assign po1013 = pi0911;// level 0
assign po1014 = pi0912;// level 0
assign po1015 = pi0914;// level 0
assign po1016 = pi0915;// level 0
assign po1017 = pi0917;// level 0
assign po1018 = pi0921;// level 0
assign po1019 = pi0922;// level 0
assign po1020 = ~w18392;// level 14
assign po1021 = w18484;// level 14
assign po1022 = pi0923;// level 0
assign po1023 = ~w18587;// level 14
assign po1024 = pi0924;// level 0
assign po1025 = w18679;// level 14
assign po1026 = ~w18696;// level 14
assign po1027 = w18726;// level 14
assign po1028 = ~w18819;// level 14
assign po1029 = w18904;// level 14
assign po1030 = pi0925;// level 0
assign po1031 = w18931;// level 14
assign po1032 = pi0919;// level 0
assign po1033 = ~w18958;// level 14
assign po1034 = w18993;// level 14
assign po1035 = w19020;// level 14
assign po1036 = ~w19051;// level 14
assign po1037 = ~w19079;// level 14
assign po1038 = pi0926;// level 0
assign po1039 = w19099;// level 14
assign po1040 = ~w19124;// level 14
assign po1041 = ~w19205;// level 14
assign po1042 = w19293;// level 14
assign po1043 = pi0927;// level 0
assign po1044 = ~w19315;// level 14
assign po1045 = w19339;// level 14
assign po1046 = w19366;// level 14
assign po1047 = w19386;// level 14
assign po1048 = w19398;// level 14
assign po1049 = w19417;// level 14
assign po1050 = ~w19447;// level 14
assign po1051 = w19470;// level 14
assign po1052 = ~w19505;// level 14
assign po1053 = w19528;// level 14
assign po1054 = w19554;// level 14
assign po1055 = w19579;// level 14
assign po1056 = ~w19601;// level 14
assign po1057 = ~w19622;// level 14
assign po1058 = pi0945;// level 0
assign po1059 = pi0967;// level 0
assign po1060 = pi0953;// level 0
assign po1061 = pi0954;// level 0
assign po1062 = pi0961;// level 0
assign po1063 = pi0968;// level 0
assign po1064 = pi0958;// level 0
assign po1065 = pi0962;// level 0
assign po1066 = pi0963;// level 0
assign po1067 = pi0972;// level 0
assign po1068 = pi0977;// level 0
assign po1069 = pi0964;// level 0
assign po1070 = pi0969;// level 0
assign po1071 = pi0970;// level 0
assign po1072 = pi0971;// level 0
assign po1073 = pi0973;// level 0
assign po1074 = pi0985;// level 0
assign po1075 = ~w19714;// level 14
assign po1076 = pi0979;// level 0
assign po1077 = pi0974;// level 0
assign po1078 = pi0975;// level 0
assign po1079 = pi0976;// level 0
assign po1080 = pi0978;// level 0
assign po1081 = pi0988;// level 0
assign po1082 = pi0981;// level 0
assign po1083 = w19815;// level 14
assign po1084 = w19920;// level 14
assign po1085 = pi0982;// level 0
assign po1086 = pi0983;// level 0
assign po1087 = pi0984;// level 0
assign po1088 = ~w20011;// level 14
assign po1089 = pi0986;// level 0
assign po1090 = pi0987;// level 0
assign po1091 = ~w20038;// level 14
assign po1092 = ~w20063;// level 14
assign po1093 = ~w20085;// level 14
assign po1094 = ~w20104;// level 14
assign po1095 = pi0989;// level 0
assign po1096 = pi0990;// level 0
assign po1097 = ~w20123;// level 14
assign po1098 = ~w20145;// level 13
assign po1099 = w20176;// level 14
assign po1100 = ~w20255;// level 14
assign po1101 = w20283;// level 14
assign po1102 = w20370;// level 14
assign po1103 = ~w20403;// level 14
assign po1104 = ~w20436;// level 14
assign po1105 = w20456;// level 14
assign po1106 = ~w20492;// level 14
assign po1107 = w20513;// level 14
assign po1108 = ~w20525;// level 14
assign po1109 = ~w20610;// level 14
assign po1110 = pi0991;// level 0
assign po1111 = w20632;// level 14
assign po1112 = w20661;// level 14
assign po1113 = w20690;// level 14
assign po1114 = ~w20717;// level 14
assign po1115 = w20743;// level 14
assign po1116 = w20825;// level 14
assign po1117 = w20846;// level 14
assign po1118 = w20882;// level 14
assign po1119 = ~w20898;// level 14
assign po1120 = ~w20918;// level 14
assign po1121 = w20938;// level 13
assign po1122 = pi0995;// level 0
assign po1123 = pi0999;// level 0
assign po1124 = pi1003;// level 0
assign po1125 = ~w21032;// level 14
assign po1126 = pi1198;// level 0
assign po1127 = w21032;// level 14
assign po1128 = pi1009;// level 0
assign po1129 = pi1013;// level 0
assign po1130 = pi1015;// level 0
assign po1131 = pi1203;// level 0
assign po1132 = w21121;// level 14
assign po1133 = ~pi1203;// level 0
assign po1134 = pi1016;// level 0
assign po1135 = pi1023;// level 0
assign po1136 = pi1022;// level 0
assign po1137 = pi1189;// level 0
assign po1138 = ~w21209;// level 13
assign po1139 = ~pi1189;// level 0
assign po1140 = pi1026;// level 0
assign po1141 = pi1031;// level 0
assign po1142 = pi1028;// level 0
assign po1143 = pi1029;// level 0
assign po1144 = pi1030;// level 0
assign po1145 = pi1195;// level 0
assign po1146 = w21231;// level 14
assign po1147 = ~pi1195;// level 0
assign po1148 = pi1032;// level 0
assign po1149 = pi1034;// level 0
assign po1150 = pi1033;// level 0
assign po1151 = w21253;// level 14
assign po1152 = pi1038;// level 0
assign po1153 = pi1197;// level 0
assign po1154 = ~w21263;// level 13
assign po1155 = ~pi1197;// level 0
assign po1156 = pi1204;// level 0
assign po1157 = ~w21373;// level 14
assign po1158 = ~pi1204;// level 0
assign po1159 = pi1043;// level 0
assign po1160 = pi1045;// level 0
assign po1161 = pi1041;// level 0
assign po1162 = pi1042;// level 0
assign po1163 = pi1044;// level 0
assign po1164 = w21408;// level 13
assign po1165 = pi1215;// level 0
assign po1166 = ~w21408;// level 13
assign po1167 = ~w21435;// level 14
assign po1168 = pi1047;// level 0
assign po1169 = pi1048;// level 0
assign po1170 = pi1185;// level 0
assign po1171 = w21528;// level 12
assign po1172 = ~pi1185;// level 0
assign po1173 = pi1049;// level 0
assign po1174 = pi1191;// level 0
assign po1175 = ~w21547;// level 13
assign po1176 = ~pi1191;// level 0
assign po1177 = pi1187;// level 0
assign po1178 = ~w21627;// level 14
assign po1179 = ~pi1187;// level 0
assign po1180 = pi1188;// level 0
assign po1181 = ~w21638;// level 14
assign po1182 = ~pi1188;// level 0
assign po1183 = pi1194;// level 0
assign po1184 = ~w21661;// level 14
assign po1185 = ~pi1194;// level 0
assign po1186 = pi1190;// level 0
assign po1187 = w21688;// level 13
assign po1188 = ~pi1190;// level 0
assign po1189 = pi1211;// level 0
assign po1190 = w21709;// level 14
assign po1191 = ~pi1211;// level 0
assign po1192 = pi1218;// level 0
assign po1193 = ~w21728;// level 14
assign po1194 = ~pi1218;// level 0
assign po1195 = pi1052;// level 0
assign po1196 = pi1051;// level 0
assign po1197 = pi1050;// level 0
assign po1198 = pi1228;// level 0
assign po1199 = ~w21746;// level 13
assign po1200 = ~pi1228;// level 0
assign po1201 = pi1053;// level 0
assign po1202 = pi1054;// level 0
assign po1203 = pi1207;// level 0
assign po1204 = ~w21826;// level 13
assign po1205 = ~pi1207;// level 0
assign po1206 = pi1199;// level 0
assign po1207 = ~w21854;// level 13
assign po1208 = ~pi1199;// level 0
assign po1209 = pi1186;// level 0
assign po1210 = ~w21882;// level 13
assign po1211 = ~pi1186;// level 0
assign po1212 = pi1196;// level 0
assign po1213 = w21906;// level 13
assign po1214 = ~pi1196;// level 0
assign po1215 = pi1205;// level 0
assign po1216 = ~w21940;// level 14
assign po1217 = ~pi1205;// level 0
assign po1218 = pi1055;// level 0
assign po1219 = pi1201;// level 0
assign po1220 = ~w22019;// level 13
assign po1221 = ~pi1201;// level 0
assign po1222 = pi1233;// level 0
assign po1223 = ~w22039;// level 12
assign po1224 = ~pi1233;// level 0
assign po1225 = pi1184;// level 0
assign po1226 = w22068;// level 14
assign po1227 = ~pi1184;// level 0
assign po1228 = w22100;// level 14
assign po1229 = pi1202;// level 0
assign po1230 = ~w22126;// level 14
assign po1231 = ~pi1202;// level 0
assign po1232 = pi1192;// level 0
assign po1233 = ~w22141;// level 14
assign po1234 = ~pi1192;// level 0
assign po1235 = ~w22162;// level 14
assign po1236 = pi1193;// level 0
assign po1237 = ~w22176;// level 14
assign po1238 = ~pi1193;// level 0
assign po1239 = pi1212;// level 0
assign po1240 = ~w22191;// level 14
assign po1241 = ~pi1212;// level 0
assign po1242 = pi1082;// level 0
assign po1243 = pi1080;// level 0
assign po1244 = pi1089;// level 0
assign po1245 = pi1074;// level 0
assign po1246 = pi1073;// level 0
assign po1247 = pi1083;// level 0
assign po1248 = pi1092;// level 0
assign po1249 = pi1099;// level 0
assign po1250 = pi1110;// level 0
assign po1251 = pi1094;// level 0
assign po1252 = pi1095;// level 0
assign po1253 = pi1098;// level 0
assign po1254 = pi1102;// level 0
assign po1255 = pi1122;// level 0
assign po1256 = pi1103;// level 0
assign po1257 = pi1104;// level 0
assign po1258 = pi1105;// level 0
assign po1259 = pi1090;// level 0
assign po1260 = pi1091;// level 0
assign po1261 = pi1109;// level 0
assign po1262 = pi1111;// level 0
assign po1263 = pi1114;// level 0
assign po1264 = pi1115;// level 0
assign po1265 = pi1116;// level 0
assign po1266 = pi1097;// level 0
assign po1267 = pi1117;// level 0
assign po1268 = pi1101;// level 0
assign po1269 = pi1100;// level 0
assign po1270 = pi1120;// level 0
assign po1271 = pi1121;// level 0
assign po1272 = pi1127;// level 0
assign po1273 = pi1128;// level 0
assign po1274 = pi1129;// level 0
assign po1275 = pi1106;// level 0
assign po1276 = pi1130;// level 0
assign po1277 = pi1131;// level 0
assign po1278 = pi1108;// level 0
assign po1279 = pi1133;// level 0
assign po1280 = pi1112;// level 0
assign po1281 = pi1113;// level 0
assign po1282 = pi1136;// level 0
assign po1283 = pi1155;// level 0
assign po1284 = pi1118;// level 0
assign po1285 = pi1119;// level 0
assign po1286 = pi1161;// level 0
assign po1287 = pi1159;// level 0
assign po1288 = pi1123;// level 0
assign po1289 = pi1124;// level 0
assign po1290 = pi1125;// level 0
assign po1291 = pi1126;// level 0
assign po1292 = pi1146;// level 0
assign po1293 = pi1150;// level 0
assign po1294 = pi1151;// level 0
assign po1295 = pi1132;// level 0
assign po1296 = pi1134;// level 0
assign po1297 = pi1135;// level 0
assign po1298 = ~pi1145;// level 0
assign po1299 = pi1173;// level 0
assign po1300 = pi1138;// level 0
assign po1301 = pi1137;// level 0
assign po1302 = pi1139;// level 0
assign po1303 = pi1140;// level 0
assign po1304 = pi1169;// level 0
assign po1305 = pi1158;// level 0
assign po1306 = pi1142;// level 0
assign po1307 = pi1143;// level 0
assign po1308 = pi1144;// level 0
assign po1309 = pi1177;// level 0
assign po1310 = pi1166;// level 0
assign po1311 = ~pi1153;// level 0
assign po1312 = pi1167;// level 0
assign po1313 = pi1147;// level 0
assign po1314 = pi1148;// level 0
assign po1315 = pi1149;// level 0
assign po1316 = w22276;// level 14
assign po1317 = ~w22371;// level 14
assign po1318 = ~pi1163;// level 0
assign po1319 = pi1152;// level 0
assign po1320 = pi1171;// level 0
assign po1321 = pi1154;// level 0
assign po1322 = pi1156;// level 0
assign po1323 = pi1157;// level 0
assign po1324 = pi1176;// level 0
assign po1325 = pi1175;// level 0
assign po1326 = pi1160;// level 0
assign po1327 = pi1162;// level 0
assign po1328 = pi1164;// level 0
assign po1329 = pi1165;// level 0
assign po1330 = pi1178;// level 0
assign po1331 = w22402;// level 14
assign po1332 = w22436;// level 14
assign po1333 = pi1168;// level 0
assign po1334 = pi1180;// level 0
assign po1335 = ~pi1174;// level 0
assign po1336 = pi1170;// level 0
assign po1337 = ~w22527;// level 14
assign po1338 = pi1172;// level 0
assign po1339 = ~w22622;// level 14
assign po1340 = w22710;// level 14
assign po1341 = w22807;// level 14
assign po1342 = ~pi1181;// level 0
assign po1343 = w22826;// level 14
assign po1344 = w22850;// level 14
assign po1345 = ~w22880;// level 14
assign po1346 = w22913;// level 14
assign po1347 = w22993;// level 14
assign po1348 = pi1179;// level 0
assign po1349 = w23021;// level 14
assign po1350 = w23103;// level 14
assign po1351 = ~w23125;// level 14
assign po1352 = ~w23159;// level 14
assign po1353 = ~w23197;// level 14
assign po1354 = ~w23222;// level 14
assign po1355 = w23252;// level 14
assign po1356 = pi1182;// level 0
assign po1357 = w23273;// level 14
assign po1358 = ~w23290;// level 14
assign po1359 = ~w23315;// level 14
assign po1360 = w23336;// level 14
assign po1361 = w23359;// level 14
assign po1362 = ~w23392;// level 14
assign po1363 = w23414;// level 14
assign po1364 = ~w23433;// level 14
assign po1365 = pi1183;// level 0
assign po1366 = ~w23456;// level 14
assign po1367 = w23479;// level 14
assign po1368 = w23500;// level 14
assign po1369 = ~w23524;// level 14
assign po1370 = pi1200;// level 0
assign po1371 = pi1206;// level 0
assign po1372 = pi1208;// level 0
assign po1373 = pi1209;// level 0
assign po1374 = pi1210;// level 0
assign po1375 = pi1216;// level 0
assign po1376 = pi1219;// level 0
assign po1377 = pi1220;// level 0
assign po1378 = pi1235;// level 0
assign po1379 = pi1226;// level 0
assign po1380 = pi1224;// level 0
assign po1381 = pi1225;// level 0
assign po1382 = pi1229;// level 0
assign po1383 = pi1230;// level 0
assign po1384 = pi1214;// level 0
assign po1385 = pi1217;// level 0
assign po1386 = w23619;// level 14
assign po1387 = pi1234;// level 0
assign po1388 = pi1236;// level 0
assign po1389 = pi1222;// level 0
assign po1390 = pi1223;// level 0
assign po1391 = pi1238;// level 0
assign po1392 = w23650;// level 14
assign po1393 = pi1239;// level 0
assign po1394 = w23673;// level 14
assign po1395 = ~w23749;// level 14
assign po1396 = w23842;// level 14
assign po1397 = pi1242;// level 0
assign po1398 = pi1243;// level 0
assign po1399 = pi1231;// level 0
assign po1400 = w23935;// level 14
assign po1401 = pi1245;// level 0
assign po1402 = w24024;// level 14
assign po1403 = w24061;// level 14
assign po1404 = pi1246;// level 0
assign po1405 = ~w24088;// level 14
assign po1406 = w24113;// level 14
assign po1407 = pi1237;// level 0
assign po1408 = w24200;// level 14
assign po1409 = ~w24227;// level 14
assign po1410 = w24245;// level 14
assign po1411 = ~w24270;// level 14
assign po1412 = w24293;// level 14
assign po1413 = pi1240;// level 0
assign po1414 = pi1241;// level 0
assign po1415 = w24319;// level 14
assign po1416 = ~w24342;// level 14
assign po1417 = w24359;// level 14
assign po1418 = pi1244;// level 0
assign po1419 = pi1247;// level 0
assign po1420 = w24431;// level 14
assign po1421 = w24460;// level 14
assign po1422 = w24481;// level 14
assign po1423 = w24504;// level 14
assign po1424 = ~w24586;// level 14
assign po1425 = w24623;// level 14
assign po1426 = ~w24644;// level 14
assign po1427 = w24670;// level 14
assign po1428 = w24696;// level 14
assign po1429 = ~w24723;// level 14
assign po1430 = w24746;// level 14
assign po1431 = w24775;// level 14
assign po1432 = w24797;// level 14
assign po1433 = w24822;// level 14
assign po1434 = pi1259;// level 0
assign po1435 = pi1271;// level 0
assign po1436 = pi1268;// level 0
assign po1437 = pi1279;// level 0
assign po1438 = pi1291;// level 0
assign po1439 = pi1275;// level 0
assign po1440 = pi1287;// level 0
assign po1441 = pi1281;// level 0
assign po1442 = pi1280;// level 0
assign po1443 = pi1299;// level 0
assign po1444 = pi1289;// level 0
assign po1445 = w24915;// level 14
assign po1446 = pi1294;// level 0
assign po1447 = pi1277;// level 0
assign po1448 = pi1295;// level 0
assign po1449 = pi1296;// level 0
assign po1450 = pi1298;// level 0
assign po1451 = pi1297;// level 0
assign po1452 = pi1290;// level 0
assign po1453 = pi1300;// level 0
assign po1454 = w25004;// level 14
assign po1455 = pi1302;// level 0
assign po1456 = pi1288;// level 0
assign po1457 = w25030;// level 14
assign po1458 = pi1293;// level 0
assign po1459 = pi1304;// level 0
assign po1460 = pi1305;// level 0
assign po1461 = ~w25124;// level 14
assign po1462 = pi1306;// level 0
assign po1463 = w25221;// level 14
assign po1464 = pi1307;// level 0
assign po1465 = ~w25312;// level 14
assign po1466 = w25407;// level 14
assign po1467 = w25447;// level 14
assign po1468 = pi1308;// level 0
assign po1469 = pi1309;// level 0
assign po1470 = pi1310;// level 0
assign po1471 = pi1301;// level 0
assign po1472 = pi1303;// level 0
assign po1473 = ~w25479;// level 14
assign po1474 = w25504;// level 14
assign po1475 = w25530;// level 14
assign po1476 = ~w25614;// level 14
assign po1477 = w25636;// level 14
assign po1478 = pi1311;// level 0
assign po1479 = ~w25657;// level 14
assign po1480 = ~w25682;// level 14
assign po1481 = ~w25714;// level 14
assign po1482 = w25740;// level 14
assign po1483 = ~w25768;// level 14
assign po1484 = w25787;// level 14
assign po1485 = w25814;// level 14
assign po1486 = ~w25910;// level 14
assign po1487 = ~w25930;// level 14
assign po1488 = ~w25954;// level 14
assign po1489 = ~w25979;// level 14
assign po1490 = w25998;// level 14
assign po1491 = ~w26019;// level 14
assign po1492 = ~w26038;// level 14
assign po1493 = ~w26064;// level 14
assign po1494 = w26087;// level 14
assign po1495 = w26107;// level 14
assign po1496 = ~w26125;// level 14
assign po1497 = w26146;// level 14
assign po1498 = pi1335;// level 0
assign po1499 = pi1334;// level 0
assign po1500 = pi1339;// level 0
assign po1501 = pi1352;// level 0
assign po1502 = pi1341;// level 0
assign po1503 = pi1350;// level 0
assign po1504 = pi1345;// level 0
assign po1505 = pi1346;// level 0
assign po1506 = pi1351;// level 0
assign po1507 = pi1353;// level 0
assign po1508 = pi1355;// level 0
assign po1509 = pi1356;// level 0
assign po1510 = pi1371;// level 0
assign po1511 = pi1357;// level 0
assign po1512 = pi1372;// level 0
assign po1513 = pi1343;// level 0
assign po1514 = pi1358;// level 0
assign po1515 = pi1360;// level 0
assign po1516 = pi1359;// level 0
assign po1517 = pi1362;// level 0
assign po1518 = pi1363;// level 0
assign po1519 = pi1364;// level 0
assign po1520 = ~w26236;// level 14
assign po1521 = w26339;// level 14
assign po1522 = pi1365;// level 0
assign po1523 = pi1367;// level 0
assign po1524 = pi1368;// level 0
assign po1525 = ~w26433;// level 14
assign po1526 = pi1369;// level 0
assign po1527 = ~w26527;// level 14
assign po1528 = pi1373;// level 0
assign po1529 = w26557;// level 14
assign po1530 = pi1361;// level 0
assign po1531 = w26647;// level 14
assign po1532 = w26725;// level 14
assign po1533 = pi1374;// level 0
assign po1534 = pi1375;// level 0
assign po1535 = pi1366;// level 0
assign po1536 = w26754;// level 14
assign po1537 = ~w26776;// level 14
assign po1538 = w26802;// level 14
assign po1539 = ~w26824;// level 14
assign po1540 = pi1370;// level 0
assign po1541 = w26865;// level 14
assign po1542 = ~w26885;// level 14
assign po1543 = w26979;// level 14
assign po1544 = w27005;// level 14
assign po1545 = w27088;// level 14
assign po1546 = w27100;// level 14
assign po1547 = ~w27125;// level 14
assign po1548 = ~w27149;// level 14
assign po1549 = ~w27180;// level 14
assign po1550 = ~w27195;// level 14
assign po1551 = w27220;// level 14
assign po1552 = w27251;// level 14
assign po1553 = ~w27275;// level 14
assign po1554 = w27297;// level 14
assign po1555 = ~w27319;// level 14
assign po1556 = ~w27341;// level 14
assign po1557 = ~w27366;// level 14
assign po1558 = w27389;// level 14
assign po1559 = ~w27411;// level 14
assign po1560 = ~w27437;// level 14
assign po1561 = ~w27453;// level 14
assign po1562 = pi1395;// level 0
assign po1563 = pi1400;// level 0
assign po1564 = pi1404;// level 0
assign po1565 = pi1415;// level 0
assign po1566 = pi1420;// level 0
assign po1567 = pi1406;// level 0
assign po1568 = pi1410;// level 0
assign po1569 = pi1411;// level 0
assign po1570 = pi1413;// level 0
assign po1571 = pi1412;// level 0
assign po1572 = pi1414;// level 0
assign po1573 = pi1416;// level 0
assign po1574 = pi1426;// level 0
assign po1575 = pi1418;// level 0
assign po1576 = pi1419;// level 0
assign po1577 = pi1421;// level 0
assign po1578 = pi1405;// level 0
assign po1579 = pi1422;// level 0
assign po1580 = pi1423;// level 0
assign po1581 = w27556;// level 14
assign po1582 = pi1424;// level 0
assign po1583 = pi1433;// level 0
assign po1584 = pi1427;// level 0
assign po1585 = pi1428;// level 0
assign po1586 = ~w27640;// level 14
assign po1587 = pi1429;// level 0
assign po1588 = pi1431;// level 0
assign po1589 = pi1432;// level 0
assign po1590 = ~w27664;// level 14
assign po1591 = w27684;// level 14
assign po1592 = w27771;// level 14
assign po1593 = pi1434;// level 0
assign po1594 = pi1435;// level 0
assign po1595 = pi1436;// level 0
assign po1596 = w27864;// level 14
assign po1597 = ~w27961;// level 14
assign po1598 = w27983;// level 14
assign po1599 = ~w28072;// level 14
assign po1600 = w28101;// level 14
assign po1601 = ~w28128;// level 14
assign po1602 = ~w28158;// level 14
assign po1603 = pi1430;// level 0
assign po1604 = ~w28182;// level 14
assign po1605 = ~w28275;// level 14
assign po1606 = ~w28297;// level 14
assign po1607 = w28318;// level 14
assign po1608 = ~w28342;// level 14
assign po1609 = w28369;// level 14
assign po1610 = ~w28389;// level 14
assign po1611 = pi1438;// level 0
assign po1612 = ~w28404;// level 14
assign po1613 = ~w28494;// level 14
assign po1614 = ~w28524;// level 14
assign po1615 = w28544;// level 14
assign po1616 = w28577;// level 14
assign po1617 = ~w28595;// level 14
assign po1618 = w28625;// level 14
assign po1619 = w28652;// level 14
assign po1620 = w28674;// level 14
assign po1621 = w28698;// level 14
assign po1622 = w28716;// level 14
assign po1623 = pi1439;// level 0
assign po1624 = w28733;// level 14
assign po1625 = w28751;// level 14
assign po1626 = pi1473;// level 0
assign po1627 = pi1464;// level 0
assign po1628 = pi1463;// level 0
assign po1629 = pi1467;// level 0
assign po1630 = pi1470;// level 0
assign po1631 = pi1469;// level 0
assign po1632 = pi1476;// level 0
assign po1633 = pi1480;// level 0
assign po1634 = pi1482;// level 0
assign po1635 = pi1475;// level 0
assign po1636 = pi1477;// level 0
assign po1637 = pi1478;// level 0
assign po1638 = pi1481;// level 0
assign po1639 = pi1483;// level 0
assign po1640 = pi1484;// level 0
assign po1641 = pi1485;// level 0
assign po1642 = pi1486;// level 0
assign po1643 = pi1487;// level 0
assign po1644 = pi1488;// level 0
assign po1645 = pi1489;// level 0
assign po1646 = pi1497;// level 0
assign po1647 = pi1490;// level 0
assign po1648 = pi1491;// level 0
assign po1649 = w28843;// level 14
assign po1650 = w28932;// level 14
assign po1651 = pi1493;// level 0
assign po1652 = pi1494;// level 0
assign po1653 = w29024;// level 14
assign po1654 = pi1495;// level 0
assign po1655 = ~w29115;// level 14
assign po1656 = w29202;// level 14
assign po1657 = pi1499;// level 0
assign po1658 = pi1500;// level 0
assign po1659 = ~w29230;// level 14
assign po1660 = pi1501;// level 0
assign po1661 = ~w29324;// level 14
assign po1662 = w29362;// level 14
assign po1663 = ~w29388;// level 14
assign po1664 = ~w29415;// level 14
assign po1665 = pi1496;// level 0
assign po1666 = w29502;// level 14
assign po1667 = w29533;// level 14
assign po1668 = w29562;// level 14
assign po1669 = w29638;// level 14
assign po1670 = ~w29682;// level 14
assign po1671 = ~w29700;// level 14
assign po1672 = w29727;// level 14
assign po1673 = w29744;// level 14
assign po1674 = w29782;// level 14
assign po1675 = w29808;// level 14
assign po1676 = ~w29825;// level 14
assign po1677 = ~w29840;// level 14
assign po1678 = pi1502;// level 0
assign po1679 = ~w29877;// level 14
assign po1680 = w29901;// level 14
assign po1681 = w29921;// level 14
assign po1682 = ~w29944;// level 14
assign po1683 = w29969;// level 14
assign po1684 = pi1503;// level 0
assign po1685 = ~w29988;// level 14
assign po1686 = ~w30013;// level 14
assign po1687 = w30035;// level 14
assign po1688 = w30050;// level 14
assign po1689 = ~w30070;// level 14
assign po1690 = pi1524;// level 0
assign po1691 = pi1528;// level 0
assign po1692 = pi1529;// level 0
assign po1693 = pi1545;// level 0
assign po1694 = pi1534;// level 0
assign po1695 = pi1535;// level 0
assign po1696 = pi1536;// level 0
assign po1697 = pi1538;// level 0
assign po1698 = pi1539;// level 0
assign po1699 = pi1544;// level 0
assign po1700 = pi1546;// level 0
assign po1701 = pi1548;// level 0
assign po1702 = pi1541;// level 0
assign po1703 = pi1551;// level 0
assign po1704 = pi1542;// level 0
assign po1705 = pi1547;// level 0
assign po1706 = pi1550;// level 0
assign po1707 = pi1549;// level 0
assign po1708 = pi1552;// level 0
assign po1709 = pi1565;// level 0
assign po1710 = ~w30168;// level 14
assign po1711 = pi1554;// level 0
assign po1712 = pi1555;// level 0
assign po1713 = pi1556;// level 0
assign po1714 = ~w30198;// level 14
assign po1715 = ~w30298;// level 14
assign po1716 = pi1564;// level 0
assign po1717 = pi1559;// level 0
assign po1718 = pi1561;// level 0
assign po1719 = pi1560;// level 0
assign po1720 = w30393;// level 14
assign po1721 = w30484;// level 14
assign po1722 = ~w30509;// level 14
assign po1723 = pi1562;// level 0
assign po1724 = w30529;// level 14
assign po1725 = w30620;// level 14
assign po1726 = pi1563;// level 0
assign po1727 = ~w30644;// level 14
assign po1728 = ~w30732;// level 14
assign po1729 = pi1558;// level 0
assign po1730 = w30770;// level 14
assign po1731 = ~w30785;// level 14
assign po1732 = ~w30815;// level 14
assign po1733 = w30901;// level 14
assign po1734 = ~w30925;// level 14
assign po1735 = w30958;// level 14
assign po1736 = w30976;// level 14
assign po1737 = w31008;// level 14
assign po1738 = ~w31026;// level 14
assign po1739 = pi1566;// level 0
assign po1740 = w31049;// level 14
assign po1741 = ~w31072;// level 15
assign po1742 = ~w31094;// level 14
assign po1743 = pi1567;// level 0
assign po1744 = w31116;// level 14
assign po1745 = w31202;// level 14
assign po1746 = w31229;// level 14
assign po1747 = w31245;// level 14
assign po1748 = ~w31266;// level 14
assign po1749 = w31286;// level 14
assign po1750 = w31306;// level 14
assign po1751 = w31332;// level 14
assign po1752 = ~w31350;// level 14
assign po1753 = ~w31373;// level 14
assign po1754 = pi1591;// level 0
assign po1755 = pi1600;// level 0
assign po1756 = pi1593;// level 0
assign po1757 = pi1598;// level 0
assign po1758 = pi1614;// level 0
assign po1759 = pi1599;// level 0
assign po1760 = pi1618;// level 0
assign po1761 = pi1603;// level 0
assign po1762 = pi1605;// level 0
assign po1763 = pi1608;// level 0
assign po1764 = pi1607;// level 0
assign po1765 = pi1609;// level 0
assign po1766 = pi1610;// level 0
assign po1767 = pi1611;// level 0
assign po1768 = pi1612;// level 0
assign po1769 = pi1615;// level 0
assign po1770 = pi1613;// level 0
assign po1771 = pi1622;// level 0
assign po1772 = pi1616;// level 0
assign po1773 = pi1617;// level 0
assign po1774 = pi1604;// level 0
assign po1775 = pi1620;// level 0
assign po1776 = pi1621;// level 0
assign po1777 = ~w31467;// level 14
assign po1778 = pi1623;// level 0
assign po1779 = w31558;// level 14
assign po1780 = pi1628;// level 0
assign po1781 = pi1626;// level 0
assign po1782 = pi1624;// level 0
assign po1783 = pi1627;// level 0
assign po1784 = w31646;// level 14
assign po1785 = w31739;// level 14
assign po1786 = ~w31821;// level 14
assign po1787 = pi1629;// level 0
assign po1788 = pi1630;// level 0
assign po1789 = w31914;// level 14
assign po1790 = w32005;// level 14
assign po1791 = ~w32029;// level 14
assign po1792 = pi1625;// level 0
assign po1793 = w32071;// level 14
assign po1794 = ~w32096;// level 14
assign po1795 = w32115;// level 14
assign po1796 = w32143;// level 14
assign po1797 = w32244;// level 14
assign po1798 = ~w32282;// level 14
assign po1799 = w32306;// level 14
assign po1800 = ~w32339;// level 14
assign po1801 = ~w32362;// level 14
assign po1802 = ~w32382;// level 14
assign po1803 = ~w32401;// level 14
assign po1804 = ~w32420;// level 14
assign po1805 = pi1631;// level 0
assign po1806 = w32436;// level 14
assign po1807 = w32467;// level 14
assign po1808 = w32493;// level 14
assign po1809 = ~w32515;// level 14
assign po1810 = w32536;// level 14
assign po1811 = w32562;// level 14
assign po1812 = ~w32581;// level 14
assign po1813 = w32602;// level 14
assign po1814 = ~w32624;// level 14
assign po1815 = w32645;// level 14
assign po1816 = w32665;// level 14
assign po1817 = w32686;// level 14
assign po1818 = pi1662;// level 0
assign po1819 = pi1672;// level 0
assign po1820 = pi1657;// level 0
assign po1821 = pi1652;// level 0
assign po1822 = pi1663;// level 0
assign po1823 = pi1664;// level 0
assign po1824 = pi1665;// level 0
assign po1825 = pi1667;// level 0
assign po1826 = pi1659;// level 0
assign po1827 = pi1661;// level 0
assign po1828 = pi1670;// level 0
assign po1829 = pi1677;// level 0
assign po1830 = pi1669;// level 0
assign po1831 = pi1676;// level 0
assign po1832 = pi1668;// level 0
assign po1833 = pi1678;// level 0
assign po1834 = pi1679;// level 0
assign po1835 = pi1690;// level 0
assign po1836 = pi1684;// level 0
assign po1837 = pi1685;// level 0
assign po1838 = ~w32776;// level 14
assign po1839 = pi1689;// level 0
assign po1840 = pi1687;// level 0
assign po1841 = pi1688;// level 0
assign po1842 = pi1675;// level 0
assign po1843 = ~w32867;// level 14
assign po1844 = pi1683;// level 0
assign po1845 = ~w32893;// level 14
assign po1846 = pi1680;// level 0
assign po1847 = w32988;// level 14
assign po1848 = w33075;// level 14
assign po1849 = ~w33112;// level 14
assign po1850 = w33137;// level 14
assign po1851 = w33161;// level 14
assign po1852 = pi1691;// level 0
assign po1853 = w33254;// level 14
assign po1854 = ~w33348;// level 14
assign po1855 = w33373;// level 15
assign po1856 = w33453;// level 14
assign po1857 = pi1686;// level 0
assign po1858 = ~w33474;// level 15
assign po1859 = pi1693;// level 0
assign po1860 = pi1694;// level 0
assign po1861 = ~w33514;// level 15
assign po1862 = w33554;// level 14
assign po1863 = w33583;// level 14
assign po1864 = ~w33611;// level 14
assign po1865 = ~w33640;// level 14
assign po1866 = w33654;// level 14
assign po1867 = pi1695;// level 0
assign po1868 = pi1692;// level 0
assign po1869 = w33674;// level 14
assign po1870 = w33695;// level 14
assign po1871 = w33729;// level 14
assign po1872 = ~w33753;// level 14
assign po1873 = w33769;// level 14
assign po1874 = ~w33791;// level 14
assign po1875 = w33814;// level 14
assign po1876 = w33898;// level 14
assign po1877 = ~w33919;// level 14
assign po1878 = ~w33937;// level 14
assign po1879 = ~w33970;// level 14
assign po1880 = ~w33992;// level 14
assign po1881 = w34014;// level 14
assign po1882 = pi1702;// level 0
assign po1883 = pi1709;// level 0
assign po1884 = pi1723;// level 0
assign po1885 = pi1724;// level 0
assign po1886 = pi1732;// level 0
assign po1887 = pi1725;// level 0
assign po1888 = ~w34107;// level 14
assign po1889 = pi1731;// level 0
assign po1890 = pi1734;// level 0
assign po1891 = pi1742;// level 0
assign po1892 = pi1736;// level 0
assign po1893 = pi1743;// level 0
assign po1894 = pi1738;// level 0
assign po1895 = w34198;// level 14
assign po1896 = pi1739;// level 0
assign po1897 = pi1744;// level 0
assign po1898 = pi1741;// level 0
assign po1899 = pi1728;// level 0
assign po1900 = pi1745;// level 0
assign po1901 = pi1746;// level 0
assign po1902 = pi1747;// level 0
assign po1903 = pi1748;// level 0
assign po1904 = pi1749;// level 0
assign po1905 = pi1755;// level 0
assign po1906 = pi1740;// level 0
assign po1907 = pi1750;// level 0
assign po1908 = pi1751;// level 0
assign po1909 = ~w34231;// level 14
assign po1910 = w34258;// level 14
assign po1911 = ~w34348;// level 14
assign po1912 = pi1752;// level 0
assign po1913 = pi1753;// level 0
assign po1914 = w34375;// level 14
assign po1915 = pi1754;// level 0
assign po1916 = pi1756;// level 0
assign po1917 = w34470;// level 14
assign po1918 = w34551;// level 14
assign po1919 = pi1757;// level 0
assign po1920 = ~w34585;// level 14
assign po1921 = pi1758;// level 0
assign po1922 = ~w34607;// level 14
assign po1923 = pi1759;// level 0
assign po1924 = ~w34704;// level 14
assign po1925 = ~w34729;// level 14
assign po1926 = w34753;// level 13
assign po1927 = w34846;// level 14
assign po1928 = w34867;// level 14
assign po1929 = w34897;// level 14
assign po1930 = w34939;// level 14
assign po1931 = ~w34966;// level 14
assign po1932 = ~w34990;// level 14
assign po1933 = ~w35027;// level 14
assign po1934 = w35049;// level 14
assign po1935 = ~w35071;// level 14
assign po1936 = ~w35090;// level 14
assign po1937 = w35115;// level 14
assign po1938 = w35194;// level 14
assign po1939 = w35226;// level 15
assign po1940 = w35253;// level 14
assign po1941 = w35272;// level 14
assign po1942 = w35289;// level 14
assign po1943 = ~w35311;// level 14
assign po1944 = ~w35332;// level 14
assign po1945 = w35353;// level 14
assign po1946 = pi1775;// level 0
assign po1947 = pi1785;// level 0
assign po1948 = pi1786;// level 0
assign po1949 = pi1787;// level 0
assign po1950 = pi1791;// level 0
assign po1951 = pi1792;// level 0
assign po1952 = pi1799;// level 0
assign po1953 = pi1794;// level 0
assign po1954 = pi1804;// level 0
assign po1955 = pi1812;// level 0
assign po1956 = pi1798;// level 0
assign po1957 = pi1800;// level 0
assign po1958 = pi1802;// level 0
assign po1959 = pi1801;// level 0
assign po1960 = pi1806;// level 0
assign po1961 = ~w35440;// level 14
assign po1962 = pi1803;// level 0
assign po1963 = pi1805;// level 0
assign po1964 = pi1807;// level 0
assign po1965 = pi1808;// level 0
assign po1966 = pi1809;// level 0
assign po1967 = pi1811;// level 0
assign po1968 = pi1813;// level 0
assign po1969 = pi1797;// level 0
assign po1970 = pi1815;// level 0
assign po1971 = w35529;// level 14
assign po1972 = ~w35561;// level 14
assign po1973 = ~w35653;// level 14
assign po1974 = pi1820;// level 0
assign po1975 = pi1816;// level 0
assign po1976 = pi1817;// level 0
assign po1977 = ~w35752;// level 14
assign po1978 = w35846;// level 14
assign po1979 = pi1818;// level 0
assign po1980 = w35872;// level 14
assign po1981 = pi1821;// level 0
assign po1982 = pi1822;// level 0
assign po1983 = ~w35898;// level 14
assign po1984 = ~w35918;// level 14
assign po1985 = w36011;// level 14
assign po1986 = ~w36105;// level 14
assign po1987 = ~w36136;// level 14
assign po1988 = w36165;// level 14
assign po1989 = w36192;// level 14
assign po1990 = w36218;// level 14
assign po1991 = w36298;// level 14
assign po1992 = ~w36321;// level 14
assign po1993 = ~w36340;// level 14
assign po1994 = ~w36370;// level 14
assign po1995 = w36394;// level 14
assign po1996 = pi1819;// level 0
assign po1997 = w36427;// level 14
assign po1998 = ~w36442;// level 14
assign po1999 = ~w36462;// level 14
assign po2000 = pi1823;// level 0
assign po2001 = ~w36484;// level 14
assign po2002 = ~w36507;// level 14
assign po2003 = ~w36532;// level 14
assign po2004 = w36567;// level 14
assign po2005 = w36594;// level 14
assign po2006 = ~w36612;// level 14
assign po2007 = w36639;// level 14
assign po2008 = ~w36657;// level 14
assign po2009 = w36681;// level 14
assign po2010 = pi1843;// level 0
assign po2011 = pi1849;// level 0
assign po2012 = pi1848;// level 0
assign po2013 = pi1855;// level 0
assign po2014 = pi1860;// level 0
assign po2015 = pi1857;// level 0
assign po2016 = pi1861;// level 0
assign po2017 = pi1856;// level 0
assign po2018 = pi1858;// level 0
assign po2019 = pi1874;// level 0
assign po2020 = pi1868;// level 0
assign po2021 = pi1862;// level 0
assign po2022 = pi1864;// level 0
assign po2023 = pi1866;// level 0
assign po2024 = pi1869;// level 0
assign po2025 = pi1854;// level 0
assign po2026 = pi1872;// level 0
assign po2027 = pi1871;// level 0
assign po2028 = pi1873;// level 0
assign po2029 = w36772;// level 14
assign po2030 = pi1875;// level 0
assign po2031 = pi1876;// level 0
assign po2032 = pi1877;// level 0
assign po2033 = pi1878;// level 0
assign po2034 = w36863;// level 14
assign po2035 = ~w36962;// level 14
assign po2036 = pi1879;// level 0
assign po2037 = pi1881;// level 0
assign po2038 = pi1882;// level 0
assign po2039 = pi1883;// level 0
assign po2040 = w37057;// level 14
assign po2041 = ~w37147;// level 14
assign po2042 = w37171;// level 14
assign po2043 = w37260;// level 14
assign po2044 = ~w37297;// level 14
assign po2045 = pi1885;// level 0
assign po2046 = ~w37332;// level 14
assign po2047 = w37428;// level 14
assign po2048 = w37459;// level 14
assign po2049 = pi1880;// level 0
assign po2050 = ~w37491;// level 14
assign po2051 = pi1886;// level 0
assign po2052 = ~w37510;// level 15
assign po2053 = pi1887;// level 0
assign po2054 = ~w37540;// level 14
assign po2055 = ~w37550;// level 14
assign po2056 = pi1884;// level 0
assign po2057 = ~w37567;// level 14
assign po2058 = ~w37589;// level 14
assign po2059 = w37611;// level 14
assign po2060 = w37633;// level 14
assign po2061 = ~w37656;// level 14
assign po2062 = w37673;// level 14
assign po2063 = ~w37686;// level 14
assign po2064 = w37707;// level 14
assign po2065 = w37752;// level 14
assign po2066 = w37770;// level 14
assign po2067 = w37796;// level 14
assign po2068 = ~w37880;// level 14
assign po2069 = ~w37899;// level 14
assign po2070 = ~w37913;// level 14
assign po2071 = ~w37950;// level 14
assign po2072 = ~w37971;// level 14
assign po2073 = ~w37988;// level 14
assign po2074 = pi1900;// level 0
assign po2075 = pi1906;// level 0
assign po2076 = pi1919;// level 0
assign po2077 = pi1920;// level 0
assign po2078 = pi1926;// level 0
assign po2079 = pi1922;// level 0
assign po2080 = pi1924;// level 0
assign po2081 = pi1923;// level 0
assign po2082 = pi1928;// level 0
assign po2083 = pi1925;// level 0
assign po2084 = pi1927;// level 0
assign po2085 = pi1929;// level 0
assign po2086 = ~w38078;// level 14
assign po2087 = pi1937;// level 0
assign po2088 = pi1932;// level 0
assign po2089 = pi1938;// level 0
assign po2090 = pi1934;// level 0
assign po2091 = pi1935;// level 0
assign po2092 = ~w38172;// level 14
assign po2093 = pi1936;// level 0
assign po2094 = pi1939;// level 0
assign po2095 = pi1940;// level 0
assign po2096 = pi1941;// level 0
assign po2097 = pi1942;// level 0
assign po2098 = pi1943;// level 0
assign po2099 = pi1944;// level 0
assign po2100 = pi1945;// level 0
assign po2101 = pi1933;// level 0
assign po2102 = pi1946;// level 0
assign po2103 = pi1947;// level 0
assign po2104 = pi1948;// level 0
assign po2105 = w38275;// level 14
assign po2106 = ~w38300;// level 14
assign po2107 = pi1949;// level 0
assign po2108 = w38330;// level 14
assign po2109 = ~w38415;// level 14
assign po2110 = w38516;// level 14
assign po2111 = w38603;// level 14
assign po2112 = w38632;// level 14
assign po2113 = w38657;// level 14
assign po2114 = w38744;// level 14
assign po2115 = ~w38762;// level 14
assign po2116 = pi1950;// level 0
assign po2117 = pi1951;// level 0
assign po2118 = ~w38796;// level 14
assign po2119 = ~w38822;// level 14
assign po2120 = ~w38837;// level 14
assign po2121 = ~w38862;// level 14
assign po2122 = w38879;// level 14
assign po2123 = w38908;// level 14
assign po2124 = ~w38934;// level 14
assign po2125 = ~w39017;// level 14
assign po2126 = ~w39042;// level 14
assign po2127 = w39082;// level 14
assign po2128 = ~w39107;// level 14
assign po2129 = w39131;// level 14
assign po2130 = w39158;// level 14
assign po2131 = w39179;// level 14
assign po2132 = w39199;// level 14
assign po2133 = ~w39215;// level 14
assign po2134 = ~w39236;// level 14
assign po2135 = ~w39253;// level 14
assign po2136 = w39278;// level 14
assign po2137 = w39298;// level 14
assign po2138 = pi1983;// level 0
assign po2139 = pi1978;// level 0
assign po2140 = pi1974;// level 0
assign po2141 = pi1990;// level 0
assign po2142 = pi1975;// level 0
assign po2143 = pi1972;// level 0
assign po2144 = pi1989;// level 0
assign po2145 = pi1982;// level 0
assign po2146 = pi1985;// level 0
assign po2147 = pi1991;// level 0
assign po2148 = pi1981;// level 0
assign po2149 = pi1997;// level 0
assign po2150 = pi1993;// level 0
assign po2151 = pi1992;// level 0
assign po2152 = pi2000;// level 0
assign po2153 = pi1999;// level 0
assign po2154 = pi2001;// level 0
assign po2155 = pi1998;// level 0
assign po2156 = pi2002;// level 0
assign po2157 = pi2005;// level 0
assign po2158 = w39390;// level 14
assign po2159 = pi2003;// level 0
assign po2160 = w39490;// level 14
assign po2161 = w39578;// level 14
assign po2162 = pi2013;// level 0
assign po2163 = pi2004;// level 0
assign po2164 = ~w39612;// level 14
assign po2165 = pi2006;// level 0
assign po2166 = pi2007;// level 0
assign po2167 = w39636;// level 14
assign po2168 = ~w39721;// level 14
assign po2169 = w39758;// level 14
assign po2170 = pi2010;// level 0
assign po2171 = w39855;// level 14
assign po2172 = pi2011;// level 0
assign po2173 = pi2012;// level 0
assign po2174 = pi2008;// level 0
assign po2175 = ~w39878;// level 14
assign po2176 = ~w39908;// level 14
assign po2177 = ~w39990;// level 14
assign po2178 = ~w40011;// level 14
assign po2179 = ~w40036;// level 14
assign po2180 = pi2015;// level 0
assign po2181 = pi2014;// level 0
assign po2182 = pi2009;// level 0
assign po2183 = ~w40060;// level 14
assign po2184 = w40098;// level 14
assign po2185 = w40176;// level 14
assign po2186 = w40217;// level 14
assign po2187 = w40241;// level 14
assign po2188 = ~w40262;// level 14
assign po2189 = w40278;// level 14
assign po2190 = ~w40358;// level 14
assign po2191 = ~w40383;// level 14
assign po2192 = ~w40411;// level 14
assign po2193 = w40435;// level 14
assign po2194 = ~w40462;// level 14
assign po2195 = w40482;// level 14
assign po2196 = w40501;// level 14
assign po2197 = w40523;// level 14
assign po2198 = w40547;// level 14
assign po2199 = w40568;// level 14
assign po2200 = w40587;// level 14
assign po2201 = w40604;// level 14
assign po2202 = pi2032;// level 0
assign po2203 = pi2043;// level 0
assign po2204 = pi2037;// level 0
assign po2205 = pi2036;// level 0
assign po2206 = pi2056;// level 0
assign po2207 = pi2045;// level 0
assign po2208 = pi2055;// level 0
assign po2209 = pi2049;// level 0
assign po2210 = pi2054;// level 0
assign po2211 = pi2052;// level 0
assign po2212 = pi2069;// level 0
assign po2213 = pi2058;// level 0
assign po2214 = pi2061;// level 0
assign po2215 = pi2059;// level 0
assign po2216 = pi2060;// level 0
assign po2217 = pi2065;// level 0
assign po2218 = w40700;// level 15
assign po2219 = pi2072;// level 0
assign po2220 = pi2074;// level 0
assign po2221 = pi2067;// level 0
assign po2222 = ~w40786;// level 14
assign po2223 = w40817;// level 14
assign po2224 = pi2066;// level 0
assign po2225 = pi2053;// level 0
assign po2226 = pi2073;// level 0
assign po2227 = pi2077;// level 0
assign po2228 = pi2068;// level 0
assign po2229 = w40907;// level 14
assign po2230 = pi2062;// level 0
assign po2231 = w40946;// level 14
assign po2232 = pi2064;// level 0
assign po2233 = pi2070;// level 0
assign po2234 = pi2075;// level 0
assign po2235 = w41038;// level 14
assign po2236 = pi2076;// level 0
assign po2237 = pi2078;// level 0
assign po2238 = w41059;// level 14
assign po2239 = ~w41100;// level 14
assign po2240 = w41128;// level 14
assign po2241 = w41215;// level 14
assign po2242 = w41238;// level 14
assign po2243 = pi2079;// level 0
assign po2244 = ~w41259;// level 14
assign po2245 = w41300;// level 14
assign po2246 = w41321;// level 14
assign po2247 = w41409;// level 14
assign po2248 = w41439;// level 14
assign po2249 = pi2071;// level 0
assign po2250 = ~w41461;// level 14
assign po2251 = ~w41490;// level 14
assign po2252 = ~w41587;// level 14
assign po2253 = ~w41606;// level 14
assign po2254 = ~w41694;// level 14
assign po2255 = w41722;// level 14
assign po2256 = ~w41743;// level 14
assign po2257 = w41768;// level 14
assign po2258 = ~w41792;// level 14
assign po2259 = ~w41820;// level 14
assign po2260 = ~w41837;// level 14
assign po2261 = ~w41856;// level 14
assign po2262 = ~w41878;// level 14
assign po2263 = w41907;// level 14
assign po2264 = ~w41928;// level 14
assign po2265 = ~w41947;// level 14
assign po2266 = pi2083;// level 0
assign po2267 = pi2089;// level 0
assign po2268 = pi2100;// level 0
assign po2269 = pi2303;// level 0
assign po2270 = w42042;// level 14
assign po2271 = ~pi2303;// level 0
assign po2272 = pi2102;// level 0
assign po2273 = pi2106;// level 0
assign po2274 = pi2107;// level 0
assign po2275 = pi2108;// level 0
assign po2276 = pi2109;// level 0
assign po2277 = pi2290;// level 0
assign po2278 = ~w42069;// level 12
assign po2279 = ~pi2290;// level 0
assign po2280 = pi2115;// level 0
assign po2281 = pi2114;// level 0
assign po2282 = pi2117;// level 0
assign po2283 = pi2110;// level 0
assign po2284 = pi2118;// level 0
assign po2285 = pi2120;// level 0
assign po2286 = pi2122;// level 0
assign po2287 = pi2111;// level 0
assign po2288 = pi2123;// level 0
assign po2289 = pi2124;// level 0
assign po2290 = pi2279;// level 0
assign po2291 = w42154;// level 14
assign po2292 = ~pi2279;// level 0
assign po2293 = pi2128;// level 0
assign po2294 = pi2302;// level 0
assign po2295 = ~w42246;// level 13
assign po2296 = ~pi2302;// level 0
assign po2297 = pi2132;// level 0
assign po2298 = pi2129;// level 0
assign po2299 = pi2133;// level 0
assign po2300 = pi2309;// level 0
assign po2301 = ~w42274;// level 13
assign po2302 = ~pi2309;// level 0
assign po2303 = pi2277;// level 0
assign po2304 = ~w42303;// level 12
assign po2305 = ~pi2277;// level 0
assign po2306 = pi2299;// level 0
assign po2307 = ~w42326;// level 14
assign po2308 = ~pi2299;// level 0
assign po2309 = w42347;// level 14
assign po2310 = ~w42434;// level 14
assign po2311 = pi2294;// level 0
assign po2312 = ~w42456;// level 14
assign po2313 = ~pi2294;// level 0
assign po2314 = pi2135;// level 0
assign po2315 = pi2136;// level 0
assign po2316 = pi2286;// level 0
assign po2317 = ~w42542;// level 14
assign po2318 = ~pi2286;// level 0
assign po2319 = pi2317;// level 0
assign po2320 = ~w42572;// level 12
assign po2321 = ~pi2317;// level 0
assign po2322 = pi2139;// level 0
assign po2323 = ~w42663;// level 14
assign po2324 = pi2285;// level 0
assign po2325 = w42663;// level 14
assign po2326 = pi2278;// level 0
assign po2327 = w42749;// level 13
assign po2328 = ~pi2278;// level 0
assign po2329 = pi2134;// level 0
assign po2330 = pi2293;// level 0
assign po2331 = w42774;// level 14
assign po2332 = ~pi2293;// level 0
assign po2333 = pi2137;// level 0
assign po2334 = pi2287;// level 0
assign po2335 = w42800;// level 13
assign po2336 = ~pi2287;// level 0
assign po2337 = w42835;// level 14
assign po2338 = pi2274;// level 0
assign po2339 = ~w42835;// level 14
assign po2340 = pi2284;// level 0
assign po2341 = ~w42860;// level 13
assign po2342 = ~pi2284;// level 0
assign po2343 = pi2141;// level 0
assign po2344 = pi2138;// level 0
assign po2345 = pi2140;// level 0
assign po2346 = w42890;// level 14
assign po2347 = pi2300;// level 0
assign po2348 = ~w42912;// level 14
assign po2349 = ~pi2300;// level 0
assign po2350 = pi2143;// level 0
assign po2351 = pi2142;// level 0
assign po2352 = w42938;// level 14
assign po2353 = pi2283;// level 0
assign po2354 = ~w43008;// level 12
assign po2355 = ~pi2283;// level 0
assign po2356 = pi2273;// level 0
assign po2357 = ~w43034;// level 14
assign po2358 = ~pi2273;// level 0
assign po2359 = pi2292;// level 0
assign po2360 = ~w43057;// level 12
assign po2361 = ~pi2292;// level 0
assign po2362 = w43075;// level 14
assign po2363 = pi2280;// level 0
assign po2364 = ~w43104;// level 14
assign po2365 = ~pi2280;// level 0
assign po2366 = w43122;// level 14
assign po2367 = w43156;// level 14
assign po2368 = ~w43175;// level 14
assign po2369 = w43202;// level 14
assign po2370 = w43223;// level 14
assign po2371 = pi2282;// level 0
assign po2372 = ~w43238;// level 13
assign po2373 = ~pi2282;// level 0
assign po2374 = pi2159;// level 0
assign po2375 = pi2162;// level 0
assign po2376 = pi2158;// level 0
assign po2377 = pi2160;// level 0
assign po2378 = pi2178;// level 0
assign po2379 = pi2164;// level 0
assign po2380 = pi2185;// level 0
assign po2381 = pi2168;// level 0
assign po2382 = pi2174;// level 0
assign po2383 = pi2176;// level 0
assign po2384 = pi2199;// level 0
assign po2385 = pi2183;// level 0
assign po2386 = pi2184;// level 0
assign po2387 = pi2182;// level 0
assign po2388 = pi2167;// level 0
assign po2389 = pi2166;// level 0
assign po2390 = pi2170;// level 0
assign po2391 = pi2192;// level 0
assign po2392 = pi2175;// level 0
assign po2393 = pi2189;// level 0
assign po2394 = pi2181;// level 0
assign po2395 = pi2196;// level 0
assign po2396 = pi2222;// level 0
assign po2397 = pi2206;// level 0
assign po2398 = pi2187;// level 0
assign po2399 = pi2209;// level 0
assign po2400 = ~pi2198;// level 0
assign po2401 = pi2210;// level 0
assign po2402 = pi2211;// level 0
assign po2403 = pi2212;// level 0
assign po2404 = pi2190;// level 0
assign po2405 = pi2227;// level 0
assign po2406 = pi2193;// level 0
assign po2407 = pi2221;// level 0
assign po2408 = pi2194;// level 0
assign po2409 = pi2215;// level 0
assign po2410 = pi2208;// level 0
assign po2411 = pi2217;// level 0
assign po2412 = pi2207;// level 0
assign po2413 = pi2202;// level 0
assign po2414 = pi2203;// level 0
assign po2415 = pi2204;// level 0
assign po2416 = pi2224;// level 0
assign po2417 = ~pi2216;// level 0
assign po2418 = pi2225;// level 0
assign po2419 = pi2214;// level 0
assign po2420 = pi2230;// level 0
assign po2421 = pi2229;// level 0
assign po2422 = pi2213;// level 0
assign po2423 = pi2233;// level 0
assign po2424 = pi2234;// level 0
assign po2425 = pi2242;// level 0
assign po2426 = pi2220;// level 0
assign po2427 = pi2243;// level 0
assign po2428 = w43323;// level 14
assign po2429 = pi2219;// level 0
assign po2430 = pi2218;// level 0
assign po2431 = pi2244;// level 0
assign po2432 = pi2223;// level 0
assign po2433 = pi2241;// level 0
assign po2434 = pi2246;// level 0
assign po2435 = pi2238;// level 0
assign po2436 = ~w43351;// level 14
assign po2437 = pi2240;// level 0
assign po2438 = pi2236;// level 0
assign po2439 = pi2228;// level 0
assign po2440 = pi2226;// level 0
assign po2441 = pi2231;// level 0
assign po2442 = pi2232;// level 0
assign po2443 = pi2254;// level 0
assign po2444 = ~pi2247;// level 0
assign po2445 = pi2235;// level 0
assign po2446 = ~w43380;// level 14
assign po2447 = ~w43397;// level 14
assign po2448 = pi2239;// level 0
assign po2449 = pi2258;// level 0
assign po2450 = pi2245;// level 0
assign po2451 = pi2237;// level 0
assign po2452 = w43480;// level 14
assign po2453 = w43517;// level 14
assign po2454 = pi2248;// level 0
assign po2455 = pi2249;// level 0
assign po2456 = pi2253;// level 0
assign po2457 = w43607;// level 14
assign po2458 = pi2251;// level 0
assign po2459 = pi2250;// level 0
assign po2460 = w43698;// level 14
assign po2461 = pi2262;// level 0
assign po2462 = pi2252;// level 0
assign po2463 = ~w43789;// level 14
assign po2464 = ~w43878;// level 14
assign po2465 = pi2255;// level 0
assign po2466 = pi2264;// level 0
assign po2467 = pi2271;// level 0
assign po2468 = pi2260;// level 0
assign po2469 = ~pi2263;// level 0
assign po2470 = ~w43902;// level 14
assign po2471 = w43935;// level 14
assign po2472 = pi2256;// level 0
assign po2473 = pi2257;// level 0
assign po2474 = pi2259;// level 0
assign po2475 = w43961;// level 14
assign po2476 = w43987;// level 14
assign po2477 = w44013;// level 14
assign po2478 = pi2266;// level 0
assign po2479 = pi2261;// level 0
assign po2480 = ~pi2269;// level 0
assign po2481 = w44031;// level 14
assign po2482 = ~w44056;// level 14
assign po2483 = w44074;// level 14
assign po2484 = w44094;// level 14
assign po2485 = w44116;// level 14
assign po2486 = pi2267;// level 0
assign po2487 = pi2268;// level 0
assign po2488 = w44197;// level 14
assign po2489 = ~pi2270;// level 0
assign po2490 = pi2265;// level 0
assign po2491 = w44218;// level 14
assign po2492 = w44257;// level 14
assign po2493 = w44275;// level 14
assign po2494 = w44355;// level 14
assign po2495 = w44387;// level 14
assign po2496 = ~w44411;// level 14
assign po2497 = w44428;// level 14
assign po2498 = ~w44461;// level 14
assign po2499 = w44479;// level 14
assign po2500 = ~w44502;// level 14
assign po2501 = w44522;// level 14
assign po2502 = pi2275;// level 0
assign po2503 = pi2295;// level 0
assign po2504 = pi2296;// level 0
assign po2505 = ~w44608;// level 14
assign po2506 = pi2304;// level 0
assign po2507 = pi2305;// level 0
assign po2508 = pi2291;// level 0
assign po2509 = pi2310;// level 0
assign po2510 = pi2312;// level 0
assign po2511 = pi2313;// level 0
assign po2512 = pi2308;// level 0
assign po2513 = pi2314;// level 0
assign po2514 = pi2301;// level 0
assign po2515 = pi2298;// level 0
assign po2516 = pi2316;// level 0
assign po2517 = pi2320;// level 0
assign po2518 = pi2307;// level 0
assign po2519 = pi2315;// level 0
assign po2520 = pi2328;// level 0
assign po2521 = w44702;// level 14
assign po2522 = pi2326;// level 0
assign po2523 = pi2324;// level 0
assign po2524 = pi2327;// level 0
assign po2525 = ~w44728;// level 14
assign po2526 = w44767;// level 14
assign po2527 = pi2322;// level 0
assign po2528 = w44859;// level 14
assign po2529 = pi2334;// level 0
assign po2530 = pi2318;// level 0
assign po2531 = ~w44943;// level 14
assign po2532 = pi2319;// level 0
assign po2533 = pi2333;// level 0
assign po2534 = w44969;// level 14
assign po2535 = w45062;// level 14
assign po2536 = pi2329;// level 0
assign po2537 = w45083;// level 14
assign po2538 = ~w45103;// level 14
assign po2539 = pi2325;// level 0
assign po2540 = w45145;// level 14
assign po2541 = pi2323;// level 0
assign po2542 = ~w45164;// level 14
assign po2543 = w45243;// level 14
assign po2544 = ~w45275;// level 14
assign po2545 = ~w45300;// level 14
assign po2546 = ~w45384;// level 14
assign po2547 = pi2332;// level 0
assign po2548 = w45422;// level 14
assign po2549 = w45450;// level 14
assign po2550 = w45471;// level 14
assign po2551 = pi2330;// level 0
assign po2552 = ~w45492;// level 14
assign po2553 = ~w45521;// level 14
assign po2554 = w45546;// level 14
assign po2555 = ~w45572;// level 14
assign po2556 = ~w45593;// level 14
assign po2557 = w45611;// level 14
assign po2558 = w45700;// level 14
assign po2559 = ~w45720;// level 14
assign po2560 = w45741;// level 13
assign po2561 = pi2335;// level 0
assign po2562 = w45756;// level 14
assign po2563 = ~w45790;// level 14
assign po2564 = w45817;// level 14
assign po2565 = w45842;// level 14
assign po2566 = pi2346;// level 0
assign po2567 = pi2360;// level 0
assign po2568 = pi2352;// level 0
assign po2569 = pi2355;// level 0
assign po2570 = pi2370;// level 0
assign po2571 = pi2364;// level 0
assign po2572 = pi2365;// level 0
assign po2573 = pi2376;// level 0
assign po2574 = pi2367;// level 0
assign po2575 = pi2366;// level 0
assign po2576 = w45932;// level 14
assign po2577 = pi2371;// level 0
assign po2578 = pi2377;// level 0
assign po2579 = pi2381;// level 0
assign po2580 = pi2385;// level 0
assign po2581 = pi2380;// level 0
assign po2582 = w45961;// level 14
assign po2583 = pi2379;// level 0
assign po2584 = pi2384;// level 0
assign po2585 = w45985;// level 14
assign po2586 = pi2383;// level 0
assign po2587 = pi2392;// level 0
assign po2588 = pi2388;// level 0
assign po2589 = pi2387;// level 0
assign po2590 = w46008;// level 14
assign po2591 = pi2389;// level 0
assign po2592 = pi2390;// level 0
assign po2593 = pi2386;// level 0
assign po2594 = ~w46095;// level 14
assign po2595 = w46184;// level 14
assign po2596 = w46270;// level 14
assign po2597 = ~w46303;// level 14
assign po2598 = pi2397;// level 0
assign po2599 = pi2394;// level 0
assign po2600 = w46405;// level 14
assign po2601 = ~w46426;// level 14
assign po2602 = pi2395;// level 0
assign po2603 = pi2393;// level 0
assign po2604 = pi2391;// level 0
assign po2605 = pi2398;// level 0
assign po2606 = w46470;// level 14
assign po2607 = w46494;// level 14
assign po2608 = pi2396;// level 0
assign po2609 = ~w46513;// level 14
assign po2610 = w46545;// level 14
assign po2611 = ~w46618;// level 14
assign po2612 = pi2399;// level 0
assign po2613 = ~w46703;// level 14
assign po2614 = ~w46727;// level 14
assign po2615 = ~w46751;// level 14
assign po2616 = ~w46840;// level 14
assign po2617 = w46866;// level 14
assign po2618 = ~w46893;// level 14
assign po2619 = ~w46931;// level 14
assign po2620 = ~w46951;// level 14
assign po2621 = w46977;// level 14
assign po2622 = w47007;// level 14
assign po2623 = ~w47027;// level 14
assign po2624 = w47048;// level 14
assign po2625 = w47073;// level 14
assign po2626 = w47097;// level 14
assign po2627 = ~w47114;// level 14
assign po2628 = ~w47141;// level 14
assign po2629 = ~w47162;// level 14
assign po2630 = pi2424;// level 0
assign po2631 = pi2417;// level 0
assign po2632 = pi2423;// level 0
assign po2633 = pi2421;// level 0
assign po2634 = pi2435;// level 0
assign po2635 = pi2426;// level 0
assign po2636 = pi2428;// level 0
assign po2637 = pi2429;// level 0
assign po2638 = pi2437;// level 0
assign po2639 = pi2439;// level 0
assign po2640 = pi2432;// level 0
assign po2641 = pi2433;// level 0
assign po2642 = pi2440;// level 0
assign po2643 = pi2434;// level 0
assign po2644 = pi2438;// level 0
assign po2645 = pi2447;// level 0
assign po2646 = pi2448;// level 0
assign po2647 = w47254;// level 14
assign po2648 = pi2444;// level 0
assign po2649 = pi2430;// level 0
assign po2650 = pi2453;// level 0
assign po2651 = ~w47290;// level 14
assign po2652 = pi2450;// level 0
assign po2653 = ~w47380;// level 14
assign po2654 = w47401;// level 14
assign po2655 = pi2452;// level 0
assign po2656 = ~w47425;// level 14
assign po2657 = pi2442;// level 0
assign po2658 = w47514;// level 14
assign po2659 = w47543;// level 14
assign po2660 = ~w47638;// level 14
assign po2661 = pi2456;// level 0
assign po2662 = w47722;// level 14
assign po2663 = ~w47747;// level 14
assign po2664 = ~w47781;// level 14
assign po2665 = ~w47801;// level 14
assign po2666 = pi2454;// level 0
assign po2667 = w47892;// level 14
assign po2668 = w47915;// level 14
assign po2669 = ~w47936;// level 14
assign po2670 = ~w47959;// level 14
assign po2671 = pi2457;// level 0
assign po2672 = w47984;// level 14
assign po2673 = pi2458;// level 0
assign po2674 = ~w48008;// level 14
assign po2675 = pi2461;// level 0
assign po2676 = pi2459;// level 0
assign po2677 = w48034;// level 14
assign po2678 = ~w48058;// level 14
assign po2679 = pi2462;// level 0
assign po2680 = ~w48081;// level 14
assign po2681 = pi2455;// level 0
assign po2682 = w48168;// level 14
assign po2683 = ~w48200;// level 14
assign po2684 = ~w48225;// level 14
assign po2685 = ~w48258;// level 14
assign po2686 = ~w48284;// level 14
assign po2687 = w48386;// level 14
assign po2688 = w48409;// level 14
assign po2689 = w48434;// level 14
assign po2690 = pi2463;// level 0
assign po2691 = ~w48449;// level 14
assign po2692 = ~w48463;// level 14
assign po2693 = ~w48484;// level 14
assign po2694 = pi2469;// level 0
assign po2695 = pi2472;// level 0
assign po2696 = pi2482;// level 0
assign po2697 = pi2493;// level 0
assign po2698 = pi2481;// level 0
assign po2699 = ~w48570;// level 14
assign po2700 = pi2499;// level 0
assign po2701 = pi2487;// level 0
assign po2702 = w48658;// level 14
assign po2703 = pi2504;// level 0
assign po2704 = ~pi2498;// level 0
assign po2705 = pi2508;// level 0
assign po2706 = pi2505;// level 0
assign po2707 = pi2510;// level 0
assign po2708 = pi2491;// level 0
assign po2709 = pi2506;// level 0
assign po2710 = pi2511;// level 0
assign po2711 = ~w48683;// level 14
assign po2712 = ~w48708;// level 14
assign po2713 = pi2512;// level 0
assign po2714 = pi2507;// level 0
assign po2715 = pi2515;// level 0
assign po2716 = pi2514;// level 0
assign po2717 = w48748;// level 14
assign po2718 = pi2518;// level 0
assign po2719 = pi2513;// level 0
assign po2720 = pi2516;// level 0
assign po2721 = w48769;// level 14
assign po2722 = pi2519;// level 0
assign po2723 = w48791;// level 14
assign po2724 = pi2526;// level 0
assign po2725 = pi2517;// level 0
assign po2726 = pi2520;// level 0
assign po2727 = pi2522;// level 0
assign po2728 = w48892;// level 14
assign po2729 = w48979;// level 14
assign po2730 = pi2523;// level 0
assign po2731 = pi2524;// level 0
assign po2732 = pi2521;// level 0
assign po2733 = pi2525;// level 0
assign po2734 = w49075;// level 14
assign po2735 = ~w49105;// level 14
assign po2736 = w49138;// level 14
assign po2737 = w49159;// level 14
assign po2738 = ~w49181;// level 14
assign po2739 = pi2527;// level 0
assign po2740 = w49203;// level 14
assign po2741 = ~w49232;// level 14
assign po2742 = w49325;// level 14
assign po2743 = w49414;// level 14
assign po2744 = w49436;// level 14
assign po2745 = w49529;// level 14
assign po2746 = ~w49552;// level 14
assign po2747 = w49573;// level 14
assign po2748 = ~w49603;// level 14
assign po2749 = ~w49620;// level 14
assign po2750 = w49648;// level 14
assign po2751 = ~w49667;// level 14
assign po2752 = ~w49686;// level 14
assign po2753 = ~w49707;// level 14
assign po2754 = ~w49726;// level 14
assign po2755 = w49751;// level 14
assign po2756 = ~w49769;// level 14
assign po2757 = w49790;// level 14
assign po2758 = pi2537;// level 0
assign po2759 = pi2564;// level 0
assign po2760 = pi2548;// level 0
assign po2761 = pi2557;// level 0
assign po2762 = pi2560;// level 0
assign po2763 = pi2554;// level 0
assign po2764 = pi2559;// level 0
assign po2765 = pi2561;// level 0
assign po2766 = pi2563;// level 0
assign po2767 = ~w49884;// level 14
assign po2768 = pi2565;// level 0
assign po2769 = pi2566;// level 0
assign po2770 = pi2569;// level 0
assign po2771 = pi2571;// level 0
assign po2772 = pi2570;// level 0
assign po2773 = pi2575;// level 0
assign po2774 = pi2558;// level 0
assign po2775 = pi2572;// level 0
assign po2776 = pi2578;// level 0
assign po2777 = pi2579;// level 0
assign po2778 = w49911;// level 14
assign po2779 = pi2587;// level 0
assign po2780 = pi2577;// level 0
assign po2781 = pi2576;// level 0
assign po2782 = pi2582;// level 0
assign po2783 = pi2580;// level 0
assign po2784 = w50003;// level 15
assign po2785 = pi2583;// level 0
assign po2786 = pi2581;// level 0
assign po2787 = w50028;// level 14
assign po2788 = ~w50056;// level 14
assign po2789 = w50146;// level 14
assign po2790 = w50246;// level 14
assign po2791 = ~w50343;// level 14
assign po2792 = pi2584;// level 0
assign po2793 = w50368;// level 14
assign po2794 = w50395;// level 14
assign po2795 = ~w50421;// level 14
assign po2796 = ~w50446;// level 14
assign po2797 = pi2585;// level 0
assign po2798 = pi2586;// level 0
assign po2799 = w50539;// level 14
assign po2800 = ~w50549;// level 14
assign po2801 = w50570;// level 14
assign po2802 = ~w50595;// level 14
assign po2803 = pi2589;// level 0
assign po2804 = pi2591;// level 0
assign po2805 = w50618;// level 14
assign po2806 = ~w50712;// level 14
assign po2807 = ~w50737;// level 14
assign po2808 = w50822;// level 14
assign po2809 = w50855;// level 14
assign po2810 = ~w50876;// level 14
assign po2811 = w50904;// level 14
assign po2812 = w50941;// level 14
assign po2813 = w50960;// level 14
assign po2814 = ~w50986;// level 14
assign po2815 = ~w51017;// level 14
assign po2816 = w51040;// level 14
assign po2817 = ~w51054;// level 14
assign po2818 = pi2590;// level 0
assign po2819 = ~w51072;// level 14
assign po2820 = ~w51096;// level 14
assign po2821 = ~w51117;// level 14
assign po2822 = pi2613;// level 0
assign po2823 = pi2610;// level 0
assign po2824 = pi2616;// level 0
assign po2825 = pi2636;// level 0
assign po2826 = pi2617;// level 0
assign po2827 = pi2630;// level 0
assign po2828 = pi2624;// level 0
assign po2829 = pi2626;// level 0
assign po2830 = pi2629;// level 0
assign po2831 = pi2638;// level 0
assign po2832 = pi2625;// level 0
assign po2833 = pi2637;// level 0
assign po2834 = pi2628;// level 0
assign po2835 = pi2631;// level 0
assign po2836 = pi2639;// level 0
assign po2837 = pi2633;// level 0
assign po2838 = pi2632;// level 0
assign po2839 = pi2634;// level 0
assign po2840 = ~w51199;// level 14
assign po2841 = pi2640;// level 0
assign po2842 = pi2644;// level 0
assign po2843 = w51238;// level 14
assign po2844 = pi2642;// level 0
assign po2845 = pi2643;// level 0
assign po2846 = ~w51263;// level 14
assign po2847 = w51358;// level 14
assign po2848 = pi2646;// level 0
assign po2849 = pi2647;// level 0
assign po2850 = pi2649;// level 0
assign po2851 = pi2650;// level 0
assign po2852 = pi2648;// level 0
assign po2853 = pi2645;// level 0
assign po2854 = ~w51453;// level 14
assign po2855 = ~w51545;// level 14
assign po2856 = w51568;// level 14
assign po2857 = pi2651;// level 0
assign po2858 = w51668;// level 14
assign po2859 = ~w51687;// level 14
assign po2860 = w51714;// level 14
assign po2861 = w51805;// level 14
assign po2862 = w51833;// level 14
assign po2863 = w51927;// level 14
assign po2864 = w51946;// level 14
assign po2865 = pi2654;// level 0
assign po2866 = ~w51966;// level 14
assign po2867 = w51996;// level 14
assign po2868 = w52020;// level 14
assign po2869 = w52047;// level 14
assign po2870 = ~w52063;// level 14
assign po2871 = pi2653;// level 0
assign po2872 = ~w52085;// level 14
assign po2873 = ~w52108;// level 14
assign po2874 = ~w52127;// level 14
assign po2875 = w52158;// level 14
assign po2876 = w52237;// level 14
assign po2877 = ~w52260;// level 14
assign po2878 = ~w52281;// level 14
assign po2879 = ~w52310;// level 14
assign po2880 = ~w52333;// level 14
assign po2881 = w52357;// level 14
assign po2882 = pi2655;// level 0
assign po2883 = w52379;// level 14
assign po2884 = ~w52400;// level 14
assign po2885 = w52423;// level 14
assign po2886 = pi2668;// level 0
assign po2887 = pi2683;// level 0
assign po2888 = pi2674;// level 0
assign po2889 = pi2694;// level 0
assign po2890 = pi2684;// level 0
assign po2891 = pi2690;// level 0
assign po2892 = pi2695;// level 0
assign po2893 = pi2692;// level 0
assign po2894 = pi2691;// level 0
assign po2895 = pi2699;// level 0
assign po2896 = pi2686;// level 0
assign po2897 = pi2702;// level 0
assign po2898 = w52512;// level 14
assign po2899 = pi2701;// level 0
assign po2900 = pi2697;// level 0
assign po2901 = pi2700;// level 0
assign po2902 = pi2703;// level 0
assign po2903 = pi2705;// level 0
assign po2904 = ~w52602;// level 14
assign po2905 = pi2709;// level 0
assign po2906 = pi2707;// level 0
assign po2907 = pi2706;// level 0
assign po2908 = pi2708;// level 0
assign po2909 = pi2713;// level 0
assign po2910 = pi2710;// level 0
assign po2911 = pi2711;// level 0
assign po2912 = pi2712;// level 0
assign po2913 = ~w52634;// level 14
assign po2914 = ~w52723;// level 14
assign po2915 = pi2718;// level 0
assign po2916 = w52750;// level 14
assign po2917 = pi2715;// level 0
assign po2918 = pi2716;// level 0
assign po2919 = pi2719;// level 0
assign po2920 = ~w52853;// level 14
assign po2921 = ~w52886;// level 14
assign po2922 = w52911;// level 14
assign po2923 = pi2704;// level 0
assign po2924 = w52996;// level 14
assign po2925 = w53011;// level 14
assign po2926 = pi2717;// level 0
assign po2927 = ~w53099;// level 14
assign po2928 = pi2714;// level 0
assign po2929 = ~w53110;// level 14
assign po2930 = w53204;// level 14
assign po2931 = w53233;// level 14
assign po2932 = ~w53256;// level 14
assign po2933 = w53270;// level 14
assign po2934 = ~w53304;// level 14
assign po2935 = w53327;// level 14
assign po2936 = ~w53354;// level 14
assign po2937 = w53386;// level 14
assign po2938 = w53409;// level 14
assign po2939 = w53433;// level 14
assign po2940 = ~w53456;// level 14
assign po2941 = ~w53473;// level 15
assign po2942 = w53554;// level 14
assign po2943 = w53570;// level 14
assign po2944 = w53590;// level 14
assign po2945 = ~w53611;// level 14
assign po2946 = ~w53634;// level 14
assign po2947 = w53665;// level 14
assign po2948 = ~w53683;// level 14
assign po2949 = w53706;// level 14
assign po2950 = pi2738;// level 0
assign po2951 = pi2741;// level 0
assign po2952 = pi2753;// level 0
assign po2953 = pi2748;// level 0
assign po2954 = pi2757;// level 0
assign po2955 = pi2759;// level 0
assign po2956 = pi2739;// level 0
assign po2957 = pi2754;// level 0
assign po2958 = pi2755;// level 0
assign po2959 = pi2758;// level 0
assign po2960 = pi2765;// level 0
assign po2961 = pi2764;// level 0
assign po2962 = pi2766;// level 0
assign po2963 = pi2760;// level 0
assign po2964 = pi2769;// level 0
assign po2965 = pi2762;// level 0
assign po2966 = pi2768;// level 0
assign po2967 = pi2761;// level 0
assign po2968 = ~w53795;// level 14
assign po2969 = w53831;// level 14
assign po2970 = pi2776;// level 0
assign po2971 = w53926;// level 14
assign po2972 = pi2772;// level 0
assign po2973 = pi2771;// level 0
assign po2974 = pi2773;// level 0
assign po2975 = pi2775;// level 0
assign po2976 = pi2777;// level 0
assign po2977 = pi2770;// level 0
assign po2978 = ~w53949;// level 14
assign po2979 = pi2779;// level 0
assign po2980 = pi2780;// level 0
assign po2981 = pi2778;// level 0
assign po2982 = pi2767;// level 0
assign po2983 = w53971;// level 14
assign po2984 = w54063;// level 14
assign po2985 = ~w54163;// level 14
assign po2986 = pi2781;// level 0
assign po2987 = ~w54186;// level 14
assign po2988 = w54271;// level 14
assign po2989 = ~w54298;// level 14
assign po2990 = ~w54390;// level 14
assign po2991 = w54423;// level 14
assign po2992 = ~w54512;// level 14
assign po2993 = pi2783;// level 0
assign po2994 = w54551;// level 14
assign po2995 = w54637;// level 14
assign po2996 = w54673;// level 14
assign po2997 = w54694;// level 14
assign po2998 = ~w54716;// level 14
assign po2999 = ~w54735;// level 14
assign po3000 = ~w54763;// level 14
assign po3001 = ~w54787;// level 14
assign po3002 = w54811;// level 14
assign po3003 = w54837;// level 14
assign po3004 = pi2782;// level 0
assign po3005 = w54877;// level 14
assign po3006 = ~w54900;// level 14
assign po3007 = ~w54919;// level 14
assign po3008 = w54940;// level 14
assign po3009 = ~w54953;// level 14
assign po3010 = w54976;// level 14
assign po3011 = ~w54999;// level 14
assign po3012 = ~w55024;// level 14
assign po3013 = ~w55045;// level 14
assign po3014 = pi2802;// level 0
assign po3015 = pi2818;// level 0
assign po3016 = pi2812;// level 0
assign po3017 = pi2817;// level 0
assign po3018 = pi2832;// level 0
assign po3019 = pi2813;// level 0
assign po3020 = pi2820;// level 0
assign po3021 = pi2822;// level 0
assign po3022 = pi2823;// level 0
assign po3023 = pi2827;// level 0
assign po3024 = pi2826;// level 0
assign po3025 = pi2821;// level 0
assign po3026 = pi2824;// level 0
assign po3027 = pi2825;// level 0
assign po3028 = pi2831;// level 0
assign po3029 = pi2835;// level 0
assign po3030 = pi2834;// level 0
assign po3031 = pi2830;// level 0
assign po3032 = w55133;// level 14
assign po3033 = pi2833;// level 0
assign po3034 = pi2819;// level 0
assign po3035 = pi2839;// level 0
assign po3036 = pi2838;// level 0
assign po3037 = pi2828;// level 0
assign po3038 = pi2836;// level 0
assign po3039 = pi2837;// level 0
assign po3040 = pi2841;// level 0
assign po3041 = pi2842;// level 0
assign po3042 = w55158;// level 14
assign po3043 = ~w55247;// level 14
assign po3044 = pi2844;// level 0
assign po3045 = pi2846;// level 0
assign po3046 = pi2845;// level 0
assign po3047 = w55335;// level 14
assign po3048 = w55371;// level 14
assign po3049 = ~w55465;// level 14
assign po3050 = w55552;// level 14
assign po3051 = w55659;// level 15
assign po3052 = ~w55741;// level 14
assign po3053 = ~w55773;// level 14
assign po3054 = ~w55794;// level 14
assign po3055 = ~w55822;// level 14
assign po3056 = w55839;// level 14
assign po3057 = ~w55869;// level 14
assign po3058 = w55886;// level 14
assign po3059 = pi2840;// level 0
assign po3060 = ~w55907;// level 14
assign po3061 = w55930;// level 14
assign po3062 = w55942;// level 14
assign po3063 = ~w55963;// level 14
assign po3064 = ~w55984;// level 14
assign po3065 = w56003;// level 14
assign po3066 = ~w56028;// level 14
assign po3067 = w56101;// level 14
assign po3068 = ~w56131;// level 14
assign po3069 = ~w56165;// level 14
assign po3070 = w56201;// level 14
assign po3071 = ~w56220;// level 14
assign po3072 = ~w56245;// level 14
assign po3073 = pi2847;// level 0
assign po3074 = ~w56268;// level 14
assign po3075 = ~w56294;// level 14
assign po3076 = w56315;// level 14
assign po3077 = ~w56338;// level 14
assign po3078 = pi2868;// level 0
assign po3079 = pi2880;// level 0
assign po3080 = pi2882;// level 0
assign po3081 = pi2879;// level 0
assign po3082 = pi2872;// level 0
assign po3083 = pi2888;// level 0
assign po3084 = pi2881;// level 0
assign po3085 = pi2890;// level 0
assign po3086 = pi2878;// level 0
assign po3087 = pi2873;// level 0
assign po3088 = pi2885;// level 0
assign po3089 = pi2891;// level 0
assign po3090 = pi2901;// level 0
assign po3091 = pi2887;// level 0
assign po3092 = pi2886;// level 0
assign po3093 = pi2892;// level 0
assign po3094 = pi2894;// level 0
assign po3095 = pi2895;// level 0
assign po3096 = pi2904;// level 0
assign po3097 = pi2899;// level 0
assign po3098 = ~w56423;// level 14
assign po3099 = pi2897;// level 0
assign po3100 = pi2900;// level 0
assign po3101 = pi2896;// level 0
assign po3102 = ~w56506;// level 14
assign po3103 = w56602;// level 14
assign po3104 = pi2905;// level 0
assign po3105 = pi2906;// level 0
assign po3106 = pi2903;// level 0
assign po3107 = pi2907;// level 0
assign po3108 = ~w56629;// level 14
assign po3109 = w56719;// level 14
assign po3110 = w56744;// level 14
assign po3111 = w56830;// level 14
assign po3112 = w56858;// level 14
assign po3113 = pi2908;// level 0
assign po3114 = pi2910;// level 0
assign po3115 = w56956;// level 14
assign po3116 = ~w56979;// level 14
assign po3117 = w57004;// level 14
assign po3118 = w57091;// level 14
assign po3119 = pi2911;// level 0
assign po3120 = w57117;// level 14
assign po3121 = w57143;// level 14
assign po3122 = ~w57182;// level 14
assign po3123 = pi2902;// level 0
assign po3124 = w57206;// level 14
assign po3125 = w57229;// level 14
assign po3126 = ~w57250;// level 14
assign po3127 = ~w57274;// level 14
assign po3128 = pi2909;// level 0
assign po3129 = ~w57294;// level 14
assign po3130 = w57312;// level 14
assign po3131 = w57343;// level 14
assign po3132 = w57381;// level 14
assign po3133 = w57457;// level 14
assign po3134 = ~w57492;// level 14
assign po3135 = ~w57524;// level 14
assign po3136 = ~w57551;// level 14
assign po3137 = w57574;// level 14
assign po3138 = w57595;// level 14
assign po3139 = ~w57614;// level 14
assign po3140 = ~w57637;// level 14
assign po3141 = ~w57657;// level 14
assign po3142 = pi2930;// level 0
assign po3143 = pi2936;// level 0
assign po3144 = pi2938;// level 0
assign po3145 = pi2944;// level 0
assign po3146 = pi2941;// level 0
assign po3147 = pi2960;// level 0
assign po3148 = pi2961;// level 0
assign po3149 = pi2946;// level 0
assign po3150 = pi2937;// level 0
assign po3151 = pi2953;// level 0
assign po3152 = pi2954;// level 0
assign po3153 = pi2962;// level 0
assign po3154 = pi2945;// level 0
assign po3155 = pi2947;// level 0
assign po3156 = pi2952;// level 0
assign po3157 = pi2966;// level 0
assign po3158 = pi2959;// level 0
assign po3159 = pi2956;// level 0
assign po3160 = w57769;// level 14
assign po3161 = pi2967;// level 0
assign po3162 = pi2957;// level 0
assign po3163 = pi2949;// level 0
assign po3164 = pi2968;// level 0
assign po3165 = pi2964;// level 0
assign po3166 = ~w57852;// level 14
assign po3167 = w57881;// level 14
assign po3168 = w57970;// level 14
assign po3169 = pi2965;// level 0
assign po3170 = pi2970;// level 0
assign po3171 = ~w57994;// level 14
assign po3172 = pi2971;// level 0
assign po3173 = pi2969;// level 0
assign po3174 = w58022;// level 14
assign po3175 = w58114;// level 15
assign po3176 = ~w58138;// level 14
assign po3177 = w58170;// level 14
assign po3178 = pi2963;// level 0
assign po3179 = w58195;// level 14
assign po3180 = pi2972;// level 0
assign po3181 = pi2973;// level 0
assign po3182 = w58285;// level 14
assign po3183 = w58312;// level 14
assign po3184 = w58325;// level 15
assign po3185 = pi2974;// level 0
assign po3186 = w58420;// level 14
assign po3187 = ~w58438;// level 14
assign po3188 = pi2975;// level 0
assign po3189 = ~w58461;// level 14
assign po3190 = ~w58480;// level 14
assign po3191 = w58564;// level 14
assign po3192 = w58597;// level 14
assign po3193 = ~w58617;// level 14
assign po3194 = ~w58648;// level 14
assign po3195 = ~w58667;// level 14
assign po3196 = w58757;// level 14
assign po3197 = w58780;// level 14
assign po3198 = ~w58812;// level 14
assign po3199 = ~w58846;// level 14
assign po3200 = ~w58866;// level 14
assign po3201 = w58885;// level 14
assign po3202 = w58900;// level 14
assign po3203 = ~w58927;// level 14
assign po3204 = w58947;// level 14
assign po3205 = ~w58970;// level 14
assign po3206 = pi3035;// level 0
assign po3207 = pi3022;// level 0
assign po3208 = pi3023;// level 0
assign po3209 = pi3048;// level 0
assign po3210 = pi3029;// level 0
assign po3211 = pi3031;// level 0
assign po3212 = pi3050;// level 0
assign po3213 = pi3021;// level 0
assign po3214 = pi3041;// level 0
assign po3215 = pi3030;// level 0
assign po3216 = pi3020;// level 0
assign po3217 = pi3014;// level 0
assign po3218 = pi3017;// level 0
assign po3219 = pi3032;// level 0
assign po3220 = pi3013;// level 0
assign po3221 = pi3025;// level 0
assign po3222 = pi3012;// level 0
assign po3223 = pi3055;// level 0
assign po3224 = pi3015;// level 0
assign po3225 = pi3034;// level 0
assign po3226 = pi3026;// level 0
assign po3227 = pi3054;// level 0
assign po3228 = pi3037;// level 0
assign po3229 = pi3036;// level 0
assign po3230 = pi3049;// level 0
assign po3231 = pi3056;// level 0
assign po3232 = pi3027;// level 0
assign po3233 = pi3024;// level 0
assign po3234 = pi3018;// level 0
assign po3235 = pi3051;// level 0
assign po3236 = pi3039;// level 0
assign po3237 = pi3019;// level 0
assign po3238 = pi3052;// level 0
assign po3239 = pi3057;// level 0
assign po3240 = pi3061;// level 0
assign po3241 = pi3067;// level 0
assign po3242 = pi3086;// level 0
assign po3243 = pi3077;// level 0
assign po3244 = pi3094;// level 0
assign po3245 = pi3080;// level 0
assign po3246 = pi3065;// level 0
assign po3247 = pi3078;// level 0
assign po3248 = pi3070;// level 0
assign po3249 = pi3093;// level 0
assign po3250 = pi3111;// level 0
assign po3251 = pi3091;// level 0
assign po3252 = pi3108;// level 0
assign po3253 = pi3079;// level 0
assign po3254 = pi3071;// level 0
assign po3255 = pi3073;// level 0
assign po3256 = pi3082;// level 0
assign po3257 = pi3088;// level 0
assign po3258 = pi3060;// level 0
assign po3259 = pi3084;// level 0
assign po3260 = pi3069;// level 0
assign po3261 = pi3104;// level 0
assign po3262 = pi3083;// level 0
assign po3263 = pi3062;// level 0
assign po3264 = pi3109;// level 0
assign po3265 = pi3074;// level 0
assign po3266 = pi3075;// level 0
assign po3267 = pi3081;// level 0
assign po3268 = pi3059;// level 0
assign po3269 = pi3076;// level 0
assign po3270 = pi3095;// level 0
assign po3271 = pi3072;// level 0
assign po3272 = pi3097;// level 0
assign po3273 = pi3101;// level 0
assign po3274 = pi3100;// level 0
assign po3275 = pi3098;// level 0
assign po3276 = pi3096;// level 0
assign po3277 = pi3099;// level 0
assign po3278 = pi3107;// level 0
assign po3279 = pi3112;// level 0
assign po3280 = pi3085;// level 0
assign po3281 = pi3090;// level 0
assign po3282 = pi3087;// level 0
assign po3283 = pi3102;// level 0
assign po3284 = pi3089;// level 0
assign po3285 = pi3110;// level 0
assign po3286 = pi3092;// level 0
assign po3287 = pi3113;// level 0
assign po3288 = pi3114;// level 0
assign po3289 = pi3122;// level 0
assign po3290 = pi3115;// level 0
assign po3291 = pi3118;// level 0
assign po3292 = pi3116;// level 0
assign po3293 = pi3124;// level 0
assign po3294 = pi3123;// level 0
assign po3295 = pi3120;// level 0
assign po3296 = pi3126;// level 0
assign po3297 = pi3119;// level 0
assign po3298 = pi3127;// level 0
assign po3299 = pi3152;// level 0
assign po3300 = pi3158;// level 0
assign po3301 = pi3141;// level 0
assign po3302 = pi3154;// level 0
assign po3303 = pi3167;// level 0
assign po3304 = pi3148;// level 0
assign po3305 = pi3146;// level 0
assign po3306 = pi3136;// level 0
assign po3307 = pi3129;// level 0
assign po3308 = pi3142;// level 0
assign po3309 = pi3147;// level 0
assign po3310 = pi3139;// level 0
assign po3311 = pi3131;// level 0
assign po3312 = pi3135;// level 0
assign po3313 = pi3155;// level 0
assign po3314 = pi3134;// level 0
assign po3315 = pi3159;// level 0
assign po3316 = pi3156;// level 0
assign po3317 = pi3133;// level 0
assign po3318 = pi3128;// level 0
assign po3319 = pi3132;// level 0
assign po3320 = pi3166;// level 0
assign po3321 = pi3170;// level 0
assign po3322 = pi3161;// level 0
assign po3323 = pi3140;// level 0
assign po3324 = pi3149;// level 0
assign po3325 = pi3168;// level 0
assign po3326 = pi3157;// level 0
assign po3327 = pi3169;// level 0
assign po3328 = pi3163;// level 0
assign po3329 = pi3117;// level 0
assign po3330 = pi3160;// level 0
assign po3331 = pi3137;// level 0
assign po3332 = pi3121;// level 0
assign po3333 = pi3125;// level 0
assign po3334 = pi3130;// level 0
assign po3335 = pi3164;// level 0
assign po3336 = pi3165;// level 0
assign po3337 = pi3150;// level 0
assign po3338 = pi3151;// level 0
assign po3339 = pi3143;// level 0
assign po3340 = pi3145;// level 0
assign po3341 = pi3144;// level 0
assign po3342 = pi3138;// level 0
assign po3343 = pi3171;// level 0
assign po3344 = pi3172;// level 0
assign po3345 = pi3176;// level 0
assign po3346 = pi3179;// level 0
assign po3347 = pi3182;// level 0
assign po3348 = pi3177;// level 0
assign po3349 = pi3181;// level 0
assign po3350 = pi3183;// level 0
assign po3351 = pi3175;// level 0
assign po3352 = pi3178;// level 0
assign po3353 = pi3162;// level 0
assign po3354 = pi3180;// level 0
assign po3355 = pi3184;// level 0
assign po3356 = pi3153;// level 0
assign po3357 = pi3188;// level 0
assign po3358 = pi3219;// level 0
assign po3359 = pi3205;// level 0
assign po3360 = pi3213;// level 0
assign po3361 = pi3221;// level 0
assign po3362 = pi3199;// level 0
assign po3363 = pi3239;// level 0
assign po3364 = pi3197;// level 0
assign po3365 = pi3223;// level 0
assign po3366 = pi3214;// level 0
assign po3367 = pi3196;// level 0
assign po3368 = pi3202;// level 0
assign po3369 = pi3208;// level 0
assign po3370 = pi3229;// level 0
assign po3371 = pi3210;// level 0
assign po3372 = pi3201;// level 0
assign po3373 = pi3234;// level 0
assign po3374 = pi3204;// level 0
assign po3375 = pi3232;// level 0
assign po3376 = pi3207;// level 0
assign po3377 = pi3226;// level 0
assign po3378 = pi3209;// level 0
assign po3379 = pi3220;// level 0
assign po3380 = pi3230;// level 0
assign po3381 = pi3211;// level 0
assign po3382 = pi3218;// level 0
assign po3383 = pi3174;// level 0
assign po3384 = pi3200;// level 0
assign po3385 = pi3212;// level 0
assign po3386 = pi3233;// level 0
assign po3387 = pi3227;// level 0
assign po3388 = pi3215;// level 0
assign po3389 = pi3222;// level 0
assign po3390 = pi3235;// level 0
assign po3391 = pi3216;// level 0
assign po3392 = pi3224;// level 0
assign po3393 = pi3217;// level 0
assign po3394 = pi3225;// level 0
assign po3395 = pi3228;// level 0
assign po3396 = pi3206;// level 0
assign po3397 = pi3238;// level 0
assign po3398 = pi3198;// level 0
assign po3399 = pi3194;// level 0
assign po3400 = pi3203;// level 0
assign po3401 = pi3250;// level 0
assign po3402 = pi3240;// level 0
assign po3403 = pi3270;// level 0
assign po3404 = pi3258;// level 0
assign po3405 = pi3257;// level 0
assign po3406 = pi3255;// level 0
assign po3407 = pi3259;// level 0
assign po3408 = pi3263;// level 0
assign po3409 = pi3253;// level 0
assign po3410 = pi3251;// level 0
assign po3411 = pi3252;// level 0
assign po3412 = pi3256;// level 0
assign po3413 = pi3254;// level 0
assign po3414 = pi3195;// level 0
assign po3415 = pi3311;// level 0
assign po3416 = pi3310;// level 0
assign po3417 = pi3267;// level 0
assign po3418 = pi3246;// level 0
assign po3419 = pi3268;// level 0
assign po3420 = pi3269;// level 0
assign po3421 = pi3266;// level 0
assign po3422 = pi3265;// level 0
assign po3423 = pi3272;// level 0
assign po3424 = pi3302;// level 0
assign po3425 = pi3294;// level 0
assign po3426 = pi3295;// level 0
assign po3427 = pi3313;// level 0
assign po3428 = pi3290;// level 0
assign po3429 = pi3287;// level 0
assign po3430 = pi3317;// level 0
assign po3431 = pi3289;// level 0
assign po3432 = pi3318;// level 0
assign po3433 = pi3316;// level 0
assign po3434 = pi3279;// level 0
assign po3435 = pi3280;// level 0
assign po3436 = pi3274;// level 0
assign po3437 = pi3304;// level 0
assign po3438 = pi3291;// level 0
assign po3439 = pi3288;// level 0
assign po3440 = pi3319;// level 0
assign po3441 = pi3277;// level 0
assign po3442 = pi3306;// level 0
assign po3443 = pi3293;// level 0
assign po3444 = pi3285;// level 0
assign po3445 = pi3303;// level 0
assign po3446 = pi3312;// level 0
assign po3447 = pi3298;// level 0
assign po3448 = pi3284;// level 0
assign po3449 = pi3286;// level 0
assign po3450 = pi3281;// level 0
assign po3451 = pi3299;// level 0
assign po3452 = pi3275;// level 0
assign po3453 = pi3276;// level 0
assign po3454 = pi3307;// level 0
assign po3455 = pi3308;// level 0
assign po3456 = pi3297;// level 0
assign po3457 = pi3292;// level 0
assign po3458 = pi3296;// level 0
assign po3459 = pi3300;// level 0
assign po3460 = pi3315;// level 0
assign po3461 = pi3314;// level 0
assign po3462 = pi3283;// level 0
assign po3463 = pi3278;// level 0
assign po3464 = pi3305;// level 0
assign po3465 = pi3282;// level 0
assign po3466 = pi3324;// level 0
assign po3467 = pi3309;// level 0
assign po3468 = pi3320;// level 0
assign po3469 = pi3301;// level 0
assign po3470 = pi3322;// level 0
assign po3471 = pi3346;// level 0
assign po3472 = pi3327;// level 0
assign po3473 = pi3332;// level 0
assign po3474 = pi3326;// level 0
assign po3475 = pi3356;// level 0
assign po3476 = pi3333;// level 0
assign po3477 = pi3330;// level 0
assign po3478 = pi3325;// level 0
assign po3479 = pi3347;// level 0
assign po3480 = pi3321;// level 0
assign po3481 = pi3345;// level 0
assign po3482 = pi3340;// level 0
assign po3483 = pi3355;// level 0
assign po3484 = pi3334;// level 0
assign po3485 = pi3352;// level 0
assign po3486 = pi3335;// level 0
assign po3487 = pi3354;// level 0
assign po3488 = pi3339;// level 0
assign po3489 = pi3338;// level 0
assign po3490 = pi3348;// level 0
assign po3491 = pi3353;// level 0
assign po3492 = pi3351;// level 0
assign po3493 = pi3341;// level 0
assign po3494 = pi3359;// level 0
assign po3495 = w59066;// level 14
assign po3496 = ~w59154;// level 14
assign po3497 = w59239;// level 14
assign po3498 = w59327;// level 14
assign po3499 = ~w59427;// level 14
assign po3500 = w59519;// level 14
assign po3501 = pi3357;// level 0
assign po3502 = ~w59548;// level 14
assign po3503 = pi3360;// level 0
assign po3504 = pi3394;// level 0
assign po3505 = pi3367;// level 0
assign po3506 = pi3365;// level 0
assign po3507 = pi3375;// level 0
assign po3508 = pi3388;// level 0
assign po3509 = pi3376;// level 0
assign po3510 = pi3383;// level 0
assign po3511 = pi3397;// level 0
assign po3512 = pi3342;// level 0
assign po3513 = pi3371;// level 0
assign po3514 = pi3392;// level 0
assign po3515 = pi3373;// level 0
assign po3516 = pi3399;// level 0
assign po3517 = pi3368;// level 0
assign po3518 = pi3363;// level 0
assign po3519 = pi3393;// level 0
assign po3520 = pi3380;// level 0
assign po3521 = pi3398;// level 0
assign po3522 = pi3336;// level 0
assign po3523 = pi3396;// level 0
assign po3524 = pi3364;// level 0
assign po3525 = pi3337;// level 0
assign po3526 = pi3385;// level 0
assign po3527 = pi3374;// level 0
assign po3528 = pi3400;// level 0
assign po3529 = pi3384;// level 0
assign po3530 = pi3377;// level 0
assign po3531 = pi3389;// level 0
assign po3532 = pi3344;// level 0
assign po3533 = pi3372;// level 0
assign po3534 = pi3390;// level 0
assign po3535 = pi3362;// level 0
assign po3536 = pi3381;// level 0
assign po3537 = pi3386;// level 0
assign po3538 = pi3343;// level 0
assign po3539 = w59583;// level 14
assign po3540 = w59669;// level 14
assign po3541 = w59698;// level 13
assign po3542 = pi3391;// level 0
assign po3543 = pi3395;// level 0
assign po3544 = w59724;// level 14
assign po3545 = pi3379;// level 0
assign po3546 = pi3382;// level 0
assign po3547 = pi3369;// level 0
assign po3548 = pi3366;// level 0
assign po3549 = pi3378;// level 0
assign po3550 = pi3370;// level 0
assign po3551 = ~pi3361;// level 0
assign po3552 = pi3402;// level 0
assign po3553 = pi3358;// level 0
assign po3554 = ~w59747;// level 14
assign po3555 = ~w59773;// level 14
assign po3556 = ~w59800;// level 14
assign po3557 = ~w59827;// level 14
assign po3558 = pi3405;// level 0
assign po3559 = pi3403;// level 0
assign po3560 = ~w59848;// level 14
assign po3561 = pi3404;// level 0
assign po3562 = w59886;// level 14
assign po3563 = pi3401;// level 0
assign po3564 = pi3406;// level 0
assign po3565 = pi3407;// level 0
assign po3566 = pi3410;// level 0
assign po3567 = pi3409;// level 0
assign po3568 = pi3416;// level 0
assign po3569 = pi3418;// level 0
assign po3570 = pi3411;// level 0
assign po3571 = pi3408;// level 0
assign po3572 = pi3415;// level 0
assign po3573 = pi3414;// level 0
assign po3574 = pi3419;// level 0
assign po3575 = pi3417;// level 0
assign po3576 = w59920;// level 14
assign po3577 = w59940;// level 14
assign po3578 = ~w59959;// level 14
assign po3579 = pi3387;// level 0
assign po3580 = pi3422;// level 0
assign po3581 = ~w59988;// level 14
assign po3582 = pi3413;// level 0
assign po3583 = w60009;// level 14
assign po3584 = pi3420;// level 0
assign po3585 = pi3412;// level 0
assign po3586 = ~w60026;// level 14
assign po3587 = w60063;// level 14
assign po3588 = w60087;// level 14
assign po3589 = ~w60163;// level 14
assign po3590 = ~w60185;// level 14
assign po3591 = pi3425;// level 0
assign po3592 = pi3430;// level 0
assign po3593 = pi3439;// level 0
assign po3594 = pi3455;// level 0
assign po3595 = pi3436;// level 0
assign po3596 = pi3438;// level 0
assign po3597 = pi3459;// level 0
assign po3598 = pi3435;// level 0
assign po3599 = pi3460;// level 0
assign po3600 = pi3449;// level 0
assign po3601 = pi3426;// level 0
assign po3602 = pi3442;// level 0
assign po3603 = pi3427;// level 0
assign po3604 = pi3437;// level 0
assign po3605 = pi3432;// level 0
assign po3606 = pi3443;// level 0
assign po3607 = pi3446;// level 0
assign po3608 = pi3444;// level 0
assign po3609 = pi3450;// level 0
assign po3610 = pi3457;// level 0
assign po3611 = pi3445;// level 0
assign po3612 = pi3440;// level 0
assign po3613 = pi3429;// level 0
assign po3614 = pi3462;// level 0
assign po3615 = pi3421;// level 0
assign po3616 = pi3456;// level 0
assign po3617 = w60210;// level 14
assign po3618 = pi3424;// level 0
assign po3619 = pi3434;// level 0
assign po3620 = pi3461;// level 0
assign po3621 = pi3453;// level 0
assign po3622 = pi3451;// level 0
assign po3623 = pi3431;// level 0
assign po3624 = pi3441;// level 0
assign po3625 = pi3448;// level 0
assign po3626 = pi3463;// level 0
assign po3627 = pi3428;// level 0
assign po3628 = pi3447;// level 0
assign po3629 = pi3433;// level 0
assign po3630 = pi3452;// level 0
assign po3631 = pi3464;// level 0
assign po3632 = pi3423;// level 0
assign po3633 = ~w60248;// level 14
assign po3634 = ~w60272;// level 14
assign po3635 = ~w60291;// level 14
assign po3636 = pi3477;// level 0
assign po3637 = pi3466;// level 0
assign po3638 = pi3474;// level 0
assign po3639 = pi3478;// level 0
assign po3640 = pi3473;// level 0
assign po3641 = pi3470;// level 0
assign po3642 = pi3467;// level 0
assign po3643 = pi3479;// level 0
assign po3644 = pi3454;// level 0
assign po3645 = pi3475;// level 0
assign po3646 = pi3472;// level 0
assign po3647 = pi3458;// level 0
assign po3648 = pi3465;// level 0
assign po3649 = pi3468;// level 0
assign po3650 = pi3476;// level 0
assign po3651 = pi3480;// level 0
assign po3652 = w60317;// level 14
assign po3653 = pi3481;// level 0
assign po3654 = pi3502;// level 0
assign po3655 = pi3519;// level 0
assign po3656 = pi3520;// level 0
assign po3657 = pi3517;// level 0
assign po3658 = pi3498;// level 0
assign po3659 = pi3522;// level 0
assign po3660 = pi3485;// level 0
assign po3661 = pi3523;// level 0
assign po3662 = pi3488;// level 0
assign po3663 = pi3515;// level 0
assign po3664 = pi3489;// level 0
assign po3665 = pi3516;// level 0
assign po3666 = pi3513;// level 0
assign po3667 = pi3503;// level 0
assign po3668 = pi3487;// level 0
assign po3669 = pi3484;// level 0
assign po3670 = pi3504;// level 0
assign po3671 = pi3496;// level 0
assign po3672 = pi3518;// level 0
assign po3673 = pi3483;// level 0
assign po3674 = pi3493;// level 0
assign po3675 = pi3492;// level 0
assign po3676 = pi3505;// level 0
assign po3677 = pi3501;// level 0
assign po3678 = pi3500;// level 0
assign po3679 = pi3495;// level 0
assign po3680 = pi3521;// level 0
assign po3681 = pi3497;// level 0
assign po3682 = pi3508;// level 0
assign po3683 = pi3494;// level 0
assign po3684 = pi3512;// level 0
assign po3685 = pi3511;// level 0
assign po3686 = pi3509;// level 0
assign po3687 = pi3469;// level 0
assign po3688 = pi3471;// level 0
assign po3689 = pi3491;// level 0
assign po3690 = pi3514;// level 0
assign po3691 = pi3507;// level 0
assign po3692 = pi3506;// level 0
assign po3693 = pi3499;// level 0
assign po3694 = pi3482;// level 0
assign po3695 = pi3537;// level 0
assign po3696 = pi3526;// level 0
assign po3697 = pi3530;// level 0
assign po3698 = pi3533;// level 0
assign po3699 = pi3486;// level 0
assign po3700 = pi3538;// level 0
assign po3701 = pi3532;// level 0
assign po3702 = pi3490;// level 0
assign po3703 = pi3525;// level 0
assign po3704 = pi3528;// level 0
assign po3705 = pi3534;// level 0
assign po3706 = pi3527;// level 0
assign po3707 = pi3531;// level 0
assign po3708 = pi3536;// level 0
assign po3709 = pi3529;// level 0
assign po3710 = pi3510;// level 0
assign po3711 = pi3539;// level 0
assign po3712 = ~pi3524;// level 0
assign po3713 = pi3553;// level 0
assign po3714 = pi3552;// level 0
assign po3715 = pi3575;// level 0
assign po3716 = pi3543;// level 0
assign po3717 = pi3549;// level 0
assign po3718 = pi3551;// level 0
assign po3719 = pi3579;// level 0
assign po3720 = pi3568;// level 0
assign po3721 = pi3545;// level 0
assign po3722 = pi3560;// level 0
assign po3723 = pi3576;// level 0
assign po3724 = pi3540;// level 0
assign po3725 = pi3565;// level 0
assign po3726 = pi3556;// level 0
assign po3727 = pi3555;// level 0
assign po3728 = pi3564;// level 0
assign po3729 = pi3566;// level 0
assign po3730 = pi3546;// level 0
assign po3731 = pi3544;// level 0
assign po3732 = pi3548;// level 0
assign po3733 = pi3571;// level 0
assign po3734 = pi3541;// level 0
assign po3735 = pi3577;// level 0
assign po3736 = pi3570;// level 0
assign po3737 = pi3550;// level 0
assign po3738 = pi3562;// level 0
assign po3739 = pi3559;// level 0
assign po3740 = pi3535;// level 0
assign po3741 = pi3580;// level 0
assign po3742 = pi3567;// level 0
assign po3743 = pi3542;// level 0
assign po3744 = pi3569;// level 0
assign po3745 = pi3547;// level 0
assign po3746 = pi3573;// level 0
assign po3747 = pi3563;// level 0
assign po3748 = pi3572;// level 0
assign po3749 = pi3554;// level 0
assign po3750 = pi3578;// level 0
assign po3751 = pi3558;// level 0
assign po3752 = pi3574;// level 0
assign po3753 = pi3561;// level 0
assign po3754 = pi3595;// level 0
assign po3755 = pi3590;// level 0
assign po3756 = pi3586;// level 0
assign po3757 = pi3587;// level 0
assign po3758 = pi3583;// level 0
assign po3759 = pi3585;// level 0
assign po3760 = pi3584;// level 0
assign po3761 = pi3593;// level 0
assign po3762 = pi3557;// level 0
assign po3763 = pi3591;// level 0
assign po3764 = pi3582;// level 0
assign po3765 = pi3594;// level 0
assign po3766 = pi3589;// level 0
assign po3767 = pi3592;// level 0
assign po3768 = pi3596;// level 0
assign po3769 = pi3581;// level 0
assign po3770 = pi3621;// level 0
assign po3771 = pi3609;// level 0
assign po3772 = pi3620;// level 0
assign po3773 = pi3627;// level 0
assign po3774 = pi3610;// level 0
assign po3775 = pi3622;// level 0
assign po3776 = pi3631;// level 0
assign po3777 = pi3600;// level 0
assign po3778 = pi3625;// level 0
assign po3779 = pi3604;// level 0
assign po3780 = pi3635;// level 0
assign po3781 = pi3617;// level 0
assign po3782 = pi3636;// level 0
assign po3783 = pi3634;// level 0
assign po3784 = pi3601;// level 0
assign po3785 = pi3599;// level 0
assign po3786 = pi3618;// level 0
assign po3787 = pi3608;// level 0
assign po3788 = pi3614;// level 0
assign po3789 = pi3613;// level 0
assign po3790 = pi3629;// level 0
assign po3791 = pi3624;// level 0
assign po3792 = pi3616;// level 0
assign po3793 = pi3619;// level 0
assign po3794 = pi3597;// level 0
assign po3795 = pi3602;// level 0
assign po3796 = pi3598;// level 0
assign po3797 = pi3588;// level 0
assign po3798 = pi3630;// level 0
assign po3799 = pi3612;// level 0
assign po3800 = pi3637;// level 0
assign po3801 = pi3628;// level 0
assign po3802 = pi3638;// level 0
assign po3803 = pi3603;// level 0
assign po3804 = pi3605;// level 0
assign po3805 = pi3632;// level 0
assign po3806 = pi3626;// level 0
assign po3807 = pi3623;// level 0
assign po3808 = pi3607;// level 0
assign po3809 = pi3633;// level 0
assign po3810 = pi3615;// level 0
assign po3811 = pi3642;// level 0
assign po3812 = pi3641;// level 0
assign po3813 = pi3649;// level 0
assign po3814 = pi3651;// level 0
assign po3815 = pi3648;// level 0
assign po3816 = pi3647;// level 0
assign po3817 = pi3650;// level 0
assign po3818 = pi3653;// level 0
assign po3819 = pi3606;// level 0
assign po3820 = pi3639;// level 0
assign po3821 = pi3611;// level 0
assign po3822 = pi3646;// level 0
assign po3823 = pi3652;// level 0
assign po3824 = pi3640;// level 0
assign po3825 = pi3643;// level 0
assign po3826 = pi3645;// level 0
assign po3827 = pi3693;// level 0
assign po3828 = pi3682;// level 0
assign po3829 = pi3658;// level 0
assign po3830 = pi3672;// level 0
assign po3831 = pi3670;// level 0
assign po3832 = pi3692;// level 0
assign po3833 = pi3664;// level 0
assign po3834 = pi3673;// level 0
assign po3835 = pi3685;// level 0
assign po3836 = pi3677;// level 0
assign po3837 = pi3675;// level 0
assign po3838 = pi3668;// level 0
assign po3839 = pi3696;// level 0
assign po3840 = pi3671;// level 0
assign po3841 = pi3667;// level 0
assign po3842 = pi3694;// level 0
assign po3843 = pi3654;// level 0
assign po3844 = pi3663;// level 0
assign po3845 = pi3698;// level 0
assign po3846 = pi3644;// level 0
assign po3847 = pi3681;// level 0
assign po3848 = pi3669;// level 0
assign po3849 = pi3690;// level 0
assign po3850 = pi3660;// level 0
assign po3851 = pi3661;// level 0
assign po3852 = pi3665;// level 0
assign po3853 = pi3662;// level 0
assign po3854 = pi3695;// level 0
assign po3855 = pi3666;// level 0
assign po3856 = pi3659;// level 0
assign po3857 = pi3678;// level 0
assign po3858 = pi3683;// level 0
assign po3859 = pi3679;// level 0
assign po3860 = pi3691;// level 0
assign po3861 = pi3676;// level 0
assign po3862 = pi3697;// level 0
assign po3863 = pi3699;// level 0
assign po3864 = pi3656;// level 0
assign po3865 = pi3680;// level 0
assign po3866 = pi3674;// level 0
assign po3867 = pi3686;// level 0
assign po3868 = pi3684;// level 0
assign po3869 = pi3687;// level 0
assign po3870 = pi3655;// level 0
assign po3871 = pi3657;// level 0
assign po3872 = ~pi3689;// level 0
assign po3873 = pi3706;// level 0
assign po3874 = pi3708;// level 0
assign po3875 = pi3701;// level 0
assign po3876 = pi3702;// level 0
assign po3877 = pi3704;// level 0
assign po3878 = pi3705;// level 0
assign po3879 = pi3700;// level 0
assign po3880 = pi3703;// level 0
assign po3881 = pi3709;// level 0
assign po3882 = pi3707;// level 0
assign po3883 = pi3688;// level 0
assign po3884 = pi3755;// level 0
assign po3885 = pi3722;// level 0
assign po3886 = pi3720;// level 0
assign po3887 = pi3733;// level 0
assign po3888 = pi3758;// level 0
assign po3889 = pi3711;// level 0
assign po3890 = pi3730;// level 0
assign po3891 = pi3732;// level 0
assign po3892 = pi3721;// level 0
assign po3893 = pi3753;// level 0
assign po3894 = pi3750;// level 0
assign po3895 = pi3745;// level 0
assign po3896 = pi3756;// level 0
assign po3897 = pi3716;// level 0
assign po3898 = pi3743;// level 0
assign po3899 = pi3723;// level 0
assign po3900 = pi3747;// level 0
assign po3901 = pi3742;// level 0
assign po3902 = pi3715;// level 0
assign po3903 = pi3734;// level 0
assign po3904 = pi3712;// level 0
assign po3905 = pi3735;// level 0
assign po3906 = pi3725;// level 0
assign po3907 = pi3726;// level 0
assign po3908 = pi3751;// level 0
assign po3909 = pi3740;// level 0
assign po3910 = pi3739;// level 0
assign po3911 = pi3714;// level 0
assign po3912 = pi3749;// level 0
assign po3913 = pi3731;// level 0
assign po3914 = pi3746;// level 0
assign po3915 = pi3717;// level 0
assign po3916 = pi3724;// level 0
assign po3917 = pi3728;// level 0
assign po3918 = pi3737;// level 0
assign po3919 = pi3738;// level 0
assign po3920 = pi3754;// level 0
assign po3921 = pi3741;// level 0
assign po3922 = pi3729;// level 0
assign po3923 = pi3713;// level 0
assign po3924 = pi3757;// level 0
assign po3925 = pi3748;// level 0
assign po3926 = pi3719;// level 0
assign po3927 = pi3718;// level 0
assign po3928 = pi3752;// level 0
assign po3929 = pi3736;// level 0
assign po3930 = pi3772;// level 0
assign po3931 = pi3769;// level 0
assign po3932 = pi3765;// level 0
assign po3933 = pi3777;// level 0
assign po3934 = pi3766;// level 0
assign po3935 = pi3768;// level 0
assign po3936 = pi3727;// level 0
assign po3937 = pi3774;// level 0
assign po3938 = pi3744;// level 0
assign po3939 = pi3773;// level 0
assign po3940 = pi3782;// level 0
assign po3941 = pi3785;// level 0
assign po3942 = pi3838;// level 0
assign po3943 = pi3820;// level 0
assign po3944 = pi3794;// level 0
assign po3945 = pi3830;// level 0
assign po3946 = pi3831;// level 0
assign po3947 = pi3799;// level 0
assign po3948 = pi3826;// level 0
assign po3949 = pi3792;// level 0
assign po3950 = pi3833;// level 0
assign po3951 = pi3811;// level 0
assign po3952 = pi3827;// level 0
assign po3953 = pi3807;// level 0
assign po3954 = pi3818;// level 0
assign po3955 = pi3822;// level 0
assign po3956 = pi3806;// level 0
assign po3957 = pi3796;// level 0
assign po3958 = pi3825;// level 0
assign po3959 = pi3788;// level 0
assign po3960 = pi3813;// level 0
assign po3961 = pi3814;// level 0
assign po3962 = pi3828;// level 0
assign po3963 = pi3804;// level 0
assign po3964 = pi3819;// level 0
assign po3965 = pi3795;// level 0
assign po3966 = pi3823;// level 0
assign po3967 = pi3791;// level 0
assign po3968 = pi3805;// level 0
assign po3969 = pi3836;// level 0
assign po3970 = pi3834;// level 0
assign po3971 = pi3784;// level 0
assign po3972 = pi3787;// level 0
assign po3973 = pi3835;// level 0
assign po3974 = pi3837;// level 0
assign po3975 = pi3829;// level 0
assign po3976 = pi3790;// level 0
assign po3977 = pi3803;// level 0
assign po3978 = pi3817;// level 0
assign po3979 = pi3832;// level 0
assign po3980 = pi3812;// level 0
assign po3981 = pi3786;// level 0
assign po3982 = pi3775;// level 0
assign po3983 = pi3802;// level 0
assign po3984 = pi3801;// level 0
assign po3985 = pi3816;// level 0
assign po3986 = pi3821;// level 0
assign po3987 = pi3808;// level 0
assign po3988 = pi3815;// level 0
assign po3989 = pi3839;// level 0
assign po3990 = pi3866;// level 0
assign po3991 = pi3840;// level 0
assign po3992 = pi3842;// level 0
assign po3993 = pi3845;// level 0
assign po3994 = pi3853;// level 0
assign po3995 = pi3797;// level 0
assign po3996 = pi3798;// level 0
assign po3997 = pi3852;// level 0
assign po3998 = pi3859;// level 0
assign po3999 = pi3858;// level 0
assign po4000 = pi3863;// level 0
assign po4001 = pi3851;// level 0
assign po4002 = pi3855;// level 0
assign po4003 = pi3854;// level 0
assign po4004 = pi3848;// level 0
assign po4005 = pi3850;// level 0
assign po4006 = pi3915;// level 0
assign po4007 = pi3793;// level 0
assign po4008 = pi3865;// level 0
assign po4009 = pi3892;// level 0
assign po4010 = pi3862;// level 0
assign po4011 = pi3861;// level 0
assign po4012 = w60415;// level 14
assign po4013 = pi3846;// level 0
assign po4014 = pi3906;// level 0
assign po4015 = pi3923;// level 0
assign po4016 = pi3888;// level 0
assign po4017 = pi3897;// level 0
assign po4018 = pi3886;// level 0
assign po4019 = pi3870;// level 0
assign po4020 = pi3879;// level 0
assign po4021 = pi3913;// level 0
assign po4022 = pi3894;// level 0
assign po4023 = pi3893;// level 0
assign po4024 = pi3890;// level 0
assign po4025 = pi3919;// level 0
assign po4026 = pi3910;// level 0
assign po4027 = pi3904;// level 0
assign po4028 = pi3905;// level 0
assign po4029 = pi3927;// level 0
assign po4030 = pi3940;// level 0
assign po4031 = pi3918;// level 0
assign po4032 = pi3887;// level 0
assign po4033 = pi3873;// level 0
assign po4034 = pi3871;// level 0
assign po4035 = pi3903;// level 0
assign po4036 = pi3911;// level 0
assign po4037 = pi3924;// level 0
assign po4038 = pi3881;// level 0
assign po4039 = pi3912;// level 0
assign po4040 = pi3930;// level 0
assign po4041 = pi3877;// level 0
assign po4042 = pi3916;// level 0
assign po4043 = pi3909;// level 0
assign po4044 = pi3900;// level 0
assign po4045 = pi3868;// level 0
assign po4046 = pi3860;// level 0
assign po4047 = pi3889;// level 0
assign po4048 = pi3901;// level 0
assign po4049 = pi3876;// level 0
assign po4050 = pi3922;// level 0
assign po4051 = pi3908;// level 0
assign po4052 = pi3882;// level 0
assign po4053 = pi3872;// level 0
assign po4054 = pi3895;// level 0
assign po4055 = pi3920;// level 0
assign po4056 = pi3874;// level 0
assign po4057 = pi3896;// level 0
assign po4058 = pi3869;// level 0
assign po4059 = pi3925;// level 0
assign po4060 = pi3880;// level 0
assign po4061 = pi3883;// level 0
assign po4062 = pi3884;// level 0
assign po4063 = pi3878;// level 0
assign po4064 = pi3907;// level 0
assign po4065 = pi3926;// level 0
assign po4066 = pi3899;// level 0
assign po4067 = pi3928;// level 0
assign po4068 = pi3891;// level 0
assign po4069 = ~w60510;// level 14
assign po4070 = w60535;// level 14
assign po4071 = pi3931;// level 0
assign po4072 = ~w60630;// level 14
assign po4073 = pi3929;// level 0
assign po4074 = pi3936;// level 0
assign po4075 = w60715;// level 14
assign po4076 = w60758;// level 14
assign po4077 = pi3935;// level 0
assign po4078 = pi3885;// level 0
assign po4079 = pi3875;// level 0
assign po4080 = pi3902;// level 0
assign po4081 = ~w60780;// level 14
assign po4082 = ~w60874;// level 14
assign po4083 = ~w60905;// level 14
assign po4084 = pi3944;// level 0
assign po4085 = pi3898;// level 0
assign po4086 = pi3943;// level 0
assign po4087 = pi3958;// level 0
assign po4088 = pi3942;// level 0
assign po4089 = pi3914;// level 0
assign po4090 = pi3941;// level 0
assign po4091 = ~w60922;// level 14
assign po4092 = w61015;// level 14
assign po4093 = w61037;// level 14
assign po4094 = pi3960;// level 0
assign po4095 = w61060;// level 14
assign po4096 = w61093;// level 14
assign po4097 = pi3939;// level 0
assign po4098 = pi3984;// level 0
assign po4099 = pi3998;// level 0
assign po4100 = w61122;// level 14
assign po4101 = pi3982;// level 0
assign po4102 = pi4007;// level 0
assign po4103 = pi4006;// level 0
assign po4104 = pi4004;// level 0
assign po4105 = w61149;// level 14
assign po4106 = pi4010;// level 0
assign po4107 = pi4018;// level 0
assign po4108 = pi4027;// level 0
assign po4109 = pi3981;// level 0
assign po4110 = pi3992;// level 0
assign po4111 = pi3983;// level 0
assign po4112 = pi4031;// level 0
assign po4113 = pi3993;// level 0
assign po4114 = pi3994;// level 0
assign po4115 = pi4019;// level 0
assign po4116 = pi4017;// level 0
assign po4117 = pi3991;// level 0
assign po4118 = pi4035;// level 0
assign po4119 = pi4009;// level 0
assign po4120 = pi3974;// level 0
assign po4121 = pi4001;// level 0
assign po4122 = w61230;// level 14
assign po4123 = pi4016;// level 0
assign po4124 = pi4026;// level 0
assign po4125 = ~w61263;// level 14
assign po4126 = pi3990;// level 0
assign po4127 = pi3999;// level 0
assign po4128 = pi3979;// level 0
assign po4129 = pi3976;// level 0
assign po4130 = pi3975;// level 0
assign po4131 = pi4013;// level 0
assign po4132 = pi4014;// level 0
assign po4133 = pi4003;// level 0
assign po4134 = pi3988;// level 0
assign po4135 = pi4012;// level 0
assign po4136 = pi3985;// level 0
assign po4137 = pi3987;// level 0
assign po4138 = pi4008;// level 0
assign po4139 = pi4015;// level 0
assign po4140 = pi4034;// level 0
assign po4141 = pi3973;// level 0
assign po4142 = w61293;// level 14
assign po4143 = pi4030;// level 0
assign po4144 = pi4005;// level 0
assign po4145 = ~w61310;// level 14
assign po4146 = pi4002;// level 0
assign po4147 = pi3972;// level 0
assign po4148 = pi4033;// level 0
assign po4149 = pi3977;// level 0
assign po4150 = pi3997;// level 0
assign po4151 = pi3989;// level 0
assign po4152 = pi3986;// level 0
assign po4153 = pi4028;// level 0
assign po4154 = pi3980;// level 0
assign po4155 = pi3995;// level 0
assign po4156 = pi3996;// level 0
assign po4157 = pi4032;// level 0
assign po4158 = pi4000;// level 0
assign po4159 = ~w61401;// level 14
assign po4160 = ~w61416;// level 14
assign po4161 = ~w61436;// level 14
assign po4162 = pi4037;// level 0
assign po4163 = pi4044;// level 0
assign po4164 = pi4042;// level 0
assign po4165 = w61475;// level 14
assign po4166 = w61492;// level 14
assign po4167 = pi4045;// level 0
assign po4168 = pi4036;// level 0
assign po4169 = w61514;// level 14
assign po4170 = w61545;// level 14
assign po4171 = pi4011;// level 0
assign po4172 = pi3978;// level 0
assign po4173 = w61569;// level 14
assign po4174 = pi4020;// level 0
assign po4175 = pi4106;// level 0
assign po4176 = pi4038;// level 0
assign po4177 = pi4097;// level 0
assign po4178 = pi4111;// level 0
assign po4179 = pi4075;// level 0
assign po4180 = pi4114;// level 0
assign po4181 = pi4100;// level 0
assign po4182 = pi4099;// level 0
assign po4183 = pi4120;// level 0
assign po4184 = pi4101;// level 0
assign po4185 = pi4110;// level 0
assign po4186 = pi4105;// level 0
assign po4187 = pi4088;// level 0
assign po4188 = ~w61592;// level 14
assign po4189 = pi4121;// level 0
assign po4190 = ~w61621;// level 14
assign po4191 = pi4122;// level 0
assign po4192 = pi4124;// level 0
assign po4193 = pi4125;// level 0
assign po4194 = pi4137;// level 0
assign po4195 = pi4123;// level 0
assign po4196 = pi4127;// level 0
assign po4197 = pi4135;// level 0
assign po4198 = pi4069;// level 0
assign po4199 = pi4104;// level 0
assign po4200 = pi4098;// level 0
assign po4201 = pi4129;// level 0
assign po4202 = ~w61638;// level 14
assign po4203 = pi4046;// level 0
assign po4204 = pi4094;// level 0
assign po4205 = pi4096;// level 0
assign po4206 = pi4066;// level 0
assign po4207 = pi4081;// level 0
assign po4208 = pi4112;// level 0
assign po4209 = pi4076;// level 0
assign po4210 = pi4062;// level 0
assign po4211 = pi4058;// level 0
assign po4212 = pi4074;// level 0
assign po4213 = pi4061;// level 0
assign po4214 = pi4092;// level 0
assign po4215 = pi4060;// level 0
assign po4216 = pi4103;// level 0
assign po4217 = pi4109;// level 0
assign po4218 = pi4115;// level 0
assign po4219 = w61656;// level 14
assign po4220 = pi4091;// level 0
assign po4221 = pi4072;// level 0
assign po4222 = pi4087;// level 0
assign po4223 = pi4116;// level 0
assign po4224 = pi4086;// level 0
assign po4225 = pi4064;// level 0
assign po4226 = pi4051;// level 0
assign po4227 = pi4070;// level 0
assign po4228 = pi4102;// level 0
assign po4229 = pi4057;// level 0
assign po4230 = pi4084;// level 0
assign po4231 = pi4052;// level 0
assign po4232 = pi4049;// level 0
assign po4233 = pi4068;// level 0
assign po4234 = pi4108;// level 0
assign po4235 = pi4113;// level 0
assign po4236 = pi4090;// level 0
assign po4237 = pi4047;// level 0
assign po4238 = pi4083;// level 0
assign po4239 = pi4050;// level 0
assign po4240 = pi4080;// level 0
assign po4241 = pi4085;// level 0
assign po4242 = pi4089;// level 0
assign po4243 = pi4053;// level 0
assign po4244 = pi4065;// level 0
assign po4245 = pi4067;// level 0
assign po4246 = pi4055;// level 0
assign po4247 = pi4056;// level 0
assign po4248 = pi4054;// level 0
assign po4249 = pi4078;// level 0
assign po4250 = pi4071;// level 0
assign po4251 = pi4190;// level 0
assign po4252 = pi4203;// level 0
assign po4253 = pi4136;// level 0
assign po4254 = pi4200;// level 0
assign po4255 = pi4159;// level 0
assign po4256 = pi4048;// level 0
assign po4257 = pi4095;// level 0
assign po4258 = pi4059;// level 0
assign po4259 = pi4169;// level 0
assign po4260 = pi4079;// level 0
assign po4261 = pi4073;// level 0
assign po4262 = pi4082;// level 0
assign po4263 = pi4077;// level 0
assign po4264 = pi4093;// level 0
assign po4265 = pi4063;// level 0
assign po4266 = pi4213;// level 0
assign po4267 = pi4215;// level 0
assign po4268 = pi4208;// level 0
assign po4269 = pi4209;// level 0
assign po4270 = pi4128;// level 0
assign po4271 = pi4207;// level 0
assign po4272 = pi4205;// level 0
assign po4273 = pi4212;// level 0
assign po4274 = pi4214;// level 0
assign po4275 = pi4206;// level 0
assign po4276 = pi4161;// level 0
assign po4277 = pi4154;// level 0
assign po4278 = pi4153;// level 0
assign po4279 = pi4142;// level 0
assign po4280 = pi4150;// level 0
assign po4281 = pi4189;// level 0
assign po4282 = pi4177;// level 0
assign po4283 = pi4155;// level 0
assign po4284 = pi4187;// level 0
assign po4285 = pi4201;// level 0
assign po4286 = pi4165;// level 0
assign po4287 = pi4174;// level 0
assign po4288 = pi4197;// level 0
assign po4289 = pi4149;// level 0
assign po4290 = pi4144;// level 0
assign po4291 = pi4172;// level 0
assign po4292 = pi4158;// level 0
assign po4293 = pi4182;// level 0
assign po4294 = pi4170;// level 0
assign po4295 = pi4185;// level 0
assign po4296 = pi4199;// level 0
assign po4297 = pi4146;// level 0
assign po4298 = pi4178;// level 0
assign po4299 = pi4220;// level 0
assign po4300 = pi4171;// level 0
assign po4301 = pi4176;// level 0
assign po4302 = pi4145;// level 0
assign po4303 = pi4167;// level 0
assign po4304 = pi4148;// level 0
assign po4305 = pi4285;// level 0
assign po4306 = pi4198;// level 0
assign po4307 = pi4162;// level 0
assign po4308 = pi4160;// level 0
assign po4309 = pi4147;// level 0
assign po4310 = pi4164;// level 0
assign po4311 = pi4166;// level 0
assign po4312 = pi4183;// level 0
assign po4313 = pi4194;// level 0
assign po4314 = pi4181;// level 0
assign po4315 = pi4152;// level 0
assign po4316 = pi4151;// level 0
assign po4317 = pi4175;// level 0
assign po4318 = pi4293;// level 0
assign po4319 = pi4140;// level 0
assign po4320 = pi4163;// level 0
assign po4321 = pi4139;// level 0
assign po4322 = pi4157;// level 0
assign po4323 = pi4195;// level 0
assign po4324 = pi4180;// level 0
assign po4325 = pi4141;// level 0
assign po4326 = pi4188;// level 0
assign po4327 = pi4246;// level 0
assign po4328 = pi4280;// level 0
assign po4329 = pi4292;// level 0
assign po4330 = pi4247;// level 0
assign po4331 = pi4211;// level 0
assign po4332 = pi4156;// level 0
assign po4333 = pi4196;// level 0
assign po4334 = pi4204;// level 0
assign po4335 = pi4249;// level 0
assign po4336 = pi4287;// level 0
assign po4337 = pi4184;// level 0
assign po4338 = pi4168;// level 0
assign po4339 = pi4143;// level 0
assign po4340 = pi4284;// level 0
assign po4341 = pi4288;// level 0
assign po4342 = pi4202;// level 0
assign po4343 = pi4173;// level 0
assign po4344 = pi4254;// level 0
assign po4345 = pi4179;// level 0
assign po4346 = pi4186;// level 0
assign po4347 = pi4279;// level 0
assign po4348 = pi4191;// level 0
assign po4349 = pi4252;// level 0
assign po4350 = pi4286;// level 0
assign po4351 = pi4228;// level 0
assign po4352 = pi4297;// level 0
assign po4353 = pi4221;// level 0
assign po4354 = pi4303;// level 0
assign po4355 = pi4294;// level 0
assign po4356 = pi4301;// level 0
assign po4357 = pi4296;// level 0
assign po4358 = pi4309;// level 0
assign po4359 = pi4308;// level 0
assign po4360 = pi4298;// level 0
assign po4361 = pi4299;// level 0
assign po4362 = pi4216;// level 0
assign po4363 = pi4300;// level 0
assign po4364 = pi4295;// level 0
assign po4365 = pi4281;// level 0
assign po4366 = pi4282;// level 0
assign po4367 = pi4302;// level 0
assign po4368 = pi4307;// level 0
assign po4369 = pi4226;// level 0
assign po4370 = pi4283;// level 0
assign po4371 = pi4225;// level 0
assign po4372 = pi4251;// level 0
assign po4373 = pi4245;// level 0
assign po4374 = pi4256;// level 0
assign po4375 = pi4255;// level 0
assign po4376 = pi4275;// level 0
assign po4377 = pi4239;// level 0
assign po4378 = pi4250;// level 0
assign po4379 = pi4274;// level 0
assign po4380 = pi4248;// level 0
assign po4381 = pi4233;// level 0
assign po4382 = pi4217;// level 0
assign po4383 = pi4231;// level 0
assign po4384 = pi4235;// level 0
assign po4385 = pi4278;// level 0
assign po4386 = pi4242;// level 0
assign po4387 = pi4229;// level 0
assign po4388 = pi4272;// level 0
assign po4389 = pi4306;// level 0
assign po4390 = pi4223;// level 0
assign po4391 = pi4289;// level 0
assign po4392 = pi4270;// level 0
assign po4393 = pi4222;// level 0
assign po4394 = pi4258;// level 0
assign po4395 = pi4224;// level 0
assign po4396 = pi4264;// level 0
assign po4397 = pi4236;// level 0
assign po4398 = pi4291;// level 0
assign po4399 = pi4379;// level 0
assign po4400 = pi4268;// level 0
assign po4401 = pi4257;// level 0
assign po4402 = pi4237;// level 0
assign po4403 = pi4262;// level 0
assign po4404 = pi4241;// level 0
assign po4405 = pi4261;// level 0
assign po4406 = pi4232;// level 0
assign po4407 = pi4263;// level 0
assign po4408 = pi4227;// level 0
assign po4409 = pi4243;// level 0
assign po4410 = pi4259;// level 0
assign po4411 = pi4219;// level 0
assign po4412 = pi4238;// level 0
assign po4413 = pi4273;// level 0
assign po4414 = pi4316;// level 0
assign po4415 = pi4230;// level 0
assign po4416 = pi4253;// level 0
assign po4417 = pi4244;// level 0
assign po4418 = pi4276;// level 0
assign po4419 = pi4218;// level 0
assign po4420 = pi4373;// level 0
assign po4421 = pi4311;// level 0
assign po4422 = pi4317;// level 0
assign po4423 = pi4375;// level 0
assign po4424 = pi4265;// level 0
assign po4425 = pi4240;// level 0
assign po4426 = pi4234;// level 0
assign po4427 = pi4290;// level 0
assign po4428 = pi4260;// level 0
assign po4429 = pi4267;// level 0
assign po4430 = pi4310;// level 0
assign po4431 = pi4269;// level 0
assign po4432 = pi4271;// level 0
assign po4433 = pi4374;// level 0
assign po4434 = pi4381;// level 0
assign po4435 = pi4397;// level 0
assign po4436 = pi4385;// level 0
assign po4437 = pi4304;// level 0
assign po4438 = pi4400;// level 0
assign po4439 = pi4380;// level 0
assign po4440 = pi4305;// level 0
assign po4441 = pi4399;// level 0
assign po4442 = pi4382;// level 0
assign po4443 = pi4393;// level 0
assign po4444 = pi4394;// level 0
assign po4445 = pi4392;// level 0
assign po4446 = pi4384;// level 0
assign po4447 = pi4338;// level 0
assign po4448 = pi4357;// level 0
assign po4449 = pi4333;// level 0
assign po4450 = pi4408;// level 0
assign po4451 = pi4490;// level 0
assign po4452 = pi4361;// level 0
assign po4453 = pi4362;// level 0
assign po4454 = pi4354;// level 0
assign po4455 = pi4345;// level 0
assign po4456 = pi4325;// level 0
assign po4457 = pi4319;// level 0
assign po4458 = pi4403;// level 0
assign po4459 = pi4363;// level 0
assign po4460 = pi4364;// level 0
assign po4461 = pi4334;// level 0
assign po4462 = pi4368;// level 0
assign po4463 = pi4340;// level 0
assign po4464 = pi4360;// level 0
assign po4465 = pi4322;// level 0
assign po4466 = pi4342;// level 0
assign po4467 = pi4366;// level 0
assign po4468 = pi4318;// level 0
assign po4469 = pi4371;// level 0
assign po4470 = pi4353;// level 0
assign po4471 = pi4356;// level 0
assign po4472 = pi4359;// level 0
assign po4473 = pi4344;// level 0
assign po4474 = pi4336;// level 0
assign po4475 = pi4335;// level 0
assign po4476 = pi4481;// level 0
assign po4477 = pi4401;// level 0
assign po4478 = pi4332;// level 0
assign po4479 = pi4396;// level 0
assign po4480 = pi4369;// level 0
assign po4481 = pi4372;// level 0
assign po4482 = pi4404;// level 0
assign po4483 = pi4330;// level 0
assign po4484 = pi4473;// level 0
assign po4485 = pi4331;// level 0
assign po4486 = pi4326;// level 0
assign po4487 = pi4337;// level 0
assign po4488 = pi4350;// level 0
assign po4489 = pi4365;// level 0
assign po4490 = pi4347;// level 0
assign po4491 = pi4358;// level 0
assign po4492 = pi4349;// level 0
assign po4493 = pi4370;// level 0
assign po4494 = pi4376;// level 0
assign po4495 = pi4355;// level 0
assign po4496 = pi4383;// level 0
assign po4497 = pi4377;// level 0
assign po4498 = pi4343;// level 0
assign po4499 = pi4315;// level 0
assign po4500 = pi4346;// level 0
assign po4501 = pi4339;// level 0
assign po4502 = pi4351;// level 0
assign po4503 = pi4367;// level 0
assign po4504 = pi4314;// level 0
assign po4505 = pi4327;// level 0
assign po4506 = pi4378;// level 0
assign po4507 = pi4446;// level 0
assign po4508 = pi4329;// level 0
assign po4509 = pi4484;// level 0
assign po4510 = pi4475;// level 0
assign po4511 = pi4413;// level 0
assign po4512 = pi4409;// level 0
assign po4513 = pi4341;// level 0
assign po4514 = pi4483;// level 0
assign po4515 = pi4402;// level 0
assign po4516 = pi4480;// level 0
assign po4517 = pi4425;// level 0
assign po4518 = pi4477;// level 0
assign po4519 = pi4328;// level 0
assign po4520 = pi4348;// level 0
assign po4521 = pi4352;// level 0
assign po4522 = pi4419;// level 0
assign po4523 = pi4482;// level 0
assign po4524 = pi4506;// level 0
assign po4525 = pi4398;// level 0
assign po4526 = pi4479;// level 0
assign po4527 = pi4485;// level 0
assign po4528 = pi4391;// level 0
assign po4529 = pi4497;// level 0
assign po4530 = pi4493;// level 0
assign po4531 = pi4505;// level 0
assign po4532 = pi4494;// level 0
assign po4533 = pi4511;// level 0
assign po4534 = pi4507;// level 0
assign po4535 = pi4491;// level 0
assign po4536 = pi4510;// level 0
assign po4537 = pi4495;// level 0
assign po4538 = pi4492;// level 0
assign po4539 = pi4509;// level 0
assign po4540 = pi4579;// level 0
assign po4541 = pi4521;// level 0
assign po4542 = pi4543;// level 0
assign po4543 = pi4542;// level 0
assign po4544 = pi4436;// level 0
assign po4545 = pi4428;// level 0
assign po4546 = pi4561;// level 0
assign po4547 = pi4489;// level 0
assign po4548 = pi4467;// level 0
assign po4549 = pi4435;// level 0
assign po4550 = pi4538;// level 0
assign po4551 = pi4544;// level 0
assign po4552 = pi4463;// level 0
assign po4553 = pi4541;// level 0
assign po4554 = pi4540;// level 0
assign po4555 = pi4486;// level 0
assign po4556 = pi4447;// level 0
assign po4557 = pi4456;// level 0
assign po4558 = pi4426;// level 0
assign po4559 = pi4437;// level 0
assign po4560 = pi4429;// level 0
assign po4561 = pi4416;// level 0
assign po4562 = pi4454;// level 0
assign po4563 = pi4452;// level 0
assign po4564 = pi4462;// level 0
assign po4565 = pi4455;// level 0
assign po4566 = pi4406;// level 0
assign po4567 = pi4469;// level 0
assign po4568 = pi4427;// level 0
assign po4569 = pi4422;// level 0
assign po4570 = pi4405;// level 0
assign po4571 = pi4464;// level 0
assign po4572 = pi4415;// level 0
assign po4573 = pi4410;// level 0
assign po4574 = pi4432;// level 0
assign po4575 = pi4430;// level 0
assign po4576 = pi4414;// level 0
assign po4577 = pi4411;// level 0
assign po4578 = pi4421;// level 0
assign po4579 = pi4448;// level 0
assign po4580 = pi4470;// level 0
assign po4581 = pi4471;// level 0
assign po4582 = pi4451;// level 0
assign po4583 = pi4444;// level 0
assign po4584 = pi4466;// level 0
assign po4585 = pi4438;// level 0
assign po4586 = pi4442;// level 0
assign po4587 = pi4412;// level 0
assign po4588 = pi4468;// level 0
assign po4589 = pi4417;// level 0
assign po4590 = pi4433;// level 0
assign po4591 = pi4418;// level 0
assign po4592 = pi4431;// level 0
assign po4593 = pi4449;// level 0
assign po4594 = pi4461;// level 0
assign po4595 = pi4420;// level 0
assign po4596 = pi4450;// level 0
assign po4597 = pi4453;// level 0
assign po4598 = pi4459;// level 0
assign po4599 = pi4465;// level 0
assign po4600 = pi4424;// level 0
assign po4601 = pi4472;// level 0
assign po4602 = pi4457;// level 0
assign po4603 = pi4508;// level 0
assign po4604 = pi4578;// level 0
assign po4605 = pi4588;// level 0
assign po4606 = pi4460;// level 0
assign po4607 = pi4441;// level 0
assign po4608 = pi4458;// level 0
assign po4609 = pi4583;// level 0
assign po4610 = pi4603;// level 0
assign po4611 = pi4590;// level 0
assign po4612 = pi4615;// level 0
assign po4613 = pi4593;// level 0
assign po4614 = pi4553;// level 0
assign po4615 = pi4607;// level 0
assign po4616 = pi4599;// level 0
assign po4617 = pi4614;// level 0
assign po4618 = pi4598;// level 0
assign po4619 = pi4592;// level 0
assign po4620 = pi4514;// level 0
assign po4621 = pi4512;// level 0
assign po4622 = pi4613;// level 0
assign po4623 = pi4619;// level 0
assign po4624 = pi4605;// level 0
assign po4625 = pi4600;// level 0
assign po4626 = pi4617;// level 0
assign po4627 = pi4611;// level 0
assign po4628 = pi4602;// level 0
assign po4629 = pi4620;// level 0
assign po4630 = pi4616;// level 0
assign po4631 = pi4692;// level 0
assign po4632 = pi4604;// level 0
assign po4633 = pi4690;// level 0
assign po4634 = pi4650;// level 0
assign po4635 = pi4527;// level 0
assign po4636 = pi4513;// level 0
assign po4637 = pi4663;// level 0
assign po4638 = pi4695;// level 0
assign po4639 = pi4691;// level 0
assign po4640 = pi4587;// level 0
assign po4641 = pi4576;// level 0
assign po4642 = pi4556;// level 0
assign po4643 = pi4612;// level 0
assign po4644 = pi4554;// level 0
assign po4645 = pi4515;// level 0
assign po4646 = pi4552;// level 0
assign po4647 = pi4571;// level 0
assign po4648 = pi4566;// level 0
assign po4649 = pi4699;// level 0
assign po4650 = pi4549;// level 0
assign po4651 = pi4545;// level 0
assign po4652 = pi4562;// level 0
assign po4653 = pi4664;// level 0
assign po4654 = pi4589;// level 0
assign po4655 = pi4685;// level 0
assign po4656 = pi4520;// level 0
assign po4657 = pi4557;// level 0
assign po4658 = pi4572;// level 0
assign po4659 = pi4581;// level 0
assign po4660 = pi4559;// level 0
assign po4661 = pi4516;// level 0
assign po4662 = pi4575;// level 0
assign po4663 = pi4582;// level 0
assign po4664 = pi4595;// level 0
assign po4665 = pi4569;// level 0
assign po4666 = pi4570;// level 0
assign po4667 = pi4535;// level 0
assign po4668 = pi4539;// level 0
assign po4669 = pi4658;// level 0
assign po4670 = pi4594;// level 0
assign po4671 = pi4550;// level 0
assign po4672 = pi4574;// level 0
assign po4673 = pi4672;// level 0
assign po4674 = pi4564;// level 0
assign po4675 = pi4669;// level 0
assign po4676 = pi4698;// level 0
assign po4677 = pi4524;// level 0
assign po4678 = pi4577;// level 0
assign po4679 = pi4565;// level 0
assign po4680 = pi4563;// level 0
assign po4681 = pi4551;// level 0
assign po4682 = pi4568;// level 0
assign po4683 = pi4525;// level 0
assign po4684 = pi4526;// level 0
assign po4685 = pi4518;// level 0
assign po4686 = pi4580;// level 0
assign po4687 = pi4519;// level 0
assign po4688 = pi4547;// level 0
assign po4689 = pi4529;// level 0
assign po4690 = pi4558;// level 0
assign po4691 = pi4586;// level 0
assign po4692 = pi4528;// level 0
assign po4693 = pi4531;// level 0
assign po4694 = pi4523;// level 0
assign po4695 = pi4567;// level 0
assign po4696 = pi4548;// level 0
assign po4697 = pi4555;// level 0
assign po4698 = pi4533;// level 0
assign po4699 = pi4517;// level 0
assign po4700 = pi4530;// level 0
assign po4701 = pi4522;// level 0
assign po4702 = pi4573;// level 0
assign po4703 = pi4654;// level 0
assign po4704 = pi4668;// level 0
assign po4705 = pi4689;// level 0
assign po4706 = pi4661;// level 0
assign po4707 = pi4606;// level 0
assign po4708 = pi4667;// level 0
assign po4709 = pi4608;// level 0
assign po4710 = pi4652;// level 0
assign po4711 = pi4623;// level 0
assign po4712 = pi4710;// level 0
assign po4713 = pi4709;// level 0
assign po4714 = pi4678;// level 0
assign po4715 = pi4618;// level 0
assign po4716 = pi4560;// level 0
assign po4717 = pi4659;// level 0
assign po4718 = pi4660;// level 0
assign po4719 = pi4711;// level 0
assign po4720 = pi4675;// level 0
assign po4721 = pi4591;// level 0
assign po4722 = pi4610;// level 0
assign po4723 = pi4718;// level 0
assign po4724 = pi4716;// level 0
assign po4725 = pi4730;// level 0
assign po4726 = pi4724;// level 0
assign po4727 = pi4735;// level 0
assign po4728 = pi4674;// level 0
assign po4729 = pi4728;// level 0
assign po4730 = pi4726;// level 0
assign po4731 = pi4719;// level 0
assign po4732 = pi4732;// level 0
assign po4733 = pi4722;// level 0
assign po4734 = pi4721;// level 0
assign po4735 = pi4609;// level 0
assign po4736 = pi4715;// level 0
assign po4737 = pi4733;// level 0
assign po4738 = pi4707;// level 0
assign po4739 = pi4734;// level 0
assign po4740 = pi4738;// level 0
assign po4741 = pi4737;// level 0
assign po4742 = pi4736;// level 0
assign po4743 = pi4697;// level 0
assign po4744 = pi4800;// level 0
assign po4745 = pi4641;// level 0
assign po4746 = pi4625;// level 0
assign po4747 = pi4643;// level 0
assign po4748 = pi4631;// level 0
assign po4749 = pi4680;// level 0
assign po4750 = pi4628;// level 0
assign po4751 = pi4754;// level 0
assign po4752 = pi4696;// level 0
assign po4753 = pi4624;// level 0
assign po4754 = pi4673;// level 0
assign po4755 = pi4653;// level 0
assign po4756 = pi4632;// level 0
assign po4757 = pi4621;// level 0
assign po4758 = pi4687;// level 0
assign po4759 = pi4636;// level 0
assign po4760 = pi4679;// level 0
assign po4761 = pi4714;// level 0
assign po4762 = pi4727;// level 0
assign po4763 = pi4644;// level 0
assign po4764 = pi4666;// level 0
assign po4765 = pi4648;// level 0
assign po4766 = pi4756;// level 0
assign po4767 = pi4665;// level 0
assign po4768 = pi4752;// level 0
assign po4769 = pi4712;// level 0
assign po4770 = pi4761;// level 0
assign po4771 = pi4759;// level 0
assign po4772 = pi4758;// level 0
assign po4773 = pi4751;// level 0
assign po4774 = pi4750;// level 0
assign po4775 = pi4703;// level 0
assign po4776 = pi4763;// level 0
assign po4777 = pi4683;// level 0
assign po4778 = pi4708;// level 0
assign po4779 = pi4713;// level 0
assign po4780 = pi4701;// level 0
assign po4781 = pi4639;// level 0
assign po4782 = pi4627;// level 0
assign po4783 = pi4780;// level 0
assign po4784 = pi4681;// level 0
assign po4785 = pi4629;// level 0
assign po4786 = pi4635;// level 0
assign po4787 = pi4676;// level 0
assign po4788 = pi4694;// level 0
assign po4789 = pi4630;// level 0
assign po4790 = pi4677;// level 0
assign po4791 = pi4781;// level 0
assign po4792 = pi4651;// level 0
assign po4793 = pi4622;// level 0
assign po4794 = pi4702;// level 0
assign po4795 = pi4626;// level 0
assign po4796 = pi4704;// level 0
assign po4797 = pi4655;// level 0
assign po4798 = pi4637;// level 0
assign po4799 = pi4640;// level 0
assign po4800 = pi4688;// level 0
assign po4801 = pi4700;// level 0
assign po4802 = pi4693;// level 0
assign po4803 = pi4671;// level 0
assign po4804 = pi4633;// level 0
assign po4805 = pi4638;// level 0
assign po4806 = pi4634;// level 0
assign po4807 = pi4649;// level 0
assign po4808 = pi4774;// level 0
assign po4809 = pi4794;// level 0
assign po4810 = pi4642;// level 0
assign po4811 = pi4684;// level 0
assign po4812 = pi4682;// level 0
assign po4813 = pi4772;// level 0
assign po4814 = pi4725;// level 0
assign po4815 = pi4670;// level 0
assign po4816 = pi4686;// level 0
assign po4817 = pi4647;// level 0
assign po4818 = pi4805;// level 0
assign po4819 = pi4705;// level 0
assign po4820 = pi4821;// level 0
assign po4821 = pi4839;// level 0
assign po4822 = pi4824;// level 0
assign po4823 = pi4731;// level 0
assign po4824 = pi4826;// level 0
assign po4825 = pi4825;// level 0
assign po4826 = pi4830;// level 0
assign po4827 = pi4723;// level 0
assign po4828 = pi4828;// level 0
assign po4829 = pi4819;// level 0
assign po4830 = pi4820;// level 0
assign po4831 = pi4823;// level 0
assign po4832 = pi4815;// level 0
assign po4833 = pi4816;// level 0
assign po4834 = pi4841;// level 0
assign po4835 = pi4844;// level 0
assign po4836 = pi4818;// level 0
assign po4837 = pi4846;// level 0
assign po4838 = pi4843;// level 0
assign po4839 = pi4817;// level 0
assign po4840 = pi4840;// level 0
assign po4841 = pi4833;// level 0
assign po4842 = pi4842;// level 0
assign po4843 = pi4834;// level 0
assign po4844 = pi4829;// level 0
assign po4845 = pi4831;// level 0
assign po4846 = pi4845;// level 0
assign po4847 = pi4849;// level 0
assign po4848 = pi4838;// level 0
assign po4849 = pi4847;// level 0
assign po4850 = pi4835;// level 0
assign po4851 = pi4770;// level 0
assign po4852 = pi4790;// level 0
assign po4853 = pi4923;// level 0
assign po4854 = pi4786;// level 0
assign po4855 = pi4788;// level 0
assign po4856 = pi4766;// level 0
assign po4857 = pi4783;// level 0
assign po4858 = pi4744;// level 0
assign po4859 = pi4777;// level 0
assign po4860 = pi4806;// level 0
assign po4861 = pi4741;// level 0
assign po4862 = pi4768;// level 0
assign po4863 = pi4739;// level 0
assign po4864 = pi4814;// level 0
assign po4865 = pi4762;// level 0
assign po4866 = pi4808;// level 0
assign po4867 = pi4775;// level 0
assign po4868 = pi4779;// level 0
assign po4869 = pi4795;// level 0
assign po4870 = pi4798;// level 0
assign po4871 = pi4753;// level 0
assign po4872 = pi4789;// level 0
assign po4873 = pi4765;// level 0
assign po4874 = pi4740;// level 0
assign po4875 = pi4873;// level 0
assign po4876 = pi4860;// level 0
assign po4877 = pi4776;// level 0
assign po4878 = pi4799;// level 0
assign po4879 = pi4797;// level 0
assign po4880 = pi4891;// level 0
assign po4881 = pi4792;// level 0
assign po4882 = pi4854;// level 0
assign po4883 = pi4745;// level 0
assign po4884 = pi4836;// level 0
assign po4885 = pi4785;// level 0
assign po4886 = pi4867;// level 0
assign po4887 = pi4858;// level 0
assign po4888 = pi4938;// level 0
assign po4889 = pi4827;// level 0
assign po4890 = pi4941;// level 0
assign po4891 = pi4862;// level 0
assign po4892 = pi4864;// level 0
assign po4893 = pi4863;// level 0
assign po4894 = pi4868;// level 0
assign po4895 = pi4859;// level 0
assign po4896 = pi4866;// level 0
assign po4897 = pi4856;// level 0
assign po4898 = pi4939;// level 0
assign po4899 = pi4942;// level 0
assign po4900 = pi4855;// level 0
assign po4901 = pi4746;// level 0
assign po4902 = pi4848;// level 0
assign po4903 = pi4769;// level 0
assign po4904 = pi4869;// level 0
assign po4905 = pi4890;// level 0
assign po4906 = pi4791;// level 0
assign po4907 = pi4793;// level 0
assign po4908 = pi4883;// level 0
assign po4909 = pi4767;// level 0
assign po4910 = pi4809;// level 0
assign po4911 = pi4812;// level 0
assign po4912 = pi4755;// level 0
assign po4913 = pi4811;// level 0
assign po4914 = pi4784;// level 0
assign po4915 = pi4943;// level 0
assign po4916 = pi4771;// level 0
assign po4917 = pi4747;// level 0
assign po4918 = pi4810;// level 0
assign po4919 = pi4881;// level 0
assign po4920 = pi4837;// level 0
assign po4921 = pi4874;// level 0
assign po4922 = pi4906;// level 0
assign po4923 = pi4796;// level 0
assign po4924 = pi4743;// level 0
assign po4925 = pi4911;// level 0
assign po4926 = pi4787;// level 0
assign po4927 = pi4801;// level 0
assign po4928 = pi4852;// level 0
assign po4929 = pi4882;// level 0
assign po4930 = pi4749;// level 0
assign po4931 = pi4742;// level 0
assign po4932 = pi4802;// level 0
assign po4933 = pi4778;// level 0
assign po4934 = pi4748;// level 0
assign po4935 = pi4807;// level 0
assign po4936 = pi4872;// level 0
assign po4937 = pi4898;// level 0
assign po4938 = pi4773;// level 0
assign po4939 = pi4876;// level 0
assign po4940 = pi4832;// level 0
assign po4941 = pi4850;// level 0
assign po4942 = pi4760;// level 0
assign po4943 = pi4813;// level 0
assign po4944 = pi4782;// level 0
assign po4945 = pi4964;// level 0
assign po4946 = pi4961;// level 0
assign po4947 = pi4950;// level 0
assign po4948 = pi4947;// level 0
assign po4949 = pi4870;// level 0
assign po4950 = pi4955;// level 0
assign po4951 = pi4865;// level 0
assign po4952 = pi4956;// level 0
assign po4953 = pi4952;// level 0
assign po4954 = pi4953;// level 0
assign po4955 = pi4954;// level 0
assign po4956 = pi4951;// level 0
assign po4957 = pi4857;// level 0
assign po4958 = pi4968;// level 0
assign po4959 = pi4871;// level 0
assign po4960 = pi4959;// level 0
assign po4961 = pi4958;// level 0
assign po4962 = pi4948;// level 0
assign po4963 = pi4957;// level 0
assign po4964 = pi4962;// level 0
assign po4965 = pi4949;// level 0
assign po4966 = pi4967;// level 0
assign po4967 = pi4963;// level 0
assign po4968 = pi4909;// level 0
assign po4969 = pi4936;// level 0
assign po4970 = pi4932;// level 0
assign po4971 = pi4908;// level 0
assign po4972 = pi4880;// level 0
assign po4973 = pi4895;// level 0
assign po4974 = pi4946;// level 0
assign po4975 = pi4878;// level 0
assign po4976 = pi4901;// level 0
assign po4977 = pi4907;// level 0
assign po4978 = pi4879;// level 0
assign po4979 = pi4851;// level 0
assign po4980 = pi4971;// level 0
assign po4981 = pi5036;// level 0
assign po4982 = pi4989;// level 0
assign po4983 = pi4886;// level 0
assign po4984 = pi5038;// level 0
assign po4985 = pi4917;// level 0
assign po4986 = pi4977;// level 0
assign po4987 = pi4975;// level 0
assign po4988 = pi4976;// level 0
assign po4989 = pi4974;// level 0
assign po4990 = pi4912;// level 0
assign po4991 = pi5042;// level 0
assign po4992 = pi4929;// level 0
assign po4993 = pi4893;// level 0
assign po4994 = pi4980;// level 0
assign po4995 = pi4920;// level 0
assign po4996 = pi4944;// level 0
assign po4997 = pi4913;// level 0
assign po4998 = pi4927;// level 0
assign po4999 = pi4925;// level 0
assign po5000 = pi4914;// level 0
assign po5001 = pi4853;// level 0
assign po5002 = pi4984;// level 0
assign po5003 = pi4889;// level 0
assign po5004 = pi4987;// level 0
assign po5005 = pi4894;// level 0
assign po5006 = pi4928;// level 0
assign po5007 = pi4904;// level 0
assign po5008 = pi4924;// level 0
assign po5009 = pi4919;// level 0
assign po5010 = pi4990;// level 0
assign po5011 = pi4988;// level 0
assign po5012 = pi4902;// level 0
assign po5013 = pi4877;// level 0
assign po5014 = pi4888;// level 0
assign po5015 = pi4900;// level 0
assign po5016 = pi4935;// level 0
assign po5017 = pi4892;// level 0
assign po5018 = pi4930;// level 0
assign po5019 = pi4915;// level 0
assign po5020 = pi4934;// level 0
assign po5021 = pi4875;// level 0
assign po5022 = pi4933;// level 0
assign po5023 = pi4905;// level 0
assign po5024 = pi5039;// level 0
assign po5025 = pi4903;// level 0
assign po5026 = pi4931;// level 0
assign po5027 = pi4921;// level 0
assign po5028 = pi4896;// level 0
assign po5029 = pi4884;// level 0
assign po5030 = pi4979;// level 0
assign po5031 = pi4916;// level 0
assign po5032 = pi4945;// level 0
assign po5033 = pi4969;// level 0
assign po5034 = pi4861;// level 0
assign po5035 = pi4937;// level 0
assign po5036 = pi4922;// level 0
assign po5037 = pi4918;// level 0
assign po5038 = pi4910;// level 0
assign po5039 = pi4885;// level 0
assign po5040 = pi4897;// level 0
assign po5041 = pi4887;// level 0
assign po5042 = pi4940;// level 0
assign po5043 = pi4899;// level 0
assign po5044 = pi4926;// level 0
assign po5045 = pi5060;// level 0
assign po5046 = pi4960;// level 0
assign po5047 = pi4966;// level 0
assign po5048 = pi5058;// level 0
assign po5049 = pi5080;// level 0
assign po5050 = pi5057;// level 0
assign po5051 = pi5065;// level 0
assign po5052 = pi5054;// level 0
assign po5053 = pi5052;// level 0
assign po5054 = pi5051;// level 0
assign po5055 = pi5055;// level 0
assign po5056 = pi5049;// level 0
assign po5057 = pi5047;// level 0
assign po5058 = pi5046;// level 0
assign po5059 = pi5082;// level 0
assign po5060 = pi5081;// level 0
assign po5061 = pi4965;// level 0
assign po5062 = pi5079;// level 0
assign po5063 = pi5068;// level 0
assign po5064 = pi5062;// level 0
assign po5065 = pi5066;// level 0
assign po5066 = pi5072;// level 0
assign po5067 = pi5078;// level 0
assign po5068 = pi5061;// level 0
assign po5069 = pi5063;// level 0
assign po5070 = pi5064;// level 0
assign po5071 = pi5075;// level 0
assign po5072 = pi5076;// level 0
assign po5073 = pi5067;// level 0
assign po5074 = pi5074;// level 0
assign po5075 = pi5083;// level 0
assign po5076 = pi5069;// level 0
assign po5077 = pi5070;// level 0
assign po5078 = pi5056;// level 0
assign po5079 = pi5071;// level 0
assign po5080 = pi5059;// level 0
assign po5081 = pi5014;// level 0
assign po5082 = pi5037;// level 0
assign po5083 = pi5040;// level 0
assign po5084 = pi5154;// level 0
assign po5085 = pi5053;// level 0
assign po5086 = pi5094;// level 0
assign po5087 = pi5093;// level 0
assign po5088 = pi5090;// level 0
assign po5089 = pi5106;// level 0
assign po5090 = pi5111;// level 0
assign po5091 = pi5114;// level 0
assign po5092 = pi5096;// level 0
assign po5093 = pi5099;// level 0
assign po5094 = pi4970;// level 0
assign po5095 = pi5108;// level 0
assign po5096 = pi5109;// level 0
assign po5097 = pi5095;// level 0
assign po5098 = pi5101;// level 0
assign po5099 = pi5091;// level 0
assign po5100 = pi5105;// level 0
assign po5101 = pi5092;// level 0
assign po5102 = pi5087;// level 0
assign po5103 = pi4978;// level 0
assign po5104 = pi5156;// level 0
assign po5105 = pi5032;// level 0
assign po5106 = pi5164;// level 0
assign po5107 = pi5017;// level 0
assign po5108 = pi4997;// level 0
assign po5109 = pi5001;// level 0
assign po5110 = pi5030;// level 0
assign po5111 = pi5112;// level 0
assign po5112 = pi5144;// level 0
assign po5113 = pi5043;// level 0
assign po5114 = pi4983;// level 0
assign po5115 = pi5031;// level 0
assign po5116 = pi5029;// level 0
assign po5117 = pi4985;// level 0
assign po5118 = pi4972;// level 0
assign po5119 = pi5022;// level 0
assign po5120 = pi5151;// level 0
assign po5121 = pi5116;// level 0
assign po5122 = pi5007;// level 0
assign po5123 = pi5104;// level 0
assign po5124 = pi4986;// level 0
assign po5125 = pi5006;// level 0
assign po5126 = pi5021;// level 0
assign po5127 = pi5008;// level 0
assign po5128 = pi5152;// level 0
assign po5129 = pi5016;// level 0
assign po5130 = pi5020;// level 0
assign po5131 = pi5010;// level 0
assign po5132 = pi4999;// level 0
assign po5133 = pi5005;// level 0
assign po5134 = pi4982;// level 0
assign po5135 = pi5041;// level 0
assign po5136 = pi5155;// level 0
assign po5137 = pi5024;// level 0
assign po5138 = pi5015;// level 0
assign po5139 = pi5117;// level 0
assign po5140 = pi5023;// level 0
assign po5141 = pi5143;// level 0
assign po5142 = pi4992;// level 0
assign po5143 = pi5044;// level 0
assign po5144 = pi4993;// level 0
assign po5145 = pi4991;// level 0
assign po5146 = pi4995;// level 0
assign po5147 = pi4981;// level 0
assign po5148 = pi5002;// level 0
assign po5149 = pi5012;// level 0
assign po5150 = pi5019;// level 0
assign po5151 = pi5004;// level 0
assign po5152 = pi4994;// level 0
assign po5153 = pi5073;// level 0
assign po5154 = pi5013;// level 0
assign po5155 = pi5018;// level 0
assign po5156 = pi5027;// level 0
assign po5157 = pi5025;// level 0
assign po5158 = pi4998;// level 0
assign po5159 = pi5009;// level 0
assign po5160 = pi5035;// level 0
assign po5161 = pi5033;// level 0
assign po5162 = pi5045;// level 0
assign po5163 = pi5028;// level 0
assign po5164 = pi4996;// level 0
assign po5165 = pi4973;// level 0
assign po5166 = pi5000;// level 0
assign po5167 = pi5150;// level 0
assign po5168 = pi5048;// level 0
assign po5169 = pi5097;// level 0
assign po5170 = pi5026;// level 0
assign po5171 = pi5107;// level 0
assign po5172 = pi5103;// level 0
assign po5173 = pi5089;// level 0
assign po5174 = pi5034;// level 0
assign po5175 = pi5011;// level 0
assign po5176 = pi5003;// level 0
assign po5177 = pi5077;// level 0
assign po5178 = pi5088;// level 0
assign po5179 = pi5185;// level 0
assign po5180 = pi5050;// level 0
assign po5181 = pi5180;// level 0
assign po5182 = pi5181;// level 0
assign po5183 = pi5179;// level 0
assign po5184 = pi5178;// level 0
assign po5185 = pi5186;// level 0
assign po5186 = pi5110;// level 0
assign po5187 = pi5194;// level 0
assign po5188 = pi5187;// level 0
assign po5189 = pi5184;// level 0
assign po5190 = pi5189;// level 0
assign po5191 = pi5190;// level 0
assign po5192 = pi5196;// level 0
assign po5193 = pi5193;// level 0
assign po5194 = pi5188;// level 0
assign po5195 = pi5182;// level 0
assign po5196 = pi5195;// level 0
assign po5197 = pi5192;// level 0
assign po5198 = pi5102;// level 0
assign po5199 = pi5211;// level 0
assign po5200 = pi5100;// level 0
assign po5201 = pi5214;// level 0
assign po5202 = pi5129;// level 0
assign po5203 = pi5175;// level 0
assign po5204 = pi5213;// level 0
assign po5205 = pi5210;// level 0
assign po5206 = pi5215;// level 0
assign po5207 = pi5208;// level 0
assign po5208 = pi5206;// level 0
assign po5209 = pi5207;// level 0
assign po5210 = pi5277;// level 0
assign po5211 = pi5177;// level 0
assign po5212 = pi5120;// level 0
assign po5213 = pi5086;// level 0
assign po5214 = pi5252;// level 0
assign po5215 = pi5165;// level 0
assign po5216 = pi5137;// level 0
assign po5217 = pi5253;// level 0
assign po5218 = pi5250;// level 0
assign po5219 = pi5204;// level 0
assign po5220 = pi5262;// level 0
assign po5221 = pi5141;// level 0
assign po5222 = pi5134;// level 0
assign po5223 = pi5124;// level 0
assign po5224 = pi5149;// level 0
assign po5225 = pi5169;// level 0
assign po5226 = pi5145;// level 0
assign po5227 = pi5133;// level 0
assign po5228 = pi5121;// level 0
assign po5229 = pi5123;// level 0
assign po5230 = pi5142;// level 0
assign po5231 = pi5172;// level 0
assign po5232 = pi5127;// level 0
assign po5233 = pi5132;// level 0
assign po5234 = pi5085;// level 0
assign po5235 = pi5167;// level 0
assign po5236 = pi5148;// level 0
assign po5237 = pi5139;// level 0
assign po5238 = pi5131;// level 0
assign po5239 = pi5115;// level 0
assign po5240 = pi5140;// level 0
assign po5241 = pi5126;// level 0
assign po5242 = pi5157;// level 0
assign po5243 = pi5138;// level 0
assign po5244 = pi5163;// level 0
assign po5245 = pi5170;// level 0
assign po5246 = pi5168;// level 0
assign po5247 = pi5176;// level 0
assign po5248 = pi5166;// level 0
assign po5249 = pi5158;// level 0
assign po5250 = pi5162;// level 0
assign po5251 = pi5147;// level 0
assign po5252 = pi5118;// level 0
assign po5253 = pi5119;// level 0
assign po5254 = pi5128;// level 0
assign po5255 = pi5084;// level 0
assign po5256 = pi5125;// level 0
assign po5257 = pi5153;// level 0
assign po5258 = pi5171;// level 0
assign po5259 = pi5159;// level 0
assign po5260 = pi5130;// level 0
assign po5261 = pi5160;// level 0
assign po5262 = pi5146;// level 0
assign po5263 = pi5136;// level 0
assign po5264 = pi5122;// level 0
assign po5265 = pi5173;// level 0
assign po5266 = pi5203;// level 0
assign po5267 = pi5278;// level 0
assign po5268 = pi5245;// level 0
assign po5269 = pi5267;// level 0
assign po5270 = pi5174;// level 0
assign po5271 = pi5135;// level 0
assign po5272 = pi5212;// level 0
assign po5273 = pi5255;// level 0
assign po5274 = pi5161;// level 0
assign po5275 = pi5113;// level 0
assign po5276 = pi5288;// level 0
assign po5277 = pi5287;// level 0
assign po5278 = pi5289;// level 0
assign po5279 = pi5297;// level 0
assign po5280 = pi5291;// level 0
assign po5281 = pi5296;// level 0
assign po5282 = pi5290;// level 0
assign po5283 = pi5283;// level 0
assign po5284 = pi5295;// level 0
assign po5285 = pi5286;// level 0
assign po5286 = pi5284;// level 0
assign po5287 = pi5285;// level 0
assign po5288 = pi5318;// level 0
assign po5289 = pi5314;// level 0
assign po5290 = pi5302;// level 0
assign po5291 = pi5303;// level 0
assign po5292 = pi5306;// level 0
assign po5293 = pi5315;// level 0
assign po5294 = pi5313;// level 0
assign po5295 = pi5316;// level 0
assign po5296 = pi5321;// level 0
assign po5297 = pi5309;// level 0
assign po5298 = pi5319;// level 0
assign po5299 = pi5325;// level 0
assign po5300 = pi5324;// level 0
assign po5301 = pi5305;// level 0
assign po5302 = pi5308;// level 0
assign po5303 = pi5299;// level 0
assign po5304 = pi5322;// level 0
assign po5305 = pi5323;// level 0
assign po5306 = pi5317;// level 0
assign po5307 = pi5312;// level 0
assign po5308 = pi5293;// level 0
assign po5309 = pi5311;// level 0
assign po5310 = pi5298;// level 0
assign po5311 = pi5281;// level 0
assign po5312 = pi5205;// level 0
assign po5313 = pi5320;// level 0
assign po5314 = pi5266;// level 0
assign po5315 = pi5220;// level 0
assign po5316 = pi5246;// level 0
assign po5317 = pi5418;// level 0
assign po5318 = pi5333;// level 0
assign po5319 = pi5310;// level 0
assign po5320 = pi5332;// level 0
assign po5321 = pi5346;// level 0
assign po5322 = pi5343;// level 0
assign po5323 = pi5378;// level 0
assign po5324 = pi5336;// level 0
assign po5325 = pi5327;// level 0
assign po5326 = pi5338;// level 0
assign po5327 = pi5337;// level 0
assign po5328 = pi5512;// level 0
assign po5329 = pi5421;// level 0
assign po5330 = pi5345;// level 0
assign po5331 = pi5344;// level 0
assign po5332 = pi5335;// level 0
assign po5333 = pi5341;// level 0
assign po5334 = pi5330;// level 0
assign po5335 = pi5422;// level 0
assign po5336 = pi5334;// level 0
assign po5337 = pi5358;// level 0
assign po5338 = pi5348;// level 0
assign po5339 = pi5340;// level 0
assign po5340 = pi5292;// level 0
assign po5341 = pi5342;// level 0
assign po5342 = pi5392;// level 0
assign po5343 = pi5224;// level 0
assign po5344 = pi5209;// level 0
assign po5345 = pi5269;// level 0
assign po5346 = pi5416;// level 0
assign po5347 = pi5403;// level 0
assign po5348 = pi5197;// level 0
assign po5349 = pi5235;// level 0
assign po5350 = pi5243;// level 0
assign po5351 = pi5272;// level 0
assign po5352 = pi5264;// level 0
assign po5353 = pi5270;// level 0
assign po5354 = pi5260;// level 0
assign po5355 = pi5247;// level 0
assign po5356 = pi5271;// level 0
assign po5357 = pi5276;// level 0
assign po5358 = pi5261;// level 0
assign po5359 = pi5241;// level 0
assign po5360 = pi5236;// level 0
assign po5361 = pi5227;// level 0
assign po5362 = pi5237;// level 0
assign po5363 = pi5225;// level 0
assign po5364 = pi5263;// level 0
assign po5365 = pi5279;// level 0
assign po5366 = pi5198;// level 0
assign po5367 = pi5244;// level 0
assign po5368 = pi5228;// level 0
assign po5369 = pi5199;// level 0
assign po5370 = pi5258;// level 0
assign po5371 = pi5239;// level 0
assign po5372 = pi5218;// level 0
assign po5373 = pi5400;// level 0
assign po5374 = pi5408;// level 0
assign po5375 = pi5221;// level 0
assign po5376 = pi5200;// level 0
assign po5377 = pi5256;// level 0
assign po5378 = pi5222;// level 0
assign po5379 = pi5232;// level 0
assign po5380 = pi5251;// level 0
assign po5381 = pi5396;// level 0
assign po5382 = pi5398;// level 0
assign po5383 = pi5273;// level 0
assign po5384 = pi5304;// level 0
assign po5385 = pi5415;// level 0
assign po5386 = pi5401;// level 0
assign po5387 = pi5275;// level 0
assign po5388 = pi5248;// level 0
assign po5389 = pi5257;// level 0
assign po5390 = pi5240;// level 0
assign po5391 = pi5249;// level 0
assign po5392 = pi5274;// level 0
assign po5393 = pi5226;// level 0
assign po5394 = pi5407;// level 0
assign po5395 = pi5259;// level 0
assign po5396 = pi5219;// level 0
assign po5397 = pi5242;// level 0
assign po5398 = pi5231;// level 0
assign po5399 = pi5268;// level 0
assign po5400 = pi5254;// level 0
assign po5401 = pi5201;// level 0
assign po5402 = pi5265;// level 0
assign po5403 = pi5234;// level 0
assign po5404 = pi5233;// level 0
assign po5405 = pi5230;// level 0
assign po5406 = pi5223;// level 0
assign po5407 = pi5229;// level 0
assign po5408 = pi5430;// level 0
assign po5409 = pi5347;// level 0
assign po5410 = pi5294;// level 0
assign po5411 = pi5429;// level 0
assign po5412 = pi5434;// level 0
assign po5413 = pi5534;// level 0
assign po5414 = pi5326;// level 0
assign po5415 = pi5439;// level 0
assign po5416 = pi5282;// level 0
assign po5417 = pi5440;// level 0
assign po5418 = pi5402;// level 0
assign po5419 = pi5438;// level 0
assign po5420 = pi5399;// level 0
assign po5421 = pi5431;// level 0
assign po5422 = pi5442;// level 0
assign po5423 = pi5328;// level 0
assign po5424 = pi5441;// level 0
assign po5425 = pi5437;// level 0
assign po5426 = pi5436;// level 0
assign po5427 = pi5371;// level 0
assign po5428 = pi5373;// level 0
assign po5429 = pi5353;// level 0
assign po5430 = pi5423;// level 0
assign po5431 = pi5381;// level 0
assign po5432 = pi5446;// level 0
assign po5433 = pi5459;// level 0
assign po5434 = pi5450;// level 0
assign po5435 = pi5455;// level 0
assign po5436 = pi5461;// level 0
assign po5437 = pi5460;// level 0
assign po5438 = pi5456;// level 0
assign po5439 = pi5506;// level 0
assign po5440 = pi5458;// level 0
assign po5441 = pi5447;// level 0
assign po5442 = pi5454;// level 0
assign po5443 = pi5464;// level 0
assign po5444 = pi5453;// level 0
assign po5445 = pi5452;// level 0
assign po5446 = pi5585;// level 0
assign po5447 = pi5475;// level 0
assign po5448 = pi5372;// level 0
assign po5449 = pi5382;// level 0
assign po5450 = pi5406;// level 0
assign po5451 = pi5388;// level 0
assign po5452 = pi5374;// level 0
assign po5453 = pi5391;// level 0
assign po5454 = pi5424;// level 0
assign po5455 = pi5375;// level 0
assign po5456 = pi5331;// level 0
assign po5457 = pi5393;// level 0
assign po5458 = pi5413;// level 0
assign po5459 = pi5370;// level 0
assign po5460 = pi5412;// level 0
assign po5461 = pi5384;// level 0
assign po5462 = pi5425;// level 0
assign po5463 = pi5410;// level 0
assign po5464 = pi5329;// level 0
assign po5465 = pi5395;// level 0
assign po5466 = pi5411;// level 0
assign po5467 = pi5380;// level 0
assign po5468 = pi5465;// level 0
assign po5469 = pi5420;// level 0
assign po5470 = pi5361;// level 0
assign po5471 = pi5419;// level 0
assign po5472 = pi5417;// level 0
assign po5473 = pi5390;// level 0
assign po5474 = pi5394;// level 0
assign po5475 = pi5510;// level 0
assign po5476 = pi5351;// level 0
assign po5477 = pi5369;// level 0
assign po5478 = pi5404;// level 0
assign po5479 = pi5354;// level 0
assign po5480 = pi5443;// level 0
assign po5481 = pi5514;// level 0
assign po5482 = pi5502;// level 0
assign po5483 = pi5509;// level 0
assign po5484 = pi5377;// level 0
assign po5485 = pi5513;// level 0
assign po5486 = pi5409;// level 0
assign po5487 = pi5389;// level 0
assign po5488 = pi5367;// level 0
assign po5489 = pi5397;// level 0
assign po5490 = pi5366;// level 0
assign po5491 = pi5386;// level 0
assign po5492 = pi5511;// level 0
assign po5493 = pi5368;// level 0
assign po5494 = pi5357;// level 0
assign po5495 = pi5364;// level 0
assign po5496 = pi5385;// level 0
assign po5497 = pi5405;// level 0
assign po5498 = pi5365;// level 0
assign po5499 = pi5387;// level 0
assign po5500 = pi5360;// level 0
assign po5501 = pi5359;// level 0
assign po5502 = pi5379;// level 0
assign po5503 = pi5383;// level 0
assign po5504 = pi5362;// level 0
assign po5505 = pi5376;// level 0
assign po5506 = pi5414;// level 0
assign po5507 = pi5339;// level 0
assign po5508 = pi5355;// level 0
assign po5509 = pi5363;// level 0
assign po5510 = pi5607;// level 0
assign po5511 = pi5584;// level 0
assign po5512 = pi5543;// level 0
assign po5513 = pi5562;// level 0
assign po5514 = pi5538;// level 0
assign po5515 = pi5537;// level 0
assign po5516 = pi5539;// level 0
assign po5517 = pi5535;// level 0
assign po5518 = pi5547;// level 0
assign po5519 = pi5548;// level 0
assign po5520 = pi5583;// level 0
assign po5521 = pi5545;// level 0
assign po5522 = pi5533;// level 0
assign po5523 = pi5560;// level 0
assign po5524 = pi5536;// level 0
assign po5525 = pi5542;// level 0
assign po5526 = pi5449;// level 0
assign po5527 = pi5552;// level 0
assign po5528 = pi5530;// level 0
assign po5529 = pi5569;// level 0
assign po5530 = pi5586;// level 0
assign po5531 = pi5587;// level 0
assign po5532 = pi5566;// level 0
assign po5533 = pi5581;// level 0
assign po5534 = pi5563;// level 0
assign po5535 = pi5564;// level 0
assign po5536 = pi5578;// level 0
assign po5537 = pi5550;// level 0
assign po5538 = pi5555;// level 0
assign po5539 = pi5574;// level 0
assign po5540 = pi5575;// level 0
assign po5541 = pi5582;// level 0
assign po5542 = pi5505;// level 0
assign po5543 = pi5553;// level 0
assign po5544 = pi5576;// level 0
assign po5545 = pi5573;// level 0
assign po5546 = pi5579;// level 0
assign po5547 = pi5554;// level 0
assign po5548 = pi5571;// level 0
assign po5549 = pi5580;// level 0
assign po5550 = pi5577;// level 0
assign po5551 = pi5559;// level 0
assign po5552 = pi5558;// level 0
assign po5553 = pi5557;// level 0
assign po5554 = pi5556;// level 0
assign po5555 = pi5568;// level 0
assign po5556 = pi5435;// level 0
assign po5557 = pi5544;// level 0
assign po5558 = pi5663;// level 0
assign po5559 = pi5527;// level 0
assign po5560 = pi5619;// level 0
assign po5561 = pi5526;// level 0
assign po5562 = ~pi5546;// level 0
assign po5563 = pi5606;// level 0
assign po5564 = pi5626;// level 0
assign po5565 = pi5608;// level 0
assign po5566 = pi5541;// level 0
assign po5567 = pi5532;// level 0
assign po5568 = pi5624;// level 0
assign po5569 = pi5630;// level 0
assign po5570 = pi5631;// level 0
assign po5571 = pi5616;// level 0
assign po5572 = pi5641;// level 0
assign po5573 = pi5662;// level 0
assign po5574 = pi5625;// level 0
assign po5575 = pi5636;// level 0
assign po5576 = pi5549;// level 0
assign po5577 = pi5668;// level 0
assign po5578 = pi5609;// level 0
assign po5579 = pi5598;// level 0
assign po5580 = pi5658;// level 0
assign po5581 = pi5504;// level 0
assign po5582 = pi5650;// level 0
assign po5583 = pi5472;// level 0
assign po5584 = pi5468;// level 0
assign po5585 = pi5665;// level 0
assign po5586 = pi5703;// level 0
assign po5587 = pi5503;// level 0
assign po5588 = pi5634;// level 0
assign po5589 = pi5491;// level 0
assign po5590 = pi5500;// level 0
assign po5591 = pi5496;// level 0
assign po5592 = pi5477;// level 0
assign po5593 = pi5525;// level 0
assign po5594 = pi5470;// level 0
assign po5595 = pi5501;// level 0
assign po5596 = pi5490;// level 0
assign po5597 = pi5489;// level 0
assign po5598 = pi5469;// level 0
assign po5599 = pi5462;// level 0
assign po5600 = pi5507;// level 0
assign po5601 = pi5520;// level 0
assign po5602 = pi5494;// level 0
assign po5603 = pi5515;// level 0
assign po5604 = pi5482;// level 0
assign po5605 = pi5480;// level 0
assign po5606 = pi5445;// level 0
assign po5607 = pi5483;// level 0
assign po5608 = pi5618;// level 0
assign po5609 = pi5516;// level 0
assign po5610 = pi5484;// level 0
assign po5611 = pi5474;// level 0
assign po5612 = pi5519;// level 0
assign po5613 = pi5528;// level 0
assign po5614 = pi5448;// level 0
assign po5615 = pi5488;// level 0
assign po5616 = pi5522;// level 0
assign po5617 = pi5485;// level 0
assign po5618 = pi5466;// level 0
assign po5619 = pi5521;// level 0
assign po5620 = pi5498;// level 0
assign po5621 = pi5495;// level 0
assign po5622 = pi5666;// level 0
assign po5623 = pi5451;// level 0
assign po5624 = pi5518;// level 0
assign po5625 = pi5486;// level 0
assign po5626 = pi5664;// level 0
assign po5627 = pi5479;// level 0
assign po5628 = pi5671;// level 0
assign po5629 = pi5561;// level 0
assign po5630 = pi5669;// level 0
assign po5631 = pi5661;// level 0
assign po5632 = pi5572;// level 0
assign po5633 = pi5677;// level 0
assign po5634 = pi5463;// level 0
assign po5635 = ~pi5567;// level 0
assign po5636 = pi5529;// level 0
assign po5637 = pi5672;// level 0
assign po5638 = pi5667;// level 0
assign po5639 = pi5492;// level 0
assign po5640 = pi5471;// level 0
assign po5641 = pi5524;// level 0
assign po5642 = pi5473;// level 0
assign po5643 = pi5481;// level 0
assign po5644 = pi5493;// level 0
assign po5645 = pi5588;// level 0
assign po5646 = pi5508;// level 0
assign po5647 = pi5478;// level 0
assign po5648 = pi5628;// level 0
assign po5649 = pi5444;// level 0
assign po5650 = pi5517;// level 0
assign po5651 = pi5633;// level 0
assign po5652 = pi5540;// level 0
assign po5653 = pi5457;// level 0
assign po5654 = pi5487;// level 0
assign po5655 = pi5476;// level 0
assign po5656 = pi5674;// level 0
assign po5657 = pi5694;// level 0
assign po5658 = pi5692;// level 0
assign po5659 = pi5687;// level 0
assign po5660 = pi5670;// level 0
assign po5661 = ~w61744;// level 14
assign po5662 = pi5693;// level 0
assign po5663 = pi5690;// level 0
assign po5664 = pi5699;// level 0
assign po5665 = pi5704;// level 0
assign po5666 = pi5698;// level 0
assign po5667 = pi5706;// level 0
assign po5668 = pi5695;// level 0
assign po5669 = pi5570;// level 0
assign po5670 = pi5565;// level 0
assign po5671 = pi5697;// level 0
assign po5672 = pi5701;// level 0
assign po5673 = pi5696;// level 0
assign po5674 = pi5591;// level 0
assign po5675 = pi5610;// level 0
assign po5676 = w61777;// level 14
assign po5677 = pi5738;// level 0
assign po5678 = pi5644;// level 0
assign po5679 = pi5747;// level 0
assign po5680 = pi5781;// level 0
assign po5681 = pi5604;// level 0
assign po5682 = pi5746;// level 0
assign po5683 = pi5741;// level 0
assign po5684 = pi5723;// level 0
assign po5685 = pi5735;// level 0
assign po5686 = pi5740;// level 0
assign po5687 = pi5680;// level 0
assign po5688 = pi5736;// level 0
assign po5689 = pi5737;// level 0
assign po5690 = pi5727;// level 0
assign po5691 = pi5734;// level 0
assign po5692 = pi5635;// level 0
assign po5693 = pi5649;// level 0
assign po5694 = pi5732;// level 0
assign po5695 = w61869;// level 14
assign po5696 = pi5657;// level 0
assign po5697 = pi5750;// level 0
assign po5698 = pi5640;// level 0
assign po5699 = pi5659;// level 0
assign po5700 = pi5652;// level 0
assign po5701 = pi5648;// level 0
assign po5702 = pi5600;// level 0
assign po5703 = pi5601;// level 0
assign po5704 = pi5681;// level 0
assign po5705 = w61962;// level 14
assign po5706 = pi5622;// level 0
assign po5707 = pi5639;// level 0
assign po5708 = pi5612;// level 0
assign po5709 = pi5593;// level 0
assign po5710 = pi5673;// level 0
assign po5711 = pi5642;// level 0
assign po5712 = pi5654;// level 0
assign po5713 = pi5637;// level 0
assign po5714 = pi5653;// level 0
assign po5715 = pi5595;// level 0
assign po5716 = pi5632;// level 0
assign po5717 = pi5660;// level 0
assign po5718 = pi5638;// level 0
assign po5719 = pi5602;// level 0
assign po5720 = pi5617;// level 0
assign po5721 = pi5597;// level 0
assign po5722 = pi5605;// level 0
assign po5723 = pi5678;// level 0
assign po5724 = pi5589;// level 0
assign po5725 = pi5623;// level 0
assign po5726 = pi5590;// level 0
assign po5727 = ~pi5684;// level 0
assign po5728 = pi5655;// level 0
assign po5729 = pi5748;// level 0
assign po5730 = pi5643;// level 0
assign po5731 = pi5682;// level 0
assign po5732 = pi5779;// level 0
assign po5733 = pi5676;// level 0
assign po5734 = pi5683;// level 0
assign po5735 = pi5700;// level 0
assign po5736 = pi5722;// level 0
assign po5737 = pi5679;// level 0
assign po5738 = pi5675;// level 0
assign po5739 = pi5784;// level 0
assign po5740 = pi5782;// level 0
assign po5741 = pi5783;// level 0
assign po5742 = w62055;// level 14
assign po5743 = pi5780;// level 0
assign po5744 = pi5785;// level 0
assign po5745 = pi5627;// level 0
assign po5746 = pi5594;// level 0
assign po5747 = pi5621;// level 0
assign po5748 = pi5645;// level 0
assign po5749 = pi5614;// level 0
assign po5750 = pi5596;// level 0
assign po5751 = pi5592;// level 0
assign po5752 = pi5651;// level 0
assign po5753 = pi5749;// level 0
assign po5754 = pi5611;// level 0
assign po5755 = pi5620;// level 0
assign po5756 = pi5615;// level 0
assign po5757 = pi5656;// level 0
assign po5758 = pi5629;// level 0
assign po5759 = pi5613;// level 0
assign po5760 = pi5814;// level 0
assign po5761 = pi5841;// level 0
assign po5762 = pi5810;// level 0
assign po5763 = pi5800;// level 0
assign po5764 = ~w62150;// level 14
assign po5765 = pi5743;// level 0
assign po5766 = pi5807;// level 0
assign po5767 = pi5811;// level 0
assign po5768 = pi5801;// level 0
assign po5769 = pi5806;// level 0
assign po5770 = pi5839;// level 0
assign po5771 = pi5812;// level 0
assign po5772 = pi5688;// level 0
assign po5773 = pi5802;// level 0
assign po5774 = pi5808;// level 0
assign po5775 = pi5794;// level 0
assign po5776 = pi5793;// level 0
assign po5777 = pi5791;// level 0
assign po5778 = pi5803;// level 0
assign po5779 = pi5797;// level 0
assign po5780 = w62183;// level 14
assign po5781 = pi5805;// level 0
assign po5782 = pi5745;// level 0
assign po5783 = pi5840;// level 0
assign po5784 = pi5824;// level 0
assign po5785 = pi5837;// level 0
assign po5786 = pi5820;// level 0
assign po5787 = pi5792;// level 0
assign po5788 = pi5829;// level 0
assign po5789 = pi5832;// level 0
assign po5790 = pi5823;// level 0
assign po5791 = pi5818;// level 0
assign po5792 = pi5804;// level 0
assign po5793 = pi5836;// level 0
assign po5794 = pi5828;// level 0
assign po5795 = pi5705;// level 0
assign po5796 = pi5830;// level 0
assign po5797 = pi5833;// level 0
assign po5798 = pi5827;// level 0
assign po5799 = pi5822;// level 0
assign po5800 = pi5702;// level 0
assign po5801 = pi5843;// level 0
assign po5802 = pi5831;// level 0
assign po5803 = pi5826;// level 0
assign po5804 = pi5825;// level 0
assign po5805 = pi5838;// level 0
assign po5806 = pi5834;// level 0
assign po5807 = pi5842;// level 0
assign po5808 = pi5817;// level 0
assign po5809 = pi5796;// level 0
assign po5810 = pi5819;// level 0
assign po5811 = pi5815;// level 0
assign po5812 = pi5821;// level 0
assign po5813 = pi5685;// level 0
assign po5814 = pi5686;// level 0
assign po5815 = w62276;// level 14
assign po5816 = ~w62314;// level 15
assign po5817 = ~w62340;// level 14
assign po5818 = pi5909;// level 0
assign po5819 = pi5708;// level 0
assign po5820 = pi5773;// level 0
assign po5821 = pi5728;// level 0
assign po5822 = pi5719;// level 0
assign po5823 = pi5761;// level 0
assign po5824 = pi5718;// level 0
assign po5825 = pi5726;// level 0
assign po5826 = pi5790;// level 0
assign po5827 = pi5721;// level 0
assign po5828 = w62355;// level 14
assign po5829 = pi5856;// level 0
assign po5830 = pi5709;// level 0
assign po5831 = pi5716;// level 0
assign po5832 = pi5768;// level 0
assign po5833 = pi5888;// level 0
assign po5834 = pi5769;// level 0
assign po5835 = pi5766;// level 0
assign po5836 = pi5884;// level 0
assign po5837 = w62444;// level 14
assign po5838 = pi5879;// level 0
assign po5839 = pi5799;// level 0
assign po5840 = pi5730;// level 0
assign po5841 = pi5714;// level 0
assign po5842 = pi5786;// level 0
assign po5843 = pi5752;// level 0
assign po5844 = pi5758;// level 0
assign po5845 = pi5755;// level 0
assign po5846 = pi5874;// level 0
assign po5847 = pi5753;// level 0
assign po5848 = pi5862;// level 0
assign po5849 = pi5871;// level 0
assign po5850 = pi5754;// level 0
assign po5851 = pi5772;// level 0
assign po5852 = pi5789;// level 0
assign po5853 = pi5707;// level 0
assign po5854 = pi5877;// level 0
assign po5855 = pi5849;// level 0
assign po5856 = pi5873;// level 0
assign po5857 = pi5765;// level 0
assign po5858 = pi5742;// level 0
assign po5859 = pi5763;// level 0
assign po5860 = pi5733;// level 0
assign po5861 = pi5844;// level 0
assign po5862 = pi5762;// level 0
assign po5863 = pi5910;// level 0
assign po5864 = pi5725;// level 0
assign po5865 = pi5757;// level 0
assign po5866 = pi5891;// level 0
assign po5867 = pi5776;// level 0
assign po5868 = pi5744;// level 0
assign po5869 = pi5777;// level 0
assign po5870 = pi5731;// level 0
assign po5871 = pi5878;// level 0
assign po5872 = pi5770;// level 0
assign po5873 = pi5712;// level 0
assign po5874 = pi5774;// level 0
assign po5875 = pi5739;// level 0
assign po5876 = pi5895;// level 0
assign po5877 = pi5798;// level 0
assign po5878 = pi5713;// level 0
assign po5879 = pi5767;// level 0
assign po5880 = ~w62476;// level 14
assign po5881 = pi5764;// level 0
assign po5882 = pi5720;// level 0
assign po5883 = pi5788;// level 0
assign po5884 = pi5724;// level 0
assign po5885 = pi5751;// level 0
assign po5886 = pi5759;// level 0
assign po5887 = pi5787;// level 0
assign po5888 = w62503;// level 14
assign po5889 = pi5717;// level 0
assign po5890 = pi5778;// level 0
assign po5891 = pi5929;// level 0
assign po5892 = pi5809;// level 0
assign po5893 = pi5921;// level 0
assign po5894 = pi5916;// level 0
assign po5895 = pi5919;// level 0
assign po5896 = ~pi5835;// level 0
assign po5897 = pi5918;// level 0
assign po5898 = pi5881;// level 0
assign po5899 = pi5920;// level 0
assign po5900 = pi5883;// level 0
assign po5901 = pi5922;// level 0
assign po5902 = pi5913;// level 0
assign po5903 = pi5710;// level 0
assign po5904 = w62531;// level 14
assign po5905 = pi5911;// level 0
assign po5906 = pi5715;// level 0
assign po5907 = pi5923;// level 0
assign po5908 = pi5771;// level 0
assign po5909 = pi5760;// level 0
assign po5910 = pi5729;// level 0
assign po5911 = pi5711;// level 0
assign po5912 = pi5775;// level 0
assign po5913 = pi5756;// level 0
assign po5914 = ~w62560;// level 14
assign po5915 = pi5944;// level 0
assign po5916 = pi5934;// level 0
assign po5917 = pi5932;// level 0
assign po5918 = pi5936;// level 0
assign po5919 = pi5813;// level 0
assign po5920 = w62637;// level 14
assign po5921 = pi5795;// level 0
assign po5922 = w62659;// level 14
assign po5923 = w62696;// level 14
assign po5924 = w62715;// level 14
assign po5925 = pi5947;// level 0
assign po5926 = pi5940;// level 0
assign po5927 = pi5942;// level 0
assign po5928 = pi5946;// level 0
assign po5929 = pi5938;// level 0
assign po5930 = pi5937;// level 0
assign po5931 = pi5943;// level 0
assign po5932 = pi5941;// level 0
assign po5933 = w62737;// level 14
assign po5934 = pi5816;// level 0
assign po5935 = pi5945;// level 0
assign po5936 = pi5948;// level 0
assign po5937 = pi5887;// level 0
assign po5938 = pi5861;// level 0
assign po5939 = pi5925;// level 0
assign po5940 = pi5889;// level 0
assign po5941 = pi5885;// level 0
assign po5942 = pi5864;// level 0
assign po5943 = pi5872;// level 0
assign po5944 = pi5869;// level 0
assign po5945 = pi5880;// level 0
assign po5946 = pi5852;// level 0
assign po5947 = pi5894;// level 0
assign po5948 = pi5846;// level 0
assign po5949 = pi5853;// level 0
assign po5950 = pi5892;// level 0
assign po5951 = pi5890;// level 0
assign po5952 = pi5951;// level 0
assign po5953 = pi5956;// level 0
assign po5954 = pi5851;// level 0
assign po5955 = pi6010;// level 0
assign po5956 = pi5845;// level 0
assign po5957 = pi6007;// level 0
assign po5958 = pi5901;// level 0
assign po5959 = pi5903;// level 0
assign po5960 = pi5899;// level 0
assign po5961 = pi5866;// level 0
assign po5962 = pi5963;// level 0
assign po5963 = pi6002;// level 0
assign po5964 = pi6016;// level 0
assign po5965 = pi5952;// level 0
assign po5966 = pi5882;// level 0
assign po5967 = pi6017;// level 0
assign po5968 = pi5931;// level 0
assign po5969 = pi5886;// level 0
assign po5970 = pi5933;// level 0
assign po5971 = pi5965;// level 0
assign po5972 = pi6011;// level 0
assign po5973 = pi5991;// level 0
assign po5974 = pi5867;// level 0
assign po5975 = pi5964;// level 0
assign po5976 = pi5960;// level 0
assign po5977 = pi6025;// level 0
assign po5978 = w62761;// level 14
assign po5979 = w62792;// level 14
assign po5980 = w62820;// level 14
assign po5981 = pi5865;// level 0
assign po5982 = pi5847;// level 0
assign po5983 = pi5855;// level 0
assign po5984 = pi5860;// level 0
assign po5985 = pi5904;// level 0
assign po5986 = pi5870;// level 0
assign po5987 = pi5930;// level 0
assign po5988 = pi5905;// level 0
assign po5989 = pi5854;// level 0
assign po5990 = pi5908;// level 0
assign po5991 = pi5897;// level 0
assign po5992 = pi5926;// level 0
assign po5993 = pi5896;// level 0
assign po5994 = pi5928;// level 0
assign po5995 = pi5848;// level 0
assign po5996 = pi5858;// level 0
assign po5997 = pi5898;// level 0
assign po5998 = pi5893;// level 0
assign po5999 = pi5914;// level 0
assign po6000 = pi5907;// level 0
assign po6001 = pi5863;// level 0
assign po6002 = pi5924;// level 0
assign po6003 = pi5900;// level 0
assign po6004 = pi5927;// level 0
assign po6005 = pi5859;// level 0
assign po6006 = pi5876;// level 0
assign po6007 = pi5850;// level 0
assign po6008 = pi5906;// level 0
assign po6009 = pi5917;// level 0
assign po6010 = pi5939;// level 0
assign po6011 = pi5950;// level 0
assign po6012 = pi6013;// level 0
assign po6013 = pi6015;// level 0
assign po6014 = pi6012;// level 0
assign po6015 = pi5915;// level 0
assign po6016 = pi5868;// level 0
assign po6017 = pi5912;// level 0
assign po6018 = pi5875;// level 0
assign po6019 = pi5857;// level 0
assign po6020 = pi5902;// level 0
assign po6021 = pi6043;// level 0
assign po6022 = pi6058;// level 0
assign po6023 = pi5935;// level 0
assign po6024 = pi6036;// level 0
assign po6025 = ~w62839;// level 14
assign po6026 = pi6050;// level 0
assign po6027 = pi6029;// level 0
assign po6028 = ~w62863;// level 14
assign po6029 = pi6042;// level 0
assign po6030 = pi6044;// level 0
assign po6031 = pi6032;// level 0
assign po6032 = pi6037;// level 0
assign po6033 = pi6068;// level 0
assign po6034 = pi6073;// level 0
assign po6035 = ~w62885;// level 14
assign po6036 = pi6047;// level 0
assign po6037 = pi6074;// level 0
assign po6038 = pi6045;// level 0
assign po6039 = pi6033;// level 0
assign po6040 = pi6030;// level 0
assign po6041 = pi6075;// level 0
assign po6042 = pi6048;// level 0
assign po6043 = w62907;// level 14
assign po6044 = pi6034;// level 0
assign po6045 = pi6038;// level 0
assign po6046 = pi6057;// level 0
assign po6047 = pi6035;// level 0
assign po6048 = pi6084;// level 0
assign po6049 = pi6041;// level 0
assign po6050 = pi6060;// level 0
assign po6051 = pi6031;// level 0
assign po6052 = pi6082;// level 0
assign po6053 = pi6071;// level 0
assign po6054 = pi6026;// level 0
assign po6055 = pi6056;// level 0
assign po6056 = pi6076;// level 0
assign po6057 = pi6078;// level 0
assign po6058 = pi6053;// level 0
assign po6059 = pi6062;// level 0
assign po6060 = pi6080;// level 0
assign po6061 = pi6066;// level 0
assign po6062 = pi6059;// level 0
assign po6063 = pi6051;// level 0
assign po6064 = pi6069;// level 0
assign po6065 = pi6063;// level 0
assign po6066 = pi6070;// level 0
assign po6067 = pi6081;// level 0
assign po6068 = pi6052;// level 0
assign po6069 = pi6046;// level 0
assign po6070 = pi6064;// level 0
assign po6071 = w62926;// level 14
assign po6072 = pi6067;// level 0
assign po6073 = pi6027;// level 0
assign po6074 = pi6139;// level 0
assign po6075 = pi6005;// level 0
assign po6076 = pi5992;// level 0
assign po6077 = pi6001;// level 0
assign po6078 = pi5969;// level 0
assign po6079 = pi6089;// level 0
assign po6080 = pi5961;// level 0
assign po6081 = pi5997;// level 0
assign po6082 = pi5987;// level 0
assign po6083 = pi6019;// level 0
assign po6084 = pi5959;// level 0
assign po6085 = pi5989;// level 0
assign po6086 = w62945;// level 15
assign po6087 = pi5966;// level 0
assign po6088 = pi6022;// level 0
assign po6089 = pi6021;// level 0
assign po6090 = pi5995;// level 0
assign po6091 = pi6024;// level 0
assign po6092 = pi6040;// level 0
assign po6093 = pi5974;// level 0
assign po6094 = pi5990;// level 0
assign po6095 = pi5970;// level 0
assign po6096 = pi5980;// level 0
assign po6097 = pi5982;// level 0
assign po6098 = pi5993;// level 0
assign po6099 = pi5958;// level 0
assign po6100 = pi5967;// level 0
assign po6101 = pi6093;// level 0
assign po6102 = pi6023;// level 0
assign po6103 = pi6094;// level 0
assign po6104 = pi6142;// level 0
assign po6105 = pi5978;// level 0
assign po6106 = pi6009;// level 0
assign po6107 = pi6079;// level 0
assign po6108 = pi6018;// level 0
assign po6109 = pi6124;// level 0
assign po6110 = pi5979;// level 0
assign po6111 = pi6121;// level 0
assign po6112 = pi6158;// level 0
assign po6113 = pi6144;// level 0
assign po6114 = pi6072;// level 0
assign po6115 = pi5976;// level 0
assign po6116 = pi5957;// level 0
assign po6117 = pi6008;// level 0
assign po6118 = w62961;// level 14
assign po6119 = pi6014;// level 0
assign po6120 = pi5994;// level 0
assign po6121 = pi6088;// level 0
assign po6122 = pi5968;// level 0
assign po6123 = pi5962;// level 0
assign po6124 = pi6003;// level 0
assign po6125 = w62983;// level 14
assign po6126 = pi5973;// level 0
assign po6127 = pi5985;// level 0
assign po6128 = pi6020;// level 0
assign po6129 = pi5984;// level 0
assign po6130 = pi5954;// level 0
assign po6131 = pi5972;// level 0
assign po6132 = pi5975;// level 0
assign po6133 = pi5971;// level 0
assign po6134 = pi5981;// level 0
assign po6135 = pi6006;// level 0
assign po6136 = pi5988;// level 0
assign po6137 = pi5999;// level 0
assign po6138 = pi5986;// level 0
assign po6139 = pi6148;// level 0
assign po6140 = pi6039;// level 0
assign po6141 = pi6159;// level 0
assign po6142 = pi5983;// level 0
assign po6143 = pi6061;// level 0
assign po6144 = pi6004;// level 0
assign po6145 = pi6150;// level 0
assign po6146 = pi6133;// level 0
assign po6147 = pi6154;// level 0
assign po6148 = pi6147;// level 0
assign po6149 = pi5949;// level 0
assign po6150 = pi6152;// level 0
assign po6151 = pi6143;// level 0
assign po6152 = pi6149;// level 0
assign po6153 = pi6151;// level 0
assign po6154 = pi5955;// level 0
assign po6155 = pi5977;// level 0
assign po6156 = pi5998;// level 0
assign po6157 = pi6000;// level 0
assign po6158 = pi5996;// level 0
assign po6159 = pi6153;// level 0
assign po6160 = pi5953;// level 0
assign po6161 = pi6146;// level 0
assign po6162 = pi6165;// level 0
assign po6163 = pi6086;// level 0
assign po6164 = pi6167;// level 0
assign po6165 = pi6166;// level 0
assign po6166 = pi6028;// level 0
assign po6167 = pi6077;// level 0
assign po6168 = pi6049;// level 0
assign po6169 = pi6055;// level 0
assign po6170 = pi6169;// level 0
assign po6171 = pi6083;// level 0
assign po6172 = pi6168;// level 0
assign po6173 = pi6174;// level 0
assign po6174 = pi6173;// level 0
assign po6175 = pi6175;// level 0
assign po6176 = pi6176;// level 0
assign po6177 = pi6065;// level 0
assign po6178 = pi6054;// level 0
assign po6179 = pi6259;// level 0
assign po6180 = pi6258;// level 0
assign po6181 = pi6256;// level 0
assign po6182 = pi6227;// level 0
assign po6183 = pi6107;// level 0
assign po6184 = pi6162;// level 0
assign po6185 = pi6120;// level 0
assign po6186 = pi6245;// level 0
assign po6187 = pi6131;// level 0
assign po6188 = pi6100;// level 0
assign po6189 = pi6110;// level 0
assign po6190 = pi6232;// level 0
assign po6191 = pi6119;// level 0
assign po6192 = pi6116;// level 0
assign po6193 = pi6234;// level 0
assign po6194 = pi6228;// level 0
assign po6195 = pi6255;// level 0
assign po6196 = pi6097;// level 0
assign po6197 = pi6108;// level 0
assign po6198 = pi6122;// level 0
assign po6199 = pi6087;// level 0
assign po6200 = pi6134;// level 0
assign po6201 = pi6125;// level 0
assign po6202 = pi6099;// level 0
assign po6203 = pi6114;// level 0
assign po6204 = pi6090;// level 0
assign po6205 = pi6104;// level 0
assign po6206 = pi6155;// level 0
assign po6207 = pi6128;// level 0
assign po6208 = pi6117;// level 0
assign po6209 = pi6130;// level 0
assign po6210 = pi6160;// level 0
assign po6211 = pi6106;// level 0
assign po6212 = pi6157;// level 0
assign po6213 = pi6109;// level 0
assign po6214 = pi6096;// level 0
assign po6215 = pi6115;// level 0
assign po6216 = pi6129;// level 0
assign po6217 = pi6127;// level 0
assign po6218 = pi6091;// level 0
assign po6219 = pi6101;// level 0
assign po6220 = pi6113;// level 0
assign po6221 = pi6244;// level 0
assign po6222 = pi6095;// level 0
assign po6223 = pi6135;// level 0
assign po6224 = pi6140;// level 0
assign po6225 = pi6103;// level 0
assign po6226 = pi6141;// level 0
assign po6227 = pi6112;// level 0
assign po6228 = pi6156;// level 0
assign po6229 = pi6098;// level 0
assign po6230 = pi6085;// level 0
assign po6231 = pi6132;// level 0
assign po6232 = pi6183;// level 0
assign po6233 = pi6138;// level 0
assign po6234 = pi6137;// level 0
assign po6235 = pi6163;// level 0
assign po6236 = pi6102;// level 0
assign po6237 = pi6242;// level 0
assign po6238 = pi6111;// level 0
assign po6239 = pi6123;// level 0
assign po6240 = pi6231;// level 0
assign po6241 = pi6179;// level 0
assign po6242 = pi6225;// level 0
assign po6243 = pi6233;// level 0
assign po6244 = pi6105;// level 0
assign po6245 = pi6257;// level 0
assign po6246 = pi6241;// level 0
assign po6247 = pi6188;// level 0
assign po6248 = pi6145;// level 0
assign po6249 = pi6092;// level 0
assign po6250 = pi6136;// level 0
assign po6251 = pi6161;// level 0
assign po6252 = pi6164;// level 0
assign po6253 = pi6118;// level 0
assign po6254 = pi6126;// level 0
assign po6255 = pi6243;// level 0
assign po6256 = pi6296;// level 0
assign po6257 = pi6311;// level 0
assign po6258 = pi6266;// level 0
assign po6259 = pi6262;// level 0
assign po6260 = pi6264;// level 0
assign po6261 = pi6260;// level 0
assign po6262 = pi6310;// level 0
assign po6263 = pi6172;// level 0
assign po6264 = pi6273;// level 0
assign po6265 = pi6281;// level 0
assign po6266 = pi6275;// level 0
assign po6267 = pi6170;// level 0
assign po6268 = pi6287;// level 0
assign po6269 = pi6240;// level 0
assign po6270 = pi6181;// level 0
assign po6271 = pi6280;// level 0
assign po6272 = pi6305;// level 0
assign po6273 = pi6279;// level 0
assign po6274 = pi6269;// level 0
assign po6275 = pi6171;// level 0
assign po6276 = pi6283;// level 0
assign po6277 = pi6246;// level 0
assign po6278 = pi6248;// level 0
assign po6279 = pi6286;// level 0
assign po6280 = pi6261;// level 0
assign po6281 = pi6289;// level 0
assign po6282 = pi6313;// level 0
assign po6283 = pi6282;// level 0
assign po6284 = pi6306;// level 0
assign po6285 = pi6277;// level 0
assign po6286 = pi6314;// level 0
assign po6287 = pi6300;// level 0
assign po6288 = pi6270;// level 0
assign po6289 = pi6285;// level 0
assign po6290 = pi6263;// level 0
assign po6291 = pi6304;// level 0
assign po6292 = pi6268;// level 0
assign po6293 = pi6288;// level 0
assign po6294 = pi6284;// level 0
assign po6295 = pi6278;// level 0
assign po6296 = pi6271;// level 0
assign po6297 = pi6290;// level 0
assign po6298 = pi6276;// level 0
assign po6299 = pi6294;// level 0
assign po6300 = pi6308;// level 0
assign po6301 = pi6292;// level 0
assign po6302 = pi6177;// level 0
assign po6303 = pi6302;// level 0
assign po6304 = pi6303;// level 0
assign po6305 = pi6301;// level 0
assign po6306 = pi6298;// level 0
assign po6307 = pi6309;// level 0
assign po6308 = pi6272;// level 0
assign po6309 = pi6247;// level 0
assign po6310 = pi6297;// level 0
assign po6311 = pi6291;// level 0
assign po6312 = pi6295;// level 0
assign po6313 = pi6293;// level 0
assign po6314 = pi6307;// level 0
assign po6315 = pi6194;// level 0
assign po6316 = pi6274;// level 0
assign po6317 = pi6199;// level 0
assign po6318 = pi6393;// level 0
assign po6319 = pi6384;// level 0
assign po6320 = pi6216;// level 0
assign po6321 = pi6250;// level 0
assign po6322 = pi6222;// level 0
assign po6323 = pi6366;// level 0
assign po6324 = pi6385;// level 0
assign po6325 = pi6226;// level 0
assign po6326 = pi6219;// level 0
assign po6327 = pi6211;// level 0
assign po6328 = pi6223;// level 0
assign po6329 = pi6193;// level 0
assign po6330 = pi6251;// level 0
assign po6331 = pi6195;// level 0
assign po6332 = pi6235;// level 0
assign po6333 = pi6205;// level 0
assign po6334 = pi6184;// level 0
assign po6335 = pi6230;// level 0
assign po6336 = pi6229;// level 0
assign po6337 = pi6237;// level 0
assign po6338 = pi6212;// level 0
assign po6339 = pi6238;// level 0
assign po6340 = pi6218;// level 0
assign po6341 = pi6224;// level 0
assign po6342 = pi6203;// level 0
assign po6343 = pi6221;// level 0
assign po6344 = pi6190;// level 0
assign po6345 = pi6239;// level 0
assign po6346 = pi6191;// level 0
assign po6347 = pi6249;// level 0
assign po6348 = pi6208;// level 0
assign po6349 = pi6186;// level 0
assign po6350 = pi6214;// level 0
assign po6351 = pi6320;// level 0
assign po6352 = pi6187;// level 0
assign po6353 = pi6196;// level 0
assign po6354 = pi6379;// level 0
assign po6355 = pi6189;// level 0
assign po6356 = pi6252;// level 0
assign po6357 = pi6207;// level 0
assign po6358 = pi6198;// level 0
assign po6359 = pi6206;// level 0
assign po6360 = pi6185;// level 0
assign po6361 = pi6180;// level 0
assign po6362 = pi6253;// level 0
assign po6363 = pi6372;// level 0
assign po6364 = pi6220;// level 0
assign po6365 = pi6200;// level 0
assign po6366 = pi6217;// level 0
assign po6367 = pi6178;// level 0
assign po6368 = pi6213;// level 0
assign po6369 = pi6392;// level 0
assign po6370 = pi6192;// level 0
assign po6371 = pi6202;// level 0
assign po6372 = pi6373;// level 0
assign po6373 = pi6367;// level 0
assign po6374 = pi6377;// level 0
assign po6375 = pi6365;// level 0
assign po6376 = pi6265;// level 0
assign po6377 = pi6374;// level 0
assign po6378 = pi6322;// level 0
assign po6379 = pi6312;// level 0
assign po6380 = ~pi6315;// level 0
assign po6381 = pi6319;// level 0
assign po6382 = pi6375;// level 0
assign po6383 = pi6369;// level 0
assign po6384 = pi6382;// level 0
assign po6385 = pi6210;// level 0
assign po6386 = pi6201;// level 0
assign po6387 = pi6182;// level 0
assign po6388 = pi6204;// level 0
assign po6389 = pi6368;// level 0
assign po6390 = pi6209;// level 0
assign po6391 = pi6197;// level 0
assign po6392 = pi6236;// level 0
assign po6393 = pi6215;// level 0
assign po6394 = pi6254;// level 0
assign po6395 = pi6381;// level 0
assign po6396 = pi6398;// level 0
assign po6397 = pi6400;// level 0
assign po6398 = pi6397;// level 0
assign po6399 = pi6402;// level 0
assign po6400 = ~pi6383;// level 0
assign po6401 = pi6267;// level 0
assign po6402 = pi6299;// level 0
assign po6403 = pi6399;// level 0
assign po6404 = pi6396;// level 0
assign po6405 = pi6395;// level 0
assign po6406 = pi6401;// level 0
assign po6407 = pi6464;// level 0
assign po6408 = pi6333;// level 0
assign po6409 = pi6407;// level 0
assign po6410 = pi6371;// level 0
assign po6411 = pi6480;// level 0
assign po6412 = pi6335;// level 0
assign po6413 = pi6469;// level 0
assign po6414 = pi6356;// level 0
assign po6415 = pi6344;// level 0
assign po6416 = pi6358;// level 0
assign po6417 = pi6359;// level 0
assign po6418 = pi6485;// level 0
assign po6419 = pi6345;// level 0
assign po6420 = pi6342;// level 0
assign po6421 = pi6350;// level 0
assign po6422 = pi6378;// level 0
assign po6423 = pi6394;// level 0
assign po6424 = pi6380;// level 0
assign po6425 = pi6326;// level 0
assign po6426 = pi6391;// level 0
assign po6427 = pi6390;// level 0
assign po6428 = pi6346;// level 0
assign po6429 = pi6351;// level 0
assign po6430 = pi6318;// level 0
assign po6431 = pi6325;// level 0
assign po6432 = pi6338;// level 0
assign po6433 = pi6364;// level 0
assign po6434 = pi6387;// level 0
assign po6435 = pi6330;// level 0
assign po6436 = pi6334;// level 0
assign po6437 = pi6389;// level 0
assign po6438 = pi6388;// level 0
assign po6439 = pi6340;// level 0
assign po6440 = pi6339;// level 0
assign po6441 = pi6341;// level 0
assign po6442 = pi6357;// level 0
assign po6443 = pi6316;// level 0
assign po6444 = pi6332;// level 0
assign po6445 = pi6353;// level 0
assign po6446 = pi6361;// level 0
assign po6447 = pi6355;// level 0
assign po6448 = pi6348;// level 0
assign po6449 = pi6354;// level 0
assign po6450 = pi6323;// level 0
assign po6451 = pi6328;// level 0
assign po6452 = pi6331;// level 0
assign po6453 = pi6349;// level 0
assign po6454 = pi6343;// level 0
assign po6455 = pi6467;// level 0
assign po6456 = pi6386;// level 0
assign po6457 = pi6483;// level 0
assign po6458 = pi6481;// level 0
assign po6459 = pi6362;// level 0
assign po6460 = pi6327;// level 0
assign po6461 = pi6419;// level 0
assign po6462 = pi6409;// level 0
assign po6463 = pi6466;// level 0
assign po6464 = pi6408;// level 0
assign po6465 = pi6317;// level 0
assign po6466 = pi6337;// level 0
assign po6467 = pi6324;// level 0
assign po6468 = pi6321;// level 0
assign po6469 = pi6363;// level 0
assign po6470 = pi6404;// level 0
assign po6471 = pi6472;// level 0
assign po6472 = pi6465;// level 0
assign po6473 = pi6468;// level 0
assign po6474 = pi6405;// level 0
assign po6475 = pi6460;// level 0
assign po6476 = pi6461;// level 0
assign po6477 = pi6421;// level 0
assign po6478 = pi6484;// level 0
assign po6479 = pi6360;// level 0
assign po6480 = pi6347;// level 0
assign po6481 = pi6336;// level 0
assign po6482 = pi6329;// level 0
assign po6483 = pi6370;// level 0
assign po6484 = pi6352;// level 0
assign po6485 = pi6463;// level 0
assign po6486 = pi6474;// level 0
assign po6487 = pi6403;// level 0
assign po6488 = pi6416;// level 0
assign po6489 = pi6376;// level 0
assign po6490 = pi6525;// level 0
assign po6491 = pi6521;// level 0
assign po6492 = pi6499;// level 0
assign po6493 = pi6517;// level 0
assign po6494 = pi6491;// level 0
assign po6495 = pi6470;// level 0
assign po6496 = pi6538;// level 0
assign po6497 = pi6495;// level 0
assign po6498 = pi6539;// level 0
assign po6499 = pi6501;// level 0
assign po6500 = pi6526;// level 0
assign po6501 = pi6536;// level 0
assign po6502 = pi6516;// level 0
assign po6503 = pi6542;// level 0
assign po6504 = pi6503;// level 0
assign po6505 = pi6537;// level 0
assign po6506 = pi6498;// level 0
assign po6507 = pi6530;// level 0
assign po6508 = pi6497;// level 0
assign po6509 = pi6500;// level 0
assign po6510 = pi6490;// level 0
assign po6511 = pi6519;// level 0
assign po6512 = pi6512;// level 0
assign po6513 = pi6507;// level 0
assign po6514 = pi6524;// level 0
assign po6515 = pi6487;// level 0
assign po6516 = pi6518;// level 0
assign po6517 = pi6520;// level 0
assign po6518 = pi6488;// level 0
assign po6519 = pi6509;// level 0
assign po6520 = pi6486;// level 0
assign po6521 = pi6515;// level 0
assign po6522 = pi6489;// level 0
assign po6523 = pi6527;// level 0
assign po6524 = pi6533;// level 0
assign po6525 = pi6529;// level 0
assign po6526 = pi6493;// level 0
assign po6527 = pi6531;// level 0
assign po6528 = pi6535;// level 0
assign po6529 = pi6508;// level 0
assign po6530 = pi6543;// level 0
assign po6531 = pi6494;// level 0
assign po6532 = pi6541;// level 0
assign po6533 = pi6514;// level 0
assign po6534 = pi6532;// level 0
assign po6535 = pi6504;// level 0
assign po6536 = pi6510;// level 0
assign po6537 = pi6496;// level 0
assign po6538 = pi6522;// level 0
assign po6539 = pi6513;// level 0
assign po6540 = pi6502;// level 0
assign po6541 = pi6540;// level 0
assign po6542 = pi6511;// level 0
assign po6543 = pi6534;// level 0
assign po6544 = pi6523;// level 0
assign po6545 = pi6528;// level 0
assign po6546 = pi6415;// level 0
assign po6547 = pi6452;// level 0
assign po6548 = pi6438;// level 0
assign po6549 = pi6546;// level 0
assign po6550 = pi6551;// level 0
assign po6551 = pi6445;// level 0
assign po6552 = pi6492;// level 0
assign po6553 = pi6475;// level 0
assign po6554 = pi6476;// level 0
assign po6555 = pi6430;// level 0
assign po6556 = pi6447;// level 0
assign po6557 = pi6434;// level 0
assign po6558 = pi6448;// level 0
assign po6559 = pi6477;// level 0
assign po6560 = pi6429;// level 0
assign po6561 = pi6424;// level 0
assign po6562 = pi6453;// level 0
assign po6563 = pi6455;// level 0
assign po6564 = pi6446;// level 0
assign po6565 = pi6482;// level 0
assign po6566 = pi6444;// level 0
assign po6567 = pi6454;// level 0
assign po6568 = pi6436;// level 0
assign po6569 = pi6457;// level 0
assign po6570 = pi6478;// level 0
assign po6571 = pi6442;// level 0
assign po6572 = pi6410;// level 0
assign po6573 = pi6450;// level 0
assign po6574 = pi6417;// level 0
assign po6575 = pi6420;// level 0
assign po6576 = pi6462;// level 0
assign po6577 = pi6458;// level 0
assign po6578 = pi6471;// level 0
assign po6579 = pi6433;// level 0
assign po6580 = pi6432;// level 0
assign po6581 = pi6473;// level 0
assign po6582 = pi6437;// level 0
assign po6583 = pi6428;// level 0
assign po6584 = pi6426;// level 0
assign po6585 = pi6479;// level 0
assign po6586 = pi6435;// level 0
assign po6587 = pi6441;// level 0
assign po6588 = pi6443;// level 0
assign po6589 = pi6413;// level 0
assign po6590 = pi6431;// level 0
assign po6591 = pi6412;// level 0
assign po6592 = pi6411;// level 0
assign po6593 = pi6406;// level 0
assign po6594 = pi6423;// level 0
assign po6595 = pi6459;// level 0
assign po6596 = pi6613;// level 0
assign po6597 = pi6606;// level 0
assign po6598 = pi6621;// level 0
assign po6599 = pi6609;// level 0
assign po6600 = pi6439;// level 0
assign po6601 = pi6414;// level 0
assign po6602 = pi6600;// level 0
assign po6603 = pi6506;// level 0
assign po6604 = pi6605;// level 0
assign po6605 = pi6607;// level 0
assign po6606 = pi6608;// level 0
assign po6607 = pi6603;// level 0
assign po6608 = pi6427;// level 0
assign po6609 = pi6577;// level 0
assign po6610 = pi6456;// level 0
assign po6611 = pi6598;// level 0
assign po6612 = pi6620;// level 0
assign po6613 = pi6555;// level 0
assign po6614 = pi6610;// level 0
assign po6615 = pi6599;// level 0
assign po6616 = pi6425;// level 0
assign po6617 = pi6619;// level 0
assign po6618 = pi6449;// level 0
assign po6619 = pi6418;// level 0
assign po6620 = pi6422;// level 0
assign po6621 = pi6451;// level 0
assign po6622 = pi6602;// level 0
assign po6623 = pi6604;// level 0
assign po6624 = pi6440;// level 0
assign po6625 = pi6544;// level 0
assign po6626 = pi6628;// level 0
assign po6627 = pi6626;// level 0
assign po6628 = pi6505;// level 0
assign po6629 = pi6627;// level 0
assign po6630 = pi6614;// level 0
assign po6631 = pi6623;// level 0
assign po6632 = pi6625;// level 0
assign po6633 = pi6629;// level 0
assign po6634 = pi6655;// level 0
assign po6635 = pi6634;// level 0
assign po6636 = pi6596;// level 0
assign po6637 = pi6637;// level 0
assign po6638 = pi6663;// level 0
assign po6639 = pi6661;// level 0
assign po6640 = pi6574;// level 0
assign po6641 = pi6553;// level 0
assign po6642 = pi6554;// level 0
assign po6643 = pi6581;// level 0
assign po6644 = pi6587;// level 0
assign po6645 = pi6569;// level 0
assign po6646 = pi6699;// level 0
assign po6647 = pi6617;// level 0
assign po6648 = pi6547;// level 0
assign po6649 = pi6676;// level 0
assign po6650 = pi6575;// level 0
assign po6651 = pi6664;// level 0
assign po6652 = pi6572;// level 0
assign po6653 = pi6582;// level 0
assign po6654 = pi6563;// level 0
assign po6655 = pi6585;// level 0
assign po6656 = pi6568;// level 0
assign po6657 = pi6584;// level 0
assign po6658 = pi6612;// level 0
assign po6659 = pi6616;// level 0
assign po6660 = pi6601;// level 0
assign po6661 = pi6590;// level 0
assign po6662 = pi6618;// level 0
assign po6663 = pi6565;// level 0
assign po6664 = pi6545;// level 0
assign po6665 = pi6611;// level 0
assign po6666 = pi6579;// level 0
assign po6667 = pi6567;// level 0
assign po6668 = pi6583;// level 0
assign po6669 = pi6566;// level 0
assign po6670 = pi6556;// level 0
assign po6671 = pi6578;// level 0
assign po6672 = pi6558;// level 0
assign po6673 = pi6562;// level 0
assign po6674 = pi6580;// level 0
assign po6675 = pi6549;// level 0
assign po6676 = pi6589;// level 0
assign po6677 = pi6595;// level 0
assign po6678 = pi6548;// level 0
assign po6679 = pi6571;// level 0
assign po6680 = pi6592;// level 0
assign po6681 = pi6560;// level 0
assign po6682 = pi6573;// level 0
assign po6683 = pi6576;// level 0
assign po6684 = pi6557;// level 0
assign po6685 = pi6597;// level 0
assign po6686 = pi6550;// level 0
assign po6687 = pi6586;// level 0
assign po6688 = pi6564;// level 0
assign po6689 = pi6671;// level 0
assign po6690 = pi6667;// level 0
assign po6691 = pi6673;// level 0
assign po6692 = pi6559;// level 0
assign po6693 = pi6658;// level 0
assign po6694 = pi6674;// level 0
assign po6695 = pi6660;// level 0
assign po6696 = pi6695;// level 0
assign po6697 = pi6693;// level 0
assign po6698 = pi6669;// level 0
assign po6699 = pi6680;// level 0
assign po6700 = pi6681;// level 0
assign po6701 = pi6552;// level 0
assign po6702 = pi6698;// level 0
assign po6703 = pi6615;// level 0
assign po6704 = pi6707;// level 0
assign po6705 = pi6591;// level 0
assign po6706 = pi6594;// level 0
assign po6707 = pi6593;// level 0
assign po6708 = pi6588;// level 0
assign po6709 = pi6570;// level 0
assign po6710 = pi6670;// level 0
assign po6711 = pi6662;// level 0
assign po6712 = pi6561;// level 0
assign po6713 = pi6632;// level 0
assign po6714 = pi6668;// level 0
assign po6715 = pi6684;// level 0
assign po6716 = pi6758;// level 0
assign po6717 = pi6749;// level 0
assign po6718 = pi6724;// level 0
assign po6719 = pi6755;// level 0
assign po6720 = pi6771;// level 0
assign po6721 = pi6672;// level 0
assign po6722 = pi6779;// level 0
assign po6723 = pi6742;// level 0
assign po6724 = pi6726;// level 0
assign po6725 = pi6763;// level 0
assign po6726 = pi6747;// level 0
assign po6727 = pi6725;// level 0
assign po6728 = pi6774;// level 0
assign po6729 = pi6766;// level 0
assign po6730 = pi6734;// level 0
assign po6731 = pi6727;// level 0
assign po6732 = pi6722;// level 0
assign po6733 = pi6736;// level 0
assign po6734 = pi6731;// level 0
assign po6735 = pi6769;// level 0
assign po6736 = pi6765;// level 0
assign po6737 = pi6730;// level 0
assign po6738 = pi6735;// level 0
assign po6739 = pi6772;// level 0
assign po6740 = pi6760;// level 0
assign po6741 = pi6741;// level 0
assign po6742 = pi6768;// level 0
assign po6743 = pi6750;// level 0
assign po6744 = pi6738;// level 0
assign po6745 = pi6761;// level 0
assign po6746 = pi6723;// level 0
assign po6747 = pi6751;// level 0
assign po6748 = pi6757;// level 0
assign po6749 = pi6743;// level 0
assign po6750 = pi6777;// level 0
assign po6751 = pi6759;// level 0
assign po6752 = pi6717;// level 0
assign po6753 = pi6720;// level 0
assign po6754 = pi6715;// level 0
assign po6755 = pi6764;// level 0
assign po6756 = pi6753;// level 0
assign po6757 = pi6773;// level 0
assign po6758 = pi6754;// level 0
assign po6759 = pi6728;// level 0
assign po6760 = pi6744;// level 0
assign po6761 = pi6718;// level 0
assign po6762 = pi6733;// level 0
assign po6763 = pi6729;// level 0
assign po6764 = pi6748;// level 0
assign po6765 = pi6622;// level 0
assign po6766 = pi6775;// level 0
assign po6767 = pi6745;// level 0
assign po6768 = pi6624;// level 0
assign po6769 = pi6752;// level 0
assign po6770 = pi6762;// level 0
assign po6771 = pi6737;// level 0
assign po6772 = pi6732;// level 0
assign po6773 = pi6767;// level 0
assign po6774 = pi6719;// level 0
assign po6775 = pi6712;// level 0
assign po6776 = pi6746;// level 0
assign po6777 = pi6665;// level 0
assign po6778 = pi6646;// level 0
assign po6779 = pi6701;// level 0
assign po6780 = pi6630;// level 0
assign po6781 = pi6799;// level 0
assign po6782 = pi6644;// level 0
assign po6783 = pi6645;// level 0
assign po6784 = pi6685;// level 0
assign po6785 = pi6828;// level 0
assign po6786 = pi6642;// level 0
assign po6787 = pi6683;// level 0
assign po6788 = pi6703;// level 0
assign po6789 = pi6638;// level 0
assign po6790 = pi6709;// level 0
assign po6791 = pi6631;// level 0
assign po6792 = pi6639;// level 0
assign po6793 = pi6678;// level 0
assign po6794 = pi6710;// level 0
assign po6795 = pi6682;// level 0
assign po6796 = pi6649;// level 0
assign po6797 = pi6675;// level 0
assign po6798 = pi6653;// level 0
assign po6799 = pi6689;// level 0
assign po6800 = pi6635;// level 0
assign po6801 = pi6659;// level 0
assign po6802 = pi6711;// level 0
assign po6803 = pi6657;// level 0
assign po6804 = pi6686;// level 0
assign po6805 = pi6690;// level 0
assign po6806 = pi6666;// level 0
assign po6807 = pi6739;// level 0
assign po6808 = pi6677;// level 0
assign po6809 = pi6643;// level 0
assign po6810 = pi6704;// level 0
assign po6811 = pi6688;// level 0
assign po6812 = pi6652;// level 0
assign po6813 = pi6708;// level 0
assign po6814 = pi6696;// level 0
assign po6815 = pi6636;// level 0
assign po6816 = pi6700;// level 0
assign po6817 = pi6647;// level 0
assign po6818 = pi6692;// level 0
assign po6819 = pi6650;// level 0
assign po6820 = pi6633;// level 0
assign po6821 = pi6640;// level 0
assign po6822 = pi6654;// level 0
assign po6823 = pi6641;// level 0
assign po6824 = pi6656;// level 0
assign po6825 = pi6651;// level 0
assign po6826 = pi6714;// level 0
assign po6827 = pi6648;// level 0
assign po6828 = pi6794;// level 0
assign po6829 = pi6839;// level 0
assign po6830 = pi6778;// level 0
assign po6831 = pi6694;// level 0
assign po6832 = pi6809;// level 0
assign po6833 = pi6721;// level 0
assign po6834 = pi6801;// level 0
assign po6835 = pi6782;// level 0
assign po6836 = pi6780;// level 0
assign po6837 = pi6827;// level 0
assign po6838 = pi6756;// level 0
assign po6839 = pi6821;// level 0
assign po6840 = pi6800;// level 0
assign po6841 = pi6691;// level 0
assign po6842 = pi6702;// level 0
assign po6843 = pi6806;// level 0
assign po6844 = pi6697;// level 0
assign po6845 = pi6679;// level 0
assign po6846 = pi6705;// level 0
assign po6847 = pi6713;// level 0
assign po6848 = pi6687;// level 0
assign po6849 = pi6706;// level 0
assign po6850 = pi6716;// level 0
assign po6851 = pi6849;// level 0
assign po6852 = pi6857;// level 0
assign po6853 = pi6859;// level 0
assign po6854 = pi6853;// level 0
assign po6855 = pi6855;// level 0
assign po6856 = pi6770;// level 0
assign po6857 = pi6740;// level 0
assign po6858 = pi6776;// level 0
assign po6859 = pi6858;// level 0
assign po6860 = pi6796;// level 0
assign po6861 = pi6824;// level 0
assign po6862 = pi6885;// level 0
assign po6863 = pi6825;// level 0
assign po6864 = pi6897;// level 0
assign po6865 = pi6836;// level 0
assign po6866 = pi6803;// level 0
assign po6867 = pi6811;// level 0
assign po6868 = pi6851;// level 0
assign po6869 = pi6843;// level 0
assign po6870 = pi6787;// level 0
assign po6871 = pi6841;// level 0
assign po6872 = pi6840;// level 0
assign po6873 = pi6845;// level 0
assign po6874 = pi6837;// level 0
assign po6875 = pi6805;// level 0
assign po6876 = pi6829;// level 0
assign po6877 = pi6790;// level 0
assign po6878 = pi6833;// level 0
assign po6879 = pi6784;// level 0
assign po6880 = pi6808;// level 0
assign po6881 = pi6817;// level 0
assign po6882 = pi6842;// level 0
assign po6883 = pi6831;// level 0
assign po6884 = pi6783;// level 0
assign po6885 = pi6864;// level 0
assign po6886 = pi6846;// level 0
assign po6887 = pi6810;// level 0
assign po6888 = pi6937;// level 0
assign po6889 = pi6834;// level 0
assign po6890 = pi6884;// level 0
assign po6891 = pi6861;// level 0
assign po6892 = pi6922;// level 0
assign po6893 = pi6870;// level 0
assign po6894 = pi6917;// level 0
assign po6895 = pi6785;// level 0
assign po6896 = pi6802;// level 0
assign po6897 = pi6905;// level 0
assign po6898 = pi6874;// level 0
assign po6899 = pi6895;// level 0
assign po6900 = pi6913;// level 0
assign po6901 = pi6860;// level 0
assign po6902 = pi6879;// level 0
assign po6903 = pi6911;// level 0
assign po6904 = pi6867;// level 0
assign po6905 = pi6820;// level 0
assign po6906 = pi6936;// level 0
assign po6907 = pi6812;// level 0
assign po6908 = pi6789;// level 0
assign po6909 = pi6832;// level 0
assign po6910 = pi6807;// level 0
assign po6911 = pi6844;// level 0
assign po6912 = pi6822;// level 0
assign po6913 = pi6835;// level 0
assign po6914 = pi6909;// level 0
assign po6915 = pi6848;// level 0
assign po6916 = pi6826;// level 0
assign po6917 = pi6823;// level 0
assign po6918 = pi6795;// level 0
assign po6919 = pi6793;// level 0
assign po6920 = pi6797;// level 0
assign po6921 = pi6818;// level 0
assign po6922 = pi6838;// level 0
assign po6923 = pi6941;// level 0
assign po6924 = pi6781;// level 0
assign po6925 = pi6854;// level 0
assign po6926 = pi6788;// level 0
assign po6927 = pi6878;// level 0
assign po6928 = pi6896;// level 0
assign po6929 = pi6889;// level 0
assign po6930 = pi6816;// level 0
assign po6931 = pi6791;// level 0
assign po6932 = pi6847;// level 0
assign po6933 = pi6792;// level 0
assign po6934 = pi6804;// level 0
assign po6935 = pi6815;// level 0
assign po6936 = pi6915;// level 0
assign po6937 = pi6866;// level 0
assign po6938 = pi6798;// level 0
assign po6939 = pi6830;// level 0
assign po6940 = pi6850;// level 0
assign po6941 = pi6786;// level 0
assign po6942 = pi6814;// level 0
assign po6943 = pi6813;// level 0
assign po6944 = pi6819;// level 0
assign po6945 = pi6947;// level 0
assign po6946 = pi6972;// level 0
assign po6947 = pi6962;// level 0
assign po6948 = pi6852;// level 0
assign po6949 = pi6993;// level 0
assign po6950 = pi6961;// level 0
assign po6951 = pi7010;// level 0
assign po6952 = pi6977;// level 0
assign po6953 = pi6945;// level 0
assign po6954 = pi6992;// level 0
assign po6955 = pi6975;// level 0
assign po6956 = pi6999;// level 0
assign po6957 = pi6963;// level 0
assign po6958 = pi6965;// level 0
assign po6959 = pi6856;// level 0
assign po6960 = pi7000;// level 0
assign po6961 = pi6998;// level 0
assign po6962 = pi6927;// level 0
assign po6963 = pi6980;// level 0
assign po6964 = pi6872;// level 0
assign po6965 = pi6971;// level 0
assign po6966 = pi6964;// level 0
assign po6967 = pi7013;// level 0
assign po6968 = ~pi6918;// level 0
assign po6969 = pi6989;// level 0
assign po6970 = pi7011;// level 0
assign po6971 = pi6957;// level 0
assign po6972 = pi6955;// level 0
assign po6973 = pi6969;// level 0
assign po6974 = pi6973;// level 0
assign po6975 = pi6987;// level 0
assign po6976 = pi6994;// level 0
assign po6977 = pi6950;// level 0
assign po6978 = pi6948;// level 0
assign po6979 = pi6968;// level 0
assign po6980 = pi6986;// level 0
assign po6981 = pi7012;// level 0
assign po6982 = pi6981;// level 0
assign po6983 = pi6956;// level 0
assign po6984 = pi6983;// level 0
assign po6985 = pi6952;// level 0
assign po6986 = pi6967;// level 0
assign po6987 = pi6979;// level 0
assign po6988 = pi6959;// level 0
assign po6989 = pi7003;// level 0
assign po6990 = pi7008;// level 0
assign po6991 = pi6988;// level 0
assign po6992 = pi7009;// level 0
assign po6993 = pi6991;// level 0
assign po6994 = pi7004;// level 0
assign po6995 = pi6997;// level 0
assign po6996 = pi6970;// level 0
assign po6997 = pi6958;// level 0
assign po6998 = pi6974;// level 0
assign po6999 = ~pi6868;// level 0
assign po7000 = pi6966;// level 0
assign po7001 = pi6985;// level 0
assign po7002 = pi6951;// level 0
assign po7003 = pi7005;// level 0
assign po7004 = pi6995;// level 0
assign po7005 = pi7002;// level 0
assign po7006 = pi6953;// level 0
assign po7007 = pi7006;// level 0
assign po7008 = pi6984;// level 0
assign po7009 = pi6946;// level 0
assign po7010 = pi7068;// level 0
assign po7011 = pi6890;// level 0
assign po7012 = pi6954;// level 0
assign po7013 = pi6914;// level 0
assign po7014 = pi6907;// level 0
assign po7015 = pi6934;// level 0
assign po7016 = pi6883;// level 0
assign po7017 = pi6899;// level 0
assign po7018 = pi6880;// level 0
assign po7019 = pi6865;// level 0
assign po7020 = pi6876;// level 0
assign po7021 = pi6904;// level 0
assign po7022 = pi6881;// level 0
assign po7023 = pi6877;// level 0
assign po7024 = pi7048;// level 0
assign po7025 = pi6921;// level 0
assign po7026 = pi6929;// level 0
assign po7027 = pi6933;// level 0
assign po7028 = pi6925;// level 0
assign po7029 = pi7001;// level 0
assign po7030 = pi7020;// level 0
assign po7031 = pi7063;// level 0
assign po7032 = pi6930;// level 0
assign po7033 = pi6894;// level 0
assign po7034 = pi6875;// level 0
assign po7035 = pi6892;// level 0
assign po7036 = pi7016;// level 0
assign po7037 = pi7073;// level 0
assign po7038 = pi6887;// level 0
assign po7039 = pi7022;// level 0
assign po7040 = pi6943;// level 0
assign po7041 = pi7028;// level 0
assign po7042 = pi6903;// level 0
assign po7043 = pi6900;// level 0
assign po7044 = pi6901;// level 0
assign po7045 = pi6908;// level 0
assign po7046 = pi6873;// level 0
assign po7047 = pi6863;// level 0
assign po7048 = pi6902;// level 0
assign po7049 = pi6926;// level 0
assign po7050 = pi6923;// level 0
assign po7051 = pi6982;// level 0
assign po7052 = pi6871;// level 0
assign po7053 = pi6893;// level 0
assign po7054 = pi6935;// level 0
assign po7055 = pi6916;// level 0
assign po7056 = pi6924;// level 0
assign po7057 = pi6960;// level 0
assign po7058 = pi7080;// level 0
assign po7059 = pi6862;// level 0
assign po7060 = pi6939;// level 0
assign po7061 = pi6919;// level 0
assign po7062 = pi6940;// level 0
assign po7063 = pi6932;// level 0
assign po7064 = pi6931;// level 0
assign po7065 = pi6891;// level 0
assign po7066 = pi6886;// level 0
assign po7067 = pi6928;// level 0
assign po7068 = pi6898;// level 0
assign po7069 = pi7018;// level 0
assign po7070 = pi6869;// level 0
assign po7071 = pi6944;// level 0
assign po7072 = pi6938;// level 0
assign po7073 = pi6912;// level 0
assign po7074 = pi7025;// level 0
assign po7075 = pi6942;// level 0
assign po7076 = pi6910;// level 0
assign po7077 = pi6906;// level 0
assign po7078 = pi6888;// level 0
assign po7079 = pi6990;// level 0
assign po7080 = pi6920;// level 0
assign po7081 = pi6882;// level 0
assign po7082 = pi7081;// level 0
assign po7083 = pi6976;// level 0
assign po7084 = pi7007;// level 0
assign po7085 = pi7083;// level 0
assign po7086 = pi7082;// level 0
assign po7087 = pi6949;// level 0
assign po7088 = pi6978;// level 0
assign po7089 = pi6996;// level 0
assign po7090 = pi7159;// level 0
assign po7091 = pi7169;// level 0
assign po7092 = pi7036;// level 0
assign po7093 = pi7069;// level 0
assign po7094 = pi7154;// level 0
assign po7095 = pi7053;// level 0
assign po7096 = pi7134;// level 0
assign po7097 = pi7151;// level 0
assign po7098 = pi7177;// level 0
assign po7099 = pi7064;// level 0
assign po7100 = pi7143;// level 0
assign po7101 = pi7062;// level 0
assign po7102 = pi7142;// level 0
assign po7103 = pi7021;// level 0
assign po7104 = pi7146;// level 0
assign po7105 = pi7035;// level 0
assign po7106 = pi7029;// level 0
assign po7107 = pi7051;// level 0
assign po7108 = pi7153;// level 0
assign po7109 = pi7117;// level 0
assign po7110 = pi7067;// level 0
assign po7111 = pi7078;// level 0
assign po7112 = pi7077;// level 0
assign po7113 = pi7060;// level 0
assign po7114 = pi7161;// level 0
assign po7115 = pi7166;// level 0
assign po7116 = pi7027;// level 0
assign po7117 = pi7026;// level 0
assign po7118 = pi7047;// level 0
assign po7119 = pi7101;// level 0
assign po7120 = pi7043;// level 0
assign po7121 = pi7033;// level 0
assign po7122 = pi7076;// level 0
assign po7123 = pi7071;// level 0
assign po7124 = pi7059;// level 0
assign po7125 = pi7158;// level 0
assign po7126 = pi7167;// level 0
assign po7127 = pi7162;// level 0
assign po7128 = pi7037;// level 0
assign po7129 = pi7057;// level 0
assign po7130 = pi7058;// level 0
assign po7131 = pi7045;// level 0
assign po7132 = pi7039;// level 0
assign po7133 = pi7044;// level 0
assign po7134 = pi7038;// level 0
assign po7135 = pi7140;// level 0
assign po7136 = pi7015;// level 0
assign po7137 = pi7041;// level 0
assign po7138 = pi7055;// level 0
assign po7139 = pi7144;// level 0
assign po7140 = pi7074;// level 0
assign po7141 = pi7145;// level 0
assign po7142 = pi7024;// level 0
assign po7143 = pi7165;// level 0
assign po7144 = pi7040;// level 0
assign po7145 = pi7148;// level 0
assign po7146 = pi7046;// level 0
assign po7147 = pi7160;// level 0
assign po7148 = pi7157;// level 0
assign po7149 = pi7052;// level 0
assign po7150 = pi7017;// level 0
assign po7151 = pi7023;// level 0
assign po7152 = pi7141;// level 0
assign po7153 = pi7049;// level 0
assign po7154 = pi7070;// level 0
assign po7155 = pi7056;// level 0
assign po7156 = pi7075;// level 0
assign po7157 = pi7135;// level 0
assign po7158 = pi7032;// level 0
assign po7159 = pi7019;// level 0
assign po7160 = pi7066;// level 0
assign po7161 = pi7050;// level 0
assign po7162 = pi7034;// level 0
assign po7163 = pi7014;// level 0
assign po7164 = pi7031;// level 0
assign po7165 = pi7079;// level 0
assign po7166 = pi7137;// level 0
assign po7167 = pi7147;// level 0
assign po7168 = pi7065;// level 0
assign po7169 = pi7054;// level 0
assign po7170 = pi7072;// level 0
assign po7171 = pi7084;// level 0
assign po7172 = pi7030;// level 0
assign po7173 = pi7042;// level 0
assign po7174 = pi7061;// level 0
assign po7175 = pi7191;// level 0
assign po7176 = pi7220;// level 0
assign po7177 = pi7183;// level 0
assign po7178 = pi7219;// level 0
assign po7179 = pi7181;// level 0
assign po7180 = pi7217;// level 0
assign po7181 = pi7199;// level 0
assign po7182 = pi7245;// level 0
assign po7183 = pi7195;// level 0
assign po7184 = pi7187;// level 0
assign po7185 = pi7182;// level 0
assign po7186 = pi7241;// level 0
assign po7187 = pi7188;// level 0
assign po7188 = pi7223;// level 0
assign po7189 = pi7197;// level 0
assign po7190 = pi7202;// level 0
assign po7191 = pi7192;// level 0
assign po7192 = pi7226;// level 0
assign po7193 = pi7118;// level 0
assign po7194 = pi7230;// level 0
assign po7195 = pi7205;// level 0
assign po7196 = pi7216;// level 0
assign po7197 = pi7208;// level 0
assign po7198 = pi7238;// level 0
assign po7199 = pi7221;// level 0
assign po7200 = pi7231;// level 0
assign po7201 = pi7218;// level 0
assign po7202 = pi7198;// level 0
assign po7203 = pi7184;// level 0
assign po7204 = pi7215;// level 0
assign po7205 = pi7225;// level 0
assign po7206 = pi7235;// level 0
assign po7207 = pi7228;// level 0
assign po7208 = pi7190;// level 0
assign po7209 = pi7196;// level 0
assign po7210 = pi7201;// level 0
assign po7211 = pi7180;// level 0
assign po7212 = pi7185;// level 0
assign po7213 = pi7200;// level 0
assign po7214 = pi7239;// level 0
assign po7215 = pi7207;// level 0
assign po7216 = pi7242;// level 0
assign po7217 = pi7098;// level 0
assign po7218 = pi7186;// level 0
assign po7219 = pi7164;// level 0
assign po7220 = pi7212;// level 0
assign po7221 = pi7138;// level 0
assign po7222 = pi7189;// level 0
assign po7223 = pi7206;// level 0
assign po7224 = pi7243;// level 0
assign po7225 = pi7155;// level 0
assign po7226 = pi7203;// level 0
assign po7227 = pi7229;// level 0
assign po7228 = pi7234;// level 0
assign po7229 = pi7150;// level 0
assign po7230 = pi7233;// level 0
assign po7231 = pi7236;// level 0
assign po7232 = pi7209;// level 0
assign po7233 = pi7213;// level 0
assign po7234 = pi7204;// level 0
assign po7235 = pi7244;// level 0
assign po7236 = pi7214;// level 0
assign po7237 = pi7237;// level 0
assign po7238 = pi7193;// level 0
assign po7239 = pi7240;// level 0
assign po7240 = pi7224;// level 0
assign po7241 = pi7136;// level 0
assign po7242 = pi7227;// level 0
assign po7243 = pi7156;// level 0
assign po7244 = pi7114;// level 0
assign po7245 = pi7102;// level 0
assign po7246 = pi7285;// level 0
assign po7247 = pi7172;// level 0
assign po7248 = pi7248;// level 0
assign po7249 = pi7116;// level 0
assign po7250 = pi7294;// level 0
assign po7251 = pi7092;// level 0
assign po7252 = pi7292;// level 0
assign po7253 = pi7091;// level 0
assign po7254 = pi7100;// level 0
assign po7255 = pi7272;// level 0
assign po7256 = pi7123;// level 0
assign po7257 = pi7128;// level 0
assign po7258 = pi7232;// level 0
assign po7259 = pi7108;// level 0
assign po7260 = pi7111;// level 0
assign po7261 = pi7095;// level 0
assign po7262 = pi7124;// level 0
assign po7263 = pi7103;// level 0
assign po7264 = pi7132;// level 0
assign po7265 = pi7130;// level 0
assign po7266 = pi7133;// level 0
assign po7267 = pi7119;// level 0
assign po7268 = pi7149;// level 0
assign po7269 = pi7121;// level 0
assign po7270 = pi7086;// level 0
assign po7271 = pi7131;// level 0
assign po7272 = pi7173;// level 0
assign po7273 = pi7104;// level 0
assign po7274 = pi7112;// level 0
assign po7275 = pi7109;// level 0
assign po7276 = pi7129;// level 0
assign po7277 = pi7097;// level 0
assign po7278 = pi7250;// level 0
assign po7279 = pi7093;// level 0
assign po7280 = pi7125;// level 0
assign po7281 = pi7105;// level 0
assign po7282 = pi7115;// level 0
assign po7283 = pi7176;// level 0
assign po7284 = pi7122;// level 0
assign po7285 = pi7152;// level 0
assign po7286 = pi7087;// level 0
assign po7287 = pi7106;// level 0
assign po7288 = pi7168;// level 0
assign po7289 = pi7178;// level 0
assign po7290 = pi7096;// level 0
assign po7291 = pi7171;// level 0
assign po7292 = pi7120;// level 0
assign po7293 = pi7246;// level 0
assign po7294 = pi7175;// level 0
assign po7295 = pi7099;// level 0
assign po7296 = pi7126;// level 0
assign po7297 = pi7110;// level 0
assign po7298 = pi7210;// level 0
assign po7299 = pi7127;// level 0
assign po7300 = pi7113;// level 0
assign po7301 = pi7089;// level 0
assign po7302 = pi7090;// level 0
assign po7303 = pi7085;// level 0
assign po7304 = pi7094;// level 0
assign po7305 = pi7139;// level 0
assign po7306 = pi7170;// level 0
assign po7307 = pi7088;// level 0
assign po7308 = pi7107;// level 0
assign po7309 = pi7174;// level 0
assign po7310 = pi7163;// level 0
assign po7311 = pi7194;// level 0
assign po7312 = pi7211;// level 0
assign po7313 = pi7222;// level 0
assign po7314 = pi7179;// level 0
assign po7315 = pi7446;// level 0
assign po7316 = pi7302;// level 0
assign po7317 = pi7282;// level 0
assign po7318 = pi7257;// level 0
assign po7319 = pi7270;// level 0
assign po7320 = pi7264;// level 0
assign po7321 = pi7283;// level 0
assign po7322 = pi7273;// level 0
assign po7323 = pi7253;// level 0
assign po7324 = pi7309;// level 0
assign po7325 = pi7254;// level 0
assign po7326 = pi7296;// level 0
assign po7327 = pi7306;// level 0
assign po7328 = pi7423;// level 0
assign po7329 = pi7262;// level 0
assign po7330 = pi7256;// level 0
assign po7331 = pi7369;// level 0
assign po7332 = pi7276;// level 0
assign po7333 = pi7281;// level 0
assign po7334 = pi7298;// level 0
assign po7335 = pi7265;// level 0
assign po7336 = pi7288;// level 0
assign po7337 = pi7252;// level 0
assign po7338 = pi7304;// level 0
assign po7339 = pi7301;// level 0
assign po7340 = pi7263;// level 0
assign po7341 = pi7277;// level 0
assign po7342 = pi7279;// level 0
assign po7343 = pi7287;// level 0
assign po7344 = pi7286;// level 0
assign po7345 = pi7259;// level 0
assign po7346 = pi7261;// level 0
assign po7347 = pi7461;// level 0
assign po7348 = pi7422;// level 0
assign po7349 = pi7268;// level 0
assign po7350 = pi7271;// level 0
assign po7351 = pi7305;// level 0
assign po7352 = pi7249;// level 0
assign po7353 = pi7295;// level 0
assign po7354 = pi7308;// level 0
assign po7355 = pi7300;// level 0
assign po7356 = pi7266;// level 0
assign po7357 = pi7255;// level 0
assign po7358 = pi7307;// level 0
assign po7359 = pi7303;// level 0
assign po7360 = pi7290;// level 0
assign po7361 = pi7274;// level 0
assign po7362 = pi7297;// level 0
assign po7363 = pi7251;// level 0
assign po7364 = pi7293;// level 0
assign po7365 = pi7462;// level 0
assign po7366 = pi7409;// level 0
assign po7367 = pi7444;// level 0
assign po7368 = pi7436;// level 0
assign po7369 = pi7278;// level 0
assign po7370 = pi7366;// level 0
assign po7371 = pi7429;// level 0
assign po7372 = pi7383;// level 0
assign po7373 = pi7411;// level 0
assign po7374 = pi7433;// level 0
assign po7375 = pi7414;// level 0
assign po7376 = pi7424;// level 0
assign po7377 = pi7415;// level 0
assign po7378 = pi7386;// level 0
assign po7379 = pi7299;// level 0
assign po7380 = pi7454;// level 0
assign po7381 = pi7428;// level 0
assign po7382 = pi7280;// level 0
assign po7383 = pi7453;// level 0
assign po7384 = pi7413;// level 0
assign po7385 = pi7421;// level 0
assign po7386 = pi7376;// level 0
assign po7387 = pi7456;// level 0
assign po7388 = pi7385;// level 0
assign po7389 = pi7410;// level 0
assign po7390 = pi7460;// level 0
assign po7391 = pi7450;// level 0
assign po7392 = pi7434;// level 0
assign po7393 = pi7425;// level 0
assign po7394 = pi7417;// level 0
assign po7395 = pi7412;// level 0
assign po7396 = pi7440;// level 0
assign po7397 = pi7426;// level 0
assign po7398 = pi7275;// level 0
assign po7399 = pi7379;// level 0
assign po7400 = pi7284;// level 0
assign po7401 = pi7269;// level 0
assign po7402 = pi7291;// level 0
assign po7403 = pi7258;// level 0
assign po7404 = pi7267;// level 0
assign po7405 = pi7247;// level 0
assign po7406 = pi7289;// level 0
assign po7407 = pi7431;// level 0
assign po7408 = pi7260;// level 0
assign po7409 = pi7335;// level 0
assign po7410 = pi7314;// level 0
assign po7411 = pi7315;// level 0
assign po7412 = pi7359;// level 0
assign po7413 = pi7320;// level 0
assign po7414 = pi7348;// level 0
assign po7415 = pi7322;// level 0
assign po7416 = pi7352;// level 0
assign po7417 = pi7344;// level 0
assign po7418 = pi7331;// level 0
assign po7419 = pi7360;// level 0
assign po7420 = pi7321;// level 0
assign po7421 = pi7333;// level 0
assign po7422 = pi7327;// level 0
assign po7423 = pi7310;// level 0
assign po7424 = pi7356;// level 0
assign po7425 = pi7345;// level 0
assign po7426 = pi7353;// level 0
assign po7427 = pi7343;// level 0
assign po7428 = pi7355;// level 0
assign po7429 = pi7324;// level 0
assign po7430 = pi7357;// level 0
assign po7431 = pi7358;// level 0
assign po7432 = pi7346;// level 0
assign po7433 = pi7329;// level 0
assign po7434 = pi7364;// level 0
assign po7435 = pi7330;// level 0
assign po7436 = pi7350;// level 0
assign po7437 = pi7319;// level 0
assign po7438 = pi7365;// level 0
assign po7439 = pi7341;// level 0
assign po7440 = pi7334;// level 0
assign po7441 = pi7323;// level 0
assign po7442 = pi7311;// level 0
assign po7443 = pi7318;// level 0
assign po7444 = pi7325;// level 0
assign po7445 = pi7354;// level 0
assign po7446 = pi7338;// level 0
assign po7447 = pi7332;// level 0
assign po7448 = pi7466;// level 0
assign po7449 = pi7351;// level 0
assign po7450 = pi7361;// level 0
assign po7451 = pi7339;// level 0
assign po7452 = pi7313;// level 0
assign po7453 = pi7347;// level 0
assign po7454 = pi7401;// level 0
assign po7455 = pi7312;// level 0
assign po7456 = pi7340;// level 0
assign po7457 = pi7349;// level 0
assign po7458 = pi7439;// level 0
assign po7459 = pi7511;// level 0
assign po7460 = pi7519;// level 0
assign po7461 = pi7522;// level 0
assign po7462 = pi7518;// level 0
assign po7463 = pi7397;// level 0
assign po7464 = pi7430;// level 0
assign po7465 = pi7396;// level 0
assign po7466 = pi7521;// level 0
assign po7467 = pi7362;// level 0
assign po7468 = pi7328;// level 0
assign po7469 = pi7317;// level 0
assign po7470 = pi7336;// level 0
assign po7471 = pi7337;// level 0
assign po7472 = pi7363;// level 0
assign po7473 = pi7342;// level 0
assign po7474 = pi7316;// level 0
assign po7475 = pi7326;// level 0
assign po7476 = pi7449;// level 0
assign po7477 = pi7464;// level 0
assign po7478 = pi7534;// level 0
assign po7479 = pi7458;// level 0
assign po7480 = pi7568;// level 0
assign po7481 = pi7371;// level 0
assign po7482 = pi7420;// level 0
assign po7483 = pi7442;// level 0
assign po7484 = pi7387;// level 0
assign po7485 = pi7378;// level 0
assign po7486 = pi7402;// level 0
assign po7487 = pi7381;// level 0
assign po7488 = pi7432;// level 0
assign po7489 = pi7373;// level 0
assign po7490 = pi7405;// level 0
assign po7491 = pi7380;// level 0
assign po7492 = pi7451;// level 0
assign po7493 = pi7445;// level 0
assign po7494 = pi7400;// level 0
assign po7495 = pi7367;// level 0
assign po7496 = pi7465;// level 0
assign po7497 = pi7416;// level 0
assign po7498 = pi7399;// level 0
assign po7499 = pi7394;// level 0
assign po7500 = pi7403;// level 0
assign po7501 = pi7408;// level 0
assign po7502 = pi7591;// level 0
assign po7503 = pi7435;// level 0
assign po7504 = pi7459;// level 0
assign po7505 = pi7447;// level 0
assign po7506 = pi7384;// level 0
assign po7507 = pi7407;// level 0
assign po7508 = pi7418;// level 0
assign po7509 = pi7463;// level 0
assign po7510 = pi7452;// level 0
assign po7511 = pi7437;// level 0
assign po7512 = pi7375;// level 0
assign po7513 = pi7393;// level 0
assign po7514 = pi7374;// level 0
assign po7515 = pi7427;// level 0
assign po7516 = pi7448;// level 0
assign po7517 = pi7398;// level 0
assign po7518 = pi7392;// level 0
assign po7519 = pi7370;// level 0
assign po7520 = pi7406;// level 0
assign po7521 = pi7441;// level 0
assign po7522 = pi7528;// level 0
assign po7523 = pi7537;// level 0
assign po7524 = pi7589;// level 0
assign po7525 = pi7438;// level 0
assign po7526 = pi7368;// level 0
assign po7527 = pi7391;// level 0
assign po7528 = pi7455;// level 0
assign po7529 = pi7377;// level 0
assign po7530 = pi7389;// level 0
assign po7531 = pi7457;// level 0
assign po7532 = pi7372;// level 0
assign po7533 = pi7404;// level 0
assign po7534 = pi7419;// level 0
assign po7535 = pi7443;// level 0
assign po7536 = pi7390;// level 0
assign po7537 = pi7395;// level 0
assign po7538 = pi7382;// level 0
assign po7539 = pi7388;// level 0
assign po7540 = pi7483;// level 0
assign po7541 = pi7474;// level 0
assign po7542 = pi7494;// level 0
assign po7543 = pi7503;// level 0
assign po7544 = pi7477;// level 0
assign po7545 = pi7491;// level 0
assign po7546 = pi7497;// level 0
assign po7547 = pi7488;// level 0
assign po7548 = pi7485;// level 0
assign po7549 = pi7484;// level 0
assign po7550 = pi7499;// level 0
assign po7551 = pi7512;// level 0
assign po7552 = pi7473;// level 0
assign po7553 = pi7505;// level 0
assign po7554 = pi7510;// level 0
assign po7555 = pi7527;// level 0
assign po7556 = pi7487;// level 0
assign po7557 = pi7472;// level 0
assign po7558 = pi7516;// level 0
assign po7559 = pi7482;// level 0
assign po7560 = pi7506;// level 0
assign po7561 = pi7523;// level 0
assign po7562 = pi7524;// level 0
assign po7563 = pi7480;// level 0
assign po7564 = pi7514;// level 0
assign po7565 = pi7504;// level 0
assign po7566 = pi7515;// level 0
assign po7567 = pi7517;// level 0
assign po7568 = pi7508;// level 0
assign po7569 = pi7509;// level 0
assign po7570 = pi7513;// level 0
assign po7571 = pi7493;// level 0
assign po7572 = pi7489;// level 0
assign po7573 = pi7475;// level 0
assign po7574 = pi7476;// level 0
assign po7575 = pi7486;// level 0
assign po7576 = pi7525;// level 0
assign po7577 = pi7496;// level 0
assign po7578 = pi7469;// level 0
assign po7579 = pi7490;// level 0
assign po7580 = pi7471;// level 0
assign po7581 = pi7502;// level 0
assign po7582 = pi7526;// level 0
assign po7583 = pi7467;// level 0
assign po7584 = pi7479;// level 0
assign po7585 = pi7495;// level 0
assign po7586 = pi7520;// level 0
assign po7587 = pi7498;// level 0
assign po7588 = pi7492;// level 0
assign po7589 = pi7468;// level 0
assign po7590 = pi7478;// level 0
assign po7591 = pi7501;// level 0
assign po7592 = pi7507;// level 0
assign po7593 = pi7470;// level 0
assign po7594 = pi7500;// level 0
assign po7595 = pi7481;// level 0
assign po7596 = pi7703;// level 0
assign po7597 = pi7555;// level 0
assign po7598 = pi7587;// level 0
assign po7599 = pi7726;// level 0
assign po7600 = pi7570;// level 0
assign po7601 = pi7564;// level 0
assign po7602 = pi7531;// level 0
assign po7603 = pi7574;// level 0
assign po7604 = pi7580;// level 0
assign po7605 = pi7538;// level 0
assign po7606 = pi7744;// level 0
assign po7607 = pi7560;// level 0
assign po7608 = pi7562;// level 0
assign po7609 = pi7674;// level 0
assign po7610 = pi7541;// level 0
assign po7611 = pi7585;// level 0
assign po7612 = pi7563;// level 0
assign po7613 = pi7711;// level 0
assign po7614 = pi7586;// level 0
assign po7615 = pi7660;// level 0
assign po7616 = pi7745;// level 0
assign po7617 = pi7567;// level 0
assign po7618 = pi7552;// level 0
assign po7619 = pi7532;// level 0
assign po7620 = pi7583;// level 0
assign po7621 = pi7565;// level 0
assign po7622 = pi7536;// level 0
assign po7623 = pi7543;// level 0
assign po7624 = pi7561;// level 0
assign po7625 = pi7571;// level 0
assign po7626 = pi7649;// level 0
assign po7627 = pi7684;// level 0
assign po7628 = pi7550;// level 0
assign po7629 = pi7549;// level 0
assign po7630 = pi7533;// level 0
assign po7631 = pi7661;// level 0
assign po7632 = pi7529;// level 0
assign po7633 = pi7539;// level 0
assign po7634 = pi7548;// level 0
assign po7635 = pi7578;// level 0
assign po7636 = pi7559;// level 0
assign po7637 = pi7545;// level 0
assign po7638 = pi7572;// level 0
assign po7639 = pi7736;// level 0
assign po7640 = pi7727;// level 0
assign po7641 = pi7648;// level 0
assign po7642 = pi7659;// level 0
assign po7643 = pi7693;// level 0
assign po7644 = pi7651;// level 0
assign po7645 = pi7668;// level 0
assign po7646 = pi7557;// level 0
assign po7647 = pi7663;// level 0
assign po7648 = pi7546;// level 0
assign po7649 = pi7576;// level 0
assign po7650 = pi7553;// level 0
assign po7651 = pi7683;// level 0
assign po7652 = pi7741;// level 0
assign po7653 = pi7590;// level 0
assign po7654 = pi7725;// level 0
assign po7655 = pi7670;// level 0
assign po7656 = pi7575;// level 0
assign po7657 = pi7653;// level 0
assign po7658 = pi7742;// level 0
assign po7659 = pi7658;// level 0
assign po7660 = pi7708;// level 0
assign po7661 = pi7739;// level 0
assign po7662 = pi7573;// level 0
assign po7663 = pi7664;// level 0
assign po7664 = pi7733;// level 0
assign po7665 = pi7558;// level 0
assign po7666 = pi7705;// level 0
assign po7667 = pi7584;// level 0
assign po7668 = pi7566;// level 0
assign po7669 = pi7689;// level 0
assign po7670 = pi7677;// level 0
assign po7671 = pi7588;// level 0
assign po7672 = pi7542;// level 0
assign po7673 = pi7530;// level 0
assign po7674 = pi7662;// level 0
assign po7675 = pi7581;// level 0
assign po7676 = pi7752;// level 0
assign po7677 = pi7544;// level 0
assign po7678 = pi7554;// level 0
assign po7679 = pi7749;// level 0
assign po7680 = pi7666;// level 0
assign po7681 = pi7577;// level 0
assign po7682 = pi7569;// level 0
assign po7683 = pi7679;// level 0
assign po7684 = pi7655;// level 0
assign po7685 = pi7582;// level 0
assign po7686 = pi7721;// level 0
assign po7687 = pi7551;// level 0
assign po7688 = pi7556;// level 0
assign po7689 = pi7547;// level 0
assign po7690 = pi7698;// level 0
assign po7691 = pi7720;// level 0
assign po7692 = pi7675;// level 0
assign po7693 = pi7540;// level 0
assign po7694 = pi7579;// level 0
assign po7695 = pi7535;// level 0
assign po7696 = pi7723;// level 0
assign po7697 = pi7634;// level 0
assign po7698 = pi7641;// level 0
assign po7699 = pi7621;// level 0
assign po7700 = pi7626;// level 0
assign po7701 = pi7645;// level 0
assign po7702 = pi7612;// level 0
assign po7703 = pi7624;// level 0
assign po7704 = pi7604;// level 0
assign po7705 = pi7628;// level 0
assign po7706 = pi7616;// level 0
assign po7707 = pi7630;// level 0
assign po7708 = pi7618;// level 0
assign po7709 = pi7633;// level 0
assign po7710 = pi7622;// level 0
assign po7711 = pi7640;// level 0
assign po7712 = pi7639;// level 0
assign po7713 = pi7593;// level 0
assign po7714 = pi7637;// level 0
assign po7715 = pi7625;// level 0
assign po7716 = pi7614;// level 0
assign po7717 = pi7608;// level 0
assign po7718 = pi7603;// level 0
assign po7719 = pi7598;// level 0
assign po7720 = pi7623;// level 0
assign po7721 = pi7611;// level 0
assign po7722 = pi7596;// level 0
assign po7723 = pi7642;// level 0
assign po7724 = pi7617;// level 0
assign po7725 = pi7632;// level 0
assign po7726 = pi7595;// level 0
assign po7727 = pi7619;// level 0
assign po7728 = pi7631;// level 0
assign po7729 = pi7635;// level 0
assign po7730 = pi7610;// level 0
assign po7731 = pi7600;// level 0
assign po7732 = pi7605;// level 0
assign po7733 = pi7644;// level 0
assign po7734 = pi7606;// level 0
assign po7735 = pi7599;// level 0
assign po7736 = pi7602;// level 0
assign po7737 = pi7646;// level 0
assign po7738 = pi7620;// level 0
assign po7739 = pi7592;// level 0
assign po7740 = pi7597;// level 0
assign po7741 = pi7686;// level 0
assign po7742 = pi7615;// level 0
assign po7743 = pi7607;// level 0
assign po7744 = pi7601;// level 0
assign po7745 = pi7594;// level 0
assign po7746 = pi7627;// level 0
assign po7747 = pi7647;// level 0
assign po7748 = pi7795;// level 0
assign po7749 = pi7811;// level 0
assign po7750 = pi7643;// level 0
assign po7751 = pi7803;// level 0
assign po7752 = pi7700;// level 0
assign po7753 = pi7609;// level 0
assign po7754 = pi7629;// level 0
assign po7755 = pi7636;// level 0
assign po7756 = pi7613;// level 0
assign po7757 = pi7638;// level 0
assign po7758 = pi7746;// level 0
assign po7759 = pi7738;// level 0
assign po7760 = pi7713;// level 0
assign po7761 = pi7716;// level 0
assign po7762 = pi7718;// level 0
assign po7763 = pi7737;// level 0
assign po7764 = pi7750;// level 0
assign po7765 = pi7728;// level 0
assign po7766 = pi7687;// level 0
assign po7767 = pi7652;// level 0
assign po7768 = pi7696;// level 0
assign po7769 = pi7680;// level 0
assign po7770 = pi7730;// level 0
assign po7771 = pi7732;// level 0
assign po7772 = pi7747;// level 0
assign po7773 = pi7734;// level 0
assign po7774 = pi7702;// level 0
assign po7775 = pi7715;// level 0
assign po7776 = pi7722;// level 0
assign po7777 = pi7740;// level 0
assign po7778 = pi7719;// level 0
assign po7779 = pi7731;// level 0
assign po7780 = pi7673;// level 0
assign po7781 = pi7690;// level 0
assign po7782 = pi7717;// level 0
assign po7783 = pi7714;// level 0
assign po7784 = pi7712;// level 0
assign po7785 = pi7697;// level 0
assign po7786 = pi7706;// level 0
assign po7787 = pi7704;// level 0
assign po7788 = pi7656;// level 0
assign po7789 = pi7709;// level 0
assign po7790 = pi7751;// level 0
assign po7791 = pi7665;// level 0
assign po7792 = pi7724;// level 0
assign po7793 = pi7688;// level 0
assign po7794 = pi7748;// level 0
assign po7795 = pi7654;// level 0
assign po7796 = pi7710;// level 0
assign po7797 = pi7676;// level 0
assign po7798 = pi7821;// level 0
assign po7799 = pi7692;// level 0
assign po7800 = pi7671;// level 0
assign po7801 = pi7743;// level 0
assign po7802 = pi7699;// level 0
assign po7803 = pi7694;// level 0
assign po7804 = pi7707;// level 0
assign po7805 = pi7817;// level 0
assign po7806 = pi7735;// level 0
assign po7807 = pi7685;// level 0
assign po7808 = pi7667;// level 0
assign po7809 = pi7657;// level 0
assign po7810 = pi7695;// level 0
assign po7811 = pi7701;// level 0
assign po7812 = pi7678;// level 0
assign po7813 = pi7682;// level 0
assign po7814 = pi7691;// level 0
assign po7815 = pi7672;// level 0
assign po7816 = pi7669;// level 0
assign po7817 = pi7729;// level 0
assign po7818 = pi7681;// level 0
assign po7819 = pi7813;// level 0
assign po7820 = pi7846;// level 0
assign po7821 = pi7650;// level 0
assign po7822 = pi7754;// level 0
assign po7823 = pi7809;// level 0
assign po7824 = pi7789;// level 0
assign po7825 = pi7775;// level 0
assign po7826 = pi7800;// level 0
assign po7827 = pi7797;// level 0
assign po7828 = pi7801;// level 0
assign po7829 = pi7804;// level 0
assign po7830 = pi7762;// level 0
assign po7831 = pi7776;// level 0
assign po7832 = pi7759;// level 0
assign po7833 = pi7771;// level 0
assign po7834 = pi7757;// level 0
assign po7835 = pi7792;// level 0
assign po7836 = pi7779;// level 0
assign po7837 = pi7778;// level 0
assign po7838 = pi7772;// level 0
assign po7839 = pi7769;// level 0
assign po7840 = pi7791;// level 0
assign po7841 = pi7785;// level 0
assign po7842 = pi7798;// level 0
assign po7843 = pi7794;// level 0
assign po7844 = pi7773;// level 0
assign po7845 = pi7787;// level 0
assign po7846 = pi7783;// level 0
assign po7847 = pi7755;// level 0
assign po7848 = pi7766;// level 0
assign po7849 = pi7781;// level 0
assign po7850 = pi7796;// level 0
assign po7851 = pi7782;// level 0
assign po7852 = pi7780;// level 0
assign po7853 = pi7802;// level 0
assign po7854 = pi7799;// level 0
assign po7855 = pi7761;// level 0
assign po7856 = pi7786;// level 0
assign po7857 = pi7764;// level 0
assign po7858 = pi7784;// level 0
assign po7859 = pi7777;// level 0
assign po7860 = pi7760;// level 0
assign po7861 = pi7810;// level 0
assign po7862 = pi7808;// level 0
assign po7863 = pi7758;// level 0
assign po7864 = pi7793;// level 0
assign po7865 = pi7770;// level 0
assign po7866 = pi7805;// level 0
assign po7867 = pi7774;// level 0
assign po7868 = pi7768;// level 0
assign po7869 = pi7788;// level 0
assign po7870 = pi7753;// level 0
assign po7871 = pi7756;// level 0
assign po7872 = pi7806;// level 0
assign po7873 = pi7807;// level 0
assign po7874 = pi7790;// level 0
assign po7875 = pi7767;// level 0
assign po7876 = pi7763;// level 0
assign po7877 = pi7765;// level 0
assign po7878 = pi7961;// level 0
assign po7879 = pi7998;// level 0
assign po7880 = pi8023;// level 0
assign po7881 = pi8005;// level 0
assign po7882 = pi7929;// level 0
assign po7883 = pi7940;// level 0
assign po7884 = pi7826;// level 0
assign po7885 = pi8001;// level 0
assign po7886 = pi7851;// level 0
assign po7887 = pi7868;// level 0
assign po7888 = pi8004;// level 0
assign po7889 = pi7991;// level 0
assign po7890 = pi8038;// level 0
assign po7891 = pi8020;// level 0
assign po7892 = pi7954;// level 0
assign po7893 = pi8017;// level 0
assign po7894 = pi8003;// level 0
assign po7895 = pi7869;// level 0
assign po7896 = pi8015;// level 0
assign po7897 = pi7838;// level 0
assign po7898 = pi7975;// level 0
assign po7899 = pi7849;// level 0
assign po7900 = pi7942;// level 0
assign po7901 = pi7866;// level 0
assign po7902 = pi7862;// level 0
assign po7903 = pi7854;// level 0
assign po7904 = pi7939;// level 0
assign po7905 = pi7999;// level 0
assign po7906 = pi7819;// level 0
assign po7907 = pi8036;// level 0
assign po7908 = pi7844;// level 0
assign po7909 = pi8033;// level 0
assign po7910 = pi7816;// level 0
assign po7911 = pi7864;// level 0
assign po7912 = pi7833;// level 0
assign po7913 = pi7971;// level 0
assign po7914 = pi7972;// level 0
assign po7915 = pi7814;// level 0
assign po7916 = pi7935;// level 0
assign po7917 = pi7870;// level 0
assign po7918 = pi7839;// level 0
assign po7919 = pi8030;// level 0
assign po7920 = pi7832;// level 0
assign po7921 = pi7858;// level 0
assign po7922 = pi7824;// level 0
assign po7923 = pi7968;// level 0
assign po7924 = pi7853;// level 0
assign po7925 = pi7836;// level 0
assign po7926 = pi7850;// level 0
assign po7927 = pi7848;// level 0
assign po7928 = pi7959;// level 0
assign po7929 = pi7837;// level 0
assign po7930 = pi8022;// level 0
assign po7931 = pi7820;// level 0
assign po7932 = pi7861;// level 0
assign po7933 = pi8016;// level 0
assign po7934 = pi7831;// level 0
assign po7935 = pi8025;// level 0
assign po7936 = pi7818;// level 0
assign po7937 = pi7842;// level 0
assign po7938 = pi7931;// level 0
assign po7939 = pi7815;// level 0
assign po7940 = pi7845;// level 0
assign po7941 = pi8011;// level 0
assign po7942 = pi7860;// level 0
assign po7943 = pi7863;// level 0
assign po7944 = pi7843;// level 0
assign po7945 = pi7827;// level 0
assign po7946 = pi7828;// level 0
assign po7947 = pi7867;// level 0
assign po7948 = pi7822;// level 0
assign po7949 = pi7865;// level 0
assign po7950 = pi7997;// level 0
assign po7951 = pi8000;// level 0
assign po7952 = pi7829;// level 0
assign po7953 = pi8034;// level 0
assign po7954 = pi7857;// level 0
assign po7955 = pi7965;// level 0
assign po7956 = pi7979;// level 0
assign po7957 = pi7946;// level 0
assign po7958 = pi7840;// level 0
assign po7959 = pi7841;// level 0
assign po7960 = pi7825;// level 0
assign po7961 = pi7852;// level 0
assign po7962 = pi7830;// level 0
assign po7963 = pi7974;// level 0
assign po7964 = pi7847;// level 0
assign po7965 = pi7855;// level 0
assign po7966 = pi7966;// level 0
assign po7967 = pi7856;// level 0
assign po7968 = pi7823;// level 0
assign po7969 = pi7957;// level 0
assign po7970 = pi7871;// level 0
assign po7971 = pi8031;// level 0
assign po7972 = pi8010;// level 0
assign po7973 = pi7812;// level 0
assign po7974 = pi7943;// level 0
assign po7975 = pi7978;// level 0
assign po7976 = pi7949;// level 0
assign po7977 = pi7834;// level 0
assign po7978 = pi7859;// level 0
assign po7979 = pi8028;// level 0
assign po7980 = pi8013;// level 0
assign po7981 = pi7835;// level 0
assign po7982 = pi7986;// level 0
assign po7983 = pi7894;// level 0
assign po7984 = pi7876;// level 0
assign po7985 = pi7874;// level 0
assign po7986 = pi7892;// level 0
assign po7987 = pi7882;// level 0
assign po7988 = pi7917;// level 0
assign po7989 = pi7907;// level 0
assign po7990 = pi7890;// level 0
assign po7991 = pi7872;// level 0
assign po7992 = pi7923;// level 0
assign po7993 = pi7902;// level 0
assign po7994 = pi7877;// level 0
assign po7995 = pi7916;// level 0
assign po7996 = pi7880;// level 0
assign po7997 = pi7881;// level 0
assign po7998 = pi7915;// level 0
assign po7999 = pi7900;// level 0
assign po8000 = pi7886;// level 0
assign po8001 = pi7908;// level 0
assign po8002 = pi7914;// level 0
assign po8003 = pi7899;// level 0
assign po8004 = pi7896;// level 0
assign po8005 = pi7924;// level 0
assign po8006 = pi7926;// level 0
assign po8007 = pi7879;// level 0
assign po8008 = pi7878;// level 0
assign po8009 = pi7912;// level 0
assign po8010 = pi7895;// level 0
assign po8011 = pi7904;// level 0
assign po8012 = pi7910;// level 0
assign po8013 = pi7898;// level 0
assign po8014 = pi7922;// level 0
assign po8015 = pi7887;// level 0
assign po8016 = pi7875;// level 0
assign po8017 = pi7903;// level 0
assign po8018 = pi7897;// level 0
assign po8019 = pi7893;// level 0
assign po8020 = pi7911;// level 0
assign po8021 = pi7883;// level 0
assign po8022 = pi7918;// level 0
assign po8023 = pi7906;// level 0
assign po8024 = pi7909;// level 0
assign po8025 = pi8039;// level 0
assign po8026 = pi7884;// level 0
assign po8027 = pi7901;// level 0
assign po8028 = pi7919;// level 0
assign po8029 = pi7873;// level 0
assign po8030 = pi7891;// level 0
assign po8031 = pi7905;// level 0
assign po8032 = pi7913;// level 0
assign po8033 = pi7952;// level 0
assign po8034 = pi7885;// level 0
assign po8035 = pi7888;// level 0
assign po8036 = pi7925;// level 0
assign po8037 = pi7921;// level 0
assign po8038 = pi7889;// level 0
assign po8039 = pi7927;// level 0
assign po8040 = pi7920;// level 0
assign po8041 = pi7963;// level 0
assign po8042 = pi8008;// level 0
assign po8043 = pi7937;// level 0
assign po8044 = pi8006;// level 0
assign po8045 = pi7984;// level 0
assign po8046 = pi7985;// level 0
assign po8047 = pi7977;// level 0
assign po8048 = pi7948;// level 0
assign po8049 = pi7969;// level 0
assign po8050 = pi7989;// level 0
assign po8051 = pi7958;// level 0
assign po8052 = pi7953;// level 0
assign po8053 = pi7973;// level 0
assign po8054 = pi7928;// level 0
assign po8055 = pi7987;// level 0
assign po8056 = pi7990;// level 0
assign po8057 = pi7947;// level 0
assign po8058 = pi7994;// level 0
assign po8059 = pi7951;// level 0
assign po8060 = pi8024;// level 0
assign po8061 = pi7992;// level 0
assign po8062 = pi7988;// level 0
assign po8063 = pi7933;// level 0
assign po8064 = pi7936;// level 0
assign po8065 = pi8027;// level 0
assign po8066 = pi8002;// level 0
assign po8067 = pi7995;// level 0
assign po8068 = pi7982;// level 0
assign po8069 = pi8029;// level 0
assign po8070 = pi8032;// level 0
assign po8071 = pi8012;// level 0
assign po8072 = pi7964;// level 0
assign po8073 = pi7932;// level 0
assign po8074 = pi7976;// level 0
assign po8075 = pi7980;// level 0
assign po8076 = pi8007;// level 0
assign po8077 = pi7930;// level 0
assign po8078 = pi7950;// level 0
assign po8079 = pi7981;// level 0
assign po8080 = pi7955;// level 0
assign po8081 = pi7962;// level 0
assign po8082 = pi7967;// level 0
assign po8083 = pi7941;// level 0
assign po8084 = pi7934;// level 0
assign po8085 = pi7993;// level 0
assign po8086 = pi7938;// level 0
assign po8087 = pi8019;// level 0
assign po8088 = pi7956;// level 0
assign po8089 = pi7945;// level 0
assign po8090 = pi8021;// level 0
assign po8091 = pi7996;// level 0
assign po8092 = pi8018;// level 0
assign po8093 = pi7983;// level 0
assign po8094 = pi8035;// level 0
assign po8095 = pi8037;// level 0
assign po8096 = pi8014;// level 0
assign po8097 = pi7970;// level 0
assign po8098 = pi8026;// level 0
assign po8099 = pi8009;// level 0
assign po8100 = pi7944;// level 0
assign po8101 = pi7960;// level 0
assign po8102 = pi8059;// level 0
assign po8103 = pi8091;// level 0
assign po8104 = pi8043;// level 0
assign po8105 = pi8071;// level 0
assign po8106 = pi8040;// level 0
assign po8107 = pi8082;// level 0
assign po8108 = pi8046;// level 0
assign po8109 = pi8053;// level 0
assign po8110 = pi8086;// level 0
assign po8111 = pi8088;// level 0
assign po8112 = pi8056;// level 0
assign po8113 = pi8070;// level 0
assign po8114 = pi8061;// level 0
assign po8115 = pi8047;// level 0
assign po8116 = pi8084;// level 0
assign po8117 = pi8054;// level 0
assign po8118 = pi8078;// level 0
assign po8119 = pi8081;// level 0
assign po8120 = pi8057;// level 0
assign po8121 = pi8063;// level 0
assign po8122 = pi8087;// level 0
assign po8123 = pi8092;// level 0
assign po8124 = pi8072;// level 0
assign po8125 = pi8068;// level 0
assign po8126 = pi8049;// level 0
assign po8127 = pi8073;// level 0
assign po8128 = pi8064;// level 0
assign po8129 = pi8058;// level 0
assign po8130 = pi8069;// level 0
assign po8131 = pi8074;// level 0
assign po8132 = pi8066;// level 0
assign po8133 = pi8055;// level 0
assign po8134 = pi8051;// level 0
assign po8135 = pi8050;// level 0
assign po8136 = pi8065;// level 0
assign po8137 = pi8042;// level 0
assign po8138 = pi8060;// level 0
assign po8139 = pi8094;// level 0
assign po8140 = pi8083;// level 0
assign po8141 = pi8044;// level 0
assign po8142 = pi8045;// level 0
assign po8143 = pi8095;// level 0
assign po8144 = pi8090;// level 0
assign po8145 = pi8089;// level 0
assign po8146 = pi8085;// level 0
assign po8147 = pi8067;// level 0
assign po8148 = pi8079;// level 0
assign po8149 = pi8052;// level 0
assign po8150 = pi8076;// level 0
assign po8151 = pi8041;// level 0
assign po8152 = pi8077;// level 0
assign po8153 = pi8048;// level 0
assign po8154 = pi8080;// level 0
assign po8155 = pi8093;// level 0
assign po8156 = pi8062;// level 0
assign po8157 = pi8075;// level 0
assign po8158 = ~w62986;// level 2
assign po8159 = ~w62989;// level 2
assign po8160 = ~w62992;// level 2
assign po8161 = ~w62995;// level 2
assign po8162 = ~w62998;// level 2
assign po8163 = ~w63001;// level 2
assign po8164 = ~w63004;// level 2
assign po8165 = ~w63007;// level 2
assign po8166 = ~w63010;// level 2
assign po8167 = ~w63013;// level 2
assign po8168 = ~w63016;// level 2
assign po8169 = ~w63019;// level 2
assign po8170 = ~w63022;// level 2
assign po8171 = ~w63025;// level 2
assign po8172 = ~w63028;// level 2
assign po8173 = ~w63031;// level 2
assign po8174 = ~w63034;// level 2
assign po8175 = ~w63037;// level 2
assign po8176 = ~w63040;// level 2
assign po8177 = ~w63043;// level 2
assign po8178 = ~w63046;// level 2
assign po8179 = ~w63049;// level 2
assign po8180 = ~w63052;// level 2
assign po8181 = ~w63055;// level 2
assign po8182 = ~w63058;// level 2
assign po8183 = ~w63061;// level 2
assign po8184 = ~w63064;// level 2
assign po8185 = ~w63067;// level 2
assign po8186 = ~w63070;// level 2
assign po8187 = ~w63073;// level 2
assign po8188 = ~w63076;// level 2
assign po8189 = ~w63079;// level 2
assign po8190 = ~w63082;// level 2
assign po8191 = ~w63085;// level 2
assign po8192 = ~w63088;// level 2
assign po8193 = ~w63091;// level 2
assign po8194 = ~w63094;// level 2
assign po8195 = ~w63097;// level 2
assign po8196 = ~w63100;// level 2
assign po8197 = ~w63103;// level 2
assign po8198 = ~w63106;// level 2
assign po8199 = ~w63109;// level 2
assign po8200 = ~w63112;// level 2
assign po8201 = ~w63115;// level 2
assign po8202 = ~w63118;// level 2
assign po8203 = ~w63121;// level 2
assign po8204 = ~w63124;// level 2
assign po8205 = ~w63127;// level 2
assign po8206 = ~w63130;// level 2
assign po8207 = ~w63133;// level 2
assign po8208 = ~w63136;// level 2
assign po8209 = ~w63139;// level 2
assign po8210 = ~w63142;// level 2
assign po8211 = ~w63145;// level 2
assign po8212 = ~w63148;// level 2
assign po8213 = ~w63151;// level 2
assign po8214 = ~w63154;// level 2
assign po8215 = ~w63157;// level 2
assign po8216 = ~w63160;// level 2
assign po8217 = ~w63163;// level 2
assign po8218 = ~w63166;// level 2
assign po8219 = ~w63169;// level 2
assign po8220 = ~w63172;// level 2
assign po8221 = ~w63175;// level 2
assign po8222 = ~w63178;// level 2
assign po8223 = ~w63181;// level 2
assign po8224 = ~w63184;// level 2
assign po8225 = ~w63187;// level 2
assign po8226 = ~w63190;// level 2
assign po8227 = ~w63193;// level 2
assign po8228 = ~w63196;// level 2
assign po8229 = ~w63199;// level 2
assign po8230 = ~w63202;// level 2
assign po8231 = ~w63205;// level 2
assign po8232 = ~w63208;// level 2
assign po8233 = ~w63211;// level 2
assign po8234 = ~w63214;// level 2
assign po8235 = ~w63217;// level 2
assign po8236 = ~w63220;// level 2
assign po8237 = ~w63223;// level 2
assign po8238 = ~w63226;// level 2
assign po8239 = ~w63229;// level 2
assign po8240 = ~w63232;// level 2
assign po8241 = ~w63235;// level 2
assign po8242 = ~w63238;// level 2
assign po8243 = ~w63241;// level 2
assign po8244 = ~w63244;// level 2
assign po8245 = ~w63247;// level 2
assign po8246 = ~w63250;// level 2
assign po8247 = ~w63253;// level 2
assign po8248 = ~w63256;// level 2
assign po8249 = ~w63259;// level 2
assign po8250 = ~w63262;// level 2
assign po8251 = ~w63265;// level 2
assign po8252 = ~w63268;// level 2
assign po8253 = ~w63271;// level 2
assign po8254 = ~w63274;// level 2
assign po8255 = ~w63277;// level 2
assign po8256 = ~w63280;// level 2
assign po8257 = ~w63283;// level 2
assign po8258 = ~w63286;// level 2
assign po8259 = ~w63289;// level 2
assign po8260 = ~w63292;// level 2
assign po8261 = ~w63295;// level 2
assign po8262 = ~w63298;// level 2
assign po8263 = ~w63301;// level 2
assign po8264 = ~w63304;// level 2
assign po8265 = ~w63307;// level 2
assign po8266 = ~w63310;// level 2
assign po8267 = ~w63313;// level 2
assign po8268 = ~w63316;// level 2
assign po8269 = ~w63319;// level 2
assign po8270 = pi8125;// level 0
assign po8271 = pi8099;// level 0
assign po8272 = pi8131;// level 0
assign po8273 = pi8096;// level 0
assign po8274 = pi8134;// level 0
assign po8275 = pi8097;// level 0
assign po8276 = pi8123;// level 0
assign po8277 = pi8145;// level 0
assign po8278 = pi8142;// level 0
assign po8279 = pi8135;// level 0
assign po8280 = pi8098;// level 0
assign po8281 = pi8103;// level 0
assign po8282 = pi8129;// level 0
assign po8283 = pi8122;// level 0
assign po8284 = pi8109;// level 0
assign po8285 = pi8149;// level 0
assign po8286 = pi8128;// level 0
assign po8287 = pi8138;// level 0
assign po8288 = pi8108;// level 0
assign po8289 = pi8100;// level 0
assign po8290 = pi8111;// level 0
assign po8291 = pi8124;// level 0
assign po8292 = pi8139;// level 0
assign po8293 = pi8116;// level 0
assign po8294 = pi8140;// level 0
assign po8295 = pi8137;// level 0
assign po8296 = pi8148;// level 0
assign po8297 = pi8120;// level 0
assign po8298 = pi8107;// level 0
assign po8299 = pi8114;// level 0
assign po8300 = pi8126;// level 0
assign po8301 = pi8102;// level 0
assign po8302 = pi8130;// level 0
assign po8303 = pi8150;// level 0
assign po8304 = pi8115;// level 0
assign po8305 = pi8112;// level 0
assign po8306 = pi8133;// level 0
assign po8307 = pi8117;// level 0
assign po8308 = pi8104;// level 0
assign po8309 = pi8143;// level 0
assign po8310 = pi8144;// level 0
assign po8311 = pi8106;// level 0
assign po8312 = pi8147;// level 0
assign po8313 = pi8118;// level 0
assign po8314 = pi8113;// level 0
assign po8315 = pi8110;// level 0
assign po8316 = pi8119;// level 0
assign po8317 = pi8151;// level 0
assign po8318 = pi8121;// level 0
assign po8319 = pi8101;// level 0
assign po8320 = pi8132;// level 0
assign po8321 = pi8141;// level 0
assign po8322 = pi8105;// level 0
assign po8323 = pi8136;// level 0
assign po8324 = pi8146;// level 0
assign po8325 = pi8127;// level 0
assign po8326 = pi8184;// level 0
assign po8327 = pi8203;// level 0
assign po8328 = pi8163;// level 0
assign po8329 = pi8205;// level 0
assign po8330 = pi8158;// level 0
assign po8331 = pi8202;// level 0
assign po8332 = pi8178;// level 0
assign po8333 = pi8177;// level 0
assign po8334 = pi8193;// level 0
assign po8335 = pi8195;// level 0
assign po8336 = pi8155;// level 0
assign po8337 = pi8179;// level 0
assign po8338 = pi8198;// level 0
assign po8339 = pi8187;// level 0
assign po8340 = pi8191;// level 0
assign po8341 = pi8156;// level 0
assign po8342 = pi8173;// level 0
assign po8343 = pi8160;// level 0
assign po8344 = pi8189;// level 0
assign po8345 = pi8152;// level 0
assign po8346 = pi8186;// level 0
assign po8347 = pi8188;// level 0
assign po8348 = pi8197;// level 0
assign po8349 = pi8196;// level 0
assign po8350 = pi8181;// level 0
assign po8351 = pi8182;// level 0
assign po8352 = pi8185;// level 0
assign po8353 = pi8183;// level 0
assign po8354 = pi8207;// level 0
assign po8355 = pi8171;// level 0
assign po8356 = pi8157;// level 0
assign po8357 = pi8167;// level 0
assign po8358 = pi8199;// level 0
assign po8359 = pi8153;// level 0
assign po8360 = pi8175;// level 0
assign po8361 = pi8154;// level 0
assign po8362 = pi8170;// level 0
assign po8363 = pi8161;// level 0
assign po8364 = pi8194;// level 0
assign po8365 = pi8166;// level 0
assign po8366 = pi8201;// level 0
assign po8367 = pi8200;// level 0
assign po8368 = pi8190;// level 0
assign po8369 = pi8164;// level 0
assign po8370 = pi8169;// level 0
assign po8371 = pi8176;// level 0
assign po8372 = pi8159;// level 0
assign po8373 = pi8165;// level 0
assign po8374 = pi8174;// level 0
assign po8375 = pi8206;// level 0
assign po8376 = pi8162;// level 0
assign po8377 = pi8204;// level 0
assign po8378 = pi8172;// level 0
assign po8379 = pi8168;// level 0
assign po8380 = pi8180;// level 0
assign po8381 = pi8192;// level 0
assign po8382 = pi8226;// level 0
assign po8383 = pi8258;// level 0
assign po8384 = pi8262;// level 0
assign po8385 = pi8221;// level 0
assign po8386 = pi8242;// level 0
assign po8387 = pi8215;// level 0
assign po8388 = pi8249;// level 0
assign po8389 = pi8240;// level 0
assign po8390 = pi8260;// level 0
assign po8391 = pi8227;// level 0
assign po8392 = pi8235;// level 0
assign po8393 = pi8231;// level 0
assign po8394 = pi8212;// level 0
assign po8395 = pi8225;// level 0
assign po8396 = pi8234;// level 0
assign po8397 = pi8255;// level 0
assign po8398 = pi8253;// level 0
assign po8399 = pi8230;// level 0
assign po8400 = pi8229;// level 0
assign po8401 = pi8236;// level 0
assign po8402 = pi8219;// level 0
assign po8403 = pi8228;// level 0
assign po8404 = pi8250;// level 0
assign po8405 = pi8224;// level 0
assign po8406 = pi8256;// level 0
assign po8407 = pi8252;// level 0
assign po8408 = pi8263;// level 0
assign po8409 = pi8237;// level 0
assign po8410 = pi8246;// level 0
assign po8411 = pi8245;// level 0
assign po8412 = pi8243;// level 0
assign po8413 = pi8217;// level 0
assign po8414 = pi8241;// level 0
assign po8415 = pi8248;// level 0
assign po8416 = pi8213;// level 0
assign po8417 = pi8216;// level 0
assign po8418 = pi8218;// level 0
assign po8419 = pi8222;// level 0
assign po8420 = pi8209;// level 0
assign po8421 = pi8211;// level 0
assign po8422 = pi8223;// level 0
assign po8423 = pi8254;// level 0
assign po8424 = pi8247;// level 0
assign po8425 = pi8208;// level 0
assign po8426 = pi8214;// level 0
assign po8427 = pi8244;// level 0
assign po8428 = pi8220;// level 0
assign po8429 = pi8257;// level 0
assign po8430 = pi8232;// level 0
assign po8431 = pi8251;// level 0
assign po8432 = pi8259;// level 0
assign po8433 = pi8239;// level 0
assign po8434 = pi8210;// level 0
assign po8435 = pi8233;// level 0
assign po8436 = pi8261;// level 0
assign po8437 = pi8238;// level 0
assign po8438 = pi8273;// level 0
assign po8439 = pi8306;// level 0
assign po8440 = pi8315;// level 0
assign po8441 = pi8311;// level 0
assign po8442 = pi8299;// level 0
assign po8443 = pi8296;// level 0
assign po8444 = pi8301;// level 0
assign po8445 = pi8295;// level 0
assign po8446 = pi8274;// level 0
assign po8447 = pi8280;// level 0
assign po8448 = pi8271;// level 0
assign po8449 = pi8310;// level 0
assign po8450 = pi8272;// level 0
assign po8451 = pi8304;// level 0
assign po8452 = pi8302;// level 0
assign po8453 = pi8282;// level 0
assign po8454 = pi8270;// level 0
assign po8455 = pi8285;// level 0
assign po8456 = pi8314;// level 0
assign po8457 = pi8313;// level 0
assign po8458 = pi8279;// level 0
assign po8459 = pi8278;// level 0
assign po8460 = pi8281;// level 0
assign po8461 = pi8275;// level 0
assign po8462 = pi8266;// level 0
assign po8463 = pi8298;// level 0
assign po8464 = pi8297;// level 0
assign po8465 = pi8303;// level 0
assign po8466 = pi8265;// level 0
assign po8467 = pi8312;// level 0
assign po8468 = pi8289;// level 0
assign po8469 = pi8309;// level 0
assign po8470 = pi8288;// level 0
assign po8471 = pi8269;// level 0
assign po8472 = pi8300;// level 0
assign po8473 = pi8284;// level 0
assign po8474 = pi8268;// level 0
assign po8475 = pi8318;// level 0
assign po8476 = pi8277;// level 0
assign po8477 = pi8292;// level 0
assign po8478 = pi8316;// level 0
assign po8479 = pi8317;// level 0
assign po8480 = pi8290;// level 0
assign po8481 = pi8286;// level 0
assign po8482 = pi8319;// level 0
assign po8483 = pi8307;// level 0
assign po8484 = pi8294;// level 0
assign po8485 = pi8293;// level 0
assign po8486 = pi8276;// level 0
assign po8487 = pi8283;// level 0
assign po8488 = pi8291;// level 0
assign po8489 = pi8308;// level 0
assign po8490 = pi8287;// level 0
assign po8491 = pi8264;// level 0
assign po8492 = pi8267;// level 0
assign po8493 = pi8305;// level 0
assign po8494 = pi8365;// level 0
assign po8495 = pi8348;// level 0
assign po8496 = pi8354;// level 0
assign po8497 = pi8341;// level 0
assign po8498 = pi8327;// level 0
assign po8499 = pi8339;// level 0
assign po8500 = pi8340;// level 0
assign po8501 = pi8331;// level 0
assign po8502 = pi8328;// level 0
assign po8503 = pi8325;// level 0
assign po8504 = pi8369;// level 0
assign po8505 = pi8371;// level 0
assign po8506 = pi8364;// level 0
assign po8507 = pi8336;// level 0
assign po8508 = pi8329;// level 0
assign po8509 = pi8338;// level 0
assign po8510 = pi8363;// level 0
assign po8511 = pi8346;// level 0
assign po8512 = pi8333;// level 0
assign po8513 = pi8361;// level 0
assign po8514 = pi8349;// level 0
assign po8515 = pi8326;// level 0
assign po8516 = pi8332;// level 0
assign po8517 = pi8356;// level 0
assign po8518 = pi8362;// level 0
assign po8519 = pi8347;// level 0
assign po8520 = pi8367;// level 0
assign po8521 = pi8352;// level 0
assign po8522 = pi8324;// level 0
assign po8523 = pi8330;// level 0
assign po8524 = pi8360;// level 0
assign po8525 = pi8322;// level 0
assign po8526 = pi8374;// level 0
assign po8527 = pi8343;// level 0
assign po8528 = pi8370;// level 0
assign po8529 = pi8337;// level 0
assign po8530 = pi8372;// level 0
assign po8531 = pi8355;// level 0
assign po8532 = pi8353;// level 0
assign po8533 = pi8345;// level 0
assign po8534 = pi8334;// level 0
assign po8535 = pi8335;// level 0
assign po8536 = pi8350;// level 0
assign po8537 = pi8359;// level 0
assign po8538 = pi8321;// level 0
assign po8539 = pi8375;// level 0
assign po8540 = pi8358;// level 0
assign po8541 = pi8351;// level 0
assign po8542 = pi8366;// level 0
assign po8543 = pi8323;// level 0
assign po8544 = pi8368;// level 0
assign po8545 = pi8342;// level 0
assign po8546 = pi8373;// level 0
assign po8547 = pi8344;// level 0
assign po8548 = pi8320;// level 0
assign po8549 = pi8357;// level 0
assign po8550 = pi8407;// level 0
assign po8551 = pi8383;// level 0
assign po8552 = pi8398;// level 0
assign po8553 = pi8418;// level 0
assign po8554 = pi8394;// level 0
assign po8555 = pi8382;// level 0
assign po8556 = pi8430;// level 0
assign po8557 = pi8409;// level 0
assign po8558 = pi8390;// level 0
assign po8559 = pi8389;// level 0
assign po8560 = pi8401;// level 0
assign po8561 = pi8406;// level 0
assign po8562 = pi8376;// level 0
assign po8563 = pi8427;// level 0
assign po8564 = pi8413;// level 0
assign po8565 = pi8379;// level 0
assign po8566 = pi8412;// level 0
assign po8567 = pi8403;// level 0
assign po8568 = pi8419;// level 0
assign po8569 = pi8391;// level 0
assign po8570 = pi8426;// level 0
assign po8571 = pi8425;// level 0
assign po8572 = pi8402;// level 0
assign po8573 = pi8414;// level 0
assign po8574 = pi8411;// level 0
assign po8575 = pi8385;// level 0
assign po8576 = pi8377;// level 0
assign po8577 = pi8395;// level 0
assign po8578 = pi8424;// level 0
assign po8579 = pi8423;// level 0
assign po8580 = pi8422;// level 0
assign po8581 = pi8408;// level 0
assign po8582 = pi8388;// level 0
assign po8583 = pi8393;// level 0
assign po8584 = pi8387;// level 0
assign po8585 = pi8392;// level 0
assign po8586 = pi8410;// level 0
assign po8587 = pi8380;// level 0
assign po8588 = pi8396;// level 0
assign po8589 = pi8421;// level 0
assign po8590 = pi8386;// level 0
assign po8591 = pi8420;// level 0
assign po8592 = pi8381;// level 0
assign po8593 = pi8384;// level 0
assign po8594 = pi8429;// level 0
assign po8595 = pi8431;// level 0
assign po8596 = pi8416;// level 0
assign po8597 = pi8397;// level 0
assign po8598 = pi8378;// level 0
assign po8599 = pi8400;// level 0
assign po8600 = pi8417;// level 0
assign po8601 = pi8399;// level 0
assign po8602 = pi8405;// level 0
assign po8603 = pi8404;// level 0
assign po8604 = pi8428;// level 0
assign po8605 = pi8415;// level 0
assign po8606 = pi8463;// level 0
assign po8607 = pi8480;// level 0
assign po8608 = pi8481;// level 0
assign po8609 = pi8456;// level 0
assign po8610 = pi8439;// level 0
assign po8611 = pi8455;// level 0
assign po8612 = pi8447;// level 0
assign po8613 = pi8451;// level 0
assign po8614 = pi8448;// level 0
assign po8615 = pi8437;// level 0
assign po8616 = pi8436;// level 0
assign po8617 = pi8457;// level 0
assign po8618 = pi8468;// level 0
assign po8619 = pi8452;// level 0
assign po8620 = pi8446;// level 0
assign po8621 = pi8469;// level 0
assign po8622 = pi8434;// level 0
assign po8623 = pi8484;// level 0
assign po8624 = pi8474;// level 0
assign po8625 = pi8473;// level 0
assign po8626 = pi8466;// level 0
assign po8627 = pi8470;// level 0
assign po8628 = pi8485;// level 0
assign po8629 = pi8433;// level 0
assign po8630 = pi8479;// level 0
assign po8631 = pi8432;// level 0
assign po8632 = pi8454;// level 0
assign po8633 = pi8453;// level 0
assign po8634 = pi8444;// level 0
assign po8635 = pi8461;// level 0
assign po8636 = pi8460;// level 0
assign po8637 = pi8482;// level 0
assign po8638 = pi8443;// level 0
assign po8639 = pi8458;// level 0
assign po8640 = pi8449;// level 0
assign po8641 = pi8467;// level 0
assign po8642 = pi8487;// level 0
assign po8643 = pi8486;// level 0
assign po8644 = pi8464;// level 0
assign po8645 = pi8478;// level 0
assign po8646 = pi8440;// level 0
assign po8647 = pi8472;// level 0
assign po8648 = pi8477;// level 0
assign po8649 = pi8476;// level 0
assign po8650 = pi8459;// level 0
assign po8651 = pi8475;// level 0
assign po8652 = pi8438;// level 0
assign po8653 = pi8462;// level 0
assign po8654 = pi8441;// level 0
assign po8655 = pi8471;// level 0
assign po8656 = pi8435;// level 0
assign po8657 = pi8483;// level 0
assign po8658 = pi8445;// level 0
assign po8659 = pi8442;// level 0
assign po8660 = pi8465;// level 0
assign po8661 = pi8450;// level 0
assign po8662 = pi8493;// level 0
assign po8663 = pi8542;// level 0
assign po8664 = pi8510;// level 0
assign po8665 = pi8512;// level 0
assign po8666 = pi8515;// level 0
assign po8667 = pi8508;// level 0
assign po8668 = pi8495;// level 0
assign po8669 = pi8524;// level 0
assign po8670 = pi8527;// level 0
assign po8671 = pi8513;// level 0
assign po8672 = pi8505;// level 0
assign po8673 = pi8517;// level 0
assign po8674 = pi8529;// level 0
assign po8675 = pi8500;// level 0
assign po8676 = pi8534;// level 0
assign po8677 = pi8525;// level 0
assign po8678 = pi8546;// level 0
assign po8679 = pi8492;// level 0
assign po8680 = pi8543;// level 0
assign po8681 = pi8537;// level 0
assign po8682 = pi8504;// level 0
assign po8683 = pi8496;// level 0
assign po8684 = pi8516;// level 0
assign po8685 = pi8545;// level 0
assign po8686 = pi8535;// level 0
assign po8687 = pi8541;// level 0
assign po8688 = pi8540;// level 0
assign po8689 = pi8532;// level 0
assign po8690 = pi8533;// level 0
assign po8691 = pi8523;// level 0
assign po8692 = pi8536;// level 0
assign po8693 = pi8498;// level 0
assign po8694 = pi8531;// level 0
assign po8695 = pi8522;// level 0
assign po8696 = pi8490;// level 0
assign po8697 = pi8502;// level 0
assign po8698 = pi8518;// level 0
assign po8699 = pi8530;// level 0
assign po8700 = pi8544;// level 0
assign po8701 = pi8521;// level 0
assign po8702 = pi8488;// level 0
assign po8703 = pi8489;// level 0
assign po8704 = pi8526;// level 0
assign po8705 = pi8501;// level 0
assign po8706 = pi8519;// level 0
assign po8707 = pi8514;// level 0
assign po8708 = pi8538;// level 0
assign po8709 = pi8497;// level 0
assign po8710 = pi8509;// level 0
assign po8711 = pi8506;// level 0
assign po8712 = pi8511;// level 0
assign po8713 = pi8499;// level 0
assign po8714 = pi8491;// level 0
assign po8715 = pi8494;// level 0
assign po8716 = pi8539;// level 0
assign po8717 = pi8507;// level 0
assign po8718 = pi8617;// level 0
assign po8719 = pi8596;// level 0
assign po8720 = pi8562;// level 0
assign po8721 = pi8604;// level 0
assign po8722 = pi8608;// level 0
assign po8723 = pi8588;// level 0
assign po8724 = pi8586;// level 0
assign po8725 = pi8618;// level 0
assign po8726 = pi8577;// level 0
assign po8727 = pi8595;// level 0
assign po8728 = pi8593;// level 0
assign po8729 = pi8574;// level 0
assign po8730 = pi8551;// level 0
assign po8731 = pi8581;// level 0
assign po8732 = pi8567;// level 0
assign po8733 = pi8742;// level 0
assign po8734 = pi8578;// level 0
assign po8735 = pi8623;// level 0
assign po8736 = pi8614;// level 0
assign po8737 = pi8611;// level 0
assign po8738 = pi8612;// level 0
assign po8739 = pi8563;// level 0
assign po8740 = pi8566;// level 0
assign po8741 = pi8589;// level 0
assign po8742 = pi8571;// level 0
assign po8743 = pi8626;// level 0
assign po8744 = pi8587;// level 0
assign po8745 = pi8552;// level 0
assign po8746 = pi8564;// level 0
assign po8747 = pi8616;// level 0
assign po8748 = pi8573;// level 0
assign po8749 = pi8610;// level 0
assign po8750 = pi8752;// level 0
assign po8751 = pi8591;// level 0
assign po8752 = pi8607;// level 0
assign po8753 = pi8620;// level 0
assign po8754 = pi8572;// level 0
assign po8755 = pi8576;// level 0
assign po8756 = pi8560;// level 0
assign po8757 = pi8584;// level 0
assign po8758 = pi8802;// level 0
assign po8759 = pi8553;// level 0
assign po8760 = pi8619;// level 0
assign po8761 = pi8598;// level 0
assign po8762 = pi8627;// level 0
assign po8763 = pi8606;// level 0
assign po8764 = pi8603;// level 0
assign po8765 = pi8555;// level 0
assign po8766 = pi8621;// level 0
assign po8767 = pi8569;// level 0
assign po8768 = pi8625;// level 0
assign po8769 = pi8558;// level 0
assign po8770 = pi8613;// level 0
assign po8771 = pi8599;// level 0
assign po8772 = pi8580;// level 0
assign po8773 = pi8565;// level 0
assign po8774 = pi8609;// level 0
assign po8775 = pi8597;// level 0
assign po8776 = pi8590;// level 0
assign po8777 = pi8748;// level 0
assign po8778 = pi8713;// level 0
assign po8779 = pi8712;// level 0
assign po8780 = pi8726;// level 0
assign po8781 = pi8687;// level 0
assign po8782 = pi8653;// level 0
assign po8783 = pi8631;// level 0
assign po8784 = pi8782;// level 0
assign po8785 = pi8661;// level 0
assign po8786 = pi8766;// level 0
assign po8787 = pi8761;// level 0
assign po8788 = pi8657;// level 0
assign po8789 = pi8803;// level 0
assign po8790 = pi8658;// level 0
assign po8791 = pi8796;// level 0
assign po8792 = pi8632;// level 0
assign po8793 = pi8683;// level 0
assign po8794 = pi8676;// level 0
assign po8795 = pi8636;// level 0
assign po8796 = pi8679;// level 0
assign po8797 = pi8643;// level 0
assign po8798 = pi8727;// level 0
assign po8799 = pi8674;// level 0
assign po8800 = pi8776;// level 0
assign po8801 = pi8656;// level 0
assign po8802 = pi8677;// level 0
assign po8803 = pi8647;// level 0
assign po8804 = pi8655;// level 0
assign po8805 = pi8781;// level 0
assign po8806 = pi8639;// level 0
assign po8807 = pi8659;// level 0
assign po8808 = pi8663;// level 0
assign po8809 = pi8717;// level 0
assign po8810 = pi8654;// level 0
assign po8811 = pi8641;// level 0
assign po8812 = pi8743;// level 0
assign po8813 = pi8719;// level 0
assign po8814 = pi8640;// level 0
assign po8815 = pi8773;// level 0
assign po8816 = pi8644;// level 0
assign po8817 = pi8637;// level 0
assign po8818 = pi8686;// level 0
assign po8819 = pi8634;// level 0
assign po8820 = pi8638;// level 0
assign po8821 = pi8672;// level 0
assign po8822 = pi8795;// level 0
assign po8823 = pi8667;// level 0
assign po8824 = pi8738;// level 0
assign po8825 = pi8645;// level 0
assign po8826 = pi8662;// level 0
assign po8827 = pi8642;// level 0
assign po8828 = pi8673;// level 0
assign po8829 = pi8664;// level 0
assign po8830 = pi8715;// level 0
assign po8831 = pi8778;// level 0
assign po8832 = pi8775;// level 0
assign po8833 = pi8652;// level 0
assign po8834 = pi8660;// level 0
assign po8835 = pi8705;// level 0
assign po8836 = pi8650;// level 0
assign po8837 = pi8630;// level 0
assign po8838 = pi8648;// level 0
assign po8839 = pi8681;// level 0
assign po8840 = pi8668;// level 0
assign po8841 = pi8670;// level 0
assign po8842 = pi8675;// level 0
assign po8843 = pi8635;// level 0
assign po8844 = pi8628;// level 0
assign po8845 = pi8750;// level 0
assign po8846 = pi8684;// level 0
assign po8847 = pi8680;// level 0
assign po8848 = pi8669;// level 0
assign po8849 = pi8646;// level 0
assign po8850 = pi8671;// level 0
assign po8851 = pi8651;// level 0
assign po8852 = pi8798;// level 0
assign po8853 = pi8682;// level 0
assign po8854 = pi8799;// level 0
assign po8855 = pi8665;// level 0
assign po8856 = pi8649;// level 0
assign po8857 = pi8666;// level 0
assign po8858 = pi8794;// level 0
assign po8859 = pi8807;// level 0
assign po8860 = pi8737;// level 0
assign po8861 = pi8732;// level 0
assign po8862 = pi8792;// level 0
assign po8863 = pi8702;// level 0
assign po8864 = pi8774;// level 0
assign po8865 = pi8791;// level 0
assign po8866 = pi8731;// level 0
assign po8867 = pi8733;// level 0
assign po8868 = pi8694;// level 0
assign po8869 = pi8756;// level 0
assign po8870 = pi8758;// level 0
assign po8871 = pi8801;// level 0
assign po8872 = pi8706;// level 0
assign po8873 = pi8711;// level 0
assign po8874 = pi8703;// level 0
assign po8875 = pi8730;// level 0
assign po8876 = pi8740;// level 0
assign po8877 = pi8800;// level 0
assign po8878 = pi8757;// level 0
assign po8879 = pi8739;// level 0
assign po8880 = pi8741;// level 0
assign po8881 = pi8699;// level 0
assign po8882 = pi8759;// level 0
assign po8883 = pi8764;// level 0
assign po8884 = pi8692;// level 0
assign po8885 = pi8690;// level 0
assign po8886 = pi8691;// level 0
assign po8887 = pi8760;// level 0
assign po8888 = pi8698;// level 0
assign po8889 = pi8700;// level 0
assign po8890 = pi8786;// level 0
assign po8891 = pi8704;// level 0
assign po8892 = pi8708;// level 0
assign po8893 = pi8785;// level 0
assign po8894 = pi8736;// level 0
assign po8895 = pi8724;// level 0
assign po8896 = pi8789;// level 0
assign po8897 = pi8805;// level 0
assign po8898 = pi8762;// level 0
assign po8899 = pi8689;// level 0
assign po8900 = pi8777;// level 0
assign po8901 = pi8745;// level 0
assign po8902 = pi8804;// level 0
assign po8903 = pi8770;// level 0
assign po8904 = pi8746;// level 0
assign po8905 = pi8707;// level 0
assign po8906 = pi8723;// level 0
assign po8907 = pi8688;// level 0
assign po8908 = pi8772;// level 0
assign po8909 = pi8735;// level 0
assign po8910 = pi8728;// level 0
assign po8911 = pi8734;// level 0
assign po8912 = pi8783;// level 0
assign po8913 = pi8769;// level 0
assign po8914 = pi8780;// level 0
assign po8915 = pi8710;// level 0
assign po8916 = pi8763;// level 0
assign po8917 = pi8806;// level 0
assign po8918 = pi8951;// level 0
assign po8919 = pi8947;// level 0
assign po8920 = pi8966;// level 0
assign po8921 = pi8941;// level 0
assign po8922 = pi8932;// level 0
assign po8923 = pi8818;// level 0
assign po8924 = pi8975;// level 0
assign po8925 = pi8834;// level 0
assign po8926 = pi8840;// level 0
assign po8927 = pi8808;// level 0
assign po8928 = pi8963;// level 0
assign po8929 = pi8958;// level 0
assign po8930 = pi8961;// level 0
assign po8931 = pi8816;// level 0
assign po8932 = pi8827;// level 0
assign po8933 = pi8979;// level 0
assign po8934 = pi8952;// level 0
assign po8935 = pi8841;// level 0
assign po8936 = pi8943;// level 0
assign po8937 = pi8971;// level 0
assign po8938 = pi8972;// level 0
assign po8939 = pi8850;// level 0
assign po8940 = pi8825;// level 0
assign po8941 = pi8956;// level 0
assign po8942 = pi8833;// level 0
assign po8943 = pi8871;// level 0
assign po8944 = pi8826;// level 0
assign po8945 = pi8823;// level 0
assign po8946 = pi8828;// level 0
assign po8947 = pi8817;// level 0
assign po8948 = pi8862;// level 0
assign po8949 = pi8815;// level 0
assign po8950 = pi8830;// level 0
assign po8951 = pi8854;// level 0
assign po8952 = pi8820;// level 0
assign po8953 = pi8939;// level 0
assign po8954 = pi8970;// level 0
assign po8955 = pi8842;// level 0
assign po8956 = pi8863;// level 0
assign po8957 = pi8851;// level 0
assign po8958 = pi8938;// level 0
assign po8959 = pi8844;// level 0
assign po8960 = pi8981;// level 0
assign po8961 = pi8967;// level 0
assign po8962 = pi8945;// level 0
assign po8963 = pi8973;// level 0
assign po8964 = pi8965;// level 0
assign po8965 = pi8937;// level 0
assign po8966 = pi8959;// level 0
assign po8967 = pi8982;// level 0
assign po8968 = pi8859;// level 0
assign po8969 = pi8968;// level 0
assign po8970 = pi8928;// level 0
assign po8971 = pi8977;// level 0
assign po8972 = pi8835;// level 0
assign po8973 = pi8855;// level 0
assign po8974 = pi8870;// level 0
assign po8975 = pi8936;// level 0
assign po8976 = pi8946;// level 0
assign po8977 = pi8866;// level 0
assign po8978 = pi8809;// level 0
assign po8979 = pi8846;// level 0
assign po8980 = pi8813;// level 0
assign po8981 = pi8810;// level 0
assign po8982 = pi8869;// level 0
assign po8983 = pi8868;// level 0
assign po8984 = pi8856;// level 0
assign po8985 = pi8824;// level 0
assign po8986 = pi8957;// level 0
assign po8987 = pi8969;// level 0
assign po8988 = pi8934;// level 0
assign po8989 = pi8935;// level 0
assign po8990 = pi8940;// level 0
assign po8991 = pi8847;// level 0
assign po8992 = pi8955;// level 0
assign po8993 = pi8933;// level 0
assign po8994 = pi8949;// level 0
assign po8995 = pi8822;// level 0
assign po8996 = pi8857;// level 0
assign po8997 = pi8858;// level 0
assign po8998 = pi8860;// level 0
assign po8999 = pi8948;// level 0
assign po9000 = pi8962;// level 0
assign po9001 = pi8832;// level 0
assign po9002 = pi8861;// level 0
assign po9003 = pi8845;// level 0
assign po9004 = pi8976;// level 0
assign po9005 = pi8837;// level 0
assign po9006 = pi8839;// level 0
assign po9007 = pi8953;// level 0
assign po9008 = pi8853;// level 0
assign po9009 = pi8814;// level 0
assign po9010 = pi8964;// level 0
assign po9011 = pi8811;// level 0
assign po9012 = pi8821;// level 0
assign po9013 = pi8942;// level 0
assign po9014 = pi8848;// level 0
assign po9015 = pi8974;// level 0
assign po9016 = pi8960;// level 0
assign po9017 = pi8864;// level 0
assign po9018 = pi8836;// level 0
assign po9019 = pi8954;// level 0
assign po9020 = pi8838;// level 0
assign po9021 = pi8930;// level 0
assign po9022 = pi8929;// level 0
assign po9023 = pi8852;// level 0
assign po9024 = pi8983;// level 0
assign po9025 = pi8829;// level 0
assign po9026 = pi8865;// level 0
assign po9027 = pi8812;// level 0
assign po9028 = pi8831;// level 0
assign po9029 = pi8819;// level 0
assign po9030 = pi8950;// level 0
assign po9031 = pi8980;// level 0
assign po9032 = pi8867;// level 0
assign po9033 = pi8843;// level 0
assign po9034 = pi8931;// level 0
assign po9035 = pi8944;// level 0
assign po9036 = pi8978;// level 0
assign po9037 = pi8849;// level 0
endmodule
