module MUL32 ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63;
  wire n130, n131, n132, n133, n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n154,
    n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
    n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234, n235, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
    n301, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n382, n383, n384, n385, n386,
    n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n560, n561, n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
    n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n914, n915, n916, n917, n918, n919,
    n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
    n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
    n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
    n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
    n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
    n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
    n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
    n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
    n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
    n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
    n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
    n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
    n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
    n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
    n2712, n2713, n2714, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
    n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
    n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
    n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
    n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
    n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
    n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
    n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
    n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
    n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
    n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
    n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
    n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
    n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
    n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
    n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
    n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
    n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
    n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
    n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
    n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
    n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
    n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
    n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
    n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
    n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
    n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
    n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
    n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
    n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
    n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
    n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
    n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
    n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
    n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5166, n5167, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
    n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
    n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
    n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
    n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
    n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
    n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
    n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
    n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
    n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
    n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
    n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
    n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
    n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
    n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
    n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
    n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
    n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
    n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
    n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
    n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
    n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
    n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
    n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5803,
    n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
    n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
    n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
    n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
    n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
    n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
    n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
    n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
    n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
    n6104, n6105, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
    n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
    n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
    n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
    n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
    n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
    n6425, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
    n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
    n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
    n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
    n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
    n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
    n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
    n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
    n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
    n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
    n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
    n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
    n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
    n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
    n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
    n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
    n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
    n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
    n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
    n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
    n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
    n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
    n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
    n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
    n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
    n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
    n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794, n7796, n7797, n7798, n7799,
    n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
    n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
    n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
    n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
    n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
    n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
    n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
    n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
    n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
    n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
    n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
    n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
    n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
    n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
    n8050, n8051, n8052, n8053, n8054, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
    n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
    n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
    n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
    n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
    n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
    n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
    n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
    n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
    n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
    n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
    n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
    n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
    n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
    n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
    n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
    n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
    n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
    n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
    n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
    n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
    n8632, n8633, n8634, n8635, n8636, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
    n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
    n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
    n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
    n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
    n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
    n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
    n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
    n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
    n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
    n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
    n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
    n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
    n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
    n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
    n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
    n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9614, n9615, n9616,
    n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
    n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
    n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
    n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
    n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
    n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
    n9797, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
    n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
    n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
    n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
    n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
    n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
    n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
    n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
    n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
    n9968, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
    n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
    n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
    n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
    n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
    n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
    n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
    n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
    n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
    n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10160, n10161,
    n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
    n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
    n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
    n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
    n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
    n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
    n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
    n10315, n10316, n10317, n10318, n10320, n10321, n10322, n10323, n10324,
    n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
    n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
    n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
    n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
    n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
    n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
    n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
    n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
    n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
    n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
    n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
    n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
    n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
    n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
    n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
    n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
    n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
    n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
    n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
    n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10798, n10799, n10801, n10802, n10803, n10804,
    n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
    n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
    n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
    n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
    n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
    n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
    n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
    n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
    n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
    n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
    n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
    n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
    n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081, n11083, n11084, n11085,
    n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
    n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
    n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
    n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
    n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
    n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
    n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
    n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
    n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
    n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
    n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
    n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
    n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
    n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
    n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
    n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
    n11485, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
    n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11622,
    n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
    n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
    n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
    n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
    n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
    n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
    n11677, n11678, n11679, n11680, n11681, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
    n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
    n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740;
  assign po00 = pi00 & pi32;
  assign n130 = pi00 & pi33;
  assign n131 = pi01 & pi32;
  assign n132 = ~n130 & n131;
  assign n133 = n130 & ~n131;
  assign po01 = n132 | n133;
  assign n135 = pi01 & ~pi32;
  assign n136 = pi02 & pi32;
  assign n137 = pi33 & ~n136;
  assign n138 = ~n135 & n137;
  assign n139 = ~pi33 & n136;
  assign n140 = ~n138 & ~n139;
  assign n141 = pi33 & ~pi34;
  assign n142 = ~pi33 & pi34;
  assign n143 = ~n141 & ~n142;
  assign n144 = pi00 & ~n143;
  assign n145 = ~n140 & n144;
  assign n146 = n140 & ~n144;
  assign n147 = ~n145 & ~n146;
  assign n148 = ~pi00 & pi33;
  assign n149 = ~n131 & n148;
  assign n150 = ~n147 & ~n149;
  assign n151 = ~n145 & n149;
  assign n152 = ~n146 & n151;
  assign po02 = ~n150 & ~n152;
  assign n154 = pi34 & ~pi35;
  assign n155 = ~pi34 & pi35;
  assign n156 = ~n154 & ~n155;
  assign n157 = pi00 & ~n141;
  assign n158 = ~n142 & n157;
  assign n159 = ~n156 & n158;
  assign n160 = pi01 & ~n143;
  assign n161 = ~n159 & ~n160;
  assign n162 = pi35 & ~n161;
  assign n163 = ~pi35 & ~n160;
  assign n164 = ~n159 & n163;
  assign n165 = pi02 & ~pi32;
  assign n166 = pi03 & pi32;
  assign n167 = pi33 & ~n166;
  assign n168 = ~n165 & n167;
  assign n169 = ~pi33 & n166;
  assign n170 = ~n168 & ~n169;
  assign n171 = ~n164 & ~n170;
  assign n172 = ~n162 & n171;
  assign n173 = ~n162 & ~n164;
  assign n174 = n170 & ~n173;
  assign n175 = ~n172 & ~n174;
  assign n176 = pi35 & ~n144;
  assign n177 = ~n145 & ~n176;
  assign n178 = ~n175 & n177;
  assign n179 = ~n172 & ~n177;
  assign n180 = ~n174 & n179;
  assign n181 = ~n178 & ~n180;
  assign n182 = ~n152 & ~n181;
  assign n183 = n152 & ~n180;
  assign n184 = ~n178 & n183;
  assign po03 = ~n182 & ~n184;
  assign n186 = ~n180 & ~n184;
  assign n187 = pi01 & ~n141;
  assign n188 = ~n142 & n187;
  assign n189 = ~n156 & n188;
  assign n190 = pi02 & ~n143;
  assign n191 = ~n189 & ~n190;
  assign n192 = pi35 & ~n191;
  assign n193 = pi35 & ~pi36;
  assign n194 = ~pi35 & pi36;
  assign n195 = ~n193 & ~n194;
  assign n196 = pi00 & ~n195;
  assign n197 = pi37 & ~n196;
  assign n198 = pi00 & ~pi37;
  assign n199 = ~n195 & n198;
  assign n200 = ~n197 & ~n199;
  assign n201 = ~pi35 & ~n190;
  assign n202 = ~n189 & n201;
  assign n203 = pi03 & ~pi32;
  assign n204 = pi04 & pi32;
  assign n205 = pi33 & ~n204;
  assign n206 = ~n203 & n205;
  assign n207 = ~pi33 & n204;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~n202 & ~n208;
  assign n210 = ~n200 & n209;
  assign n211 = ~n192 & n210;
  assign n212 = ~pi37 & ~n170;
  assign n213 = ~n164 & n212;
  assign n214 = ~n162 & n213;
  assign n215 = ~n211 & ~n214;
  assign n216 = ~n192 & ~n202;
  assign n217 = n200 & ~n208;
  assign n218 = ~n216 & n217;
  assign n219 = ~n200 & n208;
  assign n220 = ~n216 & n219;
  assign n221 = ~n218 & ~n220;
  assign n222 = n200 & n208;
  assign n223 = n216 & n222;
  assign n224 = pi37 & ~n172;
  assign n225 = ~n223 & ~n224;
  assign n226 = n221 & n225;
  assign n227 = n215 & n226;
  assign n228 = ~n211 & ~n218;
  assign n229 = ~n220 & ~n223;
  assign n230 = n228 & n229;
  assign n231 = ~n214 & ~n224;
  assign n232 = ~n230 & ~n231;
  assign n233 = ~n227 & ~n232;
  assign n234 = ~n186 & n233;
  assign n235 = n186 & ~n233;
  assign po04 = ~n234 & ~n235;
  assign n237 = pi04 & ~pi32;
  assign n238 = pi05 & pi32;
  assign n239 = pi33 & ~n238;
  assign n240 = ~n237 & n239;
  assign n241 = ~pi33 & n238;
  assign n242 = ~n240 & ~n241;
  assign n243 = pi03 & ~n143;
  assign n244 = pi02 & pi33;
  assign n245 = n154 & n244;
  assign n246 = pi02 & ~pi33;
  assign n247 = n155 & n246;
  assign n248 = ~n245 & ~n247;
  assign n249 = ~n243 & n248;
  assign n250 = pi35 & ~n249;
  assign n251 = ~pi35 & ~n245;
  assign n252 = ~n247 & n251;
  assign n253 = ~n243 & n252;
  assign n254 = ~n250 & ~n253;
  assign n255 = pi01 & ~n195;
  assign n256 = pi35 & pi36;
  assign n257 = n198 & n256;
  assign n258 = pi00 & ~pi35;
  assign n259 = ~pi36 & pi37;
  assign n260 = n258 & n259;
  assign n261 = ~n257 & ~n260;
  assign n262 = ~n255 & n261;
  assign n263 = pi37 & ~n262;
  assign n264 = ~pi37 & ~n257;
  assign n265 = ~n260 & n264;
  assign n266 = ~n255 & n265;
  assign n267 = ~n263 & ~n266;
  assign n268 = n254 & n267;
  assign n269 = ~n254 & ~n267;
  assign n270 = ~n268 & ~n269;
  assign n271 = n242 & ~n270;
  assign n272 = ~n242 & ~n268;
  assign n273 = ~n269 & n272;
  assign n274 = n200 & ~n216;
  assign n275 = ~n200 & ~n202;
  assign n276 = ~n192 & n275;
  assign n277 = n208 & ~n276;
  assign n278 = ~n274 & ~n277;
  assign n279 = ~n273 & n278;
  assign n280 = ~n271 & n279;
  assign n281 = ~n271 & ~n273;
  assign n282 = ~n278 & ~n281;
  assign n283 = ~n280 & ~n282;
  assign n284 = pi37 & ~n170;
  assign n285 = ~n164 & n284;
  assign n286 = ~n162 & n285;
  assign n287 = ~n232 & ~n286;
  assign n288 = n283 & ~n287;
  assign n289 = ~n283 & n287;
  assign n290 = n180 & ~n227;
  assign n291 = ~n232 & n290;
  assign n292 = ~n289 & n291;
  assign n293 = ~n288 & n292;
  assign n294 = ~n288 & ~n289;
  assign n295 = ~n291 & ~n294;
  assign n296 = ~n293 & ~n295;
  assign n297 = n184 & ~n227;
  assign n298 = ~n232 & n297;
  assign n299 = ~n296 & ~n298;
  assign n300 = ~n293 & n298;
  assign n301 = ~n295 & n300;
  assign po05 = ~n299 & ~n301;
  assign n303 = ~n280 & ~n288;
  assign n304 = pi37 & ~pi38;
  assign n305 = ~pi37 & pi38;
  assign n306 = ~n304 & ~n305;
  assign n307 = pi00 & ~n306;
  assign n308 = ~n242 & ~n307;
  assign n309 = ~n263 & n308;
  assign n310 = ~n266 & n309;
  assign n311 = ~n250 & n308;
  assign n312 = ~n253 & n311;
  assign n313 = ~n310 & ~n312;
  assign n314 = n242 & n307;
  assign n315 = ~n267 & n314;
  assign n316 = ~n254 & n314;
  assign n317 = ~n315 & ~n316;
  assign n318 = n313 & n317;
  assign n319 = ~n250 & ~n307;
  assign n320 = ~n253 & ~n263;
  assign n321 = ~n266 & n320;
  assign n322 = n319 & n321;
  assign n323 = ~n254 & n307;
  assign n324 = ~n267 & n323;
  assign n325 = ~n322 & ~n324;
  assign n326 = n318 & n325;
  assign n327 = pi04 & ~n143;
  assign n328 = pi03 & pi33;
  assign n329 = n154 & n328;
  assign n330 = pi03 & ~pi33;
  assign n331 = n155 & n330;
  assign n332 = ~n329 & ~n331;
  assign n333 = ~n327 & n332;
  assign n334 = pi35 & ~n333;
  assign n335 = ~pi35 & ~n329;
  assign n336 = ~n331 & n335;
  assign n337 = ~n327 & n336;
  assign n338 = ~n334 & ~n337;
  assign n339 = pi02 & ~n195;
  assign n340 = pi01 & pi35;
  assign n341 = pi36 & ~pi37;
  assign n342 = n340 & n341;
  assign n343 = pi01 & ~pi35;
  assign n344 = n259 & n343;
  assign n345 = ~n342 & ~n344;
  assign n346 = ~n339 & n345;
  assign n347 = pi37 & ~n346;
  assign n348 = ~pi37 & ~n342;
  assign n349 = ~n344 & n348;
  assign n350 = ~n339 & n349;
  assign n351 = ~n347 & ~n350;
  assign n352 = ~n338 & ~n351;
  assign n353 = n338 & n351;
  assign n354 = pi05 & ~pi32;
  assign n355 = pi06 & pi32;
  assign n356 = pi33 & ~n355;
  assign n357 = ~n354 & n356;
  assign n358 = ~pi33 & n355;
  assign n359 = ~n357 & ~n358;
  assign n360 = ~n353 & ~n359;
  assign n361 = ~n352 & n360;
  assign n362 = ~n352 & ~n353;
  assign n363 = n359 & ~n362;
  assign n364 = ~n361 & ~n363;
  assign n365 = ~n326 & n364;
  assign n366 = n326 & ~n364;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~n303 & n367;
  assign n369 = ~n280 & ~n367;
  assign n370 = ~n288 & n369;
  assign n371 = ~n368 & ~n370;
  assign n372 = ~n293 & ~n371;
  assign n373 = ~n301 & n372;
  assign n374 = n298 & ~n370;
  assign n375 = ~n293 & n374;
  assign n376 = ~n295 & ~n368;
  assign n377 = n375 & n376;
  assign n378 = n293 & ~n370;
  assign n379 = ~n368 & n378;
  assign n380 = ~n377 & ~n379;
  assign po06 = ~n373 & n380;
  assign n382 = pi39 & ~n307;
  assign n383 = ~n361 & n382;
  assign n384 = ~n363 & n383;
  assign n385 = ~n326 & n384;
  assign n386 = ~n242 & ~n269;
  assign n387 = ~n268 & ~n386;
  assign n388 = n307 & ~n387;
  assign n389 = ~n382 & ~n388;
  assign n390 = ~n365 & n389;
  assign n391 = ~n385 & ~n390;
  assign n392 = pi38 & ~pi39;
  assign n393 = ~pi38 & pi39;
  assign n394 = ~n392 & ~n393;
  assign n395 = pi00 & ~n304;
  assign n396 = ~n305 & n395;
  assign n397 = ~n394 & n396;
  assign n398 = pi01 & ~n306;
  assign n399 = ~n397 & ~n398;
  assign n400 = pi39 & ~n399;
  assign n401 = ~pi39 & ~n398;
  assign n402 = ~n397 & n401;
  assign n403 = ~n400 & ~n402;
  assign n404 = ~n352 & ~n359;
  assign n405 = ~n353 & ~n404;
  assign n406 = n403 & ~n405;
  assign n407 = ~n353 & ~n403;
  assign n408 = ~n404 & n407;
  assign n409 = pi05 & ~n143;
  assign n410 = pi04 & pi33;
  assign n411 = n154 & n410;
  assign n412 = pi04 & ~pi33;
  assign n413 = n155 & n412;
  assign n414 = ~n411 & ~n413;
  assign n415 = ~n409 & n414;
  assign n416 = pi35 & ~n415;
  assign n417 = ~pi35 & ~n411;
  assign n418 = ~n413 & n417;
  assign n419 = ~n409 & n418;
  assign n420 = ~n416 & ~n419;
  assign n421 = pi03 & ~n195;
  assign n422 = pi02 & pi35;
  assign n423 = n341 & n422;
  assign n424 = pi02 & ~pi35;
  assign n425 = n259 & n424;
  assign n426 = ~n423 & ~n425;
  assign n427 = ~n421 & n426;
  assign n428 = pi37 & ~n427;
  assign n429 = ~pi37 & ~n423;
  assign n430 = ~n425 & n429;
  assign n431 = ~n421 & n430;
  assign n432 = ~n428 & ~n431;
  assign n433 = ~n420 & ~n432;
  assign n434 = n420 & n432;
  assign n435 = pi06 & ~pi32;
  assign n436 = pi07 & pi32;
  assign n437 = pi33 & ~n436;
  assign n438 = ~n435 & n437;
  assign n439 = ~pi33 & n436;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n434 & ~n440;
  assign n442 = ~n433 & n441;
  assign n443 = ~n433 & ~n434;
  assign n444 = n440 & ~n443;
  assign n445 = ~n442 & ~n444;
  assign n446 = ~n408 & n445;
  assign n447 = ~n406 & n446;
  assign n448 = ~n406 & ~n408;
  assign n449 = ~n445 & ~n448;
  assign n450 = ~n447 & ~n449;
  assign n451 = ~n391 & n450;
  assign n452 = n391 & ~n450;
  assign n453 = ~n451 & ~n452;
  assign n454 = n283 & n367;
  assign n455 = ~n287 & n454;
  assign n456 = n280 & ~n365;
  assign n457 = ~n366 & n456;
  assign n458 = n455 & ~n457;
  assign n459 = n453 & n458;
  assign n460 = ~n451 & n457;
  assign n461 = ~n452 & ~n455;
  assign n462 = n460 & n461;
  assign n463 = ~n455 & ~n457;
  assign n464 = ~n453 & n463;
  assign n465 = ~n462 & ~n464;
  assign n466 = ~n459 & n465;
  assign n467 = n379 & ~n466;
  assign n468 = ~n379 & n466;
  assign n469 = ~n467 & ~n468;
  assign n470 = n377 & ~n469;
  assign n471 = ~n377 & ~n467;
  assign n472 = ~n468 & n471;
  assign po07 = n470 | n472;
  assign n474 = n377 & ~n468;
  assign n475 = ~n453 & n457;
  assign n476 = ~n453 & n458;
  assign n477 = ~n475 & ~n476;
  assign n478 = ~n406 & ~n447;
  assign n479 = ~n433 & ~n440;
  assign n480 = ~n434 & ~n479;
  assign n481 = pi01 & ~n304;
  assign n482 = ~n305 & n481;
  assign n483 = ~n394 & n482;
  assign n484 = pi02 & ~n306;
  assign n485 = ~n483 & ~n484;
  assign n486 = pi39 & ~n485;
  assign n487 = ~pi39 & ~n484;
  assign n488 = ~n483 & n487;
  assign n489 = pi39 & ~pi40;
  assign n490 = ~pi39 & pi40;
  assign n491 = ~n489 & ~n490;
  assign n492 = pi00 & ~n491;
  assign n493 = ~n488 & ~n492;
  assign n494 = ~n486 & n493;
  assign n495 = ~n486 & ~n488;
  assign n496 = n492 & ~n495;
  assign n497 = ~n494 & ~n496;
  assign n498 = ~n480 & ~n497;
  assign n499 = ~n434 & ~n494;
  assign n500 = ~n479 & n499;
  assign n501 = ~n496 & n500;
  assign n502 = pi06 & ~n143;
  assign n503 = pi05 & pi33;
  assign n504 = n154 & n503;
  assign n505 = pi05 & ~pi33;
  assign n506 = n155 & n505;
  assign n507 = ~n504 & ~n506;
  assign n508 = ~n502 & n507;
  assign n509 = pi35 & ~n508;
  assign n510 = ~pi35 & ~n504;
  assign n511 = ~n506 & n510;
  assign n512 = ~n502 & n511;
  assign n513 = ~n509 & ~n512;
  assign n514 = pi04 & ~n195;
  assign n515 = pi03 & pi35;
  assign n516 = n341 & n515;
  assign n517 = pi03 & ~pi35;
  assign n518 = n259 & n517;
  assign n519 = ~n516 & ~n518;
  assign n520 = ~n514 & n519;
  assign n521 = pi37 & ~n520;
  assign n522 = ~pi37 & ~n516;
  assign n523 = ~n518 & n522;
  assign n524 = ~n514 & n523;
  assign n525 = ~n521 & ~n524;
  assign n526 = ~n513 & ~n525;
  assign n527 = n513 & n525;
  assign n528 = pi07 & ~pi32;
  assign n529 = pi08 & pi32;
  assign n530 = pi33 & ~n529;
  assign n531 = ~n528 & n530;
  assign n532 = ~pi33 & n529;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~n527 & ~n533;
  assign n535 = ~n526 & n534;
  assign n536 = ~n526 & ~n527;
  assign n537 = n533 & ~n536;
  assign n538 = ~n535 & ~n537;
  assign n539 = ~n501 & n538;
  assign n540 = ~n498 & n539;
  assign n541 = ~n498 & ~n501;
  assign n542 = ~n538 & ~n541;
  assign n543 = ~n540 & ~n542;
  assign n544 = ~n478 & n543;
  assign n545 = n478 & ~n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = n391 & n450;
  assign n548 = ~n385 & ~n547;
  assign n549 = ~n546 & n548;
  assign n550 = n546 & ~n548;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~n477 & n551;
  assign n553 = n477 & ~n551;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~n467 & ~n554;
  assign n556 = ~n474 & n555;
  assign n557 = ~n467 & ~n474;
  assign n558 = n554 & ~n557;
  assign po08 = ~n556 & ~n558;
  assign n560 = ~n544 & ~n550;
  assign n561 = ~n498 & ~n540;
  assign n562 = ~n488 & n492;
  assign n563 = ~n486 & n562;
  assign n564 = pi41 & ~n492;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~n561 & ~n565;
  assign n567 = ~n498 & n565;
  assign n568 = ~n540 & n567;
  assign n569 = ~n566 & ~n568;
  assign n570 = pi40 & ~pi41;
  assign n571 = ~pi40 & pi41;
  assign n572 = ~n570 & ~n571;
  assign n573 = pi00 & ~n489;
  assign n574 = ~n490 & n573;
  assign n575 = ~n572 & n574;
  assign n576 = pi01 & ~n491;
  assign n577 = ~n575 & ~n576;
  assign n578 = pi41 & ~n577;
  assign n579 = pi02 & ~n304;
  assign n580 = ~n305 & n579;
  assign n581 = ~n394 & n580;
  assign n582 = pi03 & ~n306;
  assign n583 = ~n581 & ~n582;
  assign n584 = pi39 & ~n583;
  assign n585 = ~pi39 & ~n582;
  assign n586 = ~n581 & n585;
  assign n587 = ~pi41 & ~n576;
  assign n588 = ~n575 & n587;
  assign n589 = ~n586 & ~n588;
  assign n590 = ~n584 & n589;
  assign n591 = ~n578 & n590;
  assign n592 = ~n584 & ~n586;
  assign n593 = ~n578 & ~n588;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~n591 & ~n594;
  assign n596 = ~n526 & ~n533;
  assign n597 = ~n527 & ~n596;
  assign n598 = ~n595 & n597;
  assign n599 = n595 & ~n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = pi05 & ~n195;
  assign n602 = pi04 & pi35;
  assign n603 = n341 & n602;
  assign n604 = pi04 & ~pi35;
  assign n605 = n259 & n604;
  assign n606 = ~n603 & ~n605;
  assign n607 = ~n601 & n606;
  assign n608 = pi37 & ~n607;
  assign n609 = ~pi37 & ~n603;
  assign n610 = ~n605 & n609;
  assign n611 = ~n601 & n610;
  assign n612 = ~n608 & ~n611;
  assign n613 = pi07 & ~n143;
  assign n614 = pi06 & pi33;
  assign n615 = n154 & n614;
  assign n616 = pi06 & ~pi33;
  assign n617 = n155 & n616;
  assign n618 = ~n615 & ~n617;
  assign n619 = ~n613 & n618;
  assign n620 = pi35 & ~n619;
  assign n621 = ~pi35 & ~n615;
  assign n622 = ~n617 & n621;
  assign n623 = ~n613 & n622;
  assign n624 = ~n620 & ~n623;
  assign n625 = ~n612 & n624;
  assign n626 = n612 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = pi08 & ~pi32;
  assign n629 = pi09 & pi32;
  assign n630 = pi33 & ~n629;
  assign n631 = ~n628 & n630;
  assign n632 = ~pi33 & n629;
  assign n633 = ~n631 & ~n632;
  assign n634 = ~n627 & ~n633;
  assign n635 = ~n625 & n633;
  assign n636 = ~n626 & n635;
  assign n637 = ~n634 & ~n636;
  assign n638 = ~n600 & n637;
  assign n639 = n600 & ~n637;
  assign n640 = ~n638 & ~n639;
  assign n641 = ~n569 & n640;
  assign n642 = ~n568 & ~n640;
  assign n643 = ~n566 & n642;
  assign n644 = ~n641 & ~n643;
  assign n645 = ~n560 & n644;
  assign n646 = n475 & ~n549;
  assign n647 = ~n550 & n646;
  assign n648 = ~n645 & n647;
  assign n649 = n560 & ~n644;
  assign n650 = n476 & n551;
  assign n651 = ~n649 & ~n650;
  assign n652 = n648 & n651;
  assign n653 = ~n645 & ~n649;
  assign n654 = ~n647 & ~n650;
  assign n655 = ~n653 & n654;
  assign n656 = ~n652 & ~n655;
  assign n657 = ~n645 & n650;
  assign n658 = ~n647 & ~n649;
  assign n659 = n657 & n658;
  assign n660 = n476 & ~n550;
  assign n661 = n646 & n660;
  assign n662 = ~n653 & n661;
  assign n663 = ~n659 & ~n662;
  assign n664 = n656 & n663;
  assign n665 = n558 & ~n664;
  assign n666 = ~n558 & n664;
  assign po09 = n665 | n666;
  assign n668 = n550 & n644;
  assign n669 = ~n566 & ~n642;
  assign n670 = ~n599 & ~n637;
  assign n671 = ~n598 & ~n670;
  assign n672 = pi43 & ~n586;
  assign n673 = ~n584 & n672;
  assign n674 = n593 & n673;
  assign n675 = ~pi43 & ~n591;
  assign n676 = ~n674 & ~n675;
  assign n677 = ~n671 & ~n676;
  assign n678 = ~n598 & n676;
  assign n679 = ~n670 & n678;
  assign n680 = ~n677 & ~n679;
  assign n681 = n612 & n624;
  assign n682 = ~n634 & ~n681;
  assign n683 = pi41 & ~pi42;
  assign n684 = ~pi41 & pi42;
  assign n685 = ~n683 & ~n684;
  assign n686 = pi00 & ~n685;
  assign n687 = pi43 & ~n686;
  assign n688 = pi00 & ~pi43;
  assign n689 = ~n685 & n688;
  assign n690 = ~n687 & ~n689;
  assign n691 = pi02 & ~n491;
  assign n692 = pi01 & pi39;
  assign n693 = n570 & n692;
  assign n694 = pi01 & ~pi39;
  assign n695 = n571 & n694;
  assign n696 = ~n693 & ~n695;
  assign n697 = ~n691 & n696;
  assign n698 = pi41 & ~n697;
  assign n699 = ~pi41 & ~n693;
  assign n700 = ~n695 & n699;
  assign n701 = ~n691 & n700;
  assign n702 = ~n698 & ~n701;
  assign n703 = ~n690 & n702;
  assign n704 = n690 & ~n702;
  assign n705 = ~n703 & ~n704;
  assign n706 = pi03 & ~n304;
  assign n707 = ~n305 & n706;
  assign n708 = ~n394 & n707;
  assign n709 = pi04 & ~n306;
  assign n710 = ~n708 & ~n709;
  assign n711 = pi39 & ~n710;
  assign n712 = ~pi39 & ~n709;
  assign n713 = ~n708 & n712;
  assign n714 = ~n711 & ~n713;
  assign n715 = ~n705 & n714;
  assign n716 = n705 & ~n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = ~n682 & ~n717;
  assign n719 = n682 & n717;
  assign n720 = pi07 & ~n141;
  assign n721 = ~n142 & n720;
  assign n722 = ~n156 & n721;
  assign n723 = pi08 & ~n143;
  assign n724 = ~n722 & ~n723;
  assign n725 = pi35 & ~n724;
  assign n726 = ~pi35 & ~n723;
  assign n727 = ~n722 & n726;
  assign n728 = ~n725 & ~n727;
  assign n729 = ~n259 & ~n341;
  assign n730 = pi05 & ~n193;
  assign n731 = ~n194 & n730;
  assign n732 = ~n729 & n731;
  assign n733 = pi06 & ~n195;
  assign n734 = ~n732 & ~n733;
  assign n735 = pi37 & ~n734;
  assign n736 = ~pi37 & ~n733;
  assign n737 = ~n732 & n736;
  assign n738 = ~n735 & ~n737;
  assign n739 = ~n728 & ~n738;
  assign n740 = ~n727 & ~n737;
  assign n741 = ~n725 & n740;
  assign n742 = ~n735 & n741;
  assign n743 = pi09 & ~pi32;
  assign n744 = pi10 & pi32;
  assign n745 = pi33 & ~n744;
  assign n746 = ~n743 & n745;
  assign n747 = ~pi33 & n744;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n742 & ~n748;
  assign n750 = ~n739 & n749;
  assign n751 = ~n739 & ~n742;
  assign n752 = n748 & ~n751;
  assign n753 = ~n750 & ~n752;
  assign n754 = ~n719 & n753;
  assign n755 = ~n718 & n754;
  assign n756 = ~n718 & ~n719;
  assign n757 = ~n753 & ~n756;
  assign n758 = ~n755 & ~n757;
  assign n759 = ~n680 & ~n758;
  assign n760 = n680 & n758;
  assign n761 = ~n759 & ~n760;
  assign n762 = n669 & ~n761;
  assign n763 = ~n669 & ~n759;
  assign n764 = ~n760 & n763;
  assign n765 = n544 & ~n643;
  assign n766 = ~n641 & n765;
  assign n767 = ~n764 & n766;
  assign n768 = ~n762 & n767;
  assign n769 = ~n762 & ~n764;
  assign n770 = ~n766 & ~n769;
  assign n771 = ~n768 & ~n770;
  assign n772 = ~n668 & ~n771;
  assign n773 = n648 & ~n649;
  assign n774 = n668 & ~n768;
  assign n775 = ~n770 & n774;
  assign n776 = n773 & ~n775;
  assign n777 = ~n772 & n776;
  assign n778 = ~n772 & ~n775;
  assign n779 = ~n773 & ~n778;
  assign n780 = ~n777 & ~n779;
  assign n781 = ~n655 & ~n659;
  assign n782 = ~n662 & n781;
  assign n783 = n554 & ~n652;
  assign n784 = ~n557 & n783;
  assign n785 = n782 & n784;
  assign n786 = ~n647 & ~n653;
  assign n787 = n650 & ~n786;
  assign n788 = ~n773 & n787;
  assign n789 = ~n785 & ~n788;
  assign n790 = ~n780 & n789;
  assign n791 = n780 & ~n789;
  assign po10 = ~n790 & ~n791;
  assign n793 = ~n777 & ~n791;
  assign n794 = ~n764 & ~n768;
  assign n795 = ~n739 & ~n748;
  assign n796 = ~n742 & ~n795;
  assign n797 = pi01 & ~n685;
  assign n798 = pi41 & pi42;
  assign n799 = n688 & n798;
  assign n800 = pi00 & ~pi41;
  assign n801 = ~pi42 & pi43;
  assign n802 = n800 & n801;
  assign n803 = ~n799 & ~n802;
  assign n804 = ~n797 & n803;
  assign n805 = pi43 & ~n804;
  assign n806 = ~pi43 & ~n799;
  assign n807 = ~n802 & n806;
  assign n808 = ~n797 & n807;
  assign n809 = ~n805 & ~n808;
  assign n810 = pi03 & ~n491;
  assign n811 = pi02 & pi39;
  assign n812 = n570 & n811;
  assign n813 = pi02 & ~pi39;
  assign n814 = n571 & n813;
  assign n815 = ~n812 & ~n814;
  assign n816 = ~n810 & n815;
  assign n817 = pi41 & ~n816;
  assign n818 = ~pi41 & ~n812;
  assign n819 = ~n814 & n818;
  assign n820 = ~n810 & n819;
  assign n821 = ~n817 & ~n820;
  assign n822 = ~n809 & n821;
  assign n823 = n809 & ~n821;
  assign n824 = ~n822 & ~n823;
  assign n825 = pi04 & ~n304;
  assign n826 = ~n305 & n825;
  assign n827 = ~n394 & n826;
  assign n828 = pi05 & ~n306;
  assign n829 = ~n827 & ~n828;
  assign n830 = pi39 & ~n829;
  assign n831 = ~pi39 & ~n828;
  assign n832 = ~n827 & n831;
  assign n833 = ~n830 & ~n832;
  assign n834 = ~n824 & n833;
  assign n835 = n824 & ~n833;
  assign n836 = ~n834 & ~n835;
  assign n837 = ~n796 & n836;
  assign n838 = n796 & ~n836;
  assign n839 = ~n837 & ~n838;
  assign n840 = pi07 & ~n195;
  assign n841 = pi06 & pi35;
  assign n842 = n341 & n841;
  assign n843 = pi06 & ~pi35;
  assign n844 = n259 & n843;
  assign n845 = ~n842 & ~n844;
  assign n846 = ~n840 & n845;
  assign n847 = pi37 & ~n846;
  assign n848 = ~pi37 & ~n842;
  assign n849 = ~n844 & n848;
  assign n850 = ~n840 & n849;
  assign n851 = ~n847 & ~n850;
  assign n852 = pi09 & ~n143;
  assign n853 = pi08 & pi33;
  assign n854 = n154 & n853;
  assign n855 = pi08 & ~pi33;
  assign n856 = n155 & n855;
  assign n857 = ~n854 & ~n856;
  assign n858 = ~n852 & n857;
  assign n859 = pi35 & ~n858;
  assign n860 = ~pi35 & ~n854;
  assign n861 = ~n856 & n860;
  assign n862 = ~n852 & n861;
  assign n863 = ~n859 & ~n862;
  assign n864 = ~n851 & n863;
  assign n865 = n851 & ~n863;
  assign n866 = ~n864 & ~n865;
  assign n867 = pi10 & ~pi32;
  assign n868 = pi11 & pi32;
  assign n869 = pi33 & ~n868;
  assign n870 = ~n867 & n869;
  assign n871 = ~pi33 & n868;
  assign n872 = ~n870 & ~n871;
  assign n873 = ~n866 & ~n872;
  assign n874 = ~n864 & n872;
  assign n875 = ~n865 & n874;
  assign n876 = ~n873 & ~n875;
  assign n877 = ~n839 & n876;
  assign n878 = ~n837 & ~n876;
  assign n879 = ~n838 & n878;
  assign n880 = ~n877 & ~n879;
  assign n881 = ~n704 & ~n716;
  assign n882 = n753 & ~n881;
  assign n883 = n756 & n882;
  assign n884 = n718 & ~n881;
  assign n885 = ~n883 & ~n884;
  assign n886 = ~n718 & n881;
  assign n887 = ~n753 & n886;
  assign n888 = ~n756 & n886;
  assign n889 = ~n887 & ~n888;
  assign n890 = n885 & n889;
  assign n891 = ~n880 & n890;
  assign n892 = n880 & ~n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n674 & ~n679;
  assign n895 = ~n760 & n894;
  assign n896 = n674 & ~n679;
  assign n897 = ~n677 & n896;
  assign n898 = n758 & n897;
  assign n899 = ~n895 & ~n898;
  assign n900 = ~n893 & n899;
  assign n901 = n893 & ~n899;
  assign n902 = ~n900 & ~n901;
  assign n903 = n794 & ~n902;
  assign n904 = ~n794 & n902;
  assign n905 = n775 & ~n904;
  assign n906 = ~n903 & n905;
  assign n907 = ~n903 & ~n904;
  assign n908 = ~n775 & ~n907;
  assign n909 = ~n906 & ~n908;
  assign n910 = ~n793 & n909;
  assign n911 = ~n777 & ~n909;
  assign n912 = ~n791 & n911;
  assign po11 = ~n910 & ~n912;
  assign n914 = ~n906 & ~n910;
  assign n915 = ~n880 & ~n890;
  assign n916 = ~n718 & ~n755;
  assign n917 = n881 & ~n916;
  assign n918 = ~n915 & ~n917;
  assign n919 = n851 & n863;
  assign n920 = ~n873 & ~n919;
  assign n921 = pi02 & ~n685;
  assign n922 = pi01 & pi41;
  assign n923 = pi42 & ~pi43;
  assign n924 = n922 & n923;
  assign n925 = pi01 & ~pi41;
  assign n926 = n801 & n925;
  assign n927 = ~n924 & ~n926;
  assign n928 = ~n921 & n927;
  assign n929 = pi43 & ~n928;
  assign n930 = ~pi43 & ~n924;
  assign n931 = ~n926 & n930;
  assign n932 = ~n921 & n931;
  assign n933 = ~n929 & ~n932;
  assign n934 = pi04 & ~n491;
  assign n935 = pi03 & pi39;
  assign n936 = n570 & n935;
  assign n937 = pi03 & ~pi39;
  assign n938 = n571 & n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~n934 & n939;
  assign n941 = pi41 & ~n940;
  assign n942 = ~pi41 & ~n936;
  assign n943 = ~n938 & n942;
  assign n944 = ~n934 & n943;
  assign n945 = ~n941 & ~n944;
  assign n946 = ~n933 & n945;
  assign n947 = n933 & ~n945;
  assign n948 = ~n946 & ~n947;
  assign n949 = pi05 & ~n304;
  assign n950 = ~n305 & n949;
  assign n951 = ~n394 & n950;
  assign n952 = pi06 & ~n306;
  assign n953 = ~n951 & ~n952;
  assign n954 = pi39 & ~n953;
  assign n955 = ~pi39 & ~n952;
  assign n956 = ~n951 & n955;
  assign n957 = ~n954 & ~n956;
  assign n958 = ~n948 & n957;
  assign n959 = n948 & ~n957;
  assign n960 = ~n958 & ~n959;
  assign n961 = ~n920 & n960;
  assign n962 = n920 & ~n960;
  assign n963 = ~n961 & ~n962;
  assign n964 = pi08 & ~n195;
  assign n965 = pi07 & pi35;
  assign n966 = n341 & n965;
  assign n967 = pi07 & ~pi35;
  assign n968 = n259 & n967;
  assign n969 = ~n966 & ~n968;
  assign n970 = ~n964 & n969;
  assign n971 = pi37 & ~n970;
  assign n972 = ~pi37 & ~n966;
  assign n973 = ~n968 & n972;
  assign n974 = ~n964 & n973;
  assign n975 = ~n971 & ~n974;
  assign n976 = pi10 & ~n143;
  assign n977 = pi09 & pi33;
  assign n978 = n154 & n977;
  assign n979 = pi09 & ~pi33;
  assign n980 = n155 & n979;
  assign n981 = ~n978 & ~n980;
  assign n982 = ~n976 & n981;
  assign n983 = pi35 & ~n982;
  assign n984 = ~pi35 & ~n978;
  assign n985 = ~n980 & n984;
  assign n986 = ~n976 & n985;
  assign n987 = ~n983 & ~n986;
  assign n988 = n975 & ~n987;
  assign n989 = ~n975 & n987;
  assign n990 = pi11 & ~pi32;
  assign n991 = pi12 & pi32;
  assign n992 = pi33 & ~n991;
  assign n993 = ~n990 & n992;
  assign n994 = ~pi33 & n991;
  assign n995 = ~n993 & ~n994;
  assign n996 = ~n989 & n995;
  assign n997 = ~n988 & n996;
  assign n998 = ~n988 & ~n989;
  assign n999 = ~n995 & ~n998;
  assign n1000 = ~n997 & ~n999;
  assign n1001 = ~n963 & n1000;
  assign n1002 = ~n961 & ~n1000;
  assign n1003 = ~n962 & n1002;
  assign n1004 = ~n1001 & ~n1003;
  assign n1005 = n809 & n821;
  assign n1006 = pi43 & ~pi44;
  assign n1007 = ~pi43 & pi44;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = pi00 & ~n1008;
  assign n1010 = ~n1005 & ~n1009;
  assign n1011 = ~n834 & n1010;
  assign n1012 = ~n834 & ~n1005;
  assign n1013 = n1009 & ~n1012;
  assign n1014 = ~n1011 & ~n1013;
  assign n1015 = ~n838 & n876;
  assign n1016 = ~n837 & ~n1015;
  assign n1017 = ~n1014 & n1016;
  assign n1018 = n1014 & ~n1016;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = ~n1004 & ~n1019;
  assign n1021 = n1004 & ~n1017;
  assign n1022 = ~n1018 & n1021;
  assign n1023 = ~n1020 & ~n1022;
  assign n1024 = ~n918 & ~n1023;
  assign n1025 = n918 & n1023;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n898 & ~n900;
  assign n1028 = ~n1026 & n1027;
  assign n1029 = n1026 & ~n1027;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = ~n762 & n764;
  assign n1032 = n767 & n1031;
  assign n1033 = n902 & n1032;
  assign n1034 = ~n1030 & n1033;
  assign n1035 = n768 & n902;
  assign n1036 = ~n1028 & n1035;
  assign n1037 = n764 & ~n900;
  assign n1038 = ~n901 & n1037;
  assign n1039 = ~n1029 & ~n1038;
  assign n1040 = n1036 & n1039;
  assign n1041 = ~n1034 & ~n1040;
  assign n1042 = ~n1035 & ~n1038;
  assign n1043 = ~n1030 & n1042;
  assign n1044 = ~n1028 & n1038;
  assign n1045 = ~n1029 & ~n1035;
  assign n1046 = n1044 & n1045;
  assign n1047 = ~n1043 & ~n1046;
  assign n1048 = n1041 & n1047;
  assign n1049 = ~n914 & n1048;
  assign n1050 = ~n906 & ~n1048;
  assign n1051 = ~n910 & n1050;
  assign po12 = ~n1049 & ~n1051;
  assign n1053 = ~n906 & n1041;
  assign n1054 = n1047 & ~n1053;
  assign n1055 = n909 & n1048;
  assign n1056 = ~n793 & n1055;
  assign n1057 = ~n1054 & ~n1056;
  assign n1058 = ~n1024 & ~n1029;
  assign n1059 = ~n1004 & ~n1017;
  assign n1060 = ~n1018 & n1059;
  assign n1061 = ~n1013 & ~n1018;
  assign n1062 = ~n1060 & n1061;
  assign n1063 = ~n962 & n1000;
  assign n1064 = ~n961 & ~n1063;
  assign n1065 = n933 & n945;
  assign n1066 = pi44 & ~pi45;
  assign n1067 = ~pi44 & pi45;
  assign n1068 = ~n1066 & ~n1067;
  assign n1069 = pi00 & ~n1006;
  assign n1070 = ~n1007 & n1069;
  assign n1071 = ~n1068 & n1070;
  assign n1072 = pi01 & ~n1008;
  assign n1073 = pi00 & pi45;
  assign n1074 = ~n1008 & n1073;
  assign n1075 = ~n1072 & ~n1074;
  assign n1076 = ~n1071 & n1075;
  assign n1077 = ~n1071 & ~n1072;
  assign n1078 = n1074 & ~n1077;
  assign n1079 = ~n1076 & ~n1078;
  assign n1080 = ~n1065 & ~n1079;
  assign n1081 = ~n958 & n1080;
  assign n1082 = ~n958 & ~n1065;
  assign n1083 = n1079 & ~n1082;
  assign n1084 = ~n1081 & ~n1083;
  assign n1085 = ~n1064 & n1084;
  assign n1086 = n1064 & ~n1084;
  assign n1087 = ~n1085 & ~n1086;
  assign n1088 = pi03 & ~n685;
  assign n1089 = pi02 & pi41;
  assign n1090 = n923 & n1089;
  assign n1091 = pi02 & ~pi41;
  assign n1092 = n801 & n1091;
  assign n1093 = ~n1090 & ~n1092;
  assign n1094 = ~n1088 & n1093;
  assign n1095 = pi43 & ~n1094;
  assign n1096 = ~pi43 & ~n1090;
  assign n1097 = ~n1092 & n1096;
  assign n1098 = ~n1088 & n1097;
  assign n1099 = ~n1095 & ~n1098;
  assign n1100 = pi05 & ~n491;
  assign n1101 = pi04 & pi39;
  assign n1102 = n570 & n1101;
  assign n1103 = pi04 & ~pi39;
  assign n1104 = n571 & n1103;
  assign n1105 = ~n1102 & ~n1104;
  assign n1106 = ~n1100 & n1105;
  assign n1107 = pi41 & ~n1106;
  assign n1108 = ~pi41 & ~n1102;
  assign n1109 = ~n1104 & n1108;
  assign n1110 = ~n1100 & n1109;
  assign n1111 = ~n1107 & ~n1110;
  assign n1112 = ~n1099 & n1111;
  assign n1113 = n1099 & ~n1111;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = pi06 & ~n304;
  assign n1116 = ~n305 & n1115;
  assign n1117 = ~n394 & n1116;
  assign n1118 = pi07 & ~n306;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = pi39 & ~n1119;
  assign n1121 = ~pi39 & ~n1118;
  assign n1122 = ~n1117 & n1121;
  assign n1123 = ~n1120 & ~n1122;
  assign n1124 = ~n1114 & n1123;
  assign n1125 = n1114 & ~n1123;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = n975 & n987;
  assign n1128 = ~n999 & ~n1127;
  assign n1129 = n1126 & ~n1128;
  assign n1130 = ~n1126 & n1128;
  assign n1131 = pi08 & ~n193;
  assign n1132 = ~n194 & n1131;
  assign n1133 = ~n729 & n1132;
  assign n1134 = pi09 & ~n195;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = pi37 & ~n1135;
  assign n1137 = ~pi37 & ~n1134;
  assign n1138 = ~n1133 & n1137;
  assign n1139 = ~n1136 & ~n1138;
  assign n1140 = pi10 & ~n141;
  assign n1141 = ~n142 & n1140;
  assign n1142 = ~n156 & n1141;
  assign n1143 = pi11 & ~n143;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = pi35 & ~n1144;
  assign n1146 = ~pi35 & ~n1143;
  assign n1147 = ~n1142 & n1146;
  assign n1148 = ~n1145 & ~n1147;
  assign n1149 = ~n1139 & n1148;
  assign n1150 = n1139 & ~n1148;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = pi12 & ~pi32;
  assign n1153 = pi13 & pi32;
  assign n1154 = pi33 & ~n1153;
  assign n1155 = ~n1152 & n1154;
  assign n1156 = ~pi33 & n1153;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1151 & ~n1157;
  assign n1159 = ~n1149 & n1157;
  assign n1160 = ~n1150 & n1159;
  assign n1161 = ~n1158 & ~n1160;
  assign n1162 = ~n1130 & n1161;
  assign n1163 = ~n1129 & n1162;
  assign n1164 = ~n1129 & ~n1130;
  assign n1165 = ~n1161 & ~n1164;
  assign n1166 = ~n1163 & ~n1165;
  assign n1167 = ~n1087 & n1166;
  assign n1168 = n1087 & ~n1166;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~n1004 & n1013;
  assign n1171 = n1019 & n1170;
  assign n1172 = ~n1169 & ~n1171;
  assign n1173 = ~n1062 & n1172;
  assign n1174 = ~n1062 & ~n1171;
  assign n1175 = n1169 & ~n1174;
  assign n1176 = ~n1173 & ~n1175;
  assign n1177 = n1058 & ~n1176;
  assign n1178 = ~n1058 & n1176;
  assign n1179 = ~n1029 & n1044;
  assign n1180 = ~n1178 & n1179;
  assign n1181 = ~n1177 & n1180;
  assign n1182 = ~n1177 & ~n1178;
  assign n1183 = ~n1179 & ~n1182;
  assign n1184 = ~n1181 & ~n1183;
  assign n1185 = ~n1057 & n1184;
  assign n1186 = ~n1054 & ~n1184;
  assign n1187 = ~n1056 & n1186;
  assign po13 = ~n1185 & ~n1187;
  assign n1189 = n791 & n1184;
  assign n1190 = n1055 & n1189;
  assign n1191 = n1054 & ~n1183;
  assign n1192 = n777 & ~n906;
  assign n1193 = ~n908 & n1192;
  assign n1194 = n1048 & ~n1183;
  assign n1195 = n1193 & n1194;
  assign n1196 = ~n1181 & ~n1195;
  assign n1197 = ~n1191 & n1196;
  assign n1198 = ~n1190 & n1197;
  assign n1199 = n1024 & ~n1173;
  assign n1200 = ~n1175 & n1199;
  assign n1201 = n1099 & n1111;
  assign n1202 = ~n1124 & ~n1201;
  assign n1203 = pi01 & ~n1006;
  assign n1204 = ~n1007 & n1203;
  assign n1205 = ~n1068 & n1204;
  assign n1206 = pi02 & ~n1008;
  assign n1207 = ~n1205 & ~n1206;
  assign n1208 = pi45 & ~n1207;
  assign n1209 = ~pi45 & ~n1206;
  assign n1210 = ~n1205 & n1209;
  assign n1211 = ~n1208 & ~n1210;
  assign n1212 = pi45 & ~pi46;
  assign n1213 = ~pi45 & pi46;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = pi00 & ~n1214;
  assign n1216 = ~n1211 & n1215;
  assign n1217 = ~n1210 & ~n1215;
  assign n1218 = ~n1208 & n1217;
  assign n1219 = ~n1216 & ~n1218;
  assign n1220 = ~n1202 & ~n1219;
  assign n1221 = ~n1201 & ~n1218;
  assign n1222 = ~n1216 & n1221;
  assign n1223 = ~n1124 & n1222;
  assign n1224 = ~n1220 & ~n1223;
  assign n1225 = ~n1129 & ~n1163;
  assign n1226 = n1224 & ~n1225;
  assign n1227 = ~n1138 & ~n1147;
  assign n1228 = ~n1145 & n1227;
  assign n1229 = ~n1136 & n1228;
  assign n1230 = ~n1158 & ~n1229;
  assign n1231 = ~n801 & ~n923;
  assign n1232 = pi03 & ~n683;
  assign n1233 = ~n684 & n1232;
  assign n1234 = ~n1231 & n1233;
  assign n1235 = pi04 & ~n685;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = pi43 & ~n1236;
  assign n1238 = ~pi43 & ~n1235;
  assign n1239 = ~n1234 & n1238;
  assign n1240 = ~n1237 & ~n1239;
  assign n1241 = pi05 & ~n489;
  assign n1242 = ~n490 & n1241;
  assign n1243 = ~n572 & n1242;
  assign n1244 = pi06 & ~n491;
  assign n1245 = ~n1243 & ~n1244;
  assign n1246 = pi41 & ~n1245;
  assign n1247 = ~pi41 & ~n1244;
  assign n1248 = ~n1243 & n1247;
  assign n1249 = ~n1246 & ~n1248;
  assign n1250 = ~n1240 & n1249;
  assign n1251 = n1240 & ~n1249;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = pi07 & ~n304;
  assign n1254 = ~n305 & n1253;
  assign n1255 = ~n394 & n1254;
  assign n1256 = pi08 & ~n306;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = pi39 & ~n1257;
  assign n1259 = ~pi39 & ~n1256;
  assign n1260 = ~n1255 & n1259;
  assign n1261 = ~n1258 & ~n1260;
  assign n1262 = ~n1252 & n1261;
  assign n1263 = ~n1250 & ~n1261;
  assign n1264 = ~n1251 & n1263;
  assign n1265 = ~n1262 & ~n1264;
  assign n1266 = n1230 & ~n1265;
  assign n1267 = ~n1230 & n1265;
  assign n1268 = pi09 & ~n193;
  assign n1269 = ~n194 & n1268;
  assign n1270 = ~n729 & n1269;
  assign n1271 = pi10 & ~n195;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = pi37 & ~n1272;
  assign n1274 = ~pi37 & ~n1271;
  assign n1275 = ~n1270 & n1274;
  assign n1276 = ~n1273 & ~n1275;
  assign n1277 = pi11 & ~n141;
  assign n1278 = ~n142 & n1277;
  assign n1279 = ~n156 & n1278;
  assign n1280 = pi12 & ~n143;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = pi35 & ~n1281;
  assign n1283 = ~pi35 & ~n1280;
  assign n1284 = ~n1279 & n1283;
  assign n1285 = ~n1282 & ~n1284;
  assign n1286 = ~n1276 & n1285;
  assign n1287 = n1276 & ~n1285;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = pi13 & ~pi32;
  assign n1290 = pi14 & pi32;
  assign n1291 = pi33 & ~n1290;
  assign n1292 = ~n1289 & n1291;
  assign n1293 = ~pi33 & n1290;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n1288 & ~n1294;
  assign n1296 = ~n1286 & n1294;
  assign n1297 = ~n1287 & n1296;
  assign n1298 = ~n1295 & ~n1297;
  assign n1299 = ~n1267 & ~n1298;
  assign n1300 = ~n1266 & n1299;
  assign n1301 = ~n1129 & ~n1224;
  assign n1302 = ~n1163 & n1301;
  assign n1303 = ~n1266 & ~n1267;
  assign n1304 = n1298 & ~n1303;
  assign n1305 = ~n1302 & ~n1304;
  assign n1306 = ~n1300 & n1305;
  assign n1307 = ~n1226 & n1306;
  assign n1308 = ~n1226 & ~n1302;
  assign n1309 = ~n1300 & ~n1304;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = ~n1307 & ~n1310;
  assign n1312 = ~n1086 & n1166;
  assign n1313 = pi45 & ~n1009;
  assign n1314 = n1077 & n1313;
  assign n1315 = ~n1083 & ~n1314;
  assign n1316 = ~n1085 & ~n1315;
  assign n1317 = ~n1312 & n1316;
  assign n1318 = ~n1085 & ~n1312;
  assign n1319 = n1315 & ~n1318;
  assign n1320 = ~n1317 & ~n1319;
  assign n1321 = ~n1311 & ~n1320;
  assign n1322 = n1311 & n1320;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = ~n1171 & ~n1173;
  assign n1325 = ~n1323 & n1324;
  assign n1326 = n1323 & ~n1324;
  assign n1327 = ~n1325 & ~n1326;
  assign n1328 = ~n1200 & ~n1327;
  assign n1329 = n1200 & ~n1325;
  assign n1330 = ~n1326 & n1329;
  assign n1331 = n1029 & n1176;
  assign n1332 = ~n1330 & n1331;
  assign n1333 = ~n1328 & n1332;
  assign n1334 = ~n1328 & ~n1330;
  assign n1335 = ~n1331 & ~n1334;
  assign n1336 = ~n1333 & ~n1335;
  assign n1337 = ~n1198 & n1336;
  assign n1338 = ~n1191 & ~n1336;
  assign n1339 = n1196 & n1338;
  assign n1340 = ~n1190 & n1339;
  assign po14 = ~n1337 & ~n1340;
  assign n1342 = ~n1326 & ~n1329;
  assign n1343 = ~n1275 & ~n1284;
  assign n1344 = ~n1282 & n1343;
  assign n1345 = ~n1273 & n1344;
  assign n1346 = ~n1295 & ~n1345;
  assign n1347 = pi04 & ~n683;
  assign n1348 = ~n684 & n1347;
  assign n1349 = ~n1231 & n1348;
  assign n1350 = pi05 & ~n685;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = pi43 & ~n1351;
  assign n1353 = ~pi43 & ~n1350;
  assign n1354 = ~n1349 & n1353;
  assign n1355 = ~n1352 & ~n1354;
  assign n1356 = pi06 & ~n489;
  assign n1357 = ~n490 & n1356;
  assign n1358 = ~n572 & n1357;
  assign n1359 = pi07 & ~n491;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = pi41 & ~n1360;
  assign n1362 = ~pi41 & ~n1359;
  assign n1363 = ~n1358 & n1362;
  assign n1364 = ~n1361 & ~n1363;
  assign n1365 = ~n1355 & n1364;
  assign n1366 = n1355 & ~n1364;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = pi08 & ~n304;
  assign n1369 = ~n305 & n1368;
  assign n1370 = ~n394 & n1369;
  assign n1371 = pi09 & ~n306;
  assign n1372 = ~n1370 & ~n1371;
  assign n1373 = pi39 & ~n1372;
  assign n1374 = ~pi39 & ~n1371;
  assign n1375 = ~n1370 & n1374;
  assign n1376 = ~n1373 & ~n1375;
  assign n1377 = ~n1367 & n1376;
  assign n1378 = ~n1365 & ~n1376;
  assign n1379 = ~n1366 & n1378;
  assign n1380 = ~n1377 & ~n1379;
  assign n1381 = ~n1346 & n1380;
  assign n1382 = n1346 & ~n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = pi10 & ~n193;
  assign n1385 = ~n194 & n1384;
  assign n1386 = ~n729 & n1385;
  assign n1387 = pi11 & ~n195;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = pi37 & ~n1388;
  assign n1390 = ~pi37 & ~n1387;
  assign n1391 = ~n1386 & n1390;
  assign n1392 = ~n1389 & ~n1391;
  assign n1393 = pi12 & ~n141;
  assign n1394 = ~n142 & n1393;
  assign n1395 = ~n156 & n1394;
  assign n1396 = pi13 & ~n143;
  assign n1397 = ~n1395 & ~n1396;
  assign n1398 = pi35 & ~n1397;
  assign n1399 = ~pi35 & ~n1396;
  assign n1400 = ~n1395 & n1399;
  assign n1401 = ~n1398 & ~n1400;
  assign n1402 = ~n1392 & n1401;
  assign n1403 = n1392 & ~n1401;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = pi14 & ~pi32;
  assign n1406 = pi15 & pi32;
  assign n1407 = pi33 & ~n1406;
  assign n1408 = ~n1405 & n1407;
  assign n1409 = ~pi33 & n1406;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1404 & ~n1410;
  assign n1412 = ~n1402 & n1410;
  assign n1413 = ~n1403 & n1412;
  assign n1414 = ~n1411 & ~n1413;
  assign n1415 = ~n1383 & n1414;
  assign n1416 = ~n1381 & ~n1414;
  assign n1417 = ~n1382 & n1416;
  assign n1418 = ~n1415 & ~n1417;
  assign n1419 = ~n1239 & ~n1248;
  assign n1420 = ~n1246 & n1419;
  assign n1421 = ~n1237 & n1420;
  assign n1422 = ~n1262 & ~n1421;
  assign n1423 = pi46 & ~pi47;
  assign n1424 = ~pi46 & pi47;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = pi00 & ~n1212;
  assign n1427 = ~n1213 & n1426;
  assign n1428 = ~n1425 & n1427;
  assign n1429 = pi01 & ~n1214;
  assign n1430 = ~n1428 & ~n1429;
  assign n1431 = pi47 & ~n1430;
  assign n1432 = pi02 & ~n1006;
  assign n1433 = ~n1007 & n1432;
  assign n1434 = ~n1068 & n1433;
  assign n1435 = pi03 & ~n1008;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = pi45 & ~n1436;
  assign n1438 = ~pi45 & ~n1435;
  assign n1439 = ~n1434 & n1438;
  assign n1440 = ~pi47 & ~n1429;
  assign n1441 = ~n1428 & n1440;
  assign n1442 = ~n1439 & ~n1441;
  assign n1443 = ~n1437 & n1442;
  assign n1444 = ~n1431 & n1443;
  assign n1445 = ~n1437 & ~n1439;
  assign n1446 = ~n1431 & ~n1441;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1444 & ~n1447;
  assign n1449 = pi47 & ~n1215;
  assign n1450 = ~n1210 & n1215;
  assign n1451 = ~n1208 & n1450;
  assign n1452 = ~n1449 & ~n1451;
  assign n1453 = ~n1448 & n1452;
  assign n1454 = n1448 & ~n1452;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~n1422 & n1455;
  assign n1457 = n1422 & ~n1455;
  assign n1458 = ~n1456 & ~n1457;
  assign n1459 = ~n1266 & n1298;
  assign n1460 = ~n1267 & ~n1459;
  assign n1461 = ~n1458 & n1460;
  assign n1462 = n1458 & ~n1460;
  assign n1463 = ~n1461 & ~n1462;
  assign n1464 = ~n1418 & ~n1463;
  assign n1465 = n1418 & ~n1461;
  assign n1466 = ~n1462 & n1465;
  assign n1467 = ~n1464 & ~n1466;
  assign n1468 = ~n1226 & n1309;
  assign n1469 = ~n1302 & ~n1468;
  assign n1470 = n1220 & ~n1469;
  assign n1471 = ~n1220 & ~n1302;
  assign n1472 = ~n1468 & n1471;
  assign n1473 = ~n1470 & ~n1472;
  assign n1474 = ~n1467 & ~n1473;
  assign n1475 = n1467 & n1473;
  assign n1476 = ~n1474 & ~n1475;
  assign n1477 = ~n1315 & ~n1318;
  assign n1478 = ~n1321 & ~n1477;
  assign n1479 = ~n1476 & n1478;
  assign n1480 = n1476 & ~n1478;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = ~n1342 & n1481;
  assign n1483 = n1342 & ~n1481;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = ~n1333 & n1484;
  assign n1486 = ~n1337 & n1485;
  assign n1487 = ~n1333 & ~n1337;
  assign n1488 = ~n1484 & ~n1487;
  assign po15 = n1486 | n1488;
  assign n1490 = ~n1335 & n1485;
  assign n1491 = n1330 & n1481;
  assign n1492 = n1333 & n1484;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = ~n1490 & n1493;
  assign n1495 = ~n1181 & ~n1491;
  assign n1496 = ~n1195 & n1495;
  assign n1497 = ~n1191 & ~n1492;
  assign n1498 = n1496 & n1497;
  assign n1499 = ~n1190 & n1498;
  assign n1500 = ~n1494 & ~n1499;
  assign n1501 = n1326 & ~n1479;
  assign n1502 = ~n1480 & ~n1501;
  assign n1503 = n1220 & ~n1302;
  assign n1504 = ~n1468 & n1503;
  assign n1505 = ~n1474 & ~n1504;
  assign n1506 = n1418 & ~n1462;
  assign n1507 = ~n1461 & ~n1506;
  assign n1508 = ~n1454 & ~n1456;
  assign n1509 = pi49 & ~n1508;
  assign n1510 = ~pi49 & ~n1454;
  assign n1511 = ~n1456 & n1510;
  assign n1512 = ~n1509 & ~n1511;
  assign n1513 = ~n1507 & n1512;
  assign n1514 = ~n1391 & ~n1400;
  assign n1515 = ~n1398 & n1514;
  assign n1516 = ~n1389 & n1515;
  assign n1517 = ~n1411 & ~n1516;
  assign n1518 = pi05 & ~n683;
  assign n1519 = ~n684 & n1518;
  assign n1520 = ~n1231 & n1519;
  assign n1521 = pi06 & ~n685;
  assign n1522 = ~n1520 & ~n1521;
  assign n1523 = pi43 & ~n1522;
  assign n1524 = pi07 & ~n489;
  assign n1525 = ~n490 & n1524;
  assign n1526 = ~n572 & n1525;
  assign n1527 = pi08 & ~n491;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = pi41 & ~n1528;
  assign n1530 = ~pi41 & ~n1527;
  assign n1531 = ~n1526 & n1530;
  assign n1532 = ~pi43 & ~n1521;
  assign n1533 = ~n1520 & n1532;
  assign n1534 = ~n1531 & ~n1533;
  assign n1535 = ~n1529 & n1534;
  assign n1536 = ~n1523 & n1535;
  assign n1537 = ~n1529 & ~n1531;
  assign n1538 = ~n1523 & ~n1533;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = ~n1536 & ~n1539;
  assign n1541 = pi09 & ~n304;
  assign n1542 = ~n305 & n1541;
  assign n1543 = ~n394 & n1542;
  assign n1544 = pi10 & ~n306;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = pi39 & ~n1545;
  assign n1547 = ~pi39 & ~n1544;
  assign n1548 = ~n1543 & n1547;
  assign n1549 = ~n1546 & ~n1548;
  assign n1550 = ~n1540 & n1549;
  assign n1551 = ~n1536 & ~n1549;
  assign n1552 = ~n1539 & n1551;
  assign n1553 = ~n1550 & ~n1552;
  assign n1554 = ~n1517 & ~n1553;
  assign n1555 = n1517 & n1553;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = pi11 & ~n193;
  assign n1558 = ~n194 & n1557;
  assign n1559 = ~n729 & n1558;
  assign n1560 = pi12 & ~n195;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = pi37 & ~n1561;
  assign n1563 = ~pi37 & ~n1560;
  assign n1564 = ~n1559 & n1563;
  assign n1565 = ~n1562 & ~n1564;
  assign n1566 = pi13 & ~n141;
  assign n1567 = ~n142 & n1566;
  assign n1568 = ~n156 & n1567;
  assign n1569 = pi14 & ~n143;
  assign n1570 = ~n1568 & ~n1569;
  assign n1571 = pi35 & ~n1570;
  assign n1572 = ~pi35 & ~n1569;
  assign n1573 = ~n1568 & n1572;
  assign n1574 = ~n1571 & ~n1573;
  assign n1575 = ~n1565 & n1574;
  assign n1576 = n1565 & ~n1574;
  assign n1577 = ~n1575 & ~n1576;
  assign n1578 = pi15 & ~pi32;
  assign n1579 = pi16 & pi32;
  assign n1580 = pi33 & ~n1579;
  assign n1581 = ~n1578 & n1580;
  assign n1582 = ~pi33 & n1579;
  assign n1583 = ~n1581 & ~n1582;
  assign n1584 = ~n1577 & ~n1583;
  assign n1585 = ~n1575 & n1583;
  assign n1586 = ~n1576 & n1585;
  assign n1587 = ~n1584 & ~n1586;
  assign n1588 = ~n1556 & n1587;
  assign n1589 = ~n1554 & ~n1587;
  assign n1590 = ~n1555 & n1589;
  assign n1591 = ~n1588 & ~n1590;
  assign n1592 = ~n1382 & n1414;
  assign n1593 = ~n1381 & ~n1592;
  assign n1594 = ~n1354 & ~n1363;
  assign n1595 = ~n1361 & n1594;
  assign n1596 = ~n1352 & n1595;
  assign n1597 = ~n1377 & ~n1596;
  assign n1598 = pi01 & ~n1212;
  assign n1599 = ~n1213 & n1598;
  assign n1600 = ~n1425 & n1599;
  assign n1601 = pi02 & ~n1214;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = pi47 & ~n1602;
  assign n1604 = ~pi47 & ~n1601;
  assign n1605 = ~n1600 & n1604;
  assign n1606 = ~n1603 & ~n1605;
  assign n1607 = pi47 & ~pi48;
  assign n1608 = ~pi47 & pi48;
  assign n1609 = ~n1607 & ~n1608;
  assign n1610 = pi00 & ~n1609;
  assign n1611 = pi49 & ~n1610;
  assign n1612 = pi00 & ~pi49;
  assign n1613 = ~n1609 & n1612;
  assign n1614 = ~n1611 & ~n1613;
  assign n1615 = ~n1606 & n1614;
  assign n1616 = ~n1605 & ~n1614;
  assign n1617 = ~n1603 & n1616;
  assign n1618 = ~n1615 & ~n1617;
  assign n1619 = pi03 & ~n1006;
  assign n1620 = ~n1007 & n1619;
  assign n1621 = ~n1068 & n1620;
  assign n1622 = pi04 & ~n1008;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = pi45 & ~n1623;
  assign n1625 = ~pi45 & ~n1622;
  assign n1626 = ~n1621 & n1625;
  assign n1627 = ~n1624 & ~n1626;
  assign n1628 = ~n1444 & n1627;
  assign n1629 = ~n1618 & n1628;
  assign n1630 = n1444 & ~n1627;
  assign n1631 = ~n1618 & n1630;
  assign n1632 = ~n1629 & ~n1631;
  assign n1633 = ~n1617 & ~n1627;
  assign n1634 = ~n1444 & n1633;
  assign n1635 = ~n1615 & n1634;
  assign n1636 = ~n1617 & n1627;
  assign n1637 = n1444 & n1636;
  assign n1638 = ~n1615 & n1637;
  assign n1639 = ~n1635 & ~n1638;
  assign n1640 = n1632 & n1639;
  assign n1641 = n1597 & n1640;
  assign n1642 = ~n1597 & ~n1640;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n1593 & n1643;
  assign n1645 = n1593 & ~n1643;
  assign n1646 = ~n1644 & ~n1645;
  assign n1647 = ~n1591 & ~n1646;
  assign n1648 = n1591 & ~n1644;
  assign n1649 = ~n1645 & n1648;
  assign n1650 = ~n1647 & ~n1649;
  assign n1651 = ~n1461 & ~n1512;
  assign n1652 = ~n1506 & n1651;
  assign n1653 = ~n1650 & ~n1652;
  assign n1654 = ~n1513 & n1653;
  assign n1655 = ~n1513 & ~n1652;
  assign n1656 = n1650 & ~n1655;
  assign n1657 = ~n1654 & ~n1656;
  assign n1658 = ~n1505 & ~n1657;
  assign n1659 = n1505 & n1657;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = ~n1502 & n1660;
  assign n1662 = n1502 & ~n1660;
  assign n1663 = ~n1661 & ~n1662;
  assign n1664 = ~n1500 & n1663;
  assign n1665 = ~n1494 & ~n1663;
  assign n1666 = ~n1499 & n1665;
  assign po16 = n1664 | n1666;
  assign n1668 = n1181 & ~n1482;
  assign n1669 = ~n1483 & n1668;
  assign n1670 = n1336 & n1669;
  assign n1671 = n1493 & ~n1670;
  assign n1672 = n1663 & ~n1671;
  assign n1673 = n1184 & ~n1335;
  assign n1674 = n1663 & n1673;
  assign n1675 = n1485 & n1674;
  assign n1676 = ~n1057 & n1675;
  assign n1677 = ~n1480 & ~n1658;
  assign n1678 = ~n1659 & n1677;
  assign n1679 = n1501 & n1678;
  assign n1680 = n1480 & ~n1659;
  assign n1681 = ~n1658 & ~n1680;
  assign n1682 = ~n1461 & ~n1509;
  assign n1683 = ~n1506 & n1682;
  assign n1684 = ~n1650 & n1683;
  assign n1685 = ~n1461 & n1512;
  assign n1686 = ~n1506 & n1685;
  assign n1687 = n1509 & ~n1512;
  assign n1688 = ~n1507 & n1687;
  assign n1689 = ~n1686 & ~n1688;
  assign n1690 = ~n1684 & n1689;
  assign n1691 = n1509 & ~n1647;
  assign n1692 = ~n1649 & n1691;
  assign n1693 = n1512 & ~n1650;
  assign n1694 = ~n1692 & ~n1693;
  assign n1695 = n1690 & n1694;
  assign n1696 = ~n1564 & ~n1573;
  assign n1697 = ~n1571 & n1696;
  assign n1698 = ~n1562 & n1697;
  assign n1699 = ~n1584 & ~n1698;
  assign n1700 = pi06 & ~n683;
  assign n1701 = ~n684 & n1700;
  assign n1702 = ~n1231 & n1701;
  assign n1703 = pi07 & ~n685;
  assign n1704 = ~n1702 & ~n1703;
  assign n1705 = pi43 & ~n1704;
  assign n1706 = pi08 & ~n489;
  assign n1707 = ~n490 & n1706;
  assign n1708 = ~n572 & n1707;
  assign n1709 = pi09 & ~n491;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = pi41 & ~n1710;
  assign n1712 = ~pi41 & ~n1709;
  assign n1713 = ~n1708 & n1712;
  assign n1714 = ~pi43 & ~n1703;
  assign n1715 = ~n1702 & n1714;
  assign n1716 = ~n1713 & ~n1715;
  assign n1717 = ~n1711 & n1716;
  assign n1718 = ~n1705 & n1717;
  assign n1719 = ~n1711 & ~n1713;
  assign n1720 = ~n1705 & ~n1715;
  assign n1721 = ~n1719 & ~n1720;
  assign n1722 = ~n1718 & ~n1721;
  assign n1723 = pi10 & ~n304;
  assign n1724 = ~n305 & n1723;
  assign n1725 = ~n394 & n1724;
  assign n1726 = pi11 & ~n306;
  assign n1727 = ~n1725 & ~n1726;
  assign n1728 = pi39 & ~n1727;
  assign n1729 = ~pi39 & ~n1726;
  assign n1730 = ~n1725 & n1729;
  assign n1731 = ~n1728 & ~n1730;
  assign n1732 = ~n1722 & n1731;
  assign n1733 = ~n1718 & ~n1731;
  assign n1734 = ~n1721 & n1733;
  assign n1735 = ~n1732 & ~n1734;
  assign n1736 = ~n1699 & ~n1735;
  assign n1737 = n1699 & n1735;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = pi12 & ~n193;
  assign n1740 = ~n194 & n1739;
  assign n1741 = ~n729 & n1740;
  assign n1742 = pi13 & ~n195;
  assign n1743 = ~n1741 & ~n1742;
  assign n1744 = pi37 & ~n1743;
  assign n1745 = ~pi37 & ~n1742;
  assign n1746 = ~n1741 & n1745;
  assign n1747 = ~n1744 & ~n1746;
  assign n1748 = pi14 & ~n141;
  assign n1749 = ~n142 & n1748;
  assign n1750 = ~n156 & n1749;
  assign n1751 = pi15 & ~n143;
  assign n1752 = ~n1750 & ~n1751;
  assign n1753 = pi35 & ~n1752;
  assign n1754 = ~pi35 & ~n1751;
  assign n1755 = ~n1750 & n1754;
  assign n1756 = ~n1753 & ~n1755;
  assign n1757 = n1747 & ~n1756;
  assign n1758 = ~n1747 & n1756;
  assign n1759 = pi16 & ~pi32;
  assign n1760 = pi17 & pi32;
  assign n1761 = pi33 & ~n1760;
  assign n1762 = ~n1759 & n1761;
  assign n1763 = ~pi33 & n1760;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = ~n1758 & n1764;
  assign n1766 = ~n1757 & n1765;
  assign n1767 = ~n1757 & ~n1758;
  assign n1768 = ~n1764 & ~n1767;
  assign n1769 = ~n1766 & ~n1768;
  assign n1770 = ~n1738 & n1769;
  assign n1771 = ~n1736 & ~n1769;
  assign n1772 = ~n1737 & n1771;
  assign n1773 = ~n1770 & ~n1772;
  assign n1774 = ~n1555 & n1587;
  assign n1775 = ~n1554 & ~n1774;
  assign n1776 = ~n1615 & ~n1633;
  assign n1777 = ~n1539 & n1549;
  assign n1778 = ~n1536 & ~n1777;
  assign n1779 = ~n1776 & n1778;
  assign n1780 = pi48 & ~pi49;
  assign n1781 = ~pi48 & pi49;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = pi00 & ~n1607;
  assign n1784 = ~n1608 & n1783;
  assign n1785 = ~n1782 & n1784;
  assign n1786 = pi01 & ~n1609;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = pi49 & ~n1787;
  assign n1789 = pi02 & ~n1212;
  assign n1790 = ~n1213 & n1789;
  assign n1791 = ~n1425 & n1790;
  assign n1792 = pi03 & ~n1214;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = pi47 & ~n1793;
  assign n1795 = ~pi47 & ~n1792;
  assign n1796 = ~n1791 & n1795;
  assign n1797 = ~pi49 & ~n1786;
  assign n1798 = ~n1785 & n1797;
  assign n1799 = ~n1796 & ~n1798;
  assign n1800 = ~n1794 & n1799;
  assign n1801 = ~n1788 & n1800;
  assign n1802 = ~n1794 & ~n1796;
  assign n1803 = ~n1788 & ~n1798;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1801 & ~n1804;
  assign n1806 = pi04 & ~n1006;
  assign n1807 = ~n1007 & n1806;
  assign n1808 = ~n1068 & n1807;
  assign n1809 = pi05 & ~n1008;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = pi45 & ~n1810;
  assign n1812 = ~pi45 & ~n1809;
  assign n1813 = ~n1808 & n1812;
  assign n1814 = ~n1811 & ~n1813;
  assign n1815 = ~n1805 & n1814;
  assign n1816 = ~n1801 & ~n1814;
  assign n1817 = ~n1804 & n1816;
  assign n1818 = ~n1815 & ~n1817;
  assign n1819 = n1779 & n1818;
  assign n1820 = ~n1776 & ~n1778;
  assign n1821 = ~n1818 & n1820;
  assign n1822 = ~n1819 & ~n1821;
  assign n1823 = n1776 & ~n1815;
  assign n1824 = ~n1778 & ~n1817;
  assign n1825 = n1823 & n1824;
  assign n1826 = ~n1536 & ~n1615;
  assign n1827 = ~n1633 & n1826;
  assign n1828 = ~n1777 & n1827;
  assign n1829 = ~n1818 & n1828;
  assign n1830 = ~n1825 & ~n1829;
  assign n1831 = n1822 & n1830;
  assign n1832 = ~n1775 & n1831;
  assign n1833 = n1775 & ~n1831;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = ~n1773 & ~n1834;
  assign n1836 = n1773 & ~n1832;
  assign n1837 = ~n1833 & n1836;
  assign n1838 = ~n1835 & ~n1837;
  assign n1839 = ~n1591 & ~n1645;
  assign n1840 = ~n1618 & n1627;
  assign n1841 = ~n1615 & n1633;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = n1444 & ~n1842;
  assign n1844 = ~n1642 & ~n1843;
  assign n1845 = ~n1644 & ~n1844;
  assign n1846 = ~n1839 & n1845;
  assign n1847 = ~n1644 & ~n1839;
  assign n1848 = n1844 & ~n1847;
  assign n1849 = ~n1846 & ~n1848;
  assign n1850 = ~n1838 & ~n1849;
  assign n1851 = n1838 & n1849;
  assign n1852 = ~n1850 & ~n1851;
  assign n1853 = ~n1695 & n1852;
  assign n1854 = n1695 & ~n1852;
  assign n1855 = ~n1853 & ~n1854;
  assign n1856 = ~n1681 & n1855;
  assign n1857 = n1681 & ~n1855;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1679 & ~n1858;
  assign n1860 = ~n1676 & n1859;
  assign n1861 = ~n1672 & n1860;
  assign n1862 = ~n1676 & ~n1679;
  assign n1863 = ~n1672 & n1862;
  assign n1864 = n1858 & ~n1863;
  assign po17 = ~n1861 & ~n1864;
  assign n1866 = ~n1658 & ~n1853;
  assign n1867 = ~n1854 & n1866;
  assign n1868 = n1680 & n1867;
  assign n1869 = ~n1844 & ~n1847;
  assign n1870 = ~n1850 & ~n1869;
  assign n1871 = ~n1746 & ~n1755;
  assign n1872 = ~n1753 & n1871;
  assign n1873 = ~n1744 & n1872;
  assign n1874 = ~n1768 & ~n1873;
  assign n1875 = pi07 & ~n683;
  assign n1876 = ~n684 & n1875;
  assign n1877 = ~n1231 & n1876;
  assign n1878 = pi08 & ~n685;
  assign n1879 = ~n1877 & ~n1878;
  assign n1880 = pi43 & ~n1879;
  assign n1881 = pi09 & ~n489;
  assign n1882 = ~n490 & n1881;
  assign n1883 = ~n572 & n1882;
  assign n1884 = pi10 & ~n491;
  assign n1885 = ~n1883 & ~n1884;
  assign n1886 = pi41 & ~n1885;
  assign n1887 = ~pi41 & ~n1884;
  assign n1888 = ~n1883 & n1887;
  assign n1889 = ~pi43 & ~n1878;
  assign n1890 = ~n1877 & n1889;
  assign n1891 = ~n1888 & ~n1890;
  assign n1892 = ~n1886 & n1891;
  assign n1893 = ~n1880 & n1892;
  assign n1894 = ~n1886 & ~n1888;
  assign n1895 = ~n1880 & ~n1890;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = ~n1893 & ~n1896;
  assign n1898 = pi11 & ~n304;
  assign n1899 = ~n305 & n1898;
  assign n1900 = ~n394 & n1899;
  assign n1901 = pi12 & ~n306;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = pi39 & ~n1902;
  assign n1904 = ~pi39 & ~n1901;
  assign n1905 = ~n1900 & n1904;
  assign n1906 = ~n1903 & ~n1905;
  assign n1907 = ~n1897 & n1906;
  assign n1908 = ~n1893 & ~n1906;
  assign n1909 = ~n1896 & n1908;
  assign n1910 = ~n1907 & ~n1909;
  assign n1911 = ~n1874 & ~n1910;
  assign n1912 = n1874 & n1910;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = pi13 & ~n193;
  assign n1915 = ~n194 & n1914;
  assign n1916 = ~n729 & n1915;
  assign n1917 = pi14 & ~n195;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = pi37 & ~n1918;
  assign n1920 = ~pi37 & ~n1917;
  assign n1921 = ~n1916 & n1920;
  assign n1922 = ~n1919 & ~n1921;
  assign n1923 = pi15 & ~n141;
  assign n1924 = ~n142 & n1923;
  assign n1925 = ~n156 & n1924;
  assign n1926 = pi16 & ~n143;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = pi35 & ~n1927;
  assign n1929 = ~pi35 & ~n1926;
  assign n1930 = ~n1925 & n1929;
  assign n1931 = ~n1928 & ~n1930;
  assign n1932 = n1922 & ~n1931;
  assign n1933 = ~n1922 & n1931;
  assign n1934 = pi17 & ~pi32;
  assign n1935 = pi18 & pi32;
  assign n1936 = pi33 & ~n1935;
  assign n1937 = ~n1934 & n1936;
  assign n1938 = ~pi33 & n1935;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = ~n1933 & n1939;
  assign n1941 = ~n1932 & n1940;
  assign n1942 = ~n1932 & ~n1933;
  assign n1943 = ~n1939 & ~n1942;
  assign n1944 = ~n1941 & ~n1943;
  assign n1945 = ~n1913 & n1944;
  assign n1946 = ~n1911 & ~n1944;
  assign n1947 = ~n1912 & n1946;
  assign n1948 = ~n1945 & ~n1947;
  assign n1949 = ~n1737 & n1769;
  assign n1950 = ~n1736 & ~n1949;
  assign n1951 = pi01 & ~n1607;
  assign n1952 = ~n1608 & n1951;
  assign n1953 = ~n1782 & n1952;
  assign n1954 = pi02 & ~n1609;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = pi49 & ~n1955;
  assign n1957 = pi03 & ~n1212;
  assign n1958 = ~n1213 & n1957;
  assign n1959 = ~n1425 & n1958;
  assign n1960 = pi04 & ~n1214;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = pi47 & ~n1961;
  assign n1963 = ~pi47 & ~n1960;
  assign n1964 = ~n1959 & n1963;
  assign n1965 = ~pi49 & ~n1954;
  assign n1966 = ~n1953 & n1965;
  assign n1967 = ~n1964 & ~n1966;
  assign n1968 = ~n1962 & n1967;
  assign n1969 = ~n1956 & n1968;
  assign n1970 = ~n1962 & ~n1964;
  assign n1971 = ~n1956 & ~n1966;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1969 & ~n1972;
  assign n1974 = pi05 & ~n1006;
  assign n1975 = ~n1007 & n1974;
  assign n1976 = ~n1068 & n1975;
  assign n1977 = pi06 & ~n1008;
  assign n1978 = ~n1976 & ~n1977;
  assign n1979 = pi45 & ~n1978;
  assign n1980 = ~pi45 & ~n1977;
  assign n1981 = ~n1976 & n1980;
  assign n1982 = ~n1979 & ~n1981;
  assign n1983 = ~n1973 & n1982;
  assign n1984 = ~n1804 & n1814;
  assign n1985 = ~n1801 & ~n1984;
  assign n1986 = ~n1983 & n1985;
  assign n1987 = ~n1969 & ~n1982;
  assign n1988 = ~n1972 & n1987;
  assign n1989 = ~n1721 & n1731;
  assign n1990 = ~n1718 & ~n1989;
  assign n1991 = ~n1988 & ~n1990;
  assign n1992 = n1986 & n1991;
  assign n1993 = ~n1983 & n1990;
  assign n1994 = ~n1985 & ~n1988;
  assign n1995 = n1993 & n1994;
  assign n1996 = ~n1992 & ~n1995;
  assign n1997 = ~n1983 & ~n1988;
  assign n1998 = ~n1985 & ~n1990;
  assign n1999 = ~n1997 & n1998;
  assign n2000 = ~n1718 & ~n1801;
  assign n2001 = ~n1989 & n2000;
  assign n2002 = ~n1984 & n2001;
  assign n2003 = ~n1997 & n2002;
  assign n2004 = ~n1999 & ~n2003;
  assign n2005 = n1996 & n2004;
  assign n2006 = ~n1950 & ~n2005;
  assign n2007 = ~n1995 & ~n1999;
  assign n2008 = ~n2003 & n2007;
  assign n2009 = ~n1736 & ~n1992;
  assign n2010 = ~n1949 & n2009;
  assign n2011 = n2008 & n2010;
  assign n2012 = ~n2006 & ~n2011;
  assign n2013 = ~n1948 & ~n2012;
  assign n2014 = n1948 & ~n2006;
  assign n2015 = ~n2011 & n2014;
  assign n2016 = ~n2013 & ~n2015;
  assign n2017 = n1776 & ~n1818;
  assign n2018 = ~n1776 & ~n1815;
  assign n2019 = ~n1817 & n2018;
  assign n2020 = ~n1778 & ~n2017;
  assign n2021 = ~n2019 & n2020;
  assign n2022 = ~n2017 & ~n2021;
  assign n2023 = pi49 & ~pi50;
  assign n2024 = ~pi49 & pi50;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = pi00 & ~n2025;
  assign n2027 = ~n2022 & n2026;
  assign n2028 = ~n2017 & ~n2026;
  assign n2029 = ~n2021 & n2028;
  assign n2030 = ~n2027 & ~n2029;
  assign n2031 = ~n1773 & ~n1833;
  assign n2032 = ~n1832 & ~n2031;
  assign n2033 = ~n2030 & n2032;
  assign n2034 = n2030 & ~n2032;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = ~n2016 & ~n2035;
  assign n2037 = n2016 & ~n2033;
  assign n2038 = ~n2034 & n2037;
  assign n2039 = ~n2036 & ~n2038;
  assign n2040 = ~n1870 & ~n2039;
  assign n2041 = n1870 & n2039;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = n1509 & ~n1650;
  assign n2044 = ~n1655 & n2043;
  assign n2045 = ~n1853 & ~n2044;
  assign n2046 = n2042 & ~n2045;
  assign n2047 = ~n2042 & n2045;
  assign n2048 = n1658 & ~n1853;
  assign n2049 = ~n1854 & n2048;
  assign n2050 = ~n2047 & n2049;
  assign n2051 = ~n2046 & n2050;
  assign n2052 = ~n2046 & ~n2047;
  assign n2053 = ~n2049 & ~n2052;
  assign n2054 = ~n2051 & ~n2053;
  assign n2055 = ~n1868 & ~n2054;
  assign n2056 = ~n1864 & n2055;
  assign n2057 = n1868 & ~n2051;
  assign n2058 = ~n2053 & n2057;
  assign n2059 = n1858 & ~n2051;
  assign n2060 = ~n2053 & n2059;
  assign n2061 = ~n1863 & n2060;
  assign n2062 = ~n2058 & ~n2061;
  assign po18 = ~n2056 & n2062;
  assign n2064 = ~n1856 & n2052;
  assign n2065 = ~n1857 & n2064;
  assign n2066 = ~n1863 & n2065;
  assign n2067 = ~n2016 & ~n2033;
  assign n2068 = ~n2034 & n2067;
  assign n2069 = ~n2027 & ~n2034;
  assign n2070 = ~n2068 & n2069;
  assign n2071 = ~n2016 & n2027;
  assign n2072 = n2035 & n2071;
  assign n2073 = ~n1985 & ~n1997;
  assign n2074 = n1986 & ~n1988;
  assign n2075 = ~n1990 & ~n2074;
  assign n2076 = ~n2073 & ~n2075;
  assign n2077 = pi50 & ~pi51;
  assign n2078 = ~pi50 & pi51;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = pi00 & ~n2023;
  assign n2081 = ~n2024 & n2080;
  assign n2082 = ~n2079 & n2081;
  assign n2083 = pi01 & ~n2025;
  assign n2084 = pi00 & pi51;
  assign n2085 = ~n2025 & n2084;
  assign n2086 = ~n2083 & ~n2085;
  assign n2087 = ~n2082 & n2086;
  assign n2088 = ~n2082 & ~n2083;
  assign n2089 = n2085 & ~n2088;
  assign n2090 = ~n2087 & ~n2089;
  assign n2091 = ~n2076 & n2090;
  assign n2092 = ~n2073 & ~n2090;
  assign n2093 = ~n2075 & n2092;
  assign n2094 = ~n2091 & ~n2093;
  assign n2095 = ~n1948 & ~n2011;
  assign n2096 = ~n2006 & ~n2095;
  assign n2097 = n2094 & ~n2096;
  assign n2098 = ~n2094 & n2096;
  assign n2099 = ~n1921 & ~n1930;
  assign n2100 = ~n1928 & n2099;
  assign n2101 = ~n1919 & n2100;
  assign n2102 = ~n1943 & ~n2101;
  assign n2103 = pi08 & ~n683;
  assign n2104 = ~n684 & n2103;
  assign n2105 = ~n1231 & n2104;
  assign n2106 = pi09 & ~n685;
  assign n2107 = ~n2105 & ~n2106;
  assign n2108 = pi43 & ~n2107;
  assign n2109 = pi10 & ~n489;
  assign n2110 = ~n490 & n2109;
  assign n2111 = ~n572 & n2110;
  assign n2112 = pi11 & ~n491;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = pi41 & ~n2113;
  assign n2115 = ~pi41 & ~n2112;
  assign n2116 = ~n2111 & n2115;
  assign n2117 = ~pi43 & ~n2106;
  assign n2118 = ~n2105 & n2117;
  assign n2119 = ~n2116 & ~n2118;
  assign n2120 = ~n2114 & n2119;
  assign n2121 = ~n2108 & n2120;
  assign n2122 = ~n2114 & ~n2116;
  assign n2123 = ~n2108 & ~n2118;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = ~n2121 & ~n2124;
  assign n2126 = pi12 & ~n304;
  assign n2127 = ~n305 & n2126;
  assign n2128 = ~n394 & n2127;
  assign n2129 = pi13 & ~n306;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = pi39 & ~n2130;
  assign n2132 = ~pi39 & ~n2129;
  assign n2133 = ~n2128 & n2132;
  assign n2134 = ~n2131 & ~n2133;
  assign n2135 = ~n2125 & n2134;
  assign n2136 = ~n2121 & ~n2134;
  assign n2137 = ~n2124 & n2136;
  assign n2138 = ~n2135 & ~n2137;
  assign n2139 = ~n2102 & ~n2138;
  assign n2140 = n2102 & n2138;
  assign n2141 = ~n2139 & ~n2140;
  assign n2142 = pi14 & ~n193;
  assign n2143 = ~n194 & n2142;
  assign n2144 = ~n729 & n2143;
  assign n2145 = pi15 & ~n195;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = pi37 & ~n2146;
  assign n2148 = ~pi37 & ~n2145;
  assign n2149 = ~n2144 & n2148;
  assign n2150 = ~n2147 & ~n2149;
  assign n2151 = pi16 & ~n141;
  assign n2152 = ~n142 & n2151;
  assign n2153 = ~n156 & n2152;
  assign n2154 = pi17 & ~n143;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = pi35 & ~n2155;
  assign n2157 = ~pi35 & ~n2154;
  assign n2158 = ~n2153 & n2157;
  assign n2159 = ~n2156 & ~n2158;
  assign n2160 = ~n2150 & n2159;
  assign n2161 = n2150 & ~n2159;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = pi18 & ~pi32;
  assign n2164 = pi19 & pi32;
  assign n2165 = pi33 & ~n2164;
  assign n2166 = ~n2163 & n2165;
  assign n2167 = ~pi33 & n2164;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~n2162 & ~n2168;
  assign n2170 = ~n2160 & n2168;
  assign n2171 = ~n2161 & n2170;
  assign n2172 = ~n2169 & ~n2171;
  assign n2173 = ~n2141 & n2172;
  assign n2174 = ~n2139 & ~n2172;
  assign n2175 = ~n2140 & n2174;
  assign n2176 = ~n2173 & ~n2175;
  assign n2177 = ~n1912 & n1944;
  assign n2178 = ~n1911 & ~n2177;
  assign n2179 = pi02 & ~n1607;
  assign n2180 = ~n1608 & n2179;
  assign n2181 = ~n1782 & n2180;
  assign n2182 = pi03 & ~n1609;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = pi49 & ~n2183;
  assign n2185 = pi04 & ~n1212;
  assign n2186 = ~n1213 & n2185;
  assign n2187 = ~n1425 & n2186;
  assign n2188 = pi05 & ~n1214;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = pi47 & ~n2189;
  assign n2191 = ~pi47 & ~n2188;
  assign n2192 = ~n2187 & n2191;
  assign n2193 = ~pi49 & ~n2182;
  assign n2194 = ~n2181 & n2193;
  assign n2195 = ~n2192 & ~n2194;
  assign n2196 = ~n2190 & n2195;
  assign n2197 = ~n2184 & n2196;
  assign n2198 = ~n2190 & ~n2192;
  assign n2199 = ~n2184 & ~n2194;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = ~n2197 & ~n2200;
  assign n2202 = pi06 & ~n1006;
  assign n2203 = ~n1007 & n2202;
  assign n2204 = ~n1068 & n2203;
  assign n2205 = pi07 & ~n1008;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = pi45 & ~n2206;
  assign n2208 = ~pi45 & ~n2205;
  assign n2209 = ~n2204 & n2208;
  assign n2210 = ~n2207 & ~n2209;
  assign n2211 = ~n2201 & n2210;
  assign n2212 = ~n1972 & n1982;
  assign n2213 = ~n1969 & ~n2212;
  assign n2214 = ~n2211 & n2213;
  assign n2215 = ~n2197 & ~n2210;
  assign n2216 = ~n2200 & n2215;
  assign n2217 = ~n1896 & n1906;
  assign n2218 = ~n1893 & ~n2217;
  assign n2219 = ~n2216 & ~n2218;
  assign n2220 = n2214 & n2219;
  assign n2221 = ~n2211 & n2218;
  assign n2222 = ~n2213 & ~n2216;
  assign n2223 = n2221 & n2222;
  assign n2224 = ~n2220 & ~n2223;
  assign n2225 = ~n2211 & ~n2216;
  assign n2226 = ~n2213 & ~n2218;
  assign n2227 = ~n2225 & n2226;
  assign n2228 = ~n1893 & ~n1969;
  assign n2229 = ~n2217 & n2228;
  assign n2230 = ~n2212 & n2229;
  assign n2231 = ~n2225 & n2230;
  assign n2232 = ~n2227 & ~n2231;
  assign n2233 = n2224 & n2232;
  assign n2234 = ~n2178 & ~n2233;
  assign n2235 = ~n2223 & ~n2227;
  assign n2236 = ~n2231 & n2235;
  assign n2237 = ~n1911 & ~n2220;
  assign n2238 = ~n2177 & n2237;
  assign n2239 = n2236 & n2238;
  assign n2240 = ~n2234 & ~n2239;
  assign n2241 = ~n2176 & ~n2240;
  assign n2242 = n2176 & ~n2234;
  assign n2243 = ~n2239 & n2242;
  assign n2244 = ~n2241 & ~n2243;
  assign n2245 = ~n2098 & n2244;
  assign n2246 = ~n2097 & n2245;
  assign n2247 = ~n2097 & ~n2098;
  assign n2248 = ~n2244 & ~n2247;
  assign n2249 = ~n2246 & ~n2248;
  assign n2250 = ~n2072 & n2249;
  assign n2251 = ~n2070 & n2250;
  assign n2252 = ~n2070 & ~n2072;
  assign n2253 = ~n2249 & ~n2252;
  assign n2254 = ~n2251 & ~n2253;
  assign n2255 = ~n2040 & ~n2046;
  assign n2256 = ~n2254 & ~n2255;
  assign n2257 = ~n2040 & ~n2251;
  assign n2258 = ~n2253 & n2257;
  assign n2259 = ~n2046 & n2258;
  assign n2260 = ~n2256 & ~n2259;
  assign n2261 = ~n1868 & ~n2051;
  assign n2262 = ~n2053 & ~n2261;
  assign n2263 = ~n2260 & ~n2262;
  assign n2264 = ~n2066 & n2263;
  assign n2265 = ~n2053 & ~n2256;
  assign n2266 = ~n2259 & n2265;
  assign n2267 = ~n2261 & n2266;
  assign n2268 = n2065 & n2260;
  assign n2269 = ~n1863 & n2268;
  assign n2270 = ~n2267 & ~n2269;
  assign po19 = ~n2264 & n2270;
  assign n2272 = ~n2249 & n2252;
  assign n2273 = ~n2072 & ~n2272;
  assign n2274 = ~n2176 & ~n2239;
  assign n2275 = ~n2234 & ~n2274;
  assign n2276 = n2214 & ~n2216;
  assign n2277 = ~n2218 & ~n2276;
  assign n2278 = ~n2213 & ~n2225;
  assign n2279 = pi01 & ~n2023;
  assign n2280 = ~n2024 & n2279;
  assign n2281 = ~n2079 & n2280;
  assign n2282 = pi02 & ~n2025;
  assign n2283 = ~n2281 & ~n2282;
  assign n2284 = pi51 & ~n2283;
  assign n2285 = ~pi51 & ~n2282;
  assign n2286 = ~n2281 & n2285;
  assign n2287 = ~n2284 & ~n2286;
  assign n2288 = pi51 & ~pi52;
  assign n2289 = ~pi51 & pi52;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = pi00 & ~n2290;
  assign n2292 = ~n2287 & n2291;
  assign n2293 = ~n2286 & ~n2291;
  assign n2294 = ~n2284 & n2293;
  assign n2295 = ~n2292 & ~n2294;
  assign n2296 = pi51 & ~n2026;
  assign n2297 = n2088 & n2296;
  assign n2298 = ~n2295 & ~n2297;
  assign n2299 = ~n2294 & n2297;
  assign n2300 = ~n2292 & n2299;
  assign n2301 = ~n2298 & ~n2300;
  assign n2302 = ~n2278 & n2301;
  assign n2303 = ~n2277 & n2302;
  assign n2304 = ~n2277 & ~n2278;
  assign n2305 = ~n2301 & ~n2304;
  assign n2306 = ~n2303 & ~n2305;
  assign n2307 = ~n2275 & n2306;
  assign n2308 = n2275 & ~n2306;
  assign n2309 = ~n2307 & ~n2308;
  assign n2310 = ~n2140 & n2172;
  assign n2311 = ~n2139 & ~n2310;
  assign n2312 = pi03 & ~n1607;
  assign n2313 = ~n1608 & n2312;
  assign n2314 = ~n1782 & n2313;
  assign n2315 = pi04 & ~n1609;
  assign n2316 = ~n2314 & ~n2315;
  assign n2317 = pi49 & ~n2316;
  assign n2318 = pi05 & ~n1212;
  assign n2319 = ~n1213 & n2318;
  assign n2320 = ~n1425 & n2319;
  assign n2321 = pi06 & ~n1214;
  assign n2322 = ~n2320 & ~n2321;
  assign n2323 = pi47 & ~n2322;
  assign n2324 = ~pi47 & ~n2321;
  assign n2325 = ~n2320 & n2324;
  assign n2326 = ~pi49 & ~n2315;
  assign n2327 = ~n2314 & n2326;
  assign n2328 = ~n2325 & ~n2327;
  assign n2329 = ~n2323 & n2328;
  assign n2330 = ~n2317 & n2329;
  assign n2331 = ~n2323 & ~n2325;
  assign n2332 = ~n2317 & ~n2327;
  assign n2333 = ~n2331 & ~n2332;
  assign n2334 = ~n2330 & ~n2333;
  assign n2335 = pi07 & ~n1006;
  assign n2336 = ~n1007 & n2335;
  assign n2337 = ~n1068 & n2336;
  assign n2338 = pi08 & ~n1008;
  assign n2339 = ~n2337 & ~n2338;
  assign n2340 = pi45 & ~n2339;
  assign n2341 = ~pi45 & ~n2338;
  assign n2342 = ~n2337 & n2341;
  assign n2343 = ~n2340 & ~n2342;
  assign n2344 = ~n2334 & n2343;
  assign n2345 = ~n2200 & n2210;
  assign n2346 = ~n2197 & ~n2345;
  assign n2347 = ~n2344 & n2346;
  assign n2348 = ~n2330 & ~n2343;
  assign n2349 = ~n2333 & n2348;
  assign n2350 = ~n2124 & n2134;
  assign n2351 = ~n2121 & ~n2350;
  assign n2352 = ~n2349 & ~n2351;
  assign n2353 = n2347 & n2352;
  assign n2354 = ~n2344 & n2351;
  assign n2355 = ~n2346 & ~n2349;
  assign n2356 = n2354 & n2355;
  assign n2357 = ~n2353 & ~n2356;
  assign n2358 = ~n2344 & ~n2349;
  assign n2359 = ~n2346 & ~n2351;
  assign n2360 = ~n2358 & n2359;
  assign n2361 = ~n2121 & ~n2197;
  assign n2362 = ~n2350 & n2361;
  assign n2363 = ~n2345 & n2362;
  assign n2364 = ~n2358 & n2363;
  assign n2365 = ~n2360 & ~n2364;
  assign n2366 = n2357 & n2365;
  assign n2367 = ~n2311 & ~n2366;
  assign n2368 = ~n2149 & ~n2158;
  assign n2369 = ~n2156 & n2368;
  assign n2370 = ~n2147 & n2369;
  assign n2371 = ~n2169 & ~n2370;
  assign n2372 = pi09 & ~n683;
  assign n2373 = ~n684 & n2372;
  assign n2374 = ~n1231 & n2373;
  assign n2375 = pi10 & ~n685;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = pi43 & ~n2376;
  assign n2378 = pi11 & ~n489;
  assign n2379 = ~n490 & n2378;
  assign n2380 = ~n572 & n2379;
  assign n2381 = pi12 & ~n491;
  assign n2382 = ~n2380 & ~n2381;
  assign n2383 = pi41 & ~n2382;
  assign n2384 = ~pi41 & ~n2381;
  assign n2385 = ~n2380 & n2384;
  assign n2386 = ~pi43 & ~n2375;
  assign n2387 = ~n2374 & n2386;
  assign n2388 = ~n2385 & ~n2387;
  assign n2389 = ~n2383 & n2388;
  assign n2390 = ~n2377 & n2389;
  assign n2391 = ~n2383 & ~n2385;
  assign n2392 = ~n2377 & ~n2387;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = ~n2390 & ~n2393;
  assign n2395 = pi13 & ~n304;
  assign n2396 = ~n305 & n2395;
  assign n2397 = ~n394 & n2396;
  assign n2398 = pi14 & ~n306;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = pi39 & ~n2399;
  assign n2401 = ~pi39 & ~n2398;
  assign n2402 = ~n2397 & n2401;
  assign n2403 = ~n2400 & ~n2402;
  assign n2404 = ~n2394 & n2403;
  assign n2405 = ~n2390 & ~n2403;
  assign n2406 = ~n2393 & n2405;
  assign n2407 = ~n2404 & ~n2406;
  assign n2408 = ~n2371 & ~n2407;
  assign n2409 = n2371 & n2407;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = pi15 & ~n193;
  assign n2412 = ~n194 & n2411;
  assign n2413 = ~n729 & n2412;
  assign n2414 = pi16 & ~n195;
  assign n2415 = ~n2413 & ~n2414;
  assign n2416 = pi37 & ~n2415;
  assign n2417 = ~pi37 & ~n2414;
  assign n2418 = ~n2413 & n2417;
  assign n2419 = ~n2416 & ~n2418;
  assign n2420 = pi17 & ~n141;
  assign n2421 = ~n142 & n2420;
  assign n2422 = ~n156 & n2421;
  assign n2423 = pi18 & ~n143;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = pi35 & ~n2424;
  assign n2426 = ~pi35 & ~n2423;
  assign n2427 = ~n2422 & n2426;
  assign n2428 = ~n2425 & ~n2427;
  assign n2429 = n2419 & ~n2428;
  assign n2430 = ~n2419 & n2428;
  assign n2431 = pi19 & ~pi32;
  assign n2432 = pi20 & pi32;
  assign n2433 = pi33 & ~n2432;
  assign n2434 = ~n2431 & n2433;
  assign n2435 = ~pi33 & n2432;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = ~n2430 & n2436;
  assign n2438 = ~n2429 & n2437;
  assign n2439 = ~n2429 & ~n2430;
  assign n2440 = ~n2436 & ~n2439;
  assign n2441 = ~n2438 & ~n2440;
  assign n2442 = ~n2410 & n2441;
  assign n2443 = ~n2408 & ~n2441;
  assign n2444 = ~n2409 & n2443;
  assign n2445 = ~n2442 & ~n2444;
  assign n2446 = ~n2356 & ~n2360;
  assign n2447 = ~n2364 & n2446;
  assign n2448 = ~n2139 & ~n2353;
  assign n2449 = ~n2310 & n2448;
  assign n2450 = n2447 & n2449;
  assign n2451 = ~n2445 & ~n2450;
  assign n2452 = ~n2367 & n2451;
  assign n2453 = ~n2367 & ~n2450;
  assign n2454 = n2445 & ~n2453;
  assign n2455 = ~n2452 & ~n2454;
  assign n2456 = ~n2309 & n2455;
  assign n2457 = n2309 & ~n2455;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = ~n2097 & n2244;
  assign n2460 = ~n2098 & ~n2459;
  assign n2461 = n2091 & ~n2460;
  assign n2462 = ~n2091 & ~n2098;
  assign n2463 = ~n2459 & n2462;
  assign n2464 = ~n2461 & ~n2463;
  assign n2465 = ~n2458 & ~n2464;
  assign n2466 = n2458 & n2464;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = ~n2273 & n2467;
  assign n2469 = n2273 & ~n2467;
  assign n2470 = ~n2468 & ~n2469;
  assign n2471 = n2040 & ~n2254;
  assign n2472 = ~n2470 & n2471;
  assign n2473 = n2470 & ~n2471;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = n1663 & ~n2256;
  assign n2476 = ~n2259 & n2475;
  assign n2477 = n2065 & n2476;
  assign n2478 = n1500 & n2477;
  assign n2479 = n2046 & ~n2254;
  assign n2480 = n1679 & ~n1857;
  assign n2481 = n2064 & n2480;
  assign n2482 = ~n2262 & ~n2481;
  assign n2483 = n2260 & ~n2482;
  assign n2484 = ~n2479 & ~n2483;
  assign n2485 = ~n2478 & n2484;
  assign n2486 = ~n2474 & ~n2485;
  assign n2487 = ~n2472 & ~n2479;
  assign n2488 = ~n2473 & n2487;
  assign n2489 = ~n2483 & n2488;
  assign n2490 = ~n2478 & n2489;
  assign po20 = ~n2486 & ~n2490;
  assign n2492 = ~n2468 & n2471;
  assign n2493 = ~n2469 & n2492;
  assign n2494 = ~n2418 & ~n2427;
  assign n2495 = ~n2425 & n2494;
  assign n2496 = ~n2416 & n2495;
  assign n2497 = ~n2440 & ~n2496;
  assign n2498 = pi10 & ~n683;
  assign n2499 = ~n684 & n2498;
  assign n2500 = ~n1231 & n2499;
  assign n2501 = pi11 & ~n685;
  assign n2502 = ~n2500 & ~n2501;
  assign n2503 = pi43 & ~n2502;
  assign n2504 = pi12 & ~n489;
  assign n2505 = ~n490 & n2504;
  assign n2506 = ~n572 & n2505;
  assign n2507 = pi13 & ~n491;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = pi41 & ~n2508;
  assign n2510 = ~pi41 & ~n2507;
  assign n2511 = ~n2506 & n2510;
  assign n2512 = ~pi43 & ~n2501;
  assign n2513 = ~n2500 & n2512;
  assign n2514 = ~n2511 & ~n2513;
  assign n2515 = ~n2509 & n2514;
  assign n2516 = ~n2503 & n2515;
  assign n2517 = ~n2509 & ~n2511;
  assign n2518 = ~n2503 & ~n2513;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520 = ~n2516 & ~n2519;
  assign n2521 = pi14 & ~n304;
  assign n2522 = ~n305 & n2521;
  assign n2523 = ~n394 & n2522;
  assign n2524 = pi15 & ~n306;
  assign n2525 = ~n2523 & ~n2524;
  assign n2526 = pi39 & ~n2525;
  assign n2527 = ~pi39 & ~n2524;
  assign n2528 = ~n2523 & n2527;
  assign n2529 = ~n2526 & ~n2528;
  assign n2530 = ~n2520 & n2529;
  assign n2531 = ~n2516 & ~n2529;
  assign n2532 = ~n2519 & n2531;
  assign n2533 = ~n2530 & ~n2532;
  assign n2534 = ~n2497 & ~n2533;
  assign n2535 = n2497 & n2533;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = pi16 & ~n193;
  assign n2538 = ~n194 & n2537;
  assign n2539 = ~n729 & n2538;
  assign n2540 = pi17 & ~n195;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = pi37 & ~n2541;
  assign n2543 = ~pi37 & ~n2540;
  assign n2544 = ~n2539 & n2543;
  assign n2545 = ~n2542 & ~n2544;
  assign n2546 = pi18 & ~n141;
  assign n2547 = ~n142 & n2546;
  assign n2548 = ~n156 & n2547;
  assign n2549 = pi19 & ~n143;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = pi35 & ~n2550;
  assign n2552 = ~pi35 & ~n2549;
  assign n2553 = ~n2548 & n2552;
  assign n2554 = ~n2551 & ~n2553;
  assign n2555 = n2545 & ~n2554;
  assign n2556 = ~n2545 & n2554;
  assign n2557 = pi20 & ~pi32;
  assign n2558 = pi21 & pi32;
  assign n2559 = pi33 & ~n2558;
  assign n2560 = ~n2557 & n2559;
  assign n2561 = ~pi33 & n2558;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~n2556 & n2562;
  assign n2564 = ~n2555 & n2563;
  assign n2565 = ~n2555 & ~n2556;
  assign n2566 = ~n2562 & ~n2565;
  assign n2567 = ~n2564 & ~n2566;
  assign n2568 = ~n2536 & n2567;
  assign n2569 = ~n2534 & ~n2567;
  assign n2570 = ~n2535 & n2569;
  assign n2571 = ~n2568 & ~n2570;
  assign n2572 = ~n2409 & n2441;
  assign n2573 = ~n2408 & ~n2572;
  assign n2574 = pi04 & ~n1607;
  assign n2575 = ~n1608 & n2574;
  assign n2576 = ~n1782 & n2575;
  assign n2577 = pi05 & ~n1609;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = pi49 & ~n2578;
  assign n2580 = pi06 & ~n1212;
  assign n2581 = ~n1213 & n2580;
  assign n2582 = ~n1425 & n2581;
  assign n2583 = pi07 & ~n1214;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = pi47 & ~n2584;
  assign n2586 = ~pi47 & ~n2583;
  assign n2587 = ~n2582 & n2586;
  assign n2588 = ~pi49 & ~n2577;
  assign n2589 = ~n2576 & n2588;
  assign n2590 = ~n2587 & ~n2589;
  assign n2591 = ~n2585 & n2590;
  assign n2592 = ~n2579 & n2591;
  assign n2593 = ~n2585 & ~n2587;
  assign n2594 = ~n2579 & ~n2589;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = ~n2592 & ~n2595;
  assign n2597 = pi08 & ~n1006;
  assign n2598 = ~n1007 & n2597;
  assign n2599 = ~n1068 & n2598;
  assign n2600 = pi09 & ~n1008;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = pi45 & ~n2601;
  assign n2603 = ~pi45 & ~n2600;
  assign n2604 = ~n2599 & n2603;
  assign n2605 = ~n2602 & ~n2604;
  assign n2606 = ~n2596 & n2605;
  assign n2607 = ~n2333 & n2343;
  assign n2608 = ~n2330 & ~n2607;
  assign n2609 = ~n2606 & n2608;
  assign n2610 = ~n2592 & ~n2605;
  assign n2611 = ~n2595 & n2610;
  assign n2612 = ~n2393 & n2403;
  assign n2613 = ~n2390 & ~n2612;
  assign n2614 = ~n2611 & ~n2613;
  assign n2615 = n2609 & n2614;
  assign n2616 = ~n2606 & n2613;
  assign n2617 = ~n2608 & ~n2611;
  assign n2618 = n2616 & n2617;
  assign n2619 = ~n2615 & ~n2618;
  assign n2620 = ~n2606 & ~n2611;
  assign n2621 = ~n2608 & ~n2613;
  assign n2622 = ~n2620 & n2621;
  assign n2623 = ~n2330 & ~n2390;
  assign n2624 = ~n2612 & n2623;
  assign n2625 = ~n2607 & n2624;
  assign n2626 = ~n2620 & n2625;
  assign n2627 = ~n2622 & ~n2626;
  assign n2628 = n2619 & n2627;
  assign n2629 = ~n2573 & ~n2628;
  assign n2630 = ~n2618 & ~n2622;
  assign n2631 = ~n2626 & n2630;
  assign n2632 = ~n2408 & ~n2615;
  assign n2633 = ~n2572 & n2632;
  assign n2634 = n2631 & n2633;
  assign n2635 = ~n2629 & ~n2634;
  assign n2636 = ~n2571 & ~n2635;
  assign n2637 = n2571 & ~n2629;
  assign n2638 = ~n2634 & n2637;
  assign n2639 = ~n2636 & ~n2638;
  assign n2640 = ~n2346 & ~n2358;
  assign n2641 = n2347 & ~n2349;
  assign n2642 = ~n2351 & ~n2640;
  assign n2643 = ~n2641 & n2642;
  assign n2644 = ~n2640 & ~n2643;
  assign n2645 = pi52 & ~pi53;
  assign n2646 = ~pi52 & pi53;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = pi00 & ~n2288;
  assign n2649 = ~n2289 & n2648;
  assign n2650 = ~n2647 & n2649;
  assign n2651 = pi01 & ~n2290;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = pi53 & ~n2652;
  assign n2654 = pi02 & ~n2023;
  assign n2655 = ~n2024 & n2654;
  assign n2656 = ~n2079 & n2655;
  assign n2657 = pi03 & ~n2025;
  assign n2658 = ~n2656 & ~n2657;
  assign n2659 = pi51 & ~n2658;
  assign n2660 = ~pi51 & ~n2657;
  assign n2661 = ~n2656 & n2660;
  assign n2662 = ~pi53 & ~n2651;
  assign n2663 = ~n2650 & n2662;
  assign n2664 = ~n2661 & ~n2663;
  assign n2665 = ~n2659 & n2664;
  assign n2666 = ~n2653 & n2665;
  assign n2667 = ~n2659 & ~n2661;
  assign n2668 = ~n2653 & ~n2663;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = ~n2666 & ~n2669;
  assign n2671 = pi53 & ~n2291;
  assign n2672 = ~n2286 & n2291;
  assign n2673 = ~n2284 & n2672;
  assign n2674 = ~n2671 & ~n2673;
  assign n2675 = ~n2670 & n2674;
  assign n2676 = n2670 & ~n2674;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = ~n2644 & n2677;
  assign n2679 = ~n2640 & ~n2677;
  assign n2680 = ~n2643 & n2679;
  assign n2681 = ~n2678 & ~n2680;
  assign n2682 = ~n2367 & ~n2452;
  assign n2683 = ~n2681 & n2682;
  assign n2684 = n2681 & ~n2682;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~n2639 & ~n2685;
  assign n2687 = n2639 & ~n2683;
  assign n2688 = ~n2684 & n2687;
  assign n2689 = ~n2686 & ~n2688;
  assign n2690 = ~n2308 & n2455;
  assign n2691 = ~n2295 & n2297;
  assign n2692 = ~n2305 & ~n2691;
  assign n2693 = ~n2307 & ~n2692;
  assign n2694 = ~n2690 & n2693;
  assign n2695 = ~n2307 & ~n2690;
  assign n2696 = n2692 & ~n2695;
  assign n2697 = ~n2694 & ~n2696;
  assign n2698 = ~n2689 & ~n2697;
  assign n2699 = n2689 & n2697;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = n2091 & ~n2098;
  assign n2702 = ~n2459 & n2701;
  assign n2703 = ~n2465 & ~n2702;
  assign n2704 = n2700 & ~n2703;
  assign n2705 = ~n2700 & n2703;
  assign n2706 = n2468 & ~n2705;
  assign n2707 = ~n2704 & n2706;
  assign n2708 = ~n2704 & ~n2705;
  assign n2709 = ~n2468 & ~n2708;
  assign n2710 = ~n2707 & ~n2709;
  assign n2711 = ~n2493 & ~n2710;
  assign n2712 = ~n2486 & n2711;
  assign n2713 = ~n2486 & ~n2493;
  assign n2714 = n2710 & ~n2713;
  assign po21 = ~n2712 & ~n2714;
  assign n2716 = ~n2474 & n2710;
  assign n2717 = ~n2485 & n2716;
  assign n2718 = ~n2692 & ~n2695;
  assign n2719 = ~n2698 & ~n2718;
  assign n2720 = ~n2544 & ~n2553;
  assign n2721 = ~n2551 & n2720;
  assign n2722 = ~n2542 & n2721;
  assign n2723 = ~n2566 & ~n2722;
  assign n2724 = pi11 & ~n683;
  assign n2725 = ~n684 & n2724;
  assign n2726 = ~n1231 & n2725;
  assign n2727 = pi12 & ~n685;
  assign n2728 = ~n2726 & ~n2727;
  assign n2729 = pi43 & ~n2728;
  assign n2730 = pi13 & ~n489;
  assign n2731 = ~n490 & n2730;
  assign n2732 = ~n572 & n2731;
  assign n2733 = pi14 & ~n491;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = pi41 & ~n2734;
  assign n2736 = ~pi41 & ~n2733;
  assign n2737 = ~n2732 & n2736;
  assign n2738 = ~pi43 & ~n2727;
  assign n2739 = ~n2726 & n2738;
  assign n2740 = ~n2737 & ~n2739;
  assign n2741 = ~n2735 & n2740;
  assign n2742 = ~n2729 & n2741;
  assign n2743 = ~n2735 & ~n2737;
  assign n2744 = ~n2729 & ~n2739;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = ~n2742 & ~n2745;
  assign n2747 = pi15 & ~n304;
  assign n2748 = ~n305 & n2747;
  assign n2749 = ~n394 & n2748;
  assign n2750 = pi16 & ~n306;
  assign n2751 = ~n2749 & ~n2750;
  assign n2752 = pi39 & ~n2751;
  assign n2753 = ~pi39 & ~n2750;
  assign n2754 = ~n2749 & n2753;
  assign n2755 = ~n2752 & ~n2754;
  assign n2756 = ~n2746 & n2755;
  assign n2757 = ~n2742 & ~n2755;
  assign n2758 = ~n2745 & n2757;
  assign n2759 = ~n2756 & ~n2758;
  assign n2760 = ~n2723 & ~n2759;
  assign n2761 = n2723 & n2759;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = pi17 & ~n193;
  assign n2764 = ~n194 & n2763;
  assign n2765 = ~n729 & n2764;
  assign n2766 = pi18 & ~n195;
  assign n2767 = ~n2765 & ~n2766;
  assign n2768 = pi37 & ~n2767;
  assign n2769 = ~pi37 & ~n2766;
  assign n2770 = ~n2765 & n2769;
  assign n2771 = ~n2768 & ~n2770;
  assign n2772 = pi19 & ~n141;
  assign n2773 = ~n142 & n2772;
  assign n2774 = ~n156 & n2773;
  assign n2775 = pi20 & ~n143;
  assign n2776 = ~n2774 & ~n2775;
  assign n2777 = pi35 & ~n2776;
  assign n2778 = ~pi35 & ~n2775;
  assign n2779 = ~n2774 & n2778;
  assign n2780 = ~n2777 & ~n2779;
  assign n2781 = ~n2771 & n2780;
  assign n2782 = n2771 & ~n2780;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = pi21 & ~pi32;
  assign n2785 = pi22 & pi32;
  assign n2786 = pi33 & ~n2785;
  assign n2787 = ~n2784 & n2786;
  assign n2788 = ~pi33 & n2785;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = ~n2783 & ~n2789;
  assign n2791 = ~n2781 & n2789;
  assign n2792 = ~n2782 & n2791;
  assign n2793 = ~n2790 & ~n2792;
  assign n2794 = ~n2762 & n2793;
  assign n2795 = ~n2760 & ~n2793;
  assign n2796 = ~n2761 & n2795;
  assign n2797 = ~n2794 & ~n2796;
  assign n2798 = ~n2535 & n2567;
  assign n2799 = ~n2534 & ~n2798;
  assign n2800 = pi05 & ~n1607;
  assign n2801 = ~n1608 & n2800;
  assign n2802 = ~n1782 & n2801;
  assign n2803 = pi06 & ~n1609;
  assign n2804 = ~n2802 & ~n2803;
  assign n2805 = pi49 & ~n2804;
  assign n2806 = pi07 & ~n1212;
  assign n2807 = ~n1213 & n2806;
  assign n2808 = ~n1425 & n2807;
  assign n2809 = pi08 & ~n1214;
  assign n2810 = ~n2808 & ~n2809;
  assign n2811 = pi47 & ~n2810;
  assign n2812 = ~pi47 & ~n2809;
  assign n2813 = ~n2808 & n2812;
  assign n2814 = ~pi49 & ~n2803;
  assign n2815 = ~n2802 & n2814;
  assign n2816 = ~n2813 & ~n2815;
  assign n2817 = ~n2811 & n2816;
  assign n2818 = ~n2805 & n2817;
  assign n2819 = ~n2811 & ~n2813;
  assign n2820 = ~n2805 & ~n2815;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = ~n2818 & ~n2821;
  assign n2823 = pi09 & ~n1006;
  assign n2824 = ~n1007 & n2823;
  assign n2825 = ~n1068 & n2824;
  assign n2826 = pi10 & ~n1008;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = pi45 & ~n2827;
  assign n2829 = ~pi45 & ~n2826;
  assign n2830 = ~n2825 & n2829;
  assign n2831 = ~n2828 & ~n2830;
  assign n2832 = ~n2822 & n2831;
  assign n2833 = ~n2595 & n2605;
  assign n2834 = ~n2592 & ~n2833;
  assign n2835 = ~n2832 & n2834;
  assign n2836 = ~n2818 & ~n2831;
  assign n2837 = ~n2821 & n2836;
  assign n2838 = ~n2519 & n2529;
  assign n2839 = ~n2516 & ~n2838;
  assign n2840 = ~n2837 & ~n2839;
  assign n2841 = n2835 & n2840;
  assign n2842 = ~n2832 & n2839;
  assign n2843 = ~n2834 & ~n2837;
  assign n2844 = n2842 & n2843;
  assign n2845 = ~n2841 & ~n2844;
  assign n2846 = ~n2832 & ~n2837;
  assign n2847 = ~n2834 & ~n2839;
  assign n2848 = ~n2846 & n2847;
  assign n2849 = ~n2516 & ~n2592;
  assign n2850 = ~n2838 & n2849;
  assign n2851 = ~n2833 & n2850;
  assign n2852 = ~n2846 & n2851;
  assign n2853 = ~n2848 & ~n2852;
  assign n2854 = n2845 & n2853;
  assign n2855 = ~n2799 & ~n2854;
  assign n2856 = ~n2844 & ~n2848;
  assign n2857 = ~n2852 & n2856;
  assign n2858 = ~n2534 & ~n2841;
  assign n2859 = ~n2798 & n2858;
  assign n2860 = n2857 & n2859;
  assign n2861 = ~n2855 & ~n2860;
  assign n2862 = ~n2797 & ~n2861;
  assign n2863 = n2797 & ~n2855;
  assign n2864 = ~n2860 & n2863;
  assign n2865 = ~n2862 & ~n2864;
  assign n2866 = ~n2571 & ~n2634;
  assign n2867 = ~n2629 & ~n2866;
  assign n2868 = pi01 & ~n2288;
  assign n2869 = ~n2289 & n2868;
  assign n2870 = ~n2647 & n2869;
  assign n2871 = pi02 & ~n2290;
  assign n2872 = ~n2870 & ~n2871;
  assign n2873 = pi53 & ~n2872;
  assign n2874 = ~pi53 & ~n2871;
  assign n2875 = ~n2870 & n2874;
  assign n2876 = pi53 & ~pi54;
  assign n2877 = ~pi53 & pi54;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = pi00 & ~n2878;
  assign n2880 = pi55 & ~n2879;
  assign n2881 = pi00 & ~pi55;
  assign n2882 = ~n2878 & n2881;
  assign n2883 = ~n2880 & ~n2882;
  assign n2884 = ~n2875 & ~n2883;
  assign n2885 = ~n2873 & n2884;
  assign n2886 = ~n2873 & ~n2875;
  assign n2887 = n2883 & ~n2886;
  assign n2888 = ~n2885 & ~n2887;
  assign n2889 = pi03 & ~n2023;
  assign n2890 = ~n2024 & n2889;
  assign n2891 = ~n2079 & n2890;
  assign n2892 = pi04 & ~n2025;
  assign n2893 = ~n2891 & ~n2892;
  assign n2894 = pi51 & ~n2893;
  assign n2895 = ~pi51 & ~n2892;
  assign n2896 = ~n2891 & n2895;
  assign n2897 = ~n2894 & ~n2896;
  assign n2898 = ~n2888 & n2897;
  assign n2899 = ~n2885 & ~n2897;
  assign n2900 = ~n2887 & n2899;
  assign n2901 = ~n2898 & ~n2900;
  assign n2902 = pi55 & ~n2666;
  assign n2903 = ~pi55 & ~n2661;
  assign n2904 = ~n2659 & n2903;
  assign n2905 = n2668 & n2904;
  assign n2906 = ~n2902 & ~n2905;
  assign n2907 = ~n2901 & ~n2906;
  assign n2908 = ~n2900 & ~n2905;
  assign n2909 = ~n2902 & n2908;
  assign n2910 = ~n2898 & n2909;
  assign n2911 = ~n2676 & ~n2910;
  assign n2912 = ~n2907 & n2911;
  assign n2913 = ~n2907 & ~n2910;
  assign n2914 = n2676 & ~n2913;
  assign n2915 = ~n2608 & ~n2620;
  assign n2916 = n2609 & ~n2611;
  assign n2917 = ~n2613 & ~n2916;
  assign n2918 = ~n2915 & ~n2917;
  assign n2919 = ~n2914 & n2918;
  assign n2920 = ~n2912 & n2919;
  assign n2921 = ~n2912 & ~n2914;
  assign n2922 = ~n2918 & ~n2921;
  assign n2923 = ~n2920 & ~n2922;
  assign n2924 = ~n2867 & n2923;
  assign n2925 = n2867 & ~n2923;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = ~n2865 & ~n2926;
  assign n2928 = n2865 & ~n2924;
  assign n2929 = ~n2925 & n2928;
  assign n2930 = ~n2927 & ~n2929;
  assign n2931 = n2639 & ~n2684;
  assign n2932 = n2678 & ~n2683;
  assign n2933 = ~n2931 & n2932;
  assign n2934 = ~n2683 & ~n2931;
  assign n2935 = ~n2678 & ~n2934;
  assign n2936 = ~n2933 & ~n2935;
  assign n2937 = ~n2930 & ~n2936;
  assign n2938 = n2930 & ~n2933;
  assign n2939 = ~n2935 & n2938;
  assign n2940 = ~n2937 & ~n2939;
  assign n2941 = n2719 & n2940;
  assign n2942 = ~n2719 & ~n2940;
  assign n2943 = n2704 & ~n2942;
  assign n2944 = ~n2941 & n2943;
  assign n2945 = ~n2941 & ~n2942;
  assign n2946 = ~n2704 & ~n2945;
  assign n2947 = ~n2944 & ~n2946;
  assign n2948 = ~n2469 & n2471;
  assign n2949 = ~n2468 & ~n2948;
  assign n2950 = n2708 & ~n2949;
  assign n2951 = ~n2947 & ~n2950;
  assign n2952 = ~n2717 & n2951;
  assign n2953 = ~n2717 & ~n2950;
  assign n2954 = n2947 & ~n2953;
  assign po22 = ~n2952 & ~n2954;
  assign n2956 = ~n2797 & ~n2860;
  assign n2957 = ~n2855 & ~n2956;
  assign n2958 = pi54 & ~pi55;
  assign n2959 = ~pi54 & pi55;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = pi00 & ~n2876;
  assign n2962 = ~n2877 & n2961;
  assign n2963 = ~n2960 & n2962;
  assign n2964 = pi01 & ~n2878;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = pi55 & ~n2965;
  assign n2967 = pi02 & ~n2288;
  assign n2968 = ~n2289 & n2967;
  assign n2969 = ~n2647 & n2968;
  assign n2970 = pi03 & ~n2290;
  assign n2971 = ~n2969 & ~n2970;
  assign n2972 = pi53 & ~n2971;
  assign n2973 = ~pi53 & ~n2970;
  assign n2974 = ~n2969 & n2973;
  assign n2975 = ~pi55 & ~n2964;
  assign n2976 = ~n2963 & n2975;
  assign n2977 = ~n2974 & ~n2976;
  assign n2978 = ~n2972 & n2977;
  assign n2979 = ~n2966 & n2978;
  assign n2980 = ~n2972 & ~n2974;
  assign n2981 = ~n2966 & ~n2976;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = ~n2979 & ~n2982;
  assign n2984 = pi04 & ~n2023;
  assign n2985 = ~n2024 & n2984;
  assign n2986 = ~n2079 & n2985;
  assign n2987 = pi05 & ~n2025;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = pi51 & ~n2988;
  assign n2990 = ~pi51 & ~n2987;
  assign n2991 = ~n2986 & n2990;
  assign n2992 = ~n2989 & ~n2991;
  assign n2993 = ~n2983 & n2992;
  assign n2994 = ~n2979 & ~n2992;
  assign n2995 = ~n2982 & n2994;
  assign n2996 = ~n2993 & ~n2995;
  assign n2997 = ~n2887 & ~n2900;
  assign n2998 = ~n2996 & n2997;
  assign n2999 = n2996 & ~n2997;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = pi55 & ~n2661;
  assign n3002 = ~n2659 & n3001;
  assign n3003 = n2668 & n3002;
  assign n3004 = ~n2907 & ~n3003;
  assign n3005 = n3000 & ~n3004;
  assign n3006 = ~n3000 & n3004;
  assign n3007 = ~n2834 & ~n2846;
  assign n3008 = n2835 & ~n2837;
  assign n3009 = ~n2839 & ~n3008;
  assign n3010 = ~n3007 & ~n3009;
  assign n3011 = ~n3006 & n3010;
  assign n3012 = ~n3005 & n3011;
  assign n3013 = ~n3005 & ~n3006;
  assign n3014 = ~n3010 & ~n3013;
  assign n3015 = ~n3012 & ~n3014;
  assign n3016 = n2957 & n3015;
  assign n3017 = ~n2957 & ~n3015;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~n2761 & n2793;
  assign n3020 = ~n2760 & ~n3019;
  assign n3021 = pi06 & ~n1607;
  assign n3022 = ~n1608 & n3021;
  assign n3023 = ~n1782 & n3022;
  assign n3024 = pi07 & ~n1609;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = pi49 & ~n3025;
  assign n3027 = ~pi49 & ~n3024;
  assign n3028 = ~n3023 & n3027;
  assign n3029 = ~n3026 & ~n3028;
  assign n3030 = pi08 & ~n1212;
  assign n3031 = ~n1213 & n3030;
  assign n3032 = ~n1425 & n3031;
  assign n3033 = pi09 & ~n1214;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = pi47 & ~n3034;
  assign n3036 = ~pi47 & ~n3033;
  assign n3037 = ~n3032 & n3036;
  assign n3038 = ~n3035 & ~n3037;
  assign n3039 = n3029 & ~n3038;
  assign n3040 = pi10 & ~n1006;
  assign n3041 = ~n1007 & n3040;
  assign n3042 = ~n1068 & n3041;
  assign n3043 = pi11 & ~n1008;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = pi45 & ~n3044;
  assign n3046 = ~pi45 & ~n3043;
  assign n3047 = ~n3042 & n3046;
  assign n3048 = ~n3045 & ~n3047;
  assign n3049 = ~n3029 & n3038;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = ~n3039 & n3050;
  assign n3052 = ~n3039 & ~n3049;
  assign n3053 = n3048 & ~n3052;
  assign n3054 = ~n3051 & ~n3053;
  assign n3055 = ~n2745 & n2755;
  assign n3056 = ~n2742 & ~n3055;
  assign n3057 = ~n2821 & n2831;
  assign n3058 = ~n2818 & ~n3057;
  assign n3059 = ~n3056 & n3058;
  assign n3060 = ~n3054 & n3059;
  assign n3061 = n3056 & ~n3058;
  assign n3062 = ~n3054 & n3061;
  assign n3063 = ~n3060 & ~n3062;
  assign n3064 = ~n3056 & ~n3058;
  assign n3065 = n3054 & n3064;
  assign n3066 = ~n2742 & ~n2818;
  assign n3067 = ~n3055 & n3066;
  assign n3068 = ~n3057 & n3067;
  assign n3069 = n3054 & n3068;
  assign n3070 = ~n3065 & ~n3069;
  assign n3071 = n3063 & n3070;
  assign n3072 = ~n3020 & ~n3071;
  assign n3073 = ~n3062 & ~n3065;
  assign n3074 = ~n3069 & n3073;
  assign n3075 = ~n2760 & ~n3060;
  assign n3076 = ~n3019 & n3075;
  assign n3077 = n3074 & n3076;
  assign n3078 = pi18 & ~n193;
  assign n3079 = ~n194 & n3078;
  assign n3080 = ~n729 & n3079;
  assign n3081 = pi19 & ~n195;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = pi37 & ~n3082;
  assign n3084 = ~pi37 & ~n3081;
  assign n3085 = ~n3080 & n3084;
  assign n3086 = ~n3083 & ~n3085;
  assign n3087 = pi20 & ~n141;
  assign n3088 = ~n142 & n3087;
  assign n3089 = ~n156 & n3088;
  assign n3090 = pi21 & ~n143;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = pi35 & ~n3091;
  assign n3093 = ~pi35 & ~n3090;
  assign n3094 = ~n3089 & n3093;
  assign n3095 = ~n3092 & ~n3094;
  assign n3096 = n3086 & ~n3095;
  assign n3097 = ~n3086 & n3095;
  assign n3098 = pi22 & ~pi32;
  assign n3099 = pi23 & pi32;
  assign n3100 = pi33 & ~n3099;
  assign n3101 = ~n3098 & n3100;
  assign n3102 = ~pi33 & n3099;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n3097 & n3103;
  assign n3105 = ~n3096 & n3104;
  assign n3106 = ~n3096 & ~n3097;
  assign n3107 = ~n3103 & ~n3106;
  assign n3108 = ~n3105 & ~n3107;
  assign n3109 = pi12 & ~n683;
  assign n3110 = ~n684 & n3109;
  assign n3111 = ~n1231 & n3110;
  assign n3112 = pi13 & ~n685;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = pi43 & ~n3113;
  assign n3115 = ~pi43 & ~n3112;
  assign n3116 = ~n3111 & n3115;
  assign n3117 = ~n3114 & ~n3116;
  assign n3118 = pi14 & ~n489;
  assign n3119 = ~n490 & n3118;
  assign n3120 = ~n572 & n3119;
  assign n3121 = pi15 & ~n491;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = pi41 & ~n3122;
  assign n3124 = ~pi41 & ~n3121;
  assign n3125 = ~n3120 & n3124;
  assign n3126 = ~n3123 & ~n3125;
  assign n3127 = n3117 & ~n3126;
  assign n3128 = pi16 & ~n304;
  assign n3129 = ~n305 & n3128;
  assign n3130 = ~n394 & n3129;
  assign n3131 = pi17 & ~n306;
  assign n3132 = ~n3130 & ~n3131;
  assign n3133 = pi39 & ~n3132;
  assign n3134 = ~pi39 & ~n3131;
  assign n3135 = ~n3130 & n3134;
  assign n3136 = ~n3133 & ~n3135;
  assign n3137 = ~n3117 & n3126;
  assign n3138 = ~n3136 & ~n3137;
  assign n3139 = ~n3127 & n3138;
  assign n3140 = ~n3127 & ~n3137;
  assign n3141 = n3136 & ~n3140;
  assign n3142 = ~n3139 & ~n3141;
  assign n3143 = ~n2770 & ~n2779;
  assign n3144 = ~n2777 & n3143;
  assign n3145 = ~n2768 & n3144;
  assign n3146 = ~n2790 & ~n3145;
  assign n3147 = ~n3142 & n3146;
  assign n3148 = n3142 & ~n3146;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = ~n3108 & ~n3149;
  assign n3151 = n3108 & ~n3147;
  assign n3152 = ~n3148 & n3151;
  assign n3153 = ~n3150 & ~n3152;
  assign n3154 = ~n3077 & n3153;
  assign n3155 = ~n3072 & n3154;
  assign n3156 = ~n3072 & ~n3077;
  assign n3157 = ~n3153 & ~n3156;
  assign n3158 = ~n3155 & ~n3157;
  assign n3159 = ~n3018 & n3158;
  assign n3160 = n3018 & ~n3158;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = ~n2865 & ~n2925;
  assign n3163 = n2676 & ~n2910;
  assign n3164 = ~n2907 & n3163;
  assign n3165 = ~n2922 & ~n3164;
  assign n3166 = ~n2924 & ~n3165;
  assign n3167 = ~n3162 & n3166;
  assign n3168 = ~n2924 & ~n3162;
  assign n3169 = n3165 & ~n3168;
  assign n3170 = ~n3167 & ~n3169;
  assign n3171 = ~n3161 & ~n3170;
  assign n3172 = n3161 & n3170;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n2930 & ~n2935;
  assign n3175 = ~n2933 & ~n3174;
  assign n3176 = ~n3173 & n3175;
  assign n3177 = n3173 & ~n3175;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = n2942 & n3178;
  assign n3180 = ~n2942 & ~n3178;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~n2944 & ~n3181;
  assign n3183 = ~n2954 & n3182;
  assign n3184 = ~n2944 & ~n2954;
  assign n3185 = n3181 & ~n3184;
  assign po23 = ~n3183 & ~n3185;
  assign n3187 = n2710 & ~n3180;
  assign n3188 = ~n2474 & ~n2946;
  assign n3189 = ~n2944 & n3188;
  assign n3190 = n3187 & n3189;
  assign n3191 = ~n2270 & n3190;
  assign n3192 = n2479 & ~n2707;
  assign n3193 = ~n2709 & n3192;
  assign n3194 = n3188 & n3193;
  assign n3195 = ~n2944 & ~n2950;
  assign n3196 = ~n2946 & ~n3195;
  assign n3197 = ~n3194 & ~n3196;
  assign n3198 = ~n3180 & ~n3197;
  assign n3199 = ~n3179 & ~n3198;
  assign n3200 = ~n3191 & n3199;
  assign n3201 = ~n3165 & ~n3168;
  assign n3202 = ~n3171 & ~n3201;
  assign n3203 = ~n3072 & ~n3155;
  assign n3204 = ~n2982 & n2992;
  assign n3205 = pi55 & ~pi56;
  assign n3206 = ~pi55 & pi56;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = pi00 & ~n3207;
  assign n3209 = pi57 & ~n3208;
  assign n3210 = pi00 & ~pi57;
  assign n3211 = ~n3207 & n3210;
  assign n3212 = ~n3209 & ~n3211;
  assign n3213 = ~n2979 & ~n3212;
  assign n3214 = ~n3204 & n3213;
  assign n3215 = ~n2979 & ~n3204;
  assign n3216 = n3212 & ~n3215;
  assign n3217 = ~n3214 & ~n3216;
  assign n3218 = pi01 & ~n2876;
  assign n3219 = ~n2877 & n3218;
  assign n3220 = ~n2960 & n3219;
  assign n3221 = pi02 & ~n2878;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = pi55 & ~n3222;
  assign n3224 = pi03 & ~n2288;
  assign n3225 = ~n2289 & n3224;
  assign n3226 = ~n2647 & n3225;
  assign n3227 = pi04 & ~n2290;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = pi53 & ~n3228;
  assign n3230 = ~pi53 & ~n3227;
  assign n3231 = ~n3226 & n3230;
  assign n3232 = ~pi55 & ~n3221;
  assign n3233 = ~n3220 & n3232;
  assign n3234 = ~n3231 & ~n3233;
  assign n3235 = ~n3229 & n3234;
  assign n3236 = ~n3223 & n3235;
  assign n3237 = ~n3229 & ~n3231;
  assign n3238 = ~n3223 & ~n3233;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = ~n3236 & ~n3239;
  assign n3241 = pi05 & ~n2023;
  assign n3242 = ~n2024 & n3241;
  assign n3243 = ~n2079 & n3242;
  assign n3244 = pi06 & ~n2025;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = pi51 & ~n3245;
  assign n3247 = ~pi51 & ~n3244;
  assign n3248 = ~n3243 & n3247;
  assign n3249 = ~n3246 & ~n3248;
  assign n3250 = ~n3240 & n3249;
  assign n3251 = ~n3236 & ~n3249;
  assign n3252 = ~n3239 & n3251;
  assign n3253 = ~n3250 & ~n3252;
  assign n3254 = ~n3217 & n3253;
  assign n3255 = n3217 & ~n3253;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = n2998 & ~n3256;
  assign n3258 = ~n2998 & ~n3254;
  assign n3259 = ~n3255 & n3258;
  assign n3260 = ~n3257 & ~n3259;
  assign n3261 = n3054 & ~n3058;
  assign n3262 = ~n3054 & n3058;
  assign n3263 = ~n3056 & ~n3262;
  assign n3264 = ~n3261 & ~n3263;
  assign n3265 = ~n3260 & n3264;
  assign n3266 = ~n3257 & ~n3264;
  assign n3267 = ~n3259 & n3266;
  assign n3268 = ~n3265 & ~n3267;
  assign n3269 = n3203 & ~n3268;
  assign n3270 = ~n3085 & ~n3094;
  assign n3271 = ~n3092 & n3270;
  assign n3272 = ~n3083 & n3271;
  assign n3273 = ~n3107 & ~n3272;
  assign n3274 = pi13 & ~n683;
  assign n3275 = ~n684 & n3274;
  assign n3276 = ~n1231 & n3275;
  assign n3277 = pi14 & ~n685;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = pi43 & ~n3278;
  assign n3280 = pi15 & ~n489;
  assign n3281 = ~n490 & n3280;
  assign n3282 = ~n572 & n3281;
  assign n3283 = pi16 & ~n491;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = pi41 & ~n3284;
  assign n3286 = ~pi41 & ~n3283;
  assign n3287 = ~n3282 & n3286;
  assign n3288 = ~pi43 & ~n3277;
  assign n3289 = ~n3276 & n3288;
  assign n3290 = ~n3287 & ~n3289;
  assign n3291 = ~n3285 & n3290;
  assign n3292 = ~n3279 & n3291;
  assign n3293 = ~n3285 & ~n3287;
  assign n3294 = ~n3279 & ~n3289;
  assign n3295 = ~n3293 & ~n3294;
  assign n3296 = ~n3292 & ~n3295;
  assign n3297 = pi17 & ~n304;
  assign n3298 = ~n305 & n3297;
  assign n3299 = ~n394 & n3298;
  assign n3300 = pi18 & ~n306;
  assign n3301 = ~n3299 & ~n3300;
  assign n3302 = pi39 & ~n3301;
  assign n3303 = ~pi39 & ~n3300;
  assign n3304 = ~n3299 & n3303;
  assign n3305 = ~n3302 & ~n3304;
  assign n3306 = ~n3296 & n3305;
  assign n3307 = ~n3292 & ~n3305;
  assign n3308 = ~n3295 & n3307;
  assign n3309 = ~n3306 & ~n3308;
  assign n3310 = ~n3273 & ~n3309;
  assign n3311 = n3273 & n3309;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = pi19 & ~n193;
  assign n3314 = ~n194 & n3313;
  assign n3315 = ~n729 & n3314;
  assign n3316 = pi20 & ~n195;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = pi37 & ~n3317;
  assign n3319 = ~pi37 & ~n3316;
  assign n3320 = ~n3315 & n3319;
  assign n3321 = ~n3318 & ~n3320;
  assign n3322 = pi21 & ~n141;
  assign n3323 = ~n142 & n3322;
  assign n3324 = ~n156 & n3323;
  assign n3325 = pi22 & ~n143;
  assign n3326 = ~n3324 & ~n3325;
  assign n3327 = pi35 & ~n3326;
  assign n3328 = ~pi35 & ~n3325;
  assign n3329 = ~n3324 & n3328;
  assign n3330 = ~n3327 & ~n3329;
  assign n3331 = n3321 & ~n3330;
  assign n3332 = ~n3321 & n3330;
  assign n3333 = pi23 & ~pi32;
  assign n3334 = pi24 & pi32;
  assign n3335 = pi33 & ~n3334;
  assign n3336 = ~n3333 & n3335;
  assign n3337 = ~pi33 & n3334;
  assign n3338 = ~n3336 & ~n3337;
  assign n3339 = ~n3332 & n3338;
  assign n3340 = ~n3331 & n3339;
  assign n3341 = ~n3331 & ~n3332;
  assign n3342 = ~n3338 & ~n3341;
  assign n3343 = ~n3340 & ~n3342;
  assign n3344 = ~n3312 & n3343;
  assign n3345 = ~n3310 & ~n3343;
  assign n3346 = ~n3311 & n3345;
  assign n3347 = ~n3344 & ~n3346;
  assign n3348 = ~n3148 & ~n3152;
  assign n3349 = ~n3028 & ~n3037;
  assign n3350 = ~n3035 & n3349;
  assign n3351 = ~n3026 & n3350;
  assign n3352 = ~n3053 & ~n3351;
  assign n3353 = pi07 & ~n1607;
  assign n3354 = ~n1608 & n3353;
  assign n3355 = ~n1782 & n3354;
  assign n3356 = pi08 & ~n1609;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = pi49 & ~n3357;
  assign n3359 = pi09 & ~n1212;
  assign n3360 = ~n1213 & n3359;
  assign n3361 = ~n1425 & n3360;
  assign n3362 = pi10 & ~n1214;
  assign n3363 = ~n3361 & ~n3362;
  assign n3364 = pi47 & ~n3363;
  assign n3365 = ~pi47 & ~n3362;
  assign n3366 = ~n3361 & n3365;
  assign n3367 = ~pi49 & ~n3356;
  assign n3368 = ~n3355 & n3367;
  assign n3369 = ~n3366 & ~n3368;
  assign n3370 = ~n3364 & n3369;
  assign n3371 = ~n3358 & n3370;
  assign n3372 = ~n3364 & ~n3366;
  assign n3373 = ~n3358 & ~n3368;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = ~n3371 & ~n3374;
  assign n3376 = pi11 & ~n1006;
  assign n3377 = ~n1007 & n3376;
  assign n3378 = ~n1068 & n3377;
  assign n3379 = pi12 & ~n1008;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = pi45 & ~n3380;
  assign n3382 = ~pi45 & ~n3379;
  assign n3383 = ~n3378 & n3382;
  assign n3384 = ~n3381 & ~n3383;
  assign n3385 = ~n3375 & n3384;
  assign n3386 = ~n3371 & ~n3384;
  assign n3387 = ~n3374 & n3386;
  assign n3388 = ~n3385 & ~n3387;
  assign n3389 = n3352 & n3388;
  assign n3390 = ~n3352 & ~n3388;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = ~n3116 & ~n3125;
  assign n3393 = ~n3123 & n3392;
  assign n3394 = ~n3114 & n3393;
  assign n3395 = ~n3141 & ~n3394;
  assign n3396 = ~n3391 & n3395;
  assign n3397 = ~n3389 & ~n3395;
  assign n3398 = ~n3390 & n3397;
  assign n3399 = ~n3396 & ~n3398;
  assign n3400 = ~n3348 & n3399;
  assign n3401 = n3348 & ~n3399;
  assign n3402 = ~n3400 & ~n3401;
  assign n3403 = ~n3347 & ~n3402;
  assign n3404 = n3347 & ~n3400;
  assign n3405 = ~n3401 & n3404;
  assign n3406 = ~n3403 & ~n3405;
  assign n3407 = ~n3203 & n3268;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = ~n3269 & n3408;
  assign n3410 = ~n3269 & ~n3407;
  assign n3411 = n3406 & ~n3410;
  assign n3412 = ~n3409 & ~n3411;
  assign n3413 = ~n3017 & ~n3158;
  assign n3414 = ~n3006 & ~n3012;
  assign n3415 = ~pi57 & ~n3414;
  assign n3416 = pi57 & ~n3006;
  assign n3417 = ~n3012 & n3416;
  assign n3418 = ~n3016 & ~n3417;
  assign n3419 = ~n3415 & n3418;
  assign n3420 = ~n3413 & n3419;
  assign n3421 = ~n3415 & ~n3417;
  assign n3422 = ~n3016 & ~n3413;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = ~n3420 & ~n3423;
  assign n3425 = n3412 & n3424;
  assign n3426 = ~n3412 & ~n3424;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = n3202 & ~n3427;
  assign n3429 = ~n3202 & n3427;
  assign n3430 = n3177 & ~n3429;
  assign n3431 = ~n3428 & n3430;
  assign n3432 = ~n3428 & ~n3429;
  assign n3433 = ~n3177 & ~n3432;
  assign n3434 = ~n3431 & ~n3433;
  assign n3435 = ~n3200 & n3434;
  assign n3436 = ~n3179 & ~n3434;
  assign n3437 = ~n3198 & n3436;
  assign n3438 = ~n3191 & n3437;
  assign po24 = ~n3435 & ~n3438;
  assign n3440 = ~n2051 & ~n2058;
  assign n3441 = ~n2061 & n3440;
  assign n3442 = ~n3180 & ~n3431;
  assign n3443 = ~n3433 & n3442;
  assign n3444 = n2260 & ~n2707;
  assign n3445 = ~n2709 & ~n3179;
  assign n3446 = n3444 & n3445;
  assign n3447 = n3443 & n3446;
  assign n3448 = n3189 & n3447;
  assign n3449 = ~n3441 & n3448;
  assign n3450 = ~n3177 & ~n3179;
  assign n3451 = n3432 & ~n3450;
  assign n3452 = n3181 & n3434;
  assign n3453 = ~n3197 & n3452;
  assign n3454 = ~n3451 & ~n3453;
  assign n3455 = ~n3449 & n3454;
  assign n3456 = ~n3347 & ~n3401;
  assign n3457 = ~n3400 & ~n3456;
  assign n3458 = ~n2979 & n3212;
  assign n3459 = ~n3204 & n3458;
  assign n3460 = ~n3254 & ~n3459;
  assign n3461 = pi56 & ~pi57;
  assign n3462 = ~pi56 & pi57;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = pi00 & ~n3205;
  assign n3465 = ~n3206 & n3464;
  assign n3466 = ~n3463 & n3465;
  assign n3467 = pi01 & ~n3207;
  assign n3468 = ~n3466 & ~n3467;
  assign n3469 = pi57 & ~n3468;
  assign n3470 = ~pi57 & ~n3467;
  assign n3471 = ~n3466 & n3470;
  assign n3472 = ~n3469 & ~n3471;
  assign n3473 = ~n3239 & n3249;
  assign n3474 = ~n3236 & ~n3473;
  assign n3475 = n3472 & ~n3474;
  assign n3476 = pi02 & ~n2876;
  assign n3477 = ~n2877 & n3476;
  assign n3478 = ~n2960 & n3477;
  assign n3479 = pi03 & ~n2878;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = pi55 & ~n3480;
  assign n3482 = pi04 & ~n2288;
  assign n3483 = ~n2289 & n3482;
  assign n3484 = ~n2647 & n3483;
  assign n3485 = pi05 & ~n2290;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = pi53 & ~n3486;
  assign n3488 = ~pi53 & ~n3485;
  assign n3489 = ~n3484 & n3488;
  assign n3490 = ~pi55 & ~n3479;
  assign n3491 = ~n3478 & n3490;
  assign n3492 = ~n3489 & ~n3491;
  assign n3493 = ~n3487 & n3492;
  assign n3494 = ~n3481 & n3493;
  assign n3495 = ~n3487 & ~n3489;
  assign n3496 = ~n3481 & ~n3491;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = ~n3494 & ~n3497;
  assign n3499 = pi06 & ~n2023;
  assign n3500 = ~n2024 & n3499;
  assign n3501 = ~n2079 & n3500;
  assign n3502 = pi07 & ~n2025;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = pi51 & ~n3503;
  assign n3505 = ~pi51 & ~n3502;
  assign n3506 = ~n3501 & n3505;
  assign n3507 = ~n3504 & ~n3506;
  assign n3508 = ~n3498 & n3507;
  assign n3509 = ~n3494 & ~n3507;
  assign n3510 = ~n3497 & n3509;
  assign n3511 = ~n3508 & ~n3510;
  assign n3512 = ~n3236 & ~n3472;
  assign n3513 = ~n3473 & n3512;
  assign n3514 = ~n3511 & ~n3513;
  assign n3515 = ~n3475 & n3514;
  assign n3516 = ~n3475 & ~n3513;
  assign n3517 = n3511 & ~n3516;
  assign n3518 = ~n3515 & ~n3517;
  assign n3519 = n3460 & ~n3518;
  assign n3520 = ~n3460 & n3518;
  assign n3521 = ~n3390 & ~n3398;
  assign n3522 = ~n3520 & n3521;
  assign n3523 = ~n3519 & n3522;
  assign n3524 = ~n3519 & ~n3520;
  assign n3525 = ~n3521 & ~n3524;
  assign n3526 = ~n3523 & ~n3525;
  assign n3527 = ~n3457 & n3526;
  assign n3528 = n3457 & ~n3526;
  assign n3529 = ~n3527 & ~n3528;
  assign n3530 = ~n3311 & n3343;
  assign n3531 = ~n3310 & ~n3530;
  assign n3532 = pi08 & ~n1607;
  assign n3533 = ~n1608 & n3532;
  assign n3534 = ~n1782 & n3533;
  assign n3535 = pi09 & ~n1609;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = pi49 & ~n3536;
  assign n3538 = pi10 & ~n1212;
  assign n3539 = ~n1213 & n3538;
  assign n3540 = ~n1425 & n3539;
  assign n3541 = pi11 & ~n1214;
  assign n3542 = ~n3540 & ~n3541;
  assign n3543 = pi47 & ~n3542;
  assign n3544 = ~pi47 & ~n3541;
  assign n3545 = ~n3540 & n3544;
  assign n3546 = ~pi49 & ~n3535;
  assign n3547 = ~n3534 & n3546;
  assign n3548 = ~n3545 & ~n3547;
  assign n3549 = ~n3543 & n3548;
  assign n3550 = ~n3537 & n3549;
  assign n3551 = ~n3543 & ~n3545;
  assign n3552 = ~n3537 & ~n3547;
  assign n3553 = ~n3551 & ~n3552;
  assign n3554 = ~n3550 & ~n3553;
  assign n3555 = pi12 & ~n1006;
  assign n3556 = ~n1007 & n3555;
  assign n3557 = ~n1068 & n3556;
  assign n3558 = pi13 & ~n1008;
  assign n3559 = ~n3557 & ~n3558;
  assign n3560 = pi45 & ~n3559;
  assign n3561 = ~pi45 & ~n3558;
  assign n3562 = ~n3557 & n3561;
  assign n3563 = ~n3560 & ~n3562;
  assign n3564 = ~n3554 & n3563;
  assign n3565 = ~n3374 & n3384;
  assign n3566 = ~n3371 & ~n3565;
  assign n3567 = ~n3564 & n3566;
  assign n3568 = ~n3550 & ~n3563;
  assign n3569 = ~n3553 & n3568;
  assign n3570 = ~n3295 & n3305;
  assign n3571 = ~n3292 & ~n3570;
  assign n3572 = ~n3569 & ~n3571;
  assign n3573 = n3567 & n3572;
  assign n3574 = ~n3564 & n3571;
  assign n3575 = ~n3566 & ~n3569;
  assign n3576 = n3574 & n3575;
  assign n3577 = ~n3573 & ~n3576;
  assign n3578 = ~n3564 & ~n3569;
  assign n3579 = ~n3566 & ~n3571;
  assign n3580 = ~n3578 & n3579;
  assign n3581 = ~n3292 & ~n3371;
  assign n3582 = ~n3570 & n3581;
  assign n3583 = ~n3565 & n3582;
  assign n3584 = ~n3578 & n3583;
  assign n3585 = ~n3580 & ~n3584;
  assign n3586 = n3577 & n3585;
  assign n3587 = ~n3531 & ~n3586;
  assign n3588 = ~n3320 & ~n3329;
  assign n3589 = ~n3327 & n3588;
  assign n3590 = ~n3318 & n3589;
  assign n3591 = ~n3342 & ~n3590;
  assign n3592 = pi14 & ~n683;
  assign n3593 = ~n684 & n3592;
  assign n3594 = ~n1231 & n3593;
  assign n3595 = pi15 & ~n685;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = pi43 & ~n3596;
  assign n3598 = ~pi43 & ~n3595;
  assign n3599 = ~n3594 & n3598;
  assign n3600 = ~n3597 & ~n3599;
  assign n3601 = pi16 & ~n489;
  assign n3602 = ~n490 & n3601;
  assign n3603 = ~n572 & n3602;
  assign n3604 = pi17 & ~n491;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = pi41 & ~n3605;
  assign n3607 = ~pi41 & ~n3604;
  assign n3608 = ~n3603 & n3607;
  assign n3609 = ~n3606 & ~n3608;
  assign n3610 = ~n3600 & n3609;
  assign n3611 = n3600 & ~n3609;
  assign n3612 = ~n3610 & ~n3611;
  assign n3613 = pi18 & ~n304;
  assign n3614 = ~n305 & n3613;
  assign n3615 = ~n394 & n3614;
  assign n3616 = pi19 & ~n306;
  assign n3617 = ~n3615 & ~n3616;
  assign n3618 = pi39 & ~n3617;
  assign n3619 = ~pi39 & ~n3616;
  assign n3620 = ~n3615 & n3619;
  assign n3621 = ~n3618 & ~n3620;
  assign n3622 = ~n3612 & n3621;
  assign n3623 = ~n3610 & ~n3621;
  assign n3624 = ~n3611 & n3623;
  assign n3625 = ~n3622 & ~n3624;
  assign n3626 = ~n3591 & n3625;
  assign n3627 = n3591 & ~n3625;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = pi22 & ~n141;
  assign n3630 = ~n142 & n3629;
  assign n3631 = ~n156 & n3630;
  assign n3632 = pi23 & ~n143;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = pi35 & ~n3633;
  assign n3635 = ~pi35 & ~n3632;
  assign n3636 = ~n3631 & n3635;
  assign n3637 = ~n3634 & ~n3636;
  assign n3638 = pi20 & ~n193;
  assign n3639 = ~n194 & n3638;
  assign n3640 = ~n729 & n3639;
  assign n3641 = pi21 & ~n195;
  assign n3642 = ~n3640 & ~n3641;
  assign n3643 = pi37 & ~n3642;
  assign n3644 = ~pi37 & ~n3641;
  assign n3645 = ~n3640 & n3644;
  assign n3646 = ~n3643 & ~n3645;
  assign n3647 = ~n3637 & ~n3646;
  assign n3648 = ~n3636 & ~n3645;
  assign n3649 = ~n3634 & n3648;
  assign n3650 = ~n3643 & n3649;
  assign n3651 = pi24 & ~pi32;
  assign n3652 = pi25 & pi32;
  assign n3653 = pi33 & ~n3652;
  assign n3654 = ~n3651 & n3653;
  assign n3655 = ~pi33 & n3652;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = ~n3650 & ~n3656;
  assign n3658 = ~n3647 & n3657;
  assign n3659 = ~n3647 & ~n3650;
  assign n3660 = n3656 & ~n3659;
  assign n3661 = ~n3658 & ~n3660;
  assign n3662 = ~n3628 & n3661;
  assign n3663 = ~n3626 & ~n3661;
  assign n3664 = ~n3627 & n3663;
  assign n3665 = ~n3662 & ~n3664;
  assign n3666 = ~n3576 & ~n3580;
  assign n3667 = ~n3584 & n3666;
  assign n3668 = ~n3310 & ~n3573;
  assign n3669 = ~n3530 & n3668;
  assign n3670 = n3667 & n3669;
  assign n3671 = ~n3665 & ~n3670;
  assign n3672 = ~n3587 & n3671;
  assign n3673 = ~n3587 & ~n3670;
  assign n3674 = n3665 & ~n3673;
  assign n3675 = ~n3672 & ~n3674;
  assign n3676 = ~n3529 & n3675;
  assign n3677 = ~n3527 & ~n3675;
  assign n3678 = ~n3528 & n3677;
  assign n3679 = ~n3676 & ~n3678;
  assign n3680 = ~n3257 & ~n3267;
  assign n3681 = ~n3406 & ~n3680;
  assign n3682 = n3410 & n3681;
  assign n3683 = n3407 & ~n3680;
  assign n3684 = ~n3682 & ~n3683;
  assign n3685 = ~n3407 & n3680;
  assign n3686 = ~n3410 & n3685;
  assign n3687 = ~n3403 & n3680;
  assign n3688 = ~n3405 & n3687;
  assign n3689 = ~n3407 & n3688;
  assign n3690 = ~n3686 & ~n3689;
  assign n3691 = n3684 & n3690;
  assign n3692 = ~n3679 & ~n3691;
  assign n3693 = n3679 & n3691;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = ~n3417 & ~n3420;
  assign n3696 = ~n3425 & n3695;
  assign n3697 = ~n3409 & n3417;
  assign n3698 = ~n3411 & ~n3420;
  assign n3699 = ~n3423 & n3698;
  assign n3700 = n3697 & n3699;
  assign n3701 = ~n3696 & ~n3700;
  assign n3702 = n3694 & ~n3701;
  assign n3703 = ~n3694 & n3701;
  assign n3704 = n3429 & ~n3703;
  assign n3705 = ~n3702 & n3704;
  assign n3706 = ~n3702 & ~n3703;
  assign n3707 = ~n3429 & ~n3706;
  assign n3708 = ~n3705 & ~n3707;
  assign n3709 = ~n3455 & n3708;
  assign n3710 = ~n3451 & ~n3708;
  assign n3711 = ~n3453 & n3710;
  assign n3712 = ~n3449 & n3711;
  assign po25 = ~n3709 & ~n3712;
  assign n3714 = ~n2267 & ~n2479;
  assign n3715 = ~n2269 & n3714;
  assign n3716 = n2947 & n3708;
  assign n3717 = n2716 & n3452;
  assign n3718 = n3716 & n3717;
  assign n3719 = ~n3715 & n3718;
  assign n3720 = n2944 & n3452;
  assign n3721 = ~n3451 & ~n3705;
  assign n3722 = ~n3720 & n3721;
  assign n3723 = ~n3707 & ~n3722;
  assign n3724 = ~n2946 & ~n3705;
  assign n3725 = ~n3707 & n3724;
  assign n3726 = ~n2944 & n2950;
  assign n3727 = n3452 & n3726;
  assign n3728 = n3725 & n3727;
  assign n3729 = ~n3407 & ~n3409;
  assign n3730 = ~n3680 & ~n3729;
  assign n3731 = ~n3679 & n3691;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = ~n3647 & ~n3656;
  assign n3734 = ~n3650 & ~n3733;
  assign n3735 = pi18 & ~n491;
  assign n3736 = pi17 & pi39;
  assign n3737 = n570 & n3736;
  assign n3738 = pi17 & ~pi39;
  assign n3739 = n571 & n3738;
  assign n3740 = ~n3737 & ~n3739;
  assign n3741 = ~n3735 & n3740;
  assign n3742 = pi41 & ~n3741;
  assign n3743 = ~pi41 & ~n3737;
  assign n3744 = ~n3739 & n3743;
  assign n3745 = ~n3735 & n3744;
  assign n3746 = ~n3742 & ~n3745;
  assign n3747 = pi16 & ~n685;
  assign n3748 = pi15 & pi41;
  assign n3749 = n923 & n3748;
  assign n3750 = pi15 & ~pi41;
  assign n3751 = n801 & n3750;
  assign n3752 = ~n3749 & ~n3751;
  assign n3753 = ~n3747 & n3752;
  assign n3754 = pi43 & ~n3753;
  assign n3755 = ~pi43 & ~n3749;
  assign n3756 = ~n3751 & n3755;
  assign n3757 = ~n3747 & n3756;
  assign n3758 = ~n3754 & ~n3757;
  assign n3759 = n3746 & n3758;
  assign n3760 = ~n3746 & ~n3758;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = pi19 & ~n304;
  assign n3763 = ~n305 & n3762;
  assign n3764 = ~n394 & n3763;
  assign n3765 = pi20 & ~n306;
  assign n3766 = ~n3764 & ~n3765;
  assign n3767 = pi39 & ~n3766;
  assign n3768 = ~pi39 & ~n3765;
  assign n3769 = ~n3764 & n3768;
  assign n3770 = ~n3767 & ~n3769;
  assign n3771 = ~n3761 & n3770;
  assign n3772 = n3761 & ~n3770;
  assign n3773 = ~n3771 & ~n3772;
  assign n3774 = ~n3734 & ~n3773;
  assign n3775 = n3734 & n3773;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = pi22 & ~n195;
  assign n3778 = pi21 & pi35;
  assign n3779 = n341 & n3778;
  assign n3780 = pi21 & ~pi35;
  assign n3781 = n259 & n3780;
  assign n3782 = ~n3779 & ~n3781;
  assign n3783 = ~n3777 & n3782;
  assign n3784 = pi37 & ~n3783;
  assign n3785 = ~pi37 & ~n3779;
  assign n3786 = ~n3781 & n3785;
  assign n3787 = ~n3777 & n3786;
  assign n3788 = ~n3784 & ~n3787;
  assign n3789 = pi24 & ~n143;
  assign n3790 = pi23 & pi33;
  assign n3791 = n154 & n3790;
  assign n3792 = pi23 & ~pi33;
  assign n3793 = n155 & n3792;
  assign n3794 = ~n3791 & ~n3793;
  assign n3795 = ~n3789 & n3794;
  assign n3796 = pi35 & ~n3795;
  assign n3797 = ~pi35 & ~n3791;
  assign n3798 = ~n3793 & n3797;
  assign n3799 = ~n3789 & n3798;
  assign n3800 = ~n3796 & ~n3799;
  assign n3801 = n3788 & ~n3800;
  assign n3802 = ~n3788 & n3800;
  assign n3803 = pi25 & ~pi32;
  assign n3804 = pi26 & pi32;
  assign n3805 = pi33 & ~n3804;
  assign n3806 = ~n3803 & n3805;
  assign n3807 = ~pi33 & n3804;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = ~n3802 & n3808;
  assign n3810 = ~n3801 & n3809;
  assign n3811 = ~n3801 & ~n3802;
  assign n3812 = ~n3808 & ~n3811;
  assign n3813 = ~n3810 & ~n3812;
  assign n3814 = ~n3776 & n3813;
  assign n3815 = ~n3774 & ~n3813;
  assign n3816 = ~n3775 & n3815;
  assign n3817 = ~n3814 & ~n3816;
  assign n3818 = ~n3627 & n3661;
  assign n3819 = ~n3626 & ~n3818;
  assign n3820 = ~n3553 & n3563;
  assign n3821 = ~n3550 & ~n3820;
  assign n3822 = pi12 & ~n1214;
  assign n3823 = pi11 & pi45;
  assign n3824 = n1423 & n3823;
  assign n3825 = pi11 & ~pi45;
  assign n3826 = n1424 & n3825;
  assign n3827 = ~n3824 & ~n3826;
  assign n3828 = ~n3822 & n3827;
  assign n3829 = pi47 & ~n3828;
  assign n3830 = ~pi47 & ~n3824;
  assign n3831 = ~n3826 & n3830;
  assign n3832 = ~n3822 & n3831;
  assign n3833 = ~n3829 & ~n3832;
  assign n3834 = pi10 & ~n1609;
  assign n3835 = pi09 & pi47;
  assign n3836 = n1780 & n3835;
  assign n3837 = pi09 & ~pi47;
  assign n3838 = n1781 & n3837;
  assign n3839 = ~n3836 & ~n3838;
  assign n3840 = ~n3834 & n3839;
  assign n3841 = pi49 & ~n3840;
  assign n3842 = ~pi49 & ~n3836;
  assign n3843 = ~n3838 & n3842;
  assign n3844 = ~n3834 & n3843;
  assign n3845 = ~n3841 & ~n3844;
  assign n3846 = n3833 & n3845;
  assign n3847 = ~n3833 & ~n3845;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = pi13 & ~n1006;
  assign n3850 = ~n1007 & n3849;
  assign n3851 = ~n1068 & n3850;
  assign n3852 = pi14 & ~n1008;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = pi45 & ~n3853;
  assign n3855 = ~pi45 & ~n3852;
  assign n3856 = ~n3851 & n3855;
  assign n3857 = ~n3854 & ~n3856;
  assign n3858 = ~n3848 & n3857;
  assign n3859 = n3848 & ~n3857;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = n3821 & n3860;
  assign n3862 = ~n3821 & ~n3860;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~n3599 & ~n3608;
  assign n3865 = ~n3606 & n3864;
  assign n3866 = ~n3597 & n3865;
  assign n3867 = ~n3622 & ~n3866;
  assign n3868 = ~n3863 & n3867;
  assign n3869 = n3863 & ~n3867;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = ~n3819 & n3870;
  assign n3872 = n3819 & ~n3870;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = ~n3817 & ~n3873;
  assign n3875 = n3817 & ~n3871;
  assign n3876 = ~n3872 & n3875;
  assign n3877 = ~n3874 & ~n3876;
  assign n3878 = ~n3587 & ~n3672;
  assign n3879 = pi06 & ~n2290;
  assign n3880 = pi05 & pi51;
  assign n3881 = n2645 & n3880;
  assign n3882 = pi05 & ~pi51;
  assign n3883 = n2646 & n3882;
  assign n3884 = ~n3881 & ~n3883;
  assign n3885 = ~n3879 & n3884;
  assign n3886 = pi53 & ~n3885;
  assign n3887 = ~pi53 & ~n3881;
  assign n3888 = ~n3883 & n3887;
  assign n3889 = ~n3879 & n3888;
  assign n3890 = ~n3886 & ~n3889;
  assign n3891 = pi04 & ~n2878;
  assign n3892 = pi03 & pi53;
  assign n3893 = n2958 & n3892;
  assign n3894 = pi03 & ~pi53;
  assign n3895 = n2959 & n3894;
  assign n3896 = ~n3893 & ~n3895;
  assign n3897 = ~n3891 & n3896;
  assign n3898 = pi55 & ~n3897;
  assign n3899 = ~pi55 & ~n3893;
  assign n3900 = ~n3895 & n3899;
  assign n3901 = ~n3891 & n3900;
  assign n3902 = ~n3898 & ~n3901;
  assign n3903 = n3890 & n3902;
  assign n3904 = ~n3890 & ~n3902;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = pi07 & ~n2023;
  assign n3907 = ~n2024 & n3906;
  assign n3908 = ~n2079 & n3907;
  assign n3909 = pi08 & ~n2025;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = pi51 & ~n3910;
  assign n3912 = ~pi51 & ~n3909;
  assign n3913 = ~n3908 & n3912;
  assign n3914 = ~n3911 & ~n3913;
  assign n3915 = ~n3905 & n3914;
  assign n3916 = n3905 & ~n3914;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = ~n3497 & n3507;
  assign n3919 = ~n3494 & ~n3918;
  assign n3920 = pi01 & ~n3205;
  assign n3921 = ~n3206 & n3920;
  assign n3922 = ~n3463 & n3921;
  assign n3923 = pi02 & ~n3207;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = pi57 & ~n3924;
  assign n3926 = ~pi57 & ~n3923;
  assign n3927 = ~n3922 & n3926;
  assign n3928 = ~n3925 & ~n3927;
  assign n3929 = ~n3919 & n3928;
  assign n3930 = ~n3494 & ~n3928;
  assign n3931 = ~n3918 & n3930;
  assign n3932 = ~n3929 & ~n3931;
  assign n3933 = ~n3917 & ~n3932;
  assign n3934 = n3917 & ~n3931;
  assign n3935 = ~n3929 & n3934;
  assign n3936 = ~n3475 & ~n3935;
  assign n3937 = ~n3515 & n3936;
  assign n3938 = ~n3933 & n3937;
  assign n3939 = ~n3475 & ~n3515;
  assign n3940 = ~n3933 & ~n3935;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3938 & ~n3941;
  assign n3943 = ~n3566 & ~n3578;
  assign n3944 = n3567 & ~n3569;
  assign n3945 = ~n3571 & ~n3944;
  assign n3946 = ~n3943 & ~n3945;
  assign n3947 = ~n3942 & n3946;
  assign n3948 = ~n3938 & ~n3946;
  assign n3949 = ~n3941 & n3948;
  assign n3950 = ~n3947 & ~n3949;
  assign n3951 = ~n3878 & n3950;
  assign n3952 = n3878 & ~n3950;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3877 & ~n3953;
  assign n3955 = n3877 & ~n3951;
  assign n3956 = ~n3952 & n3955;
  assign n3957 = ~n3954 & ~n3956;
  assign n3958 = n3460 & n3518;
  assign n3959 = pi57 & ~pi58;
  assign n3960 = ~pi57 & pi58;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = pi00 & ~n3961;
  assign n3963 = ~n3958 & ~n3962;
  assign n3964 = ~n3525 & n3963;
  assign n3965 = ~n3525 & ~n3958;
  assign n3966 = n3962 & ~n3965;
  assign n3967 = ~n3964 & ~n3966;
  assign n3968 = ~n3528 & n3675;
  assign n3969 = ~n3527 & ~n3968;
  assign n3970 = ~n3967 & n3969;
  assign n3971 = n3967 & ~n3969;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n3957 & ~n3972;
  assign n3974 = n3957 & ~n3970;
  assign n3975 = ~n3971 & n3974;
  assign n3976 = ~n3973 & ~n3975;
  assign n3977 = ~n3732 & ~n3976;
  assign n3978 = n3732 & n3976;
  assign n3979 = ~n3977 & ~n3978;
  assign n3980 = ~n3700 & ~n3703;
  assign n3981 = ~n3979 & n3980;
  assign n3982 = n3979 & ~n3980;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n3728 & ~n3983;
  assign n3985 = ~n3723 & n3984;
  assign n3986 = ~n3719 & n3985;
  assign n3987 = ~n3723 & ~n3728;
  assign n3988 = ~n3719 & n3987;
  assign n3989 = n3983 & ~n3988;
  assign po26 = ~n3986 & ~n3989;
  assign n3991 = ~n2485 & n3718;
  assign n3992 = n3987 & ~n3991;
  assign n3993 = ~n3981 & ~n3992;
  assign n3994 = ~n3982 & ~n3993;
  assign n3995 = ~n3966 & ~n3969;
  assign n3996 = ~n3957 & n3995;
  assign n3997 = ~n3527 & n3966;
  assign n3998 = ~n3968 & n3997;
  assign n3999 = ~n3967 & n3998;
  assign n4000 = ~n3971 & ~n3999;
  assign n4001 = ~n3996 & n4000;
  assign n4002 = ~n3954 & n3966;
  assign n4003 = ~n3956 & n4002;
  assign n4004 = ~n3957 & n3967;
  assign n4005 = ~n4003 & ~n4004;
  assign n4006 = n4001 & n4005;
  assign n4007 = ~n3817 & ~n3872;
  assign n4008 = ~n3871 & ~n4007;
  assign n4009 = ~n3904 & n3914;
  assign n4010 = pi02 & ~n3205;
  assign n4011 = ~n3206 & n4010;
  assign n4012 = ~n3463 & n4011;
  assign n4013 = pi03 & ~n3207;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = pi57 & ~n4014;
  assign n4016 = ~pi57 & ~n4013;
  assign n4017 = ~n4012 & n4016;
  assign n4018 = ~n4015 & ~n4017;
  assign n4019 = ~n3903 & ~n4018;
  assign n4020 = ~n4009 & n4019;
  assign n4021 = ~n3903 & ~n4009;
  assign n4022 = n4018 & ~n4021;
  assign n4023 = ~n4020 & ~n4022;
  assign n4024 = pi07 & ~n2290;
  assign n4025 = pi06 & pi51;
  assign n4026 = n2645 & n4025;
  assign n4027 = pi06 & ~pi51;
  assign n4028 = n2646 & n4027;
  assign n4029 = ~n4026 & ~n4028;
  assign n4030 = ~n4024 & n4029;
  assign n4031 = pi53 & ~n4030;
  assign n4032 = ~pi53 & ~n4026;
  assign n4033 = ~n4028 & n4032;
  assign n4034 = ~n4024 & n4033;
  assign n4035 = ~n4031 & ~n4034;
  assign n4036 = pi05 & ~n2878;
  assign n4037 = pi04 & pi53;
  assign n4038 = n2958 & n4037;
  assign n4039 = pi04 & ~pi53;
  assign n4040 = n2959 & n4039;
  assign n4041 = ~n4038 & ~n4040;
  assign n4042 = ~n4036 & n4041;
  assign n4043 = pi55 & ~n4042;
  assign n4044 = ~pi55 & ~n4038;
  assign n4045 = ~n4040 & n4044;
  assign n4046 = ~n4036 & n4045;
  assign n4047 = ~n4043 & ~n4046;
  assign n4048 = n4035 & n4047;
  assign n4049 = ~n4035 & ~n4047;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = pi08 & ~n2023;
  assign n4052 = ~n2024 & n4051;
  assign n4053 = ~n2079 & n4052;
  assign n4054 = pi09 & ~n2025;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = pi51 & ~n4055;
  assign n4057 = ~pi51 & ~n4054;
  assign n4058 = ~n4053 & n4057;
  assign n4059 = ~n4056 & ~n4058;
  assign n4060 = ~n4050 & n4059;
  assign n4061 = n4050 & ~n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = ~n4023 & n4062;
  assign n4064 = n4023 & ~n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~n3917 & ~n3931;
  assign n4067 = ~n3929 & ~n4066;
  assign n4068 = ~n4065 & n4067;
  assign n4069 = n4065 & ~n4067;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = ~n3862 & ~n3869;
  assign n4072 = ~n4070 & n4071;
  assign n4073 = n4070 & ~n4071;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = ~n4008 & n4074;
  assign n4076 = n4008 & ~n4074;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = pi13 & ~n1214;
  assign n4079 = pi12 & pi45;
  assign n4080 = n1423 & n4079;
  assign n4081 = pi12 & ~pi45;
  assign n4082 = n1424 & n4081;
  assign n4083 = ~n4080 & ~n4082;
  assign n4084 = ~n4078 & n4083;
  assign n4085 = pi47 & ~n4084;
  assign n4086 = ~pi47 & ~n4080;
  assign n4087 = ~n4082 & n4086;
  assign n4088 = ~n4078 & n4087;
  assign n4089 = ~n4085 & ~n4088;
  assign n4090 = pi11 & ~n1609;
  assign n4091 = pi10 & pi47;
  assign n4092 = n1780 & n4091;
  assign n4093 = pi10 & ~pi47;
  assign n4094 = n1781 & n4093;
  assign n4095 = ~n4092 & ~n4094;
  assign n4096 = ~n4090 & n4095;
  assign n4097 = pi49 & ~n4096;
  assign n4098 = ~pi49 & ~n4092;
  assign n4099 = ~n4094 & n4098;
  assign n4100 = ~n4090 & n4099;
  assign n4101 = ~n4097 & ~n4100;
  assign n4102 = n4089 & n4101;
  assign n4103 = ~n4089 & ~n4101;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = pi14 & ~n1006;
  assign n4106 = ~n1007 & n4105;
  assign n4107 = ~n1068 & n4106;
  assign n4108 = pi15 & ~n1008;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = pi45 & ~n4109;
  assign n4111 = ~pi45 & ~n4108;
  assign n4112 = ~n4107 & n4111;
  assign n4113 = ~n4110 & ~n4112;
  assign n4114 = ~n4104 & n4113;
  assign n4115 = n4104 & ~n4113;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = ~n3847 & n3857;
  assign n4118 = ~n3760 & n3770;
  assign n4119 = ~n3759 & ~n3846;
  assign n4120 = ~n4118 & n4119;
  assign n4121 = ~n4117 & n4120;
  assign n4122 = ~n4116 & n4121;
  assign n4123 = ~n3759 & ~n4118;
  assign n4124 = ~n4114 & n4123;
  assign n4125 = ~n3846 & ~n4117;
  assign n4126 = ~n4115 & ~n4125;
  assign n4127 = n4124 & n4126;
  assign n4128 = ~n4123 & ~n4125;
  assign n4129 = ~n4116 & n4128;
  assign n4130 = ~n4127 & ~n4129;
  assign n4131 = ~n4122 & n4130;
  assign n4132 = ~n3775 & n3813;
  assign n4133 = ~n4114 & n4125;
  assign n4134 = ~n4115 & ~n4123;
  assign n4135 = n4133 & n4134;
  assign n4136 = ~n3774 & ~n4135;
  assign n4137 = ~n4132 & n4136;
  assign n4138 = n4131 & n4137;
  assign n4139 = ~n3774 & ~n4132;
  assign n4140 = ~n4127 & ~n4135;
  assign n4141 = ~n4122 & ~n4129;
  assign n4142 = n4140 & n4141;
  assign n4143 = ~n4139 & ~n4142;
  assign n4144 = ~n4138 & ~n4143;
  assign n4145 = n3788 & n3800;
  assign n4146 = ~n3812 & ~n4145;
  assign n4147 = pi19 & ~n491;
  assign n4148 = pi18 & pi39;
  assign n4149 = n570 & n4148;
  assign n4150 = pi18 & ~pi39;
  assign n4151 = n571 & n4150;
  assign n4152 = ~n4149 & ~n4151;
  assign n4153 = ~n4147 & n4152;
  assign n4154 = pi41 & ~n4153;
  assign n4155 = ~pi41 & ~n4149;
  assign n4156 = ~n4151 & n4155;
  assign n4157 = ~n4147 & n4156;
  assign n4158 = ~n4154 & ~n4157;
  assign n4159 = pi17 & ~n685;
  assign n4160 = pi16 & pi41;
  assign n4161 = n923 & n4160;
  assign n4162 = pi16 & ~pi41;
  assign n4163 = n801 & n4162;
  assign n4164 = ~n4161 & ~n4163;
  assign n4165 = ~n4159 & n4164;
  assign n4166 = pi43 & ~n4165;
  assign n4167 = ~pi43 & ~n4161;
  assign n4168 = ~n4163 & n4167;
  assign n4169 = ~n4159 & n4168;
  assign n4170 = ~n4166 & ~n4169;
  assign n4171 = n4158 & n4170;
  assign n4172 = ~n4158 & ~n4170;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = pi20 & ~n304;
  assign n4175 = ~n305 & n4174;
  assign n4176 = ~n394 & n4175;
  assign n4177 = pi21 & ~n306;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = pi39 & ~n4178;
  assign n4180 = ~pi39 & ~n4177;
  assign n4181 = ~n4176 & n4180;
  assign n4182 = ~n4179 & ~n4181;
  assign n4183 = ~n4173 & n4182;
  assign n4184 = n4173 & ~n4182;
  assign n4185 = ~n4183 & ~n4184;
  assign n4186 = ~n4146 & ~n4185;
  assign n4187 = n4146 & n4185;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = pi22 & ~n193;
  assign n4190 = ~n194 & n4189;
  assign n4191 = ~n729 & n4190;
  assign n4192 = pi23 & ~n195;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = pi37 & ~n4193;
  assign n4195 = ~pi37 & ~n4192;
  assign n4196 = ~n4191 & n4195;
  assign n4197 = ~n4194 & ~n4196;
  assign n4198 = pi24 & ~n141;
  assign n4199 = ~n142 & n4198;
  assign n4200 = ~n156 & n4199;
  assign n4201 = pi25 & ~n143;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = pi35 & ~n4202;
  assign n4204 = ~pi35 & ~n4201;
  assign n4205 = ~n4200 & n4204;
  assign n4206 = ~n4203 & ~n4205;
  assign n4207 = n4197 & ~n4206;
  assign n4208 = ~n4197 & n4206;
  assign n4209 = pi26 & ~pi32;
  assign n4210 = pi27 & pi32;
  assign n4211 = pi33 & ~n4210;
  assign n4212 = ~n4209 & n4211;
  assign n4213 = ~pi33 & n4210;
  assign n4214 = ~n4212 & ~n4213;
  assign n4215 = ~n4208 & n4214;
  assign n4216 = ~n4207 & n4215;
  assign n4217 = ~n4207 & ~n4208;
  assign n4218 = ~n4214 & ~n4217;
  assign n4219 = ~n4216 & ~n4218;
  assign n4220 = ~n4188 & n4219;
  assign n4221 = n4188 & ~n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = ~n4144 & n4222;
  assign n4224 = n4144 & ~n4222;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = ~n4077 & n4225;
  assign n4227 = ~n4075 & ~n4225;
  assign n4228 = ~n4076 & n4227;
  assign n4229 = ~n4226 & ~n4228;
  assign n4230 = ~n3941 & ~n3949;
  assign n4231 = pi58 & ~pi59;
  assign n4232 = ~pi58 & pi59;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = pi00 & ~n3959;
  assign n4235 = ~n3960 & n4234;
  assign n4236 = ~n4233 & n4235;
  assign n4237 = pi01 & ~n3961;
  assign n4238 = pi00 & pi59;
  assign n4239 = ~n3961 & n4238;
  assign n4240 = ~n4237 & ~n4239;
  assign n4241 = ~n4236 & n4240;
  assign n4242 = ~n4236 & ~n4237;
  assign n4243 = n4239 & ~n4242;
  assign n4244 = ~n4241 & ~n4243;
  assign n4245 = ~n4230 & n4244;
  assign n4246 = ~n3941 & ~n4244;
  assign n4247 = ~n3949 & n4246;
  assign n4248 = ~n4245 & ~n4247;
  assign n4249 = ~n3877 & ~n3952;
  assign n4250 = ~n3951 & ~n4249;
  assign n4251 = ~n4248 & n4250;
  assign n4252 = n4248 & ~n4250;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~n4229 & ~n4253;
  assign n4255 = n4229 & ~n4251;
  assign n4256 = ~n4252 & n4255;
  assign n4257 = ~n4254 & ~n4256;
  assign n4258 = ~n4006 & n4257;
  assign n4259 = n4006 & ~n4257;
  assign n4260 = ~n4258 & ~n4259;
  assign n4261 = n3977 & ~n4260;
  assign n4262 = ~n3977 & ~n4258;
  assign n4263 = ~n4259 & n4262;
  assign n4264 = ~n4261 & ~n4263;
  assign n4265 = ~n3994 & n4264;
  assign n4266 = ~n3982 & ~n4264;
  assign n4267 = ~n3993 & n4266;
  assign po27 = ~n4265 & ~n4267;
  assign n4269 = ~n3977 & ~n3982;
  assign n4270 = ~n4260 & ~n4269;
  assign n4271 = n3983 & n4264;
  assign n4272 = ~n3992 & n4271;
  assign n4273 = ~n4270 & ~n4272;
  assign n4274 = ~n3957 & n3966;
  assign n4275 = n3972 & n4274;
  assign n4276 = ~n4006 & ~n4257;
  assign n4277 = ~n4275 & ~n4276;
  assign n4278 = ~n4196 & ~n4205;
  assign n4279 = ~n4203 & n4278;
  assign n4280 = ~n4194 & n4279;
  assign n4281 = ~n4218 & ~n4280;
  assign n4282 = pi17 & ~n683;
  assign n4283 = ~n684 & n4282;
  assign n4284 = ~n1231 & n4283;
  assign n4285 = pi18 & ~n685;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = pi43 & ~n4286;
  assign n4288 = pi19 & ~n489;
  assign n4289 = ~n490 & n4288;
  assign n4290 = ~n572 & n4289;
  assign n4291 = pi20 & ~n491;
  assign n4292 = ~n4290 & ~n4291;
  assign n4293 = pi41 & ~n4292;
  assign n4294 = ~pi41 & ~n4291;
  assign n4295 = ~n4290 & n4294;
  assign n4296 = ~pi43 & ~n4285;
  assign n4297 = ~n4284 & n4296;
  assign n4298 = ~n4295 & ~n4297;
  assign n4299 = ~n4293 & n4298;
  assign n4300 = ~n4287 & n4299;
  assign n4301 = ~n4293 & ~n4295;
  assign n4302 = ~n4287 & ~n4297;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = ~n4300 & ~n4303;
  assign n4305 = pi21 & ~n304;
  assign n4306 = ~n305 & n4305;
  assign n4307 = ~n394 & n4306;
  assign n4308 = pi22 & ~n306;
  assign n4309 = ~n4307 & ~n4308;
  assign n4310 = pi39 & ~n4309;
  assign n4311 = ~pi39 & ~n4308;
  assign n4312 = ~n4307 & n4311;
  assign n4313 = ~n4310 & ~n4312;
  assign n4314 = ~n4304 & n4313;
  assign n4315 = ~n4300 & ~n4313;
  assign n4316 = ~n4303 & n4315;
  assign n4317 = ~n4314 & ~n4316;
  assign n4318 = ~n4281 & ~n4317;
  assign n4319 = n4281 & n4317;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = pi23 & ~n193;
  assign n4322 = ~n194 & n4321;
  assign n4323 = ~n729 & n4322;
  assign n4324 = pi24 & ~n195;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = pi37 & ~n4325;
  assign n4327 = ~pi37 & ~n4324;
  assign n4328 = ~n4323 & n4327;
  assign n4329 = ~n4326 & ~n4328;
  assign n4330 = pi25 & ~n141;
  assign n4331 = ~n142 & n4330;
  assign n4332 = ~n156 & n4331;
  assign n4333 = pi26 & ~n143;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = pi35 & ~n4334;
  assign n4336 = ~pi35 & ~n4333;
  assign n4337 = ~n4332 & n4336;
  assign n4338 = ~n4335 & ~n4337;
  assign n4339 = ~n4329 & n4338;
  assign n4340 = n4329 & ~n4338;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = pi27 & ~pi32;
  assign n4343 = pi28 & pi32;
  assign n4344 = pi33 & ~n4343;
  assign n4345 = ~n4342 & n4344;
  assign n4346 = ~pi33 & n4343;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = ~n4341 & ~n4347;
  assign n4349 = ~n4339 & n4347;
  assign n4350 = ~n4340 & n4349;
  assign n4351 = ~n4348 & ~n4350;
  assign n4352 = ~n4320 & n4351;
  assign n4353 = ~n4318 & ~n4351;
  assign n4354 = ~n4319 & n4353;
  assign n4355 = ~n4352 & ~n4354;
  assign n4356 = pi12 & ~n1609;
  assign n4357 = pi11 & pi47;
  assign n4358 = n1780 & n4357;
  assign n4359 = pi11 & ~pi47;
  assign n4360 = n1781 & n4359;
  assign n4361 = ~n4358 & ~n4360;
  assign n4362 = ~n4356 & n4361;
  assign n4363 = pi49 & ~n4362;
  assign n4364 = ~pi49 & ~n4358;
  assign n4365 = ~n4360 & n4364;
  assign n4366 = ~n4356 & n4365;
  assign n4367 = ~n4363 & ~n4366;
  assign n4368 = pi14 & ~n1214;
  assign n4369 = pi13 & pi45;
  assign n4370 = n1423 & n4369;
  assign n4371 = pi13 & ~pi45;
  assign n4372 = n1424 & n4371;
  assign n4373 = ~n4370 & ~n4372;
  assign n4374 = ~n4368 & n4373;
  assign n4375 = pi47 & ~n4374;
  assign n4376 = ~pi47 & ~n4370;
  assign n4377 = ~n4372 & n4376;
  assign n4378 = ~n4368 & n4377;
  assign n4379 = ~n4375 & ~n4378;
  assign n4380 = ~n4367 & n4379;
  assign n4381 = n4367 & ~n4379;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = pi15 & ~n1006;
  assign n4384 = ~n1007 & n4383;
  assign n4385 = ~n1068 & n4384;
  assign n4386 = pi16 & ~n1008;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = pi45 & ~n4387;
  assign n4389 = ~pi45 & ~n4386;
  assign n4390 = ~n4385 & n4389;
  assign n4391 = ~n4388 & ~n4390;
  assign n4392 = ~n4382 & n4391;
  assign n4393 = n4382 & ~n4391;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = ~n4103 & n4113;
  assign n4396 = ~n4172 & n4182;
  assign n4397 = ~n4102 & ~n4171;
  assign n4398 = ~n4396 & n4397;
  assign n4399 = ~n4395 & n4398;
  assign n4400 = n4394 & n4399;
  assign n4401 = ~n4171 & ~n4396;
  assign n4402 = ~n4102 & ~n4395;
  assign n4403 = n4401 & ~n4402;
  assign n4404 = ~n4394 & n4403;
  assign n4405 = ~n4401 & ~n4402;
  assign n4406 = n4394 & n4405;
  assign n4407 = ~n4404 & ~n4406;
  assign n4408 = ~n4400 & n4407;
  assign n4409 = ~n4187 & n4219;
  assign n4410 = ~n4401 & n4402;
  assign n4411 = ~n4394 & n4410;
  assign n4412 = ~n4186 & ~n4411;
  assign n4413 = ~n4409 & n4412;
  assign n4414 = n4408 & n4413;
  assign n4415 = ~n4186 & ~n4409;
  assign n4416 = ~n4404 & ~n4411;
  assign n4417 = ~n4400 & ~n4406;
  assign n4418 = n4416 & n4417;
  assign n4419 = ~n4415 & ~n4418;
  assign n4420 = ~n4414 & ~n4419;
  assign n4421 = ~n4355 & ~n4420;
  assign n4422 = n4355 & n4420;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = ~n4143 & ~n4224;
  assign n4425 = ~n4022 & ~n4064;
  assign n4426 = pi03 & ~n3205;
  assign n4427 = ~n3206 & n4426;
  assign n4428 = ~n3463 & n4427;
  assign n4429 = pi04 & ~n3207;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = pi57 & ~n4430;
  assign n4432 = ~pi57 & ~n4429;
  assign n4433 = ~n4428 & n4432;
  assign n4434 = ~n4431 & ~n4433;
  assign n4435 = ~n4049 & n4059;
  assign n4436 = ~n4048 & ~n4435;
  assign n4437 = n4434 & ~n4436;
  assign n4438 = pi08 & ~n2290;
  assign n4439 = pi07 & pi51;
  assign n4440 = n2645 & n4439;
  assign n4441 = pi07 & ~pi51;
  assign n4442 = n2646 & n4441;
  assign n4443 = ~n4440 & ~n4442;
  assign n4444 = ~n4438 & n4443;
  assign n4445 = pi53 & ~n4444;
  assign n4446 = ~pi53 & ~n4440;
  assign n4447 = ~n4442 & n4446;
  assign n4448 = ~n4438 & n4447;
  assign n4449 = ~n4445 & ~n4448;
  assign n4450 = pi06 & ~n2878;
  assign n4451 = pi05 & pi53;
  assign n4452 = n2958 & n4451;
  assign n4453 = pi05 & ~pi53;
  assign n4454 = n2959 & n4453;
  assign n4455 = ~n4452 & ~n4454;
  assign n4456 = ~n4450 & n4455;
  assign n4457 = pi55 & ~n4456;
  assign n4458 = ~pi55 & ~n4452;
  assign n4459 = ~n4454 & n4458;
  assign n4460 = ~n4450 & n4459;
  assign n4461 = ~n4457 & ~n4460;
  assign n4462 = n4449 & n4461;
  assign n4463 = ~n4449 & ~n4461;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = pi09 & ~n2023;
  assign n4466 = ~n2024 & n4465;
  assign n4467 = ~n2079 & n4466;
  assign n4468 = pi10 & ~n2025;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = pi51 & ~n4469;
  assign n4471 = ~pi51 & ~n4468;
  assign n4472 = ~n4467 & n4471;
  assign n4473 = ~n4470 & ~n4472;
  assign n4474 = ~n4464 & n4473;
  assign n4475 = n4464 & ~n4473;
  assign n4476 = ~n4474 & ~n4475;
  assign n4477 = ~n4048 & ~n4434;
  assign n4478 = ~n4435 & n4477;
  assign n4479 = ~n4476 & ~n4478;
  assign n4480 = ~n4437 & n4479;
  assign n4481 = ~n4437 & ~n4478;
  assign n4482 = n4476 & ~n4481;
  assign n4483 = ~n4480 & ~n4482;
  assign n4484 = ~n4425 & n4483;
  assign n4485 = n4425 & ~n4483;
  assign n4486 = ~n4484 & ~n4485;
  assign n4487 = ~n4116 & ~n4125;
  assign n4488 = ~n4115 & n4133;
  assign n4489 = ~n4123 & ~n4488;
  assign n4490 = ~n4487 & ~n4489;
  assign n4491 = ~n4486 & n4490;
  assign n4492 = ~n4484 & ~n4490;
  assign n4493 = ~n4485 & n4492;
  assign n4494 = ~n4491 & ~n4493;
  assign n4495 = ~n4424 & n4494;
  assign n4496 = n4424 & ~n4494;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = ~n4423 & ~n4497;
  assign n4499 = n4423 & ~n4495;
  assign n4500 = ~n4496 & n4499;
  assign n4501 = ~n4498 & ~n4500;
  assign n4502 = ~n4076 & n4225;
  assign n4503 = ~n4075 & ~n4502;
  assign n4504 = pi01 & ~n3959;
  assign n4505 = ~n3960 & n4504;
  assign n4506 = ~n4233 & n4505;
  assign n4507 = pi02 & ~n3961;
  assign n4508 = ~n4506 & ~n4507;
  assign n4509 = pi59 & ~n4508;
  assign n4510 = ~pi59 & ~n4507;
  assign n4511 = ~n4506 & n4510;
  assign n4512 = ~n4509 & ~n4511;
  assign n4513 = pi59 & ~pi60;
  assign n4514 = ~pi59 & pi60;
  assign n4515 = ~n4513 & ~n4514;
  assign n4516 = pi00 & ~n4515;
  assign n4517 = ~n4512 & n4516;
  assign n4518 = ~n4511 & ~n4516;
  assign n4519 = ~n4509 & n4518;
  assign n4520 = ~n4517 & ~n4519;
  assign n4521 = pi59 & ~n3962;
  assign n4522 = n4242 & n4521;
  assign n4523 = ~n4520 & ~n4522;
  assign n4524 = ~n4519 & n4522;
  assign n4525 = ~n4517 & n4524;
  assign n4526 = ~n4523 & ~n4525;
  assign n4527 = ~n4069 & n4526;
  assign n4528 = ~n4073 & n4527;
  assign n4529 = ~n4069 & ~n4073;
  assign n4530 = ~n4526 & ~n4529;
  assign n4531 = ~n4528 & ~n4530;
  assign n4532 = ~n4503 & n4531;
  assign n4533 = n4503 & ~n4531;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n4501 & ~n4534;
  assign n4536 = n4501 & ~n4532;
  assign n4537 = ~n4533 & n4536;
  assign n4538 = ~n4535 & ~n4537;
  assign n4539 = n4229 & ~n4252;
  assign n4540 = n4245 & ~n4251;
  assign n4541 = ~n4539 & n4540;
  assign n4542 = ~n4251 & ~n4539;
  assign n4543 = ~n4245 & ~n4542;
  assign n4544 = ~n4541 & ~n4543;
  assign n4545 = ~n4538 & ~n4544;
  assign n4546 = n4538 & ~n4541;
  assign n4547 = ~n4543 & n4546;
  assign n4548 = ~n4545 & ~n4547;
  assign n4549 = ~n4277 & ~n4548;
  assign n4550 = n4277 & n4548;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = ~n4273 & n4551;
  assign n4553 = ~n4270 & ~n4551;
  assign n4554 = ~n4272 & n4553;
  assign po28 = ~n4552 & ~n4554;
  assign n4556 = n3705 & ~n3981;
  assign n4557 = ~n3982 & ~n4261;
  assign n4558 = ~n4263 & n4557;
  assign n4559 = n4556 & n4558;
  assign n4560 = ~n4270 & ~n4549;
  assign n4561 = ~n4559 & n4560;
  assign n4562 = ~n4550 & ~n4561;
  assign n4563 = n2947 & n3452;
  assign n4564 = ~n2953 & n4563;
  assign n4565 = ~n3451 & ~n3720;
  assign n4566 = ~n4564 & n4565;
  assign n4567 = n3708 & ~n4549;
  assign n4568 = ~n4550 & n4567;
  assign n4569 = n4271 & n4568;
  assign n4570 = ~n4566 & n4569;
  assign n4571 = ~n4562 & ~n4570;
  assign n4572 = ~n4423 & ~n4496;
  assign n4573 = ~n4485 & ~n4490;
  assign n4574 = ~n4484 & ~n4573;
  assign n4575 = pi60 & ~pi61;
  assign n4576 = ~pi60 & pi61;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = pi00 & ~n4513;
  assign n4579 = ~n4514 & n4578;
  assign n4580 = ~n4577 & n4579;
  assign n4581 = pi01 & ~n4515;
  assign n4582 = ~n4580 & ~n4581;
  assign n4583 = pi61 & ~n4582;
  assign n4584 = pi02 & ~n3959;
  assign n4585 = ~n3960 & n4584;
  assign n4586 = ~n4233 & n4585;
  assign n4587 = pi03 & ~n3961;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = pi59 & ~n4588;
  assign n4590 = ~pi59 & ~n4587;
  assign n4591 = ~n4586 & n4590;
  assign n4592 = ~pi61 & ~n4581;
  assign n4593 = ~n4580 & n4592;
  assign n4594 = ~n4591 & ~n4593;
  assign n4595 = ~n4589 & n4594;
  assign n4596 = ~n4583 & n4595;
  assign n4597 = ~n4589 & ~n4591;
  assign n4598 = ~n4583 & ~n4593;
  assign n4599 = ~n4597 & ~n4598;
  assign n4600 = ~n4596 & ~n4599;
  assign n4601 = pi61 & ~n4516;
  assign n4602 = ~n4511 & n4516;
  assign n4603 = ~n4509 & n4602;
  assign n4604 = ~n4601 & ~n4603;
  assign n4605 = ~n4600 & n4604;
  assign n4606 = n4600 & ~n4604;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4574 & n4607;
  assign n4609 = ~n4484 & ~n4607;
  assign n4610 = ~n4573 & n4609;
  assign n4611 = ~n4608 & ~n4610;
  assign n4612 = ~n4495 & ~n4611;
  assign n4613 = ~n4572 & n4612;
  assign n4614 = ~n4495 & ~n4572;
  assign n4615 = n4611 & ~n4614;
  assign n4616 = ~n4613 & ~n4615;
  assign n4617 = ~n4463 & n4473;
  assign n4618 = pi04 & ~n3205;
  assign n4619 = ~n3206 & n4618;
  assign n4620 = ~n3463 & n4619;
  assign n4621 = pi05 & ~n3207;
  assign n4622 = ~n4620 & ~n4621;
  assign n4623 = pi57 & ~n4622;
  assign n4624 = ~pi57 & ~n4621;
  assign n4625 = ~n4620 & n4624;
  assign n4626 = ~n4623 & ~n4625;
  assign n4627 = ~n4462 & ~n4626;
  assign n4628 = ~n4617 & n4627;
  assign n4629 = ~n4462 & ~n4617;
  assign n4630 = n4626 & ~n4629;
  assign n4631 = ~n4628 & ~n4630;
  assign n4632 = pi06 & ~n2876;
  assign n4633 = ~n2877 & n4632;
  assign n4634 = ~n2960 & n4633;
  assign n4635 = pi07 & ~n2878;
  assign n4636 = ~n4634 & ~n4635;
  assign n4637 = pi55 & ~n4636;
  assign n4638 = pi08 & ~n2288;
  assign n4639 = ~n2289 & n4638;
  assign n4640 = ~n2647 & n4639;
  assign n4641 = pi09 & ~n2290;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = pi53 & ~n4642;
  assign n4644 = ~pi53 & ~n4641;
  assign n4645 = ~n4640 & n4644;
  assign n4646 = ~pi55 & ~n4635;
  assign n4647 = ~n4634 & n4646;
  assign n4648 = ~n4645 & ~n4647;
  assign n4649 = ~n4643 & n4648;
  assign n4650 = ~n4637 & n4649;
  assign n4651 = ~n4643 & ~n4645;
  assign n4652 = ~n4637 & ~n4647;
  assign n4653 = ~n4651 & ~n4652;
  assign n4654 = ~n4650 & ~n4653;
  assign n4655 = pi10 & ~n2023;
  assign n4656 = ~n2024 & n4655;
  assign n4657 = ~n2079 & n4656;
  assign n4658 = pi11 & ~n2025;
  assign n4659 = ~n4657 & ~n4658;
  assign n4660 = pi51 & ~n4659;
  assign n4661 = ~pi51 & ~n4658;
  assign n4662 = ~n4657 & n4661;
  assign n4663 = ~n4660 & ~n4662;
  assign n4664 = ~n4654 & n4663;
  assign n4665 = ~n4650 & ~n4663;
  assign n4666 = ~n4653 & n4665;
  assign n4667 = ~n4664 & ~n4666;
  assign n4668 = ~n4631 & n4667;
  assign n4669 = n4631 & ~n4667;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = ~n4437 & ~n4480;
  assign n4672 = ~n4670 & n4671;
  assign n4673 = n4670 & ~n4671;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = n4394 & ~n4402;
  assign n4676 = ~n4394 & n4402;
  assign n4677 = ~n4401 & ~n4676;
  assign n4678 = ~n4675 & ~n4677;
  assign n4679 = ~n4674 & n4678;
  assign n4680 = ~n4672 & ~n4678;
  assign n4681 = ~n4673 & n4680;
  assign n4682 = ~n4679 & ~n4681;
  assign n4683 = ~n4355 & n4420;
  assign n4684 = ~n4419 & ~n4683;
  assign n4685 = n4682 & ~n4684;
  assign n4686 = ~n4682 & n4684;
  assign n4687 = pi12 & ~n1607;
  assign n4688 = ~n1608 & n4687;
  assign n4689 = ~n1782 & n4688;
  assign n4690 = pi13 & ~n1609;
  assign n4691 = ~n4689 & ~n4690;
  assign n4692 = pi49 & ~n4691;
  assign n4693 = pi14 & ~n1212;
  assign n4694 = ~n1213 & n4693;
  assign n4695 = ~n1425 & n4694;
  assign n4696 = pi15 & ~n1214;
  assign n4697 = ~n4695 & ~n4696;
  assign n4698 = pi47 & ~n4697;
  assign n4699 = ~pi47 & ~n4696;
  assign n4700 = ~n4695 & n4699;
  assign n4701 = ~pi49 & ~n4690;
  assign n4702 = ~n4689 & n4701;
  assign n4703 = ~n4700 & ~n4702;
  assign n4704 = ~n4698 & n4703;
  assign n4705 = ~n4692 & n4704;
  assign n4706 = ~n4698 & ~n4700;
  assign n4707 = ~n4692 & ~n4702;
  assign n4708 = ~n4706 & ~n4707;
  assign n4709 = ~n4705 & ~n4708;
  assign n4710 = pi16 & ~n1006;
  assign n4711 = ~n1007 & n4710;
  assign n4712 = ~n1068 & n4711;
  assign n4713 = pi17 & ~n1008;
  assign n4714 = ~n4712 & ~n4713;
  assign n4715 = pi45 & ~n4714;
  assign n4716 = ~pi45 & ~n4713;
  assign n4717 = ~n4712 & n4716;
  assign n4718 = ~n4715 & ~n4717;
  assign n4719 = ~n4709 & n4718;
  assign n4720 = ~n4705 & ~n4718;
  assign n4721 = ~n4708 & n4720;
  assign n4722 = ~n4719 & ~n4721;
  assign n4723 = ~n4303 & n4313;
  assign n4724 = n4367 & n4379;
  assign n4725 = ~n4300 & ~n4724;
  assign n4726 = ~n4392 & n4725;
  assign n4727 = ~n4723 & n4726;
  assign n4728 = ~n4722 & n4727;
  assign n4729 = ~n4300 & ~n4723;
  assign n4730 = ~n4719 & n4729;
  assign n4731 = ~n4392 & ~n4724;
  assign n4732 = ~n4721 & ~n4731;
  assign n4733 = n4730 & n4732;
  assign n4734 = ~n4729 & ~n4731;
  assign n4735 = ~n4722 & n4734;
  assign n4736 = ~n4733 & ~n4735;
  assign n4737 = ~n4728 & n4736;
  assign n4738 = ~n4319 & n4351;
  assign n4739 = ~n4719 & n4731;
  assign n4740 = ~n4721 & ~n4729;
  assign n4741 = n4739 & n4740;
  assign n4742 = ~n4318 & ~n4741;
  assign n4743 = ~n4738 & n4742;
  assign n4744 = n4737 & n4743;
  assign n4745 = ~n4318 & ~n4738;
  assign n4746 = ~n4733 & ~n4741;
  assign n4747 = ~n4728 & ~n4735;
  assign n4748 = n4746 & n4747;
  assign n4749 = ~n4745 & ~n4748;
  assign n4750 = ~n4744 & ~n4749;
  assign n4751 = ~n4328 & ~n4337;
  assign n4752 = ~n4335 & n4751;
  assign n4753 = ~n4326 & n4752;
  assign n4754 = ~n4348 & ~n4753;
  assign n4755 = pi18 & ~n683;
  assign n4756 = ~n684 & n4755;
  assign n4757 = ~n1231 & n4756;
  assign n4758 = pi19 & ~n685;
  assign n4759 = ~n4757 & ~n4758;
  assign n4760 = pi43 & ~n4759;
  assign n4761 = pi20 & ~n489;
  assign n4762 = ~n490 & n4761;
  assign n4763 = ~n572 & n4762;
  assign n4764 = pi21 & ~n491;
  assign n4765 = ~n4763 & ~n4764;
  assign n4766 = pi41 & ~n4765;
  assign n4767 = ~pi41 & ~n4764;
  assign n4768 = ~n4763 & n4767;
  assign n4769 = ~pi43 & ~n4758;
  assign n4770 = ~n4757 & n4769;
  assign n4771 = ~n4768 & ~n4770;
  assign n4772 = ~n4766 & n4771;
  assign n4773 = ~n4760 & n4772;
  assign n4774 = ~n4766 & ~n4768;
  assign n4775 = ~n4760 & ~n4770;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = ~n4773 & ~n4776;
  assign n4778 = pi22 & ~n304;
  assign n4779 = ~n305 & n4778;
  assign n4780 = ~n394 & n4779;
  assign n4781 = pi23 & ~n306;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = pi39 & ~n4782;
  assign n4784 = ~pi39 & ~n4781;
  assign n4785 = ~n4780 & n4784;
  assign n4786 = ~n4783 & ~n4785;
  assign n4787 = ~n4777 & n4786;
  assign n4788 = ~n4773 & ~n4786;
  assign n4789 = ~n4776 & n4788;
  assign n4790 = ~n4787 & ~n4789;
  assign n4791 = ~n4754 & ~n4790;
  assign n4792 = n4754 & n4790;
  assign n4793 = ~n4791 & ~n4792;
  assign n4794 = pi24 & ~n193;
  assign n4795 = ~n194 & n4794;
  assign n4796 = ~n729 & n4795;
  assign n4797 = pi25 & ~n195;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = pi37 & ~n4798;
  assign n4800 = ~pi37 & ~n4797;
  assign n4801 = ~n4796 & n4800;
  assign n4802 = ~n4799 & ~n4801;
  assign n4803 = pi26 & ~n141;
  assign n4804 = ~n142 & n4803;
  assign n4805 = ~n156 & n4804;
  assign n4806 = pi27 & ~n143;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = pi35 & ~n4807;
  assign n4809 = ~pi35 & ~n4806;
  assign n4810 = ~n4805 & n4809;
  assign n4811 = ~n4808 & ~n4810;
  assign n4812 = n4802 & ~n4811;
  assign n4813 = ~n4802 & n4811;
  assign n4814 = pi28 & ~pi32;
  assign n4815 = pi29 & pi32;
  assign n4816 = pi33 & ~n4815;
  assign n4817 = ~n4814 & n4816;
  assign n4818 = ~pi33 & n4815;
  assign n4819 = ~n4817 & ~n4818;
  assign n4820 = ~n4813 & n4819;
  assign n4821 = ~n4812 & n4820;
  assign n4822 = ~n4812 & ~n4813;
  assign n4823 = ~n4819 & ~n4822;
  assign n4824 = ~n4821 & ~n4823;
  assign n4825 = ~n4793 & n4824;
  assign n4826 = ~n4791 & ~n4824;
  assign n4827 = ~n4792 & n4826;
  assign n4828 = ~n4825 & ~n4827;
  assign n4829 = ~n4750 & n4828;
  assign n4830 = n4750 & ~n4828;
  assign n4831 = ~n4829 & ~n4830;
  assign n4832 = ~n4686 & n4831;
  assign n4833 = ~n4685 & n4832;
  assign n4834 = ~n4685 & ~n4686;
  assign n4835 = ~n4831 & ~n4834;
  assign n4836 = ~n4833 & ~n4835;
  assign n4837 = ~n4616 & n4836;
  assign n4838 = n4616 & ~n4836;
  assign n4839 = ~n4837 & ~n4838;
  assign n4840 = ~n4501 & ~n4533;
  assign n4841 = ~n4520 & n4522;
  assign n4842 = ~n4530 & ~n4841;
  assign n4843 = ~n4532 & ~n4842;
  assign n4844 = ~n4840 & n4843;
  assign n4845 = ~n4532 & ~n4840;
  assign n4846 = n4842 & ~n4845;
  assign n4847 = ~n4844 & ~n4846;
  assign n4848 = ~n4839 & ~n4847;
  assign n4849 = n4839 & n4847;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4538 & ~n4543;
  assign n4852 = ~n4541 & ~n4851;
  assign n4853 = ~n4850 & n4852;
  assign n4854 = n4850 & ~n4852;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = ~n4571 & n4855;
  assign n4857 = ~n4562 & ~n4855;
  assign n4858 = ~n4570 & n4857;
  assign po29 = ~n4856 & ~n4858;
  assign n4860 = n2716 & n4563;
  assign n4861 = ~n2270 & n4860;
  assign n4862 = n3454 & ~n4562;
  assign n4863 = ~n4861 & n4862;
  assign n4864 = ~n4562 & ~n4569;
  assign n4865 = ~n4853 & ~n4864;
  assign n4866 = ~n4863 & n4865;
  assign n4867 = ~n4854 & ~n4866;
  assign n4868 = ~n4842 & ~n4845;
  assign n4869 = ~n4848 & ~n4868;
  assign n4870 = ~n4749 & ~n4830;
  assign n4871 = ~n4653 & n4663;
  assign n4872 = pi05 & ~n3205;
  assign n4873 = ~n3206 & n4872;
  assign n4874 = ~n3463 & n4873;
  assign n4875 = pi06 & ~n3207;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = pi57 & ~n4876;
  assign n4878 = ~pi57 & ~n4875;
  assign n4879 = ~n4874 & n4878;
  assign n4880 = ~n4877 & ~n4879;
  assign n4881 = ~n4650 & ~n4880;
  assign n4882 = ~n4871 & n4881;
  assign n4883 = ~n4650 & ~n4871;
  assign n4884 = n4880 & ~n4883;
  assign n4885 = ~n4882 & ~n4884;
  assign n4886 = pi07 & ~n2876;
  assign n4887 = ~n2877 & n4886;
  assign n4888 = ~n2960 & n4887;
  assign n4889 = pi08 & ~n2878;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = pi55 & ~n4890;
  assign n4892 = pi09 & ~n2288;
  assign n4893 = ~n2289 & n4892;
  assign n4894 = ~n2647 & n4893;
  assign n4895 = pi10 & ~n2290;
  assign n4896 = ~n4894 & ~n4895;
  assign n4897 = pi53 & ~n4896;
  assign n4898 = ~pi53 & ~n4895;
  assign n4899 = ~n4894 & n4898;
  assign n4900 = ~pi55 & ~n4889;
  assign n4901 = ~n4888 & n4900;
  assign n4902 = ~n4899 & ~n4901;
  assign n4903 = ~n4897 & n4902;
  assign n4904 = ~n4891 & n4903;
  assign n4905 = ~n4897 & ~n4899;
  assign n4906 = ~n4891 & ~n4901;
  assign n4907 = ~n4905 & ~n4906;
  assign n4908 = ~n4904 & ~n4907;
  assign n4909 = pi11 & ~n2023;
  assign n4910 = ~n2024 & n4909;
  assign n4911 = ~n2079 & n4910;
  assign n4912 = pi12 & ~n2025;
  assign n4913 = ~n4911 & ~n4912;
  assign n4914 = pi51 & ~n4913;
  assign n4915 = ~pi51 & ~n4912;
  assign n4916 = ~n4911 & n4915;
  assign n4917 = ~n4914 & ~n4916;
  assign n4918 = ~n4908 & n4917;
  assign n4919 = ~n4904 & ~n4917;
  assign n4920 = ~n4907 & n4919;
  assign n4921 = ~n4918 & ~n4920;
  assign n4922 = n4885 & ~n4921;
  assign n4923 = ~n4630 & ~n4669;
  assign n4924 = ~n4885 & n4921;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = ~n4922 & n4925;
  assign n4927 = ~n4922 & ~n4924;
  assign n4928 = n4923 & ~n4927;
  assign n4929 = ~n4926 & ~n4928;
  assign n4930 = ~n4722 & ~n4731;
  assign n4931 = ~n4721 & n4739;
  assign n4932 = ~n4729 & ~n4931;
  assign n4933 = ~n4930 & ~n4932;
  assign n4934 = ~n4929 & n4933;
  assign n4935 = ~n4926 & ~n4933;
  assign n4936 = ~n4928 & n4935;
  assign n4937 = ~n4934 & ~n4936;
  assign n4938 = ~n4870 & n4937;
  assign n4939 = n4870 & ~n4937;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = pi13 & ~n1607;
  assign n4942 = ~n1608 & n4941;
  assign n4943 = ~n1782 & n4942;
  assign n4944 = pi14 & ~n1609;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = pi49 & ~n4945;
  assign n4947 = pi15 & ~n1212;
  assign n4948 = ~n1213 & n4947;
  assign n4949 = ~n1425 & n4948;
  assign n4950 = pi16 & ~n1214;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = pi47 & ~n4951;
  assign n4953 = ~pi47 & ~n4950;
  assign n4954 = ~n4949 & n4953;
  assign n4955 = ~pi49 & ~n4944;
  assign n4956 = ~n4943 & n4955;
  assign n4957 = ~n4954 & ~n4956;
  assign n4958 = ~n4952 & n4957;
  assign n4959 = ~n4946 & n4958;
  assign n4960 = ~n4952 & ~n4954;
  assign n4961 = ~n4946 & ~n4956;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = ~n4959 & ~n4962;
  assign n4964 = pi17 & ~n1006;
  assign n4965 = ~n1007 & n4964;
  assign n4966 = ~n1068 & n4965;
  assign n4967 = pi18 & ~n1008;
  assign n4968 = ~n4966 & ~n4967;
  assign n4969 = pi45 & ~n4968;
  assign n4970 = ~pi45 & ~n4967;
  assign n4971 = ~n4966 & n4970;
  assign n4972 = ~n4969 & ~n4971;
  assign n4973 = ~n4963 & n4972;
  assign n4974 = ~n4959 & ~n4972;
  assign n4975 = ~n4962 & n4974;
  assign n4976 = ~n4973 & ~n4975;
  assign n4977 = ~n4708 & n4718;
  assign n4978 = ~n4776 & n4786;
  assign n4979 = ~n4705 & ~n4773;
  assign n4980 = ~n4978 & n4979;
  assign n4981 = ~n4977 & n4980;
  assign n4982 = ~n4976 & n4981;
  assign n4983 = ~n4773 & ~n4978;
  assign n4984 = ~n4973 & n4983;
  assign n4985 = ~n4705 & ~n4977;
  assign n4986 = ~n4975 & ~n4985;
  assign n4987 = n4984 & n4986;
  assign n4988 = ~n4983 & ~n4985;
  assign n4989 = ~n4976 & n4988;
  assign n4990 = ~n4987 & ~n4989;
  assign n4991 = ~n4982 & n4990;
  assign n4992 = ~n4792 & n4824;
  assign n4993 = ~n4973 & n4985;
  assign n4994 = ~n4975 & ~n4983;
  assign n4995 = n4993 & n4994;
  assign n4996 = ~n4791 & ~n4995;
  assign n4997 = ~n4992 & n4996;
  assign n4998 = n4991 & n4997;
  assign n4999 = ~n4791 & ~n4992;
  assign n5000 = ~n4987 & ~n4995;
  assign n5001 = ~n4982 & ~n4989;
  assign n5002 = n5000 & n5001;
  assign n5003 = ~n4999 & ~n5002;
  assign n5004 = ~n4998 & ~n5003;
  assign n5005 = ~n4801 & ~n4810;
  assign n5006 = ~n4808 & n5005;
  assign n5007 = ~n4799 & n5006;
  assign n5008 = ~n4823 & ~n5007;
  assign n5009 = pi19 & ~n683;
  assign n5010 = ~n684 & n5009;
  assign n5011 = ~n1231 & n5010;
  assign n5012 = pi20 & ~n685;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = pi43 & ~n5013;
  assign n5015 = pi21 & ~n489;
  assign n5016 = ~n490 & n5015;
  assign n5017 = ~n572 & n5016;
  assign n5018 = pi22 & ~n491;
  assign n5019 = ~n5017 & ~n5018;
  assign n5020 = pi41 & ~n5019;
  assign n5021 = ~pi41 & ~n5018;
  assign n5022 = ~n5017 & n5021;
  assign n5023 = ~pi43 & ~n5012;
  assign n5024 = ~n5011 & n5023;
  assign n5025 = ~n5022 & ~n5024;
  assign n5026 = ~n5020 & n5025;
  assign n5027 = ~n5014 & n5026;
  assign n5028 = ~n5020 & ~n5022;
  assign n5029 = ~n5014 & ~n5024;
  assign n5030 = ~n5028 & ~n5029;
  assign n5031 = ~n5027 & ~n5030;
  assign n5032 = pi23 & ~n304;
  assign n5033 = ~n305 & n5032;
  assign n5034 = ~n394 & n5033;
  assign n5035 = pi24 & ~n306;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = pi39 & ~n5036;
  assign n5038 = ~pi39 & ~n5035;
  assign n5039 = ~n5034 & n5038;
  assign n5040 = ~n5037 & ~n5039;
  assign n5041 = ~n5031 & n5040;
  assign n5042 = ~n5027 & ~n5040;
  assign n5043 = ~n5030 & n5042;
  assign n5044 = ~n5041 & ~n5043;
  assign n5045 = ~n5008 & ~n5044;
  assign n5046 = n5008 & n5044;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = pi25 & ~n193;
  assign n5049 = ~n194 & n5048;
  assign n5050 = ~n729 & n5049;
  assign n5051 = pi26 & ~n195;
  assign n5052 = ~n5050 & ~n5051;
  assign n5053 = pi37 & ~n5052;
  assign n5054 = ~pi37 & ~n5051;
  assign n5055 = ~n5050 & n5054;
  assign n5056 = ~n5053 & ~n5055;
  assign n5057 = pi27 & ~n141;
  assign n5058 = ~n142 & n5057;
  assign n5059 = ~n156 & n5058;
  assign n5060 = pi28 & ~n143;
  assign n5061 = ~n5059 & ~n5060;
  assign n5062 = pi35 & ~n5061;
  assign n5063 = ~pi35 & ~n5060;
  assign n5064 = ~n5059 & n5063;
  assign n5065 = ~n5062 & ~n5064;
  assign n5066 = n5056 & ~n5065;
  assign n5067 = ~n5056 & n5065;
  assign n5068 = pi29 & ~pi32;
  assign n5069 = pi30 & pi32;
  assign n5070 = pi33 & ~n5069;
  assign n5071 = ~n5068 & n5070;
  assign n5072 = ~pi33 & n5069;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = ~n5067 & n5073;
  assign n5075 = ~n5066 & n5074;
  assign n5076 = ~n5066 & ~n5067;
  assign n5077 = ~n5073 & ~n5076;
  assign n5078 = ~n5075 & ~n5077;
  assign n5079 = ~n5047 & n5078;
  assign n5080 = ~n5045 & ~n5078;
  assign n5081 = ~n5046 & n5080;
  assign n5082 = ~n5079 & ~n5081;
  assign n5083 = ~n5004 & n5082;
  assign n5084 = n5004 & ~n5082;
  assign n5085 = ~n5083 & ~n5084;
  assign n5086 = ~n4940 & n5085;
  assign n5087 = ~n4938 & ~n5085;
  assign n5088 = ~n4939 & n5087;
  assign n5089 = ~n5086 & ~n5088;
  assign n5090 = ~n4685 & ~n4833;
  assign n5091 = pi61 & ~pi62;
  assign n5092 = ~pi61 & pi62;
  assign n5093 = ~n5091 & ~n5092;
  assign n5094 = pi00 & ~n5093;
  assign n5095 = pi63 & ~n5094;
  assign n5096 = pi00 & ~pi63;
  assign n5097 = ~n5093 & n5096;
  assign n5098 = ~n5095 & ~n5097;
  assign n5099 = pi01 & ~n4513;
  assign n5100 = ~n4514 & n5099;
  assign n5101 = ~n4577 & n5100;
  assign n5102 = pi02 & ~n4515;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = pi61 & ~n5103;
  assign n5105 = ~pi61 & ~n5102;
  assign n5106 = ~n5101 & n5105;
  assign n5107 = ~n5104 & ~n5106;
  assign n5108 = n5098 & ~n5107;
  assign n5109 = pi03 & ~n3959;
  assign n5110 = ~n3960 & n5109;
  assign n5111 = ~n4233 & n5110;
  assign n5112 = pi04 & ~n3961;
  assign n5113 = ~n5111 & ~n5112;
  assign n5114 = pi59 & ~n5113;
  assign n5115 = ~pi59 & ~n5112;
  assign n5116 = ~n5111 & n5115;
  assign n5117 = ~n5114 & ~n5116;
  assign n5118 = ~n5098 & ~n5106;
  assign n5119 = ~n5104 & n5118;
  assign n5120 = ~n5117 & ~n5119;
  assign n5121 = ~n5108 & n5120;
  assign n5122 = ~n5108 & ~n5119;
  assign n5123 = n5117 & ~n5122;
  assign n5124 = ~n5121 & ~n5123;
  assign n5125 = pi63 & ~n4596;
  assign n5126 = ~pi63 & ~n4591;
  assign n5127 = ~n4589 & n5126;
  assign n5128 = n4598 & n5127;
  assign n5129 = ~n5125 & ~n5128;
  assign n5130 = n5124 & n5129;
  assign n5131 = ~n5124 & ~n5129;
  assign n5132 = ~n4606 & ~n5131;
  assign n5133 = ~n5130 & n5132;
  assign n5134 = ~n5130 & ~n5131;
  assign n5135 = n4606 & ~n5134;
  assign n5136 = ~n4673 & ~n5135;
  assign n5137 = ~n5133 & n5136;
  assign n5138 = ~n4681 & n5137;
  assign n5139 = ~n4673 & ~n4681;
  assign n5140 = ~n5133 & ~n5135;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = ~n5138 & ~n5141;
  assign n5143 = ~n5090 & n5142;
  assign n5144 = ~n4685 & ~n5142;
  assign n5145 = ~n4833 & n5144;
  assign n5146 = ~n5143 & ~n5145;
  assign n5147 = ~n5089 & ~n5146;
  assign n5148 = n5089 & n5146;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = ~n4615 & ~n4836;
  assign n5151 = ~n4613 & ~n5150;
  assign n5152 = n4608 & ~n5151;
  assign n5153 = ~n4608 & ~n4613;
  assign n5154 = ~n5150 & n5153;
  assign n5155 = ~n5152 & ~n5154;
  assign n5156 = ~n5149 & ~n5155;
  assign n5157 = n5149 & n5155;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = ~n4869 & n5158;
  assign n5160 = n4869 & ~n5158;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = ~n4867 & n5161;
  assign n5163 = ~n4854 & ~n5161;
  assign n5164 = ~n4866 & n5163;
  assign po30 = ~n5162 & ~n5164;
  assign n5166 = n4855 & n5161;
  assign n5167 = n4271 & n5166;
  assign n5168 = n4568 & n5167;
  assign n5169 = ~n3455 & n5168;
  assign n5170 = ~n4550 & n5166;
  assign n5171 = ~n4561 & n5170;
  assign n5172 = ~n4854 & ~n5159;
  assign n5173 = ~n5160 & ~n5172;
  assign n5174 = ~n4928 & ~n4933;
  assign n5175 = ~n4926 & ~n5174;
  assign n5176 = pi62 & ~pi63;
  assign n5177 = ~pi62 & pi63;
  assign n5178 = ~n5176 & ~n5177;
  assign n5179 = pi00 & ~n5091;
  assign n5180 = ~n5092 & n5179;
  assign n5181 = ~n5178 & n5180;
  assign n5182 = pi01 & ~n5093;
  assign n5183 = ~n5181 & ~n5182;
  assign n5184 = pi63 & ~n5183;
  assign n5185 = ~pi63 & ~n5182;
  assign n5186 = ~n5181 & n5185;
  assign n5187 = ~n5184 & ~n5186;
  assign n5188 = pi02 & ~n4513;
  assign n5189 = ~n4514 & n5188;
  assign n5190 = ~n4577 & n5189;
  assign n5191 = pi03 & ~n4515;
  assign n5192 = ~n5190 & ~n5191;
  assign n5193 = pi61 & ~n5192;
  assign n5194 = ~pi61 & ~n5191;
  assign n5195 = ~n5190 & n5194;
  assign n5196 = ~n5193 & ~n5195;
  assign n5197 = n5187 & ~n5196;
  assign n5198 = ~n5187 & n5196;
  assign n5199 = pi04 & ~n3959;
  assign n5200 = ~n3960 & n5199;
  assign n5201 = ~n4233 & n5200;
  assign n5202 = pi05 & ~n3961;
  assign n5203 = ~n5201 & ~n5202;
  assign n5204 = pi59 & ~n5203;
  assign n5205 = ~pi59 & ~n5202;
  assign n5206 = ~n5201 & n5205;
  assign n5207 = ~n5204 & ~n5206;
  assign n5208 = ~n5198 & ~n5207;
  assign n5209 = ~n5197 & n5208;
  assign n5210 = ~n5197 & ~n5198;
  assign n5211 = n5207 & ~n5210;
  assign n5212 = ~n5108 & ~n5121;
  assign n5213 = ~n5211 & n5212;
  assign n5214 = ~n5209 & n5213;
  assign n5215 = ~n5209 & ~n5211;
  assign n5216 = ~n5212 & ~n5215;
  assign n5217 = ~n5214 & ~n5216;
  assign n5218 = pi63 & ~n4591;
  assign n5219 = ~n4589 & n5218;
  assign n5220 = n4598 & n5219;
  assign n5221 = ~n5131 & ~n5220;
  assign n5222 = ~n5217 & n5221;
  assign n5223 = n5217 & ~n5221;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5175 & n5224;
  assign n5226 = ~n4926 & ~n5224;
  assign n5227 = ~n5174 & n5226;
  assign n5228 = ~n5225 & ~n5227;
  assign n5229 = ~n4939 & n5085;
  assign n5230 = ~n4938 & ~n5229;
  assign n5231 = n5228 & ~n5230;
  assign n5232 = ~n5003 & ~n5084;
  assign n5233 = ~n4884 & ~n4922;
  assign n5234 = pi06 & ~n3205;
  assign n5235 = ~n3206 & n5234;
  assign n5236 = ~n3463 & n5235;
  assign n5237 = pi07 & ~n3207;
  assign n5238 = ~n5236 & ~n5237;
  assign n5239 = pi57 & ~n5238;
  assign n5240 = ~pi57 & ~n5237;
  assign n5241 = ~n5236 & n5240;
  assign n5242 = ~n5239 & ~n5241;
  assign n5243 = ~n4907 & n4917;
  assign n5244 = ~n4904 & ~n5243;
  assign n5245 = n5242 & ~n5244;
  assign n5246 = pi08 & ~n2876;
  assign n5247 = ~n2877 & n5246;
  assign n5248 = ~n2960 & n5247;
  assign n5249 = pi09 & ~n2878;
  assign n5250 = ~n5248 & ~n5249;
  assign n5251 = pi55 & ~n5250;
  assign n5252 = pi10 & ~n2288;
  assign n5253 = ~n2289 & n5252;
  assign n5254 = ~n2647 & n5253;
  assign n5255 = pi11 & ~n2290;
  assign n5256 = ~n5254 & ~n5255;
  assign n5257 = pi53 & ~n5256;
  assign n5258 = ~pi53 & ~n5255;
  assign n5259 = ~n5254 & n5258;
  assign n5260 = ~pi55 & ~n5249;
  assign n5261 = ~n5248 & n5260;
  assign n5262 = ~n5259 & ~n5261;
  assign n5263 = ~n5257 & n5262;
  assign n5264 = ~n5251 & n5263;
  assign n5265 = ~n5257 & ~n5259;
  assign n5266 = ~n5251 & ~n5261;
  assign n5267 = ~n5265 & ~n5266;
  assign n5268 = ~n5264 & ~n5267;
  assign n5269 = pi12 & ~n2023;
  assign n5270 = ~n2024 & n5269;
  assign n5271 = ~n2079 & n5270;
  assign n5272 = pi13 & ~n2025;
  assign n5273 = ~n5271 & ~n5272;
  assign n5274 = pi51 & ~n5273;
  assign n5275 = ~pi51 & ~n5272;
  assign n5276 = ~n5271 & n5275;
  assign n5277 = ~n5274 & ~n5276;
  assign n5278 = ~n5268 & n5277;
  assign n5279 = ~n5264 & ~n5277;
  assign n5280 = ~n5267 & n5279;
  assign n5281 = ~n5278 & ~n5280;
  assign n5282 = ~n4904 & ~n5242;
  assign n5283 = ~n5243 & n5282;
  assign n5284 = ~n5281 & ~n5283;
  assign n5285 = ~n5245 & n5284;
  assign n5286 = ~n5245 & ~n5283;
  assign n5287 = n5281 & ~n5286;
  assign n5288 = ~n5285 & ~n5287;
  assign n5289 = ~n5233 & n5288;
  assign n5290 = n5233 & ~n5288;
  assign n5291 = ~n5289 & ~n5290;
  assign n5292 = ~n4976 & ~n4985;
  assign n5293 = ~n4975 & n4993;
  assign n5294 = ~n4983 & ~n5293;
  assign n5295 = ~n5292 & ~n5294;
  assign n5296 = ~n5291 & n5295;
  assign n5297 = ~n5289 & ~n5295;
  assign n5298 = ~n5290 & n5297;
  assign n5299 = ~n5296 & ~n5298;
  assign n5300 = n5232 & ~n5299;
  assign n5301 = ~n5232 & n5299;
  assign n5302 = ~n5046 & n5078;
  assign n5303 = ~n5045 & ~n5302;
  assign n5304 = pi14 & ~n1607;
  assign n5305 = ~n1608 & n5304;
  assign n5306 = ~n1782 & n5305;
  assign n5307 = pi15 & ~n1609;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = pi49 & ~n5308;
  assign n5310 = pi16 & ~n1212;
  assign n5311 = ~n1213 & n5310;
  assign n5312 = ~n1425 & n5311;
  assign n5313 = pi17 & ~n1214;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = pi47 & ~n5314;
  assign n5316 = ~pi47 & ~n5313;
  assign n5317 = ~n5312 & n5316;
  assign n5318 = ~pi49 & ~n5307;
  assign n5319 = ~n5306 & n5318;
  assign n5320 = ~n5317 & ~n5319;
  assign n5321 = ~n5315 & n5320;
  assign n5322 = ~n5309 & n5321;
  assign n5323 = ~n5315 & ~n5317;
  assign n5324 = ~n5309 & ~n5319;
  assign n5325 = ~n5323 & ~n5324;
  assign n5326 = ~n5322 & ~n5325;
  assign n5327 = pi18 & ~n1006;
  assign n5328 = ~n1007 & n5327;
  assign n5329 = ~n1068 & n5328;
  assign n5330 = pi19 & ~n1008;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = pi45 & ~n5331;
  assign n5333 = ~pi45 & ~n5330;
  assign n5334 = ~n5329 & n5333;
  assign n5335 = ~n5332 & ~n5334;
  assign n5336 = ~n5326 & n5335;
  assign n5337 = ~n4962 & n4972;
  assign n5338 = ~n4959 & ~n5337;
  assign n5339 = ~n5336 & n5338;
  assign n5340 = ~n5322 & ~n5335;
  assign n5341 = ~n5325 & n5340;
  assign n5342 = ~n5030 & n5040;
  assign n5343 = ~n5027 & ~n5342;
  assign n5344 = ~n5341 & ~n5343;
  assign n5345 = n5339 & n5344;
  assign n5346 = ~n5336 & n5343;
  assign n5347 = ~n5338 & ~n5341;
  assign n5348 = n5346 & n5347;
  assign n5349 = ~n5345 & ~n5348;
  assign n5350 = ~n5336 & ~n5341;
  assign n5351 = ~n5338 & ~n5343;
  assign n5352 = ~n5350 & n5351;
  assign n5353 = ~n4959 & ~n5027;
  assign n5354 = ~n5342 & n5353;
  assign n5355 = ~n5337 & n5354;
  assign n5356 = ~n5350 & n5355;
  assign n5357 = ~n5352 & ~n5356;
  assign n5358 = n5349 & n5357;
  assign n5359 = ~n5303 & ~n5358;
  assign n5360 = ~n5055 & ~n5064;
  assign n5361 = ~n5062 & n5360;
  assign n5362 = ~n5053 & n5361;
  assign n5363 = ~n5077 & ~n5362;
  assign n5364 = pi20 & ~n683;
  assign n5365 = ~n684 & n5364;
  assign n5366 = ~n1231 & n5365;
  assign n5367 = pi21 & ~n685;
  assign n5368 = ~n5366 & ~n5367;
  assign n5369 = pi43 & ~n5368;
  assign n5370 = pi22 & ~n489;
  assign n5371 = ~n490 & n5370;
  assign n5372 = ~n572 & n5371;
  assign n5373 = pi23 & ~n491;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = pi41 & ~n5374;
  assign n5376 = ~pi41 & ~n5373;
  assign n5377 = ~n5372 & n5376;
  assign n5378 = ~pi43 & ~n5367;
  assign n5379 = ~n5366 & n5378;
  assign n5380 = ~n5377 & ~n5379;
  assign n5381 = ~n5375 & n5380;
  assign n5382 = ~n5369 & n5381;
  assign n5383 = ~n5375 & ~n5377;
  assign n5384 = ~n5369 & ~n5379;
  assign n5385 = ~n5383 & ~n5384;
  assign n5386 = ~n5382 & ~n5385;
  assign n5387 = pi24 & ~n304;
  assign n5388 = ~n305 & n5387;
  assign n5389 = ~n394 & n5388;
  assign n5390 = pi25 & ~n306;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = pi39 & ~n5391;
  assign n5393 = ~pi39 & ~n5390;
  assign n5394 = ~n5389 & n5393;
  assign n5395 = ~n5392 & ~n5394;
  assign n5396 = ~n5386 & n5395;
  assign n5397 = ~n5382 & ~n5395;
  assign n5398 = ~n5385 & n5397;
  assign n5399 = ~n5396 & ~n5398;
  assign n5400 = ~n5363 & ~n5399;
  assign n5401 = n5363 & n5399;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = pi26 & ~n193;
  assign n5404 = ~n194 & n5403;
  assign n5405 = ~n729 & n5404;
  assign n5406 = pi27 & ~n195;
  assign n5407 = ~n5405 & ~n5406;
  assign n5408 = pi37 & ~n5407;
  assign n5409 = ~pi37 & ~n5406;
  assign n5410 = ~n5405 & n5409;
  assign n5411 = ~n5408 & ~n5410;
  assign n5412 = pi28 & ~n141;
  assign n5413 = ~n142 & n5412;
  assign n5414 = ~n156 & n5413;
  assign n5415 = pi29 & ~n143;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = pi35 & ~n5416;
  assign n5418 = ~pi35 & ~n5415;
  assign n5419 = ~n5414 & n5418;
  assign n5420 = ~n5417 & ~n5419;
  assign n5421 = ~n5411 & n5420;
  assign n5422 = n5411 & ~n5420;
  assign n5423 = ~n5421 & ~n5422;
  assign n5424 = pi30 & ~pi32;
  assign n5425 = pi33 & n5424;
  assign n5426 = pi31 & pi32;
  assign n5427 = ~pi33 & n5426;
  assign n5428 = ~pi32 & pi33;
  assign n5429 = ~pi31 & pi33;
  assign n5430 = ~n5428 & ~n5429;
  assign n5431 = ~n5427 & n5430;
  assign n5432 = ~n5425 & ~n5431;
  assign n5433 = ~n5423 & n5432;
  assign n5434 = ~n5421 & ~n5432;
  assign n5435 = ~n5422 & n5434;
  assign n5436 = ~n5433 & ~n5435;
  assign n5437 = ~n5402 & n5436;
  assign n5438 = ~n5400 & ~n5436;
  assign n5439 = ~n5401 & n5438;
  assign n5440 = ~n5437 & ~n5439;
  assign n5441 = ~n5348 & ~n5352;
  assign n5442 = ~n5356 & n5441;
  assign n5443 = ~n5045 & ~n5345;
  assign n5444 = ~n5302 & n5443;
  assign n5445 = n5442 & n5444;
  assign n5446 = ~n5440 & ~n5445;
  assign n5447 = ~n5359 & n5446;
  assign n5448 = ~n5359 & ~n5445;
  assign n5449 = n5440 & ~n5448;
  assign n5450 = ~n5447 & ~n5449;
  assign n5451 = ~n5301 & ~n5450;
  assign n5452 = ~n5300 & n5451;
  assign n5453 = ~n4938 & ~n5228;
  assign n5454 = ~n5229 & n5453;
  assign n5455 = ~n5300 & ~n5301;
  assign n5456 = n5450 & ~n5455;
  assign n5457 = ~n5454 & ~n5456;
  assign n5458 = ~n5452 & n5457;
  assign n5459 = ~n5231 & n5458;
  assign n5460 = ~n5231 & ~n5454;
  assign n5461 = ~n5452 & ~n5456;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = ~n5459 & ~n5462;
  assign n5464 = ~n5089 & ~n5145;
  assign n5465 = n4606 & ~n5131;
  assign n5466 = ~n5130 & n5465;
  assign n5467 = ~n5141 & ~n5466;
  assign n5468 = ~n5143 & ~n5467;
  assign n5469 = ~n5464 & n5468;
  assign n5470 = ~n5143 & ~n5464;
  assign n5471 = n5467 & ~n5470;
  assign n5472 = ~n5469 & ~n5471;
  assign n5473 = ~n5463 & ~n5472;
  assign n5474 = n5463 & n5472;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = n4608 & ~n4613;
  assign n5477 = ~n5150 & n5476;
  assign n5478 = ~n5156 & ~n5477;
  assign n5479 = ~n5475 & n5478;
  assign n5480 = n5475 & ~n5478;
  assign n5481 = ~n5479 & ~n5480;
  assign n5482 = ~n5173 & ~n5481;
  assign n5483 = ~n5171 & n5482;
  assign n5484 = ~n5169 & n5483;
  assign n5485 = ~n5171 & ~n5173;
  assign n5486 = ~n5169 & n5485;
  assign n5487 = n5481 & ~n5486;
  assign po31 = ~n5484 & ~n5487;
  assign n5489 = n3454 & ~n4861;
  assign n5490 = ~n4550 & ~n5479;
  assign n5491 = ~n5480 & n5490;
  assign n5492 = n4271 & n4567;
  assign n5493 = n5166 & n5492;
  assign n5494 = n5491 & n5493;
  assign n5495 = ~n5489 & n5494;
  assign n5496 = ~n4270 & ~n4559;
  assign n5497 = n4551 & n5481;
  assign n5498 = n5166 & n5497;
  assign n5499 = ~n5496 & n5498;
  assign n5500 = n4549 & n5166;
  assign n5501 = ~n5173 & ~n5480;
  assign n5502 = ~n5500 & n5501;
  assign n5503 = ~n5479 & ~n5502;
  assign n5504 = ~n5499 & ~n5503;
  assign n5505 = ~n5495 & n5504;
  assign n5506 = ~n5467 & ~n5470;
  assign n5507 = ~n5473 & ~n5506;
  assign n5508 = ~n5231 & n5461;
  assign n5509 = ~n5454 & ~n5508;
  assign n5510 = ~n5223 & ~n5225;
  assign n5511 = ~n5509 & n5510;
  assign n5512 = ~n5359 & ~n5447;
  assign n5513 = ~n5245 & ~n5285;
  assign n5514 = pi07 & ~n3205;
  assign n5515 = ~n3206 & n5514;
  assign n5516 = ~n3463 & n5515;
  assign n5517 = pi08 & ~n3207;
  assign n5518 = ~n5516 & ~n5517;
  assign n5519 = pi57 & ~n5518;
  assign n5520 = ~pi57 & ~n5517;
  assign n5521 = ~n5516 & n5520;
  assign n5522 = ~n5519 & ~n5521;
  assign n5523 = ~n5267 & n5277;
  assign n5524 = ~n5264 & ~n5523;
  assign n5525 = n5522 & ~n5524;
  assign n5526 = pi09 & ~n2876;
  assign n5527 = ~n2877 & n5526;
  assign n5528 = ~n2960 & n5527;
  assign n5529 = pi10 & ~n2878;
  assign n5530 = ~n5528 & ~n5529;
  assign n5531 = pi55 & ~n5530;
  assign n5532 = pi11 & ~n2288;
  assign n5533 = ~n2289 & n5532;
  assign n5534 = ~n2647 & n5533;
  assign n5535 = pi12 & ~n2290;
  assign n5536 = ~n5534 & ~n5535;
  assign n5537 = pi53 & ~n5536;
  assign n5538 = ~pi53 & ~n5535;
  assign n5539 = ~n5534 & n5538;
  assign n5540 = ~pi55 & ~n5529;
  assign n5541 = ~n5528 & n5540;
  assign n5542 = ~n5539 & ~n5541;
  assign n5543 = ~n5537 & n5542;
  assign n5544 = ~n5531 & n5543;
  assign n5545 = ~n5537 & ~n5539;
  assign n5546 = ~n5531 & ~n5541;
  assign n5547 = ~n5545 & ~n5546;
  assign n5548 = ~n5544 & ~n5547;
  assign n5549 = pi13 & ~n2023;
  assign n5550 = ~n2024 & n5549;
  assign n5551 = ~n2079 & n5550;
  assign n5552 = pi14 & ~n2025;
  assign n5553 = ~n5551 & ~n5552;
  assign n5554 = pi51 & ~n5553;
  assign n5555 = ~pi51 & ~n5552;
  assign n5556 = ~n5551 & n5555;
  assign n5557 = ~n5554 & ~n5556;
  assign n5558 = ~n5548 & n5557;
  assign n5559 = ~n5544 & ~n5557;
  assign n5560 = ~n5547 & n5559;
  assign n5561 = ~n5558 & ~n5560;
  assign n5562 = ~n5264 & ~n5522;
  assign n5563 = ~n5523 & n5562;
  assign n5564 = ~n5561 & ~n5563;
  assign n5565 = ~n5525 & n5564;
  assign n5566 = ~n5525 & ~n5563;
  assign n5567 = n5561 & ~n5566;
  assign n5568 = ~n5565 & ~n5567;
  assign n5569 = ~n5513 & n5568;
  assign n5570 = n5513 & ~n5568;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = ~n5338 & ~n5350;
  assign n5573 = n5339 & ~n5341;
  assign n5574 = ~n5343 & ~n5573;
  assign n5575 = ~n5572 & ~n5574;
  assign n5576 = ~n5571 & n5575;
  assign n5577 = ~n5569 & ~n5575;
  assign n5578 = ~n5570 & n5577;
  assign n5579 = ~n5576 & ~n5578;
  assign n5580 = ~n5512 & n5579;
  assign n5581 = n5512 & ~n5579;
  assign n5582 = ~n5580 & ~n5581;
  assign n5583 = ~n5401 & n5436;
  assign n5584 = ~n5400 & ~n5583;
  assign n5585 = pi15 & ~n1607;
  assign n5586 = ~n1608 & n5585;
  assign n5587 = ~n1782 & n5586;
  assign n5588 = pi16 & ~n1609;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = pi49 & ~n5589;
  assign n5591 = pi17 & ~n1212;
  assign n5592 = ~n1213 & n5591;
  assign n5593 = ~n1425 & n5592;
  assign n5594 = pi18 & ~n1214;
  assign n5595 = ~n5593 & ~n5594;
  assign n5596 = pi47 & ~n5595;
  assign n5597 = ~pi47 & ~n5594;
  assign n5598 = ~n5593 & n5597;
  assign n5599 = ~pi49 & ~n5588;
  assign n5600 = ~n5587 & n5599;
  assign n5601 = ~n5598 & ~n5600;
  assign n5602 = ~n5596 & n5601;
  assign n5603 = ~n5590 & n5602;
  assign n5604 = ~n5596 & ~n5598;
  assign n5605 = ~n5590 & ~n5600;
  assign n5606 = ~n5604 & ~n5605;
  assign n5607 = ~n5603 & ~n5606;
  assign n5608 = pi19 & ~n1006;
  assign n5609 = ~n1007 & n5608;
  assign n5610 = ~n1068 & n5609;
  assign n5611 = pi20 & ~n1008;
  assign n5612 = ~n5610 & ~n5611;
  assign n5613 = pi45 & ~n5612;
  assign n5614 = ~pi45 & ~n5611;
  assign n5615 = ~n5610 & n5614;
  assign n5616 = ~n5613 & ~n5615;
  assign n5617 = ~n5607 & n5616;
  assign n5618 = ~n5325 & n5335;
  assign n5619 = ~n5322 & ~n5618;
  assign n5620 = ~n5617 & n5619;
  assign n5621 = ~n5603 & ~n5616;
  assign n5622 = ~n5606 & n5621;
  assign n5623 = ~n5385 & n5395;
  assign n5624 = ~n5382 & ~n5623;
  assign n5625 = ~n5622 & ~n5624;
  assign n5626 = n5620 & n5625;
  assign n5627 = ~n5617 & n5624;
  assign n5628 = ~n5619 & ~n5622;
  assign n5629 = n5627 & n5628;
  assign n5630 = ~n5626 & ~n5629;
  assign n5631 = ~n5617 & ~n5622;
  assign n5632 = ~n5619 & ~n5624;
  assign n5633 = ~n5631 & n5632;
  assign n5634 = ~n5322 & ~n5382;
  assign n5635 = ~n5623 & n5634;
  assign n5636 = ~n5618 & n5635;
  assign n5637 = ~n5631 & n5636;
  assign n5638 = ~n5633 & ~n5637;
  assign n5639 = n5630 & n5638;
  assign n5640 = ~n5584 & ~n5639;
  assign n5641 = ~n5410 & ~n5419;
  assign n5642 = ~n5417 & n5641;
  assign n5643 = ~n5408 & n5642;
  assign n5644 = ~n5433 & ~n5643;
  assign n5645 = pi21 & ~n683;
  assign n5646 = ~n684 & n5645;
  assign n5647 = ~n1231 & n5646;
  assign n5648 = pi22 & ~n685;
  assign n5649 = ~n5647 & ~n5648;
  assign n5650 = pi43 & ~n5649;
  assign n5651 = pi23 & ~n489;
  assign n5652 = ~n490 & n5651;
  assign n5653 = ~n572 & n5652;
  assign n5654 = pi24 & ~n491;
  assign n5655 = ~n5653 & ~n5654;
  assign n5656 = pi41 & ~n5655;
  assign n5657 = ~pi41 & ~n5654;
  assign n5658 = ~n5653 & n5657;
  assign n5659 = ~pi43 & ~n5648;
  assign n5660 = ~n5647 & n5659;
  assign n5661 = ~n5658 & ~n5660;
  assign n5662 = ~n5656 & n5661;
  assign n5663 = ~n5650 & n5662;
  assign n5664 = ~n5656 & ~n5658;
  assign n5665 = ~n5650 & ~n5660;
  assign n5666 = ~n5664 & ~n5665;
  assign n5667 = ~n5663 & ~n5666;
  assign n5668 = pi25 & ~n304;
  assign n5669 = ~n305 & n5668;
  assign n5670 = ~n394 & n5669;
  assign n5671 = pi26 & ~n306;
  assign n5672 = ~n5670 & ~n5671;
  assign n5673 = pi39 & ~n5672;
  assign n5674 = ~pi39 & ~n5671;
  assign n5675 = ~n5670 & n5674;
  assign n5676 = ~n5673 & ~n5675;
  assign n5677 = ~n5667 & n5676;
  assign n5678 = ~n5663 & ~n5676;
  assign n5679 = ~n5666 & n5678;
  assign n5680 = ~n5677 & ~n5679;
  assign n5681 = ~n5644 & ~n5680;
  assign n5682 = n5644 & n5680;
  assign n5683 = ~n5681 & ~n5682;
  assign n5684 = pi27 & ~n193;
  assign n5685 = ~n194 & n5684;
  assign n5686 = ~n729 & n5685;
  assign n5687 = pi28 & ~n195;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = pi37 & ~n5688;
  assign n5690 = ~pi37 & ~n5687;
  assign n5691 = ~n5686 & n5690;
  assign n5692 = ~n5689 & ~n5691;
  assign n5693 = pi29 & ~n141;
  assign n5694 = ~n142 & n5693;
  assign n5695 = ~n156 & n5694;
  assign n5696 = pi30 & ~n143;
  assign n5697 = ~n5695 & ~n5696;
  assign n5698 = pi35 & ~n5697;
  assign n5699 = ~pi35 & ~n5696;
  assign n5700 = ~n5695 & n5699;
  assign n5701 = ~n5698 & ~n5700;
  assign n5702 = n5692 & ~n5701;
  assign n5703 = ~n5427 & ~n5429;
  assign n5704 = ~n5692 & n5701;
  assign n5705 = ~n5703 & ~n5704;
  assign n5706 = ~n5702 & n5705;
  assign n5707 = ~n5702 & ~n5704;
  assign n5708 = n5703 & ~n5707;
  assign n5709 = ~n5706 & ~n5708;
  assign n5710 = ~n5683 & n5709;
  assign n5711 = ~n5681 & ~n5709;
  assign n5712 = ~n5682 & n5711;
  assign n5713 = ~n5710 & ~n5712;
  assign n5714 = ~n5629 & ~n5633;
  assign n5715 = ~n5637 & n5714;
  assign n5716 = ~n5400 & ~n5626;
  assign n5717 = ~n5583 & n5716;
  assign n5718 = n5715 & n5717;
  assign n5719 = ~n5713 & ~n5718;
  assign n5720 = ~n5640 & n5719;
  assign n5721 = ~n5640 & ~n5718;
  assign n5722 = n5713 & ~n5721;
  assign n5723 = ~n5720 & ~n5722;
  assign n5724 = ~n5582 & n5723;
  assign n5725 = ~n5580 & ~n5723;
  assign n5726 = ~n5581 & n5725;
  assign n5727 = ~n5724 & ~n5726;
  assign n5728 = ~n5300 & n5450;
  assign n5729 = ~n5301 & ~n5728;
  assign n5730 = ~n5290 & ~n5295;
  assign n5731 = ~n5186 & ~n5195;
  assign n5732 = ~n5193 & n5731;
  assign n5733 = ~n5184 & n5732;
  assign n5734 = ~n5211 & ~n5733;
  assign n5735 = pi01 & ~n5091;
  assign n5736 = ~n5092 & n5735;
  assign n5737 = ~n5178 & n5736;
  assign n5738 = pi02 & ~n5093;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = pi63 & ~n5739;
  assign n5741 = ~pi63 & ~n5738;
  assign n5742 = ~n5737 & n5741;
  assign n5743 = ~n5740 & ~n5742;
  assign n5744 = pi03 & ~n4513;
  assign n5745 = ~n4514 & n5744;
  assign n5746 = ~n4577 & n5745;
  assign n5747 = pi04 & ~n4515;
  assign n5748 = ~n5746 & ~n5747;
  assign n5749 = pi61 & ~n5748;
  assign n5750 = ~pi61 & ~n5747;
  assign n5751 = ~n5746 & n5750;
  assign n5752 = ~n5749 & ~n5751;
  assign n5753 = ~n5743 & n5752;
  assign n5754 = n5743 & ~n5752;
  assign n5755 = ~n5753 & ~n5754;
  assign n5756 = pi05 & ~n3959;
  assign n5757 = ~n3960 & n5756;
  assign n5758 = ~n4233 & n5757;
  assign n5759 = pi06 & ~n3961;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = pi59 & ~n5760;
  assign n5762 = ~pi59 & ~n5759;
  assign n5763 = ~n5758 & n5762;
  assign n5764 = ~n5761 & ~n5763;
  assign n5765 = ~n5755 & n5764;
  assign n5766 = ~n5753 & ~n5764;
  assign n5767 = ~n5754 & n5766;
  assign n5768 = ~n5765 & ~n5767;
  assign n5769 = ~n5734 & n5768;
  assign n5770 = n5734 & ~n5768;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = n5214 & ~n5771;
  assign n5773 = ~n5214 & ~n5769;
  assign n5774 = ~n5770 & n5773;
  assign n5775 = ~n5772 & ~n5774;
  assign n5776 = ~n5289 & ~n5775;
  assign n5777 = ~n5730 & n5776;
  assign n5778 = ~n5289 & ~n5730;
  assign n5779 = n5775 & ~n5778;
  assign n5780 = ~n5777 & ~n5779;
  assign n5781 = ~n5729 & n5780;
  assign n5782 = ~n5301 & ~n5780;
  assign n5783 = ~n5728 & n5782;
  assign n5784 = ~n5781 & ~n5783;
  assign n5785 = ~n5727 & ~n5784;
  assign n5786 = n5727 & n5784;
  assign n5787 = ~n5785 & ~n5786;
  assign n5788 = ~n5454 & ~n5510;
  assign n5789 = ~n5508 & n5788;
  assign n5790 = ~n5787 & ~n5789;
  assign n5791 = ~n5511 & n5790;
  assign n5792 = ~n5511 & ~n5789;
  assign n5793 = n5787 & ~n5792;
  assign n5794 = ~n5791 & ~n5793;
  assign n5795 = ~n5507 & n5794;
  assign n5796 = n5507 & ~n5794;
  assign n5797 = ~n5795 & ~n5796;
  assign n5798 = ~n5505 & n5797;
  assign n5799 = ~n5499 & ~n5797;
  assign n5800 = ~n5503 & n5799;
  assign n5801 = ~n5495 & n5800;
  assign po32 = ~n5798 & ~n5801;
  assign n5803 = n5167 & n5497;
  assign n5804 = ~n3992 & n5803;
  assign n5805 = ~n4269 & ~n5480;
  assign n5806 = n5490 & n5805;
  assign n5807 = ~n5160 & n5172;
  assign n5808 = ~n4260 & ~n4853;
  assign n5809 = ~n4549 & n5808;
  assign n5810 = n5807 & n5809;
  assign n5811 = n5806 & n5810;
  assign n5812 = ~n5503 & ~n5811;
  assign n5813 = ~n5804 & n5812;
  assign n5814 = ~n5796 & ~n5813;
  assign n5815 = ~n5795 & ~n5814;
  assign n5816 = ~n5640 & ~n5720;
  assign n5817 = ~n5525 & ~n5565;
  assign n5818 = pi08 & ~n3205;
  assign n5819 = ~n3206 & n5818;
  assign n5820 = ~n3463 & n5819;
  assign n5821 = pi09 & ~n3207;
  assign n5822 = ~n5820 & ~n5821;
  assign n5823 = pi57 & ~n5822;
  assign n5824 = ~pi57 & ~n5821;
  assign n5825 = ~n5820 & n5824;
  assign n5826 = ~n5823 & ~n5825;
  assign n5827 = ~n5547 & n5557;
  assign n5828 = ~n5544 & ~n5827;
  assign n5829 = n5826 & ~n5828;
  assign n5830 = pi10 & ~n2876;
  assign n5831 = ~n2877 & n5830;
  assign n5832 = ~n2960 & n5831;
  assign n5833 = pi11 & ~n2878;
  assign n5834 = ~n5832 & ~n5833;
  assign n5835 = pi55 & ~n5834;
  assign n5836 = pi12 & ~n2288;
  assign n5837 = ~n2289 & n5836;
  assign n5838 = ~n2647 & n5837;
  assign n5839 = pi13 & ~n2290;
  assign n5840 = ~n5838 & ~n5839;
  assign n5841 = pi53 & ~n5840;
  assign n5842 = ~pi53 & ~n5839;
  assign n5843 = ~n5838 & n5842;
  assign n5844 = ~pi55 & ~n5833;
  assign n5845 = ~n5832 & n5844;
  assign n5846 = ~n5843 & ~n5845;
  assign n5847 = ~n5841 & n5846;
  assign n5848 = ~n5835 & n5847;
  assign n5849 = ~n5841 & ~n5843;
  assign n5850 = ~n5835 & ~n5845;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = ~n5848 & ~n5851;
  assign n5853 = pi14 & ~n2023;
  assign n5854 = ~n2024 & n5853;
  assign n5855 = ~n2079 & n5854;
  assign n5856 = pi15 & ~n2025;
  assign n5857 = ~n5855 & ~n5856;
  assign n5858 = pi51 & ~n5857;
  assign n5859 = ~pi51 & ~n5856;
  assign n5860 = ~n5855 & n5859;
  assign n5861 = ~n5858 & ~n5860;
  assign n5862 = ~n5852 & n5861;
  assign n5863 = ~n5848 & ~n5861;
  assign n5864 = ~n5851 & n5863;
  assign n5865 = ~n5862 & ~n5864;
  assign n5866 = ~n5544 & ~n5826;
  assign n5867 = ~n5827 & n5866;
  assign n5868 = ~n5865 & ~n5867;
  assign n5869 = ~n5829 & n5868;
  assign n5870 = ~n5829 & ~n5867;
  assign n5871 = n5865 & ~n5870;
  assign n5872 = ~n5869 & ~n5871;
  assign n5873 = ~n5817 & n5872;
  assign n5874 = n5817 & ~n5872;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n5619 & ~n5631;
  assign n5877 = n5620 & ~n5622;
  assign n5878 = ~n5624 & ~n5877;
  assign n5879 = ~n5876 & ~n5878;
  assign n5880 = ~n5875 & n5879;
  assign n5881 = ~n5873 & ~n5879;
  assign n5882 = ~n5874 & n5881;
  assign n5883 = ~n5880 & ~n5882;
  assign n5884 = ~n5816 & n5883;
  assign n5885 = n5816 & ~n5883;
  assign n5886 = ~n5884 & ~n5885;
  assign n5887 = ~n5682 & n5709;
  assign n5888 = ~n5681 & ~n5887;
  assign n5889 = pi16 & ~n1607;
  assign n5890 = ~n1608 & n5889;
  assign n5891 = ~n1782 & n5890;
  assign n5892 = pi17 & ~n1609;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = pi49 & ~n5893;
  assign n5895 = pi18 & ~n1212;
  assign n5896 = ~n1213 & n5895;
  assign n5897 = ~n1425 & n5896;
  assign n5898 = pi19 & ~n1214;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = pi47 & ~n5899;
  assign n5901 = ~pi47 & ~n5898;
  assign n5902 = ~n5897 & n5901;
  assign n5903 = ~pi49 & ~n5892;
  assign n5904 = ~n5891 & n5903;
  assign n5905 = ~n5902 & ~n5904;
  assign n5906 = ~n5900 & n5905;
  assign n5907 = ~n5894 & n5906;
  assign n5908 = ~n5900 & ~n5902;
  assign n5909 = ~n5894 & ~n5904;
  assign n5910 = ~n5908 & ~n5909;
  assign n5911 = ~n5907 & ~n5910;
  assign n5912 = pi20 & ~n1006;
  assign n5913 = ~n1007 & n5912;
  assign n5914 = ~n1068 & n5913;
  assign n5915 = pi21 & ~n1008;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = pi45 & ~n5916;
  assign n5918 = ~pi45 & ~n5915;
  assign n5919 = ~n5914 & n5918;
  assign n5920 = ~n5917 & ~n5919;
  assign n5921 = ~n5911 & n5920;
  assign n5922 = ~n5606 & n5616;
  assign n5923 = ~n5603 & ~n5922;
  assign n5924 = ~n5921 & n5923;
  assign n5925 = ~n5907 & ~n5920;
  assign n5926 = ~n5910 & n5925;
  assign n5927 = ~n5666 & n5676;
  assign n5928 = ~n5663 & ~n5927;
  assign n5929 = ~n5926 & ~n5928;
  assign n5930 = n5924 & n5929;
  assign n5931 = ~n5921 & n5928;
  assign n5932 = ~n5923 & ~n5926;
  assign n5933 = n5931 & n5932;
  assign n5934 = ~n5930 & ~n5933;
  assign n5935 = ~n5921 & ~n5926;
  assign n5936 = ~n5923 & ~n5928;
  assign n5937 = ~n5935 & n5936;
  assign n5938 = ~n5603 & ~n5663;
  assign n5939 = ~n5927 & n5938;
  assign n5940 = ~n5922 & n5939;
  assign n5941 = ~n5935 & n5940;
  assign n5942 = ~n5937 & ~n5941;
  assign n5943 = n5934 & n5942;
  assign n5944 = ~n5888 & ~n5943;
  assign n5945 = ~n5933 & ~n5937;
  assign n5946 = ~n5941 & n5945;
  assign n5947 = ~n5681 & ~n5930;
  assign n5948 = ~n5887 & n5947;
  assign n5949 = n5946 & n5948;
  assign n5950 = ~n5691 & ~n5700;
  assign n5951 = ~n5698 & n5950;
  assign n5952 = ~n5689 & n5951;
  assign n5953 = ~n5708 & ~n5952;
  assign n5954 = pi22 & ~n683;
  assign n5955 = ~n684 & n5954;
  assign n5956 = ~n1231 & n5955;
  assign n5957 = pi23 & ~n685;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = pi43 & ~n5958;
  assign n5960 = pi24 & ~n489;
  assign n5961 = ~n490 & n5960;
  assign n5962 = ~n572 & n5961;
  assign n5963 = pi25 & ~n491;
  assign n5964 = ~n5962 & ~n5963;
  assign n5965 = pi41 & ~n5964;
  assign n5966 = ~pi41 & ~n5963;
  assign n5967 = ~n5962 & n5966;
  assign n5968 = ~pi43 & ~n5957;
  assign n5969 = ~n5956 & n5968;
  assign n5970 = ~n5967 & ~n5969;
  assign n5971 = ~n5965 & n5970;
  assign n5972 = ~n5959 & n5971;
  assign n5973 = ~n5965 & ~n5967;
  assign n5974 = ~n5959 & ~n5969;
  assign n5975 = ~n5973 & ~n5974;
  assign n5976 = ~n5972 & ~n5975;
  assign n5977 = pi26 & ~n304;
  assign n5978 = ~n305 & n5977;
  assign n5979 = ~n394 & n5978;
  assign n5980 = pi27 & ~n306;
  assign n5981 = ~n5979 & ~n5980;
  assign n5982 = pi39 & ~n5981;
  assign n5983 = ~pi39 & ~n5980;
  assign n5984 = ~n5979 & n5983;
  assign n5985 = ~n5982 & ~n5984;
  assign n5986 = ~n5976 & n5985;
  assign n5987 = ~n5972 & ~n5985;
  assign n5988 = ~n5975 & n5987;
  assign n5989 = ~n5986 & ~n5988;
  assign n5990 = n5953 & n5989;
  assign n5991 = ~n5953 & ~n5989;
  assign n5992 = pi30 & ~n141;
  assign n5993 = ~n142 & n5992;
  assign n5994 = ~n156 & n5993;
  assign n5995 = pi31 & ~n143;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = pi35 & ~n5996;
  assign n5998 = pi28 & ~n193;
  assign n5999 = ~n194 & n5998;
  assign n6000 = ~n729 & n5999;
  assign n6001 = pi29 & ~n195;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = pi37 & ~n6002;
  assign n6004 = ~pi37 & ~n6001;
  assign n6005 = ~n6000 & n6004;
  assign n6006 = ~pi35 & ~n5995;
  assign n6007 = ~n5994 & n6006;
  assign n6008 = ~n6005 & ~n6007;
  assign n6009 = ~n6003 & n6008;
  assign n6010 = ~n5997 & n6009;
  assign n6011 = ~n6003 & ~n6005;
  assign n6012 = ~n5997 & ~n6007;
  assign n6013 = ~n6011 & ~n6012;
  assign n6014 = ~n6010 & ~n6013;
  assign n6015 = ~n5991 & ~n6014;
  assign n6016 = ~n5990 & n6015;
  assign n6017 = ~n5990 & ~n5991;
  assign n6018 = n6014 & ~n6017;
  assign n6019 = ~n6016 & ~n6018;
  assign n6020 = ~n5949 & n6019;
  assign n6021 = ~n5944 & n6020;
  assign n6022 = ~n5944 & ~n5949;
  assign n6023 = ~n6019 & ~n6022;
  assign n6024 = ~n6021 & ~n6023;
  assign n6025 = ~n5886 & n6024;
  assign n6026 = ~n5884 & ~n6024;
  assign n6027 = ~n5885 & n6026;
  assign n6028 = ~n6025 & ~n6027;
  assign n6029 = ~n5581 & n5723;
  assign n6030 = ~n5570 & ~n5575;
  assign n6031 = ~n5569 & ~n6030;
  assign n6032 = ~n5742 & ~n5751;
  assign n6033 = ~n5749 & n6032;
  assign n6034 = ~n5740 & n6033;
  assign n6035 = ~n5765 & ~n6034;
  assign n6036 = pi02 & ~n5091;
  assign n6037 = ~n5092 & n6036;
  assign n6038 = ~n5178 & n6037;
  assign n6039 = pi03 & ~n5093;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = pi63 & ~n6040;
  assign n6042 = ~pi63 & ~n6039;
  assign n6043 = ~n6038 & n6042;
  assign n6044 = ~n6041 & ~n6043;
  assign n6045 = pi04 & ~n4513;
  assign n6046 = ~n4514 & n6045;
  assign n6047 = ~n4577 & n6046;
  assign n6048 = pi05 & ~n4515;
  assign n6049 = ~n6047 & ~n6048;
  assign n6050 = pi61 & ~n6049;
  assign n6051 = ~pi61 & ~n6048;
  assign n6052 = ~n6047 & n6051;
  assign n6053 = ~n6050 & ~n6052;
  assign n6054 = ~n6044 & n6053;
  assign n6055 = n6044 & ~n6053;
  assign n6056 = ~n6054 & ~n6055;
  assign n6057 = pi06 & ~n3959;
  assign n6058 = ~n3960 & n6057;
  assign n6059 = ~n4233 & n6058;
  assign n6060 = pi07 & ~n3961;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = pi59 & ~n6061;
  assign n6063 = ~pi59 & ~n6060;
  assign n6064 = ~n6059 & n6063;
  assign n6065 = ~n6062 & ~n6064;
  assign n6066 = ~n6056 & n6065;
  assign n6067 = ~n6054 & ~n6065;
  assign n6068 = ~n6055 & n6067;
  assign n6069 = ~n6066 & ~n6068;
  assign n6070 = ~n6035 & n6069;
  assign n6071 = n6035 & ~n6069;
  assign n6072 = ~n6070 & ~n6071;
  assign n6073 = n5770 & ~n6072;
  assign n6074 = ~n5770 & ~n6070;
  assign n6075 = ~n6071 & n6074;
  assign n6076 = ~n6073 & ~n6075;
  assign n6077 = ~n6031 & n6076;
  assign n6078 = ~n5569 & ~n6076;
  assign n6079 = ~n6030 & n6078;
  assign n6080 = ~n6077 & ~n6079;
  assign n6081 = ~n5580 & ~n6080;
  assign n6082 = ~n6029 & n6081;
  assign n6083 = ~n5580 & ~n6029;
  assign n6084 = n6080 & ~n6083;
  assign n6085 = ~n6082 & ~n6084;
  assign n6086 = ~n6028 & ~n6085;
  assign n6087 = n6028 & n6085;
  assign n6088 = ~n6086 & ~n6087;
  assign n6089 = ~n5727 & ~n5783;
  assign n6090 = ~n5772 & ~n5779;
  assign n6091 = ~n5781 & ~n6090;
  assign n6092 = ~n6089 & n6091;
  assign n6093 = ~n5781 & ~n6089;
  assign n6094 = n6090 & ~n6093;
  assign n6095 = ~n6092 & ~n6094;
  assign n6096 = ~n6088 & ~n6095;
  assign n6097 = n6088 & n6095;
  assign n6098 = ~n6096 & ~n6097;
  assign n6099 = ~n5789 & ~n5791;
  assign n6100 = ~n6098 & n6099;
  assign n6101 = n6098 & ~n6099;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = ~n5815 & n6102;
  assign n6104 = ~n5795 & ~n6102;
  assign n6105 = ~n5814 & n6104;
  assign po33 = ~n6103 & ~n6105;
  assign n6107 = ~n3707 & ~n3981;
  assign n6108 = ~n3982 & n6107;
  assign n6109 = n2710 & ~n2944;
  assign n6110 = n3724 & n6109;
  assign n6111 = n3452 & n6110;
  assign n6112 = n6108 & n6111;
  assign n6113 = ~n2713 & n6112;
  assign n6114 = n2707 & ~n3179;
  assign n6115 = ~n2944 & n6114;
  assign n6116 = n3443 & n6115;
  assign n6117 = n3725 & n6116;
  assign n6118 = ~n3982 & ~n6117;
  assign n6119 = ~n3723 & n6118;
  assign n6120 = ~n3981 & ~n6119;
  assign n6121 = ~n4261 & ~n6120;
  assign n6122 = ~n6113 & n6121;
  assign n6123 = ~n5796 & ~n6100;
  assign n6124 = ~n6101 & n6123;
  assign n6125 = ~n5480 & ~n5795;
  assign n6126 = n5490 & n6125;
  assign n6127 = ~n4263 & ~n4853;
  assign n6128 = ~n4549 & n6127;
  assign n6129 = n5807 & n6128;
  assign n6130 = n6126 & n6129;
  assign n6131 = n6124 & n6130;
  assign n6132 = ~n6122 & n6131;
  assign n6133 = ~n5795 & ~n6101;
  assign n6134 = ~n6100 & ~n6133;
  assign n6135 = ~n5479 & ~n5795;
  assign n6136 = n6124 & n6135;
  assign n6137 = ~n5502 & n6136;
  assign n6138 = ~n6134 & ~n6137;
  assign n6139 = ~n6132 & n6138;
  assign n6140 = ~n5885 & n6024;
  assign n6141 = ~n5884 & ~n6140;
  assign n6142 = ~n5874 & ~n5879;
  assign n6143 = ~n6043 & ~n6052;
  assign n6144 = ~n6050 & n6143;
  assign n6145 = ~n6041 & n6144;
  assign n6146 = ~n6066 & ~n6145;
  assign n6147 = pi03 & ~n5091;
  assign n6148 = ~n5092 & n6147;
  assign n6149 = ~n5178 & n6148;
  assign n6150 = pi04 & ~n5093;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = pi63 & ~n6151;
  assign n6153 = ~pi63 & ~n6150;
  assign n6154 = ~n6149 & n6153;
  assign n6155 = ~n6152 & ~n6154;
  assign n6156 = pi05 & ~n4513;
  assign n6157 = ~n4514 & n6156;
  assign n6158 = ~n4577 & n6157;
  assign n6159 = pi06 & ~n4515;
  assign n6160 = ~n6158 & ~n6159;
  assign n6161 = pi61 & ~n6160;
  assign n6162 = ~pi61 & ~n6159;
  assign n6163 = ~n6158 & n6162;
  assign n6164 = ~n6161 & ~n6163;
  assign n6165 = ~n6155 & n6164;
  assign n6166 = n6155 & ~n6164;
  assign n6167 = ~n6165 & ~n6166;
  assign n6168 = pi07 & ~n3959;
  assign n6169 = ~n3960 & n6168;
  assign n6170 = ~n4233 & n6169;
  assign n6171 = pi08 & ~n3961;
  assign n6172 = ~n6170 & ~n6171;
  assign n6173 = pi59 & ~n6172;
  assign n6174 = ~pi59 & ~n6171;
  assign n6175 = ~n6170 & n6174;
  assign n6176 = ~n6173 & ~n6175;
  assign n6177 = ~n6167 & n6176;
  assign n6178 = ~n6165 & ~n6176;
  assign n6179 = ~n6166 & n6178;
  assign n6180 = ~n6177 & ~n6179;
  assign n6181 = ~n6146 & n6180;
  assign n6182 = n6146 & ~n6180;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = n6070 & ~n6183;
  assign n6185 = ~n6070 & ~n6181;
  assign n6186 = ~n6182 & n6185;
  assign n6187 = ~n6184 & ~n6186;
  assign n6188 = ~n5873 & n6187;
  assign n6189 = ~n6142 & n6188;
  assign n6190 = ~n5873 & ~n6142;
  assign n6191 = ~n6187 & ~n6190;
  assign n6192 = ~n6189 & ~n6191;
  assign n6193 = ~n6141 & n6192;
  assign n6194 = pi17 & ~n1607;
  assign n6195 = ~n1608 & n6194;
  assign n6196 = ~n1782 & n6195;
  assign n6197 = pi18 & ~n1609;
  assign n6198 = ~n6196 & ~n6197;
  assign n6199 = pi49 & ~n6198;
  assign n6200 = pi19 & ~n1212;
  assign n6201 = ~n1213 & n6200;
  assign n6202 = ~n1425 & n6201;
  assign n6203 = pi20 & ~n1214;
  assign n6204 = ~n6202 & ~n6203;
  assign n6205 = pi47 & ~n6204;
  assign n6206 = ~pi47 & ~n6203;
  assign n6207 = ~n6202 & n6206;
  assign n6208 = ~pi49 & ~n6197;
  assign n6209 = ~n6196 & n6208;
  assign n6210 = ~n6207 & ~n6209;
  assign n6211 = ~n6205 & n6210;
  assign n6212 = ~n6199 & n6211;
  assign n6213 = ~n6205 & ~n6207;
  assign n6214 = ~n6199 & ~n6209;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = ~n6212 & ~n6215;
  assign n6217 = pi21 & ~n1006;
  assign n6218 = ~n1007 & n6217;
  assign n6219 = ~n1068 & n6218;
  assign n6220 = pi22 & ~n1008;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = pi45 & ~n6221;
  assign n6223 = ~pi45 & ~n6220;
  assign n6224 = ~n6219 & n6223;
  assign n6225 = ~n6222 & ~n6224;
  assign n6226 = ~n6216 & n6225;
  assign n6227 = ~n6212 & ~n6225;
  assign n6228 = ~n6215 & n6227;
  assign n6229 = ~n6226 & ~n6228;
  assign n6230 = ~n5910 & n5920;
  assign n6231 = ~n5975 & n5985;
  assign n6232 = ~n5907 & ~n5972;
  assign n6233 = ~n6231 & n6232;
  assign n6234 = ~n6230 & n6233;
  assign n6235 = ~n6229 & n6234;
  assign n6236 = ~n5972 & ~n6231;
  assign n6237 = ~n6226 & n6236;
  assign n6238 = ~n5907 & ~n6230;
  assign n6239 = ~n6228 & ~n6238;
  assign n6240 = n6237 & n6239;
  assign n6241 = ~n6236 & ~n6238;
  assign n6242 = ~n6229 & n6241;
  assign n6243 = ~n6240 & ~n6242;
  assign n6244 = ~n6235 & n6243;
  assign n6245 = ~n5990 & ~n6014;
  assign n6246 = ~n6226 & n6238;
  assign n6247 = ~n6228 & ~n6236;
  assign n6248 = n6246 & n6247;
  assign n6249 = ~n5991 & ~n6248;
  assign n6250 = ~n6245 & n6249;
  assign n6251 = n6244 & n6250;
  assign n6252 = ~n5991 & ~n6245;
  assign n6253 = ~n6240 & ~n6248;
  assign n6254 = ~n6235 & ~n6242;
  assign n6255 = n6253 & n6254;
  assign n6256 = ~n6252 & ~n6255;
  assign n6257 = pi23 & ~n683;
  assign n6258 = ~n684 & n6257;
  assign n6259 = ~n1231 & n6258;
  assign n6260 = pi24 & ~n685;
  assign n6261 = ~n6259 & ~n6260;
  assign n6262 = pi43 & ~n6261;
  assign n6263 = pi25 & ~n489;
  assign n6264 = ~n490 & n6263;
  assign n6265 = ~n572 & n6264;
  assign n6266 = pi26 & ~n491;
  assign n6267 = ~n6265 & ~n6266;
  assign n6268 = pi41 & ~n6267;
  assign n6269 = ~pi41 & ~n6266;
  assign n6270 = ~n6265 & n6269;
  assign n6271 = ~pi43 & ~n6260;
  assign n6272 = ~n6259 & n6271;
  assign n6273 = ~n6270 & ~n6272;
  assign n6274 = ~n6268 & n6273;
  assign n6275 = ~n6262 & n6274;
  assign n6276 = ~n6268 & ~n6270;
  assign n6277 = ~n6262 & ~n6272;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = ~n6275 & ~n6278;
  assign n6280 = pi27 & ~n304;
  assign n6281 = ~n305 & n6280;
  assign n6282 = ~n394 & n6281;
  assign n6283 = pi28 & ~n306;
  assign n6284 = ~n6282 & ~n6283;
  assign n6285 = pi39 & ~n6284;
  assign n6286 = ~pi39 & ~n6283;
  assign n6287 = ~n6282 & n6286;
  assign n6288 = ~n6285 & ~n6287;
  assign n6289 = ~n6279 & n6288;
  assign n6290 = ~n6275 & ~n6288;
  assign n6291 = ~n6278 & n6290;
  assign n6292 = ~n6289 & ~n6291;
  assign n6293 = ~n6013 & ~n6292;
  assign n6294 = n6013 & ~n6289;
  assign n6295 = ~n6291 & n6294;
  assign n6296 = n143 & n156;
  assign n6297 = pi31 & pi35;
  assign n6298 = ~n6296 & n6297;
  assign n6299 = pi31 & ~n6296;
  assign n6300 = ~pi35 & ~n6299;
  assign n6301 = ~n6298 & ~n6300;
  assign n6302 = pi29 & ~n193;
  assign n6303 = ~n194 & n6302;
  assign n6304 = ~n729 & n6303;
  assign n6305 = pi30 & ~n195;
  assign n6306 = ~n6304 & ~n6305;
  assign n6307 = pi37 & ~n6306;
  assign n6308 = ~pi37 & ~n6305;
  assign n6309 = ~n6304 & n6308;
  assign n6310 = ~n6307 & ~n6309;
  assign n6311 = ~n6301 & n6310;
  assign n6312 = n6301 & ~n6310;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = ~n6295 & ~n6313;
  assign n6315 = ~n6293 & n6314;
  assign n6316 = ~n6293 & ~n6295;
  assign n6317 = n6313 & ~n6316;
  assign n6318 = ~n6315 & ~n6317;
  assign n6319 = ~n6256 & n6318;
  assign n6320 = ~n6251 & n6319;
  assign n6321 = ~n6251 & ~n6256;
  assign n6322 = ~n6318 & ~n6321;
  assign n6323 = ~n6320 & ~n6322;
  assign n6324 = ~n5944 & ~n6021;
  assign n6325 = ~n5829 & ~n5869;
  assign n6326 = pi09 & ~n3205;
  assign n6327 = ~n3206 & n6326;
  assign n6328 = ~n3463 & n6327;
  assign n6329 = pi10 & ~n3207;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = pi57 & ~n6330;
  assign n6332 = ~pi57 & ~n6329;
  assign n6333 = ~n6328 & n6332;
  assign n6334 = ~n6331 & ~n6333;
  assign n6335 = ~n5851 & n5861;
  assign n6336 = ~n5848 & ~n6335;
  assign n6337 = n6334 & ~n6336;
  assign n6338 = pi11 & ~n2876;
  assign n6339 = ~n2877 & n6338;
  assign n6340 = ~n2960 & n6339;
  assign n6341 = pi12 & ~n2878;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = pi55 & ~n6342;
  assign n6344 = pi13 & ~n2288;
  assign n6345 = ~n2289 & n6344;
  assign n6346 = ~n2647 & n6345;
  assign n6347 = pi14 & ~n2290;
  assign n6348 = ~n6346 & ~n6347;
  assign n6349 = pi53 & ~n6348;
  assign n6350 = ~pi53 & ~n6347;
  assign n6351 = ~n6346 & n6350;
  assign n6352 = ~pi55 & ~n6341;
  assign n6353 = ~n6340 & n6352;
  assign n6354 = ~n6351 & ~n6353;
  assign n6355 = ~n6349 & n6354;
  assign n6356 = ~n6343 & n6355;
  assign n6357 = ~n6349 & ~n6351;
  assign n6358 = ~n6343 & ~n6353;
  assign n6359 = ~n6357 & ~n6358;
  assign n6360 = ~n6356 & ~n6359;
  assign n6361 = pi15 & ~n2023;
  assign n6362 = ~n2024 & n6361;
  assign n6363 = ~n2079 & n6362;
  assign n6364 = pi16 & ~n2025;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = pi51 & ~n6365;
  assign n6367 = ~pi51 & ~n6364;
  assign n6368 = ~n6363 & n6367;
  assign n6369 = ~n6366 & ~n6368;
  assign n6370 = ~n6360 & n6369;
  assign n6371 = ~n6356 & ~n6369;
  assign n6372 = ~n6359 & n6371;
  assign n6373 = ~n6370 & ~n6372;
  assign n6374 = ~n5848 & ~n6334;
  assign n6375 = ~n6335 & n6374;
  assign n6376 = ~n6373 & ~n6375;
  assign n6377 = ~n6337 & n6376;
  assign n6378 = ~n6337 & ~n6375;
  assign n6379 = n6373 & ~n6378;
  assign n6380 = ~n6377 & ~n6379;
  assign n6381 = ~n6325 & n6380;
  assign n6382 = n6325 & ~n6380;
  assign n6383 = ~n6381 & ~n6382;
  assign n6384 = ~n5923 & ~n5935;
  assign n6385 = n5924 & ~n5926;
  assign n6386 = ~n5928 & ~n6385;
  assign n6387 = ~n6384 & ~n6386;
  assign n6388 = ~n6383 & n6387;
  assign n6389 = ~n6381 & ~n6387;
  assign n6390 = ~n6382 & n6389;
  assign n6391 = ~n6388 & ~n6390;
  assign n6392 = ~n6324 & n6391;
  assign n6393 = n6324 & ~n6391;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = ~n6323 & ~n6394;
  assign n6396 = ~n5884 & ~n6192;
  assign n6397 = ~n6140 & n6396;
  assign n6398 = n6323 & ~n6392;
  assign n6399 = ~n6393 & n6398;
  assign n6400 = ~n6397 & ~n6399;
  assign n6401 = ~n6395 & n6400;
  assign n6402 = ~n6193 & n6401;
  assign n6403 = ~n6193 & ~n6397;
  assign n6404 = ~n6395 & ~n6399;
  assign n6405 = ~n6403 & ~n6404;
  assign n6406 = ~n6402 & ~n6405;
  assign n6407 = n6028 & ~n6084;
  assign n6408 = ~n6082 & ~n6407;
  assign n6409 = ~n6075 & ~n6077;
  assign n6410 = ~n6408 & n6409;
  assign n6411 = ~n6082 & ~n6409;
  assign n6412 = ~n6407 & n6411;
  assign n6413 = ~n6410 & ~n6412;
  assign n6414 = ~n6406 & n6413;
  assign n6415 = n6406 & ~n6413;
  assign n6416 = ~n6414 & ~n6415;
  assign n6417 = ~n6090 & ~n6093;
  assign n6418 = ~n6096 & ~n6417;
  assign n6419 = ~n6416 & n6418;
  assign n6420 = n6416 & ~n6418;
  assign n6421 = ~n6419 & ~n6420;
  assign n6422 = ~n6139 & n6421;
  assign n6423 = ~n6134 & ~n6421;
  assign n6424 = ~n6137 & n6423;
  assign n6425 = ~n6132 & n6424;
  assign po34 = ~n6422 & ~n6425;
  assign n6427 = n6102 & n6421;
  assign n6428 = n5481 & n5797;
  assign n6429 = n4551 & n5166;
  assign n6430 = n6428 & n6429;
  assign n6431 = n6427 & n6430;
  assign n6432 = ~n4273 & n6431;
  assign n6433 = ~n6138 & ~n6419;
  assign n6434 = ~n6420 & ~n6433;
  assign n6435 = ~n6432 & n6434;
  assign n6436 = ~n6412 & ~n6414;
  assign n6437 = ~n6382 & ~n6387;
  assign n6438 = ~n6154 & ~n6163;
  assign n6439 = ~n6161 & n6438;
  assign n6440 = ~n6152 & n6439;
  assign n6441 = ~n6177 & ~n6440;
  assign n6442 = pi04 & ~n5091;
  assign n6443 = ~n5092 & n6442;
  assign n6444 = ~n5178 & n6443;
  assign n6445 = pi05 & ~n5093;
  assign n6446 = ~n6444 & ~n6445;
  assign n6447 = pi63 & ~n6446;
  assign n6448 = ~pi63 & ~n6445;
  assign n6449 = ~n6444 & n6448;
  assign n6450 = ~n6447 & ~n6449;
  assign n6451 = pi06 & ~n4513;
  assign n6452 = ~n4514 & n6451;
  assign n6453 = ~n4577 & n6452;
  assign n6454 = pi07 & ~n4515;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = pi61 & ~n6455;
  assign n6457 = ~pi61 & ~n6454;
  assign n6458 = ~n6453 & n6457;
  assign n6459 = ~n6456 & ~n6458;
  assign n6460 = ~n6450 & n6459;
  assign n6461 = n6450 & ~n6459;
  assign n6462 = ~n6460 & ~n6461;
  assign n6463 = pi08 & ~n3959;
  assign n6464 = ~n3960 & n6463;
  assign n6465 = ~n4233 & n6464;
  assign n6466 = pi09 & ~n3961;
  assign n6467 = ~n6465 & ~n6466;
  assign n6468 = pi59 & ~n6467;
  assign n6469 = ~pi59 & ~n6466;
  assign n6470 = ~n6465 & n6469;
  assign n6471 = ~n6468 & ~n6470;
  assign n6472 = ~n6462 & n6471;
  assign n6473 = ~n6460 & ~n6471;
  assign n6474 = ~n6461 & n6473;
  assign n6475 = ~n6472 & ~n6474;
  assign n6476 = ~n6441 & n6475;
  assign n6477 = n6441 & ~n6475;
  assign n6478 = ~n6476 & ~n6477;
  assign n6479 = n6181 & ~n6478;
  assign n6480 = ~n6181 & ~n6476;
  assign n6481 = ~n6477 & n6480;
  assign n6482 = ~n6479 & ~n6481;
  assign n6483 = ~n6381 & n6482;
  assign n6484 = ~n6437 & n6483;
  assign n6485 = ~n6381 & ~n6437;
  assign n6486 = ~n6482 & ~n6485;
  assign n6487 = ~n6484 & ~n6486;
  assign n6488 = ~n6323 & ~n6393;
  assign n6489 = ~n6392 & ~n6488;
  assign n6490 = n6487 & ~n6489;
  assign n6491 = ~n6392 & ~n6487;
  assign n6492 = ~n6488 & n6491;
  assign n6493 = ~n6337 & ~n6377;
  assign n6494 = pi10 & ~n3205;
  assign n6495 = ~n3206 & n6494;
  assign n6496 = ~n3463 & n6495;
  assign n6497 = pi11 & ~n3207;
  assign n6498 = ~n6496 & ~n6497;
  assign n6499 = pi57 & ~n6498;
  assign n6500 = ~pi57 & ~n6497;
  assign n6501 = ~n6496 & n6500;
  assign n6502 = ~n6499 & ~n6501;
  assign n6503 = ~n6359 & n6369;
  assign n6504 = ~n6356 & ~n6503;
  assign n6505 = n6502 & ~n6504;
  assign n6506 = pi12 & ~n2876;
  assign n6507 = ~n2877 & n6506;
  assign n6508 = ~n2960 & n6507;
  assign n6509 = pi13 & ~n2878;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = pi55 & ~n6510;
  assign n6512 = pi14 & ~n2288;
  assign n6513 = ~n2289 & n6512;
  assign n6514 = ~n2647 & n6513;
  assign n6515 = pi15 & ~n2290;
  assign n6516 = ~n6514 & ~n6515;
  assign n6517 = pi53 & ~n6516;
  assign n6518 = ~pi53 & ~n6515;
  assign n6519 = ~n6514 & n6518;
  assign n6520 = ~pi55 & ~n6509;
  assign n6521 = ~n6508 & n6520;
  assign n6522 = ~n6519 & ~n6521;
  assign n6523 = ~n6517 & n6522;
  assign n6524 = ~n6511 & n6523;
  assign n6525 = ~n6517 & ~n6519;
  assign n6526 = ~n6511 & ~n6521;
  assign n6527 = ~n6525 & ~n6526;
  assign n6528 = ~n6524 & ~n6527;
  assign n6529 = pi16 & ~n2023;
  assign n6530 = ~n2024 & n6529;
  assign n6531 = ~n2079 & n6530;
  assign n6532 = pi17 & ~n2025;
  assign n6533 = ~n6531 & ~n6532;
  assign n6534 = pi51 & ~n6533;
  assign n6535 = ~pi51 & ~n6532;
  assign n6536 = ~n6531 & n6535;
  assign n6537 = ~n6534 & ~n6536;
  assign n6538 = ~n6528 & n6537;
  assign n6539 = ~n6524 & ~n6537;
  assign n6540 = ~n6527 & n6539;
  assign n6541 = ~n6538 & ~n6540;
  assign n6542 = ~n6356 & ~n6502;
  assign n6543 = ~n6503 & n6542;
  assign n6544 = ~n6541 & ~n6543;
  assign n6545 = ~n6505 & n6544;
  assign n6546 = ~n6505 & ~n6543;
  assign n6547 = n6541 & ~n6546;
  assign n6548 = ~n6545 & ~n6547;
  assign n6549 = ~n6493 & n6548;
  assign n6550 = n6493 & ~n6548;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = ~n6229 & ~n6238;
  assign n6553 = ~n6228 & n6246;
  assign n6554 = ~n6236 & ~n6553;
  assign n6555 = ~n6552 & ~n6554;
  assign n6556 = ~n6551 & n6555;
  assign n6557 = ~n6549 & ~n6555;
  assign n6558 = ~n6550 & n6557;
  assign n6559 = ~n6556 & ~n6558;
  assign n6560 = pi18 & ~n1607;
  assign n6561 = ~n1608 & n6560;
  assign n6562 = ~n1782 & n6561;
  assign n6563 = pi19 & ~n1609;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = pi49 & ~n6564;
  assign n6566 = pi20 & ~n1212;
  assign n6567 = ~n1213 & n6566;
  assign n6568 = ~n1425 & n6567;
  assign n6569 = pi21 & ~n1214;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = pi47 & ~n6570;
  assign n6572 = ~pi47 & ~n6569;
  assign n6573 = ~n6568 & n6572;
  assign n6574 = ~pi49 & ~n6563;
  assign n6575 = ~n6562 & n6574;
  assign n6576 = ~n6573 & ~n6575;
  assign n6577 = ~n6571 & n6576;
  assign n6578 = ~n6565 & n6577;
  assign n6579 = ~n6571 & ~n6573;
  assign n6580 = ~n6565 & ~n6575;
  assign n6581 = ~n6579 & ~n6580;
  assign n6582 = ~n6578 & ~n6581;
  assign n6583 = pi22 & ~n1006;
  assign n6584 = ~n1007 & n6583;
  assign n6585 = ~n1068 & n6584;
  assign n6586 = pi23 & ~n1008;
  assign n6587 = ~n6585 & ~n6586;
  assign n6588 = pi45 & ~n6587;
  assign n6589 = ~pi45 & ~n6586;
  assign n6590 = ~n6585 & n6589;
  assign n6591 = ~n6588 & ~n6590;
  assign n6592 = ~n6582 & n6591;
  assign n6593 = ~n6215 & n6225;
  assign n6594 = ~n6212 & ~n6593;
  assign n6595 = ~n6592 & n6594;
  assign n6596 = ~n6578 & ~n6591;
  assign n6597 = ~n6581 & n6596;
  assign n6598 = ~n6278 & n6288;
  assign n6599 = ~n6275 & ~n6598;
  assign n6600 = ~n6597 & ~n6599;
  assign n6601 = n6595 & n6600;
  assign n6602 = ~n6592 & n6599;
  assign n6603 = ~n6594 & ~n6597;
  assign n6604 = n6602 & n6603;
  assign n6605 = ~n6601 & ~n6604;
  assign n6606 = ~n6592 & ~n6597;
  assign n6607 = ~n6594 & ~n6599;
  assign n6608 = ~n6606 & n6607;
  assign n6609 = ~n6212 & ~n6275;
  assign n6610 = ~n6598 & n6609;
  assign n6611 = ~n6593 & n6610;
  assign n6612 = ~n6606 & n6611;
  assign n6613 = ~n6608 & ~n6612;
  assign n6614 = n6605 & n6613;
  assign n6615 = ~n6278 & ~n6311;
  assign n6616 = ~n6312 & n6615;
  assign n6617 = n6290 & n6616;
  assign n6618 = n6288 & ~n6311;
  assign n6619 = ~n6312 & n6618;
  assign n6620 = ~n6279 & n6619;
  assign n6621 = ~n6617 & ~n6620;
  assign n6622 = ~n6013 & ~n6278;
  assign n6623 = n6290 & n6622;
  assign n6624 = ~n6013 & ~n6311;
  assign n6625 = ~n6312 & n6624;
  assign n6626 = ~n6013 & n6288;
  assign n6627 = ~n6279 & n6626;
  assign n6628 = ~n6625 & ~n6627;
  assign n6629 = ~n6623 & n6628;
  assign n6630 = n6621 & n6629;
  assign n6631 = pi24 & ~n683;
  assign n6632 = ~n684 & n6631;
  assign n6633 = ~n1231 & n6632;
  assign n6634 = pi25 & ~n685;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = pi43 & ~n6635;
  assign n6637 = pi26 & ~n489;
  assign n6638 = ~n490 & n6637;
  assign n6639 = ~n572 & n6638;
  assign n6640 = pi27 & ~n491;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = pi41 & ~n6641;
  assign n6643 = ~pi41 & ~n6640;
  assign n6644 = ~n6639 & n6643;
  assign n6645 = ~pi43 & ~n6634;
  assign n6646 = ~n6633 & n6645;
  assign n6647 = ~n6644 & ~n6646;
  assign n6648 = ~n6642 & n6647;
  assign n6649 = ~n6636 & n6648;
  assign n6650 = ~n6642 & ~n6644;
  assign n6651 = ~n6636 & ~n6646;
  assign n6652 = ~n6650 & ~n6651;
  assign n6653 = ~n6649 & ~n6652;
  assign n6654 = pi30 & ~n193;
  assign n6655 = ~n194 & n6654;
  assign n6656 = ~n729 & n6655;
  assign n6657 = pi31 & ~n195;
  assign n6658 = ~n6656 & ~n6657;
  assign n6659 = pi37 & ~n6658;
  assign n6660 = ~pi37 & ~n6657;
  assign n6661 = ~n6656 & n6660;
  assign n6662 = ~n6659 & ~n6661;
  assign n6663 = pi28 & ~n304;
  assign n6664 = ~n305 & n6663;
  assign n6665 = ~n394 & n6664;
  assign n6666 = pi29 & ~n306;
  assign n6667 = ~n6665 & ~n6666;
  assign n6668 = pi39 & ~n6667;
  assign n6669 = ~pi39 & ~n6666;
  assign n6670 = ~n6665 & n6669;
  assign n6671 = ~n6668 & ~n6670;
  assign n6672 = ~n6662 & ~n6671;
  assign n6673 = n6311 & n6672;
  assign n6674 = ~n6653 & n6673;
  assign n6675 = n6662 & ~n6671;
  assign n6676 = ~n6311 & n6675;
  assign n6677 = ~n6653 & n6676;
  assign n6678 = ~n6674 & ~n6677;
  assign n6679 = ~n6662 & n6671;
  assign n6680 = ~n6311 & n6679;
  assign n6681 = ~n6653 & n6680;
  assign n6682 = ~n6309 & ~n6661;
  assign n6683 = ~n6307 & n6682;
  assign n6684 = ~n6301 & ~n6659;
  assign n6685 = n6683 & n6684;
  assign n6686 = n6671 & n6685;
  assign n6687 = ~n6653 & n6686;
  assign n6688 = ~n6681 & ~n6687;
  assign n6689 = n6678 & n6688;
  assign n6690 = ~n6311 & n6672;
  assign n6691 = n6653 & n6690;
  assign n6692 = ~n6671 & n6685;
  assign n6693 = n6653 & n6692;
  assign n6694 = ~n6691 & ~n6693;
  assign n6695 = ~n6309 & ~n6670;
  assign n6696 = ~n6307 & n6695;
  assign n6697 = ~n6301 & ~n6668;
  assign n6698 = n6696 & n6697;
  assign n6699 = ~n6662 & n6698;
  assign n6700 = n6653 & n6699;
  assign n6701 = ~n6661 & ~n6670;
  assign n6702 = ~n6659 & n6701;
  assign n6703 = ~n6668 & n6702;
  assign n6704 = ~n6311 & n6703;
  assign n6705 = n6653 & n6704;
  assign n6706 = ~n6700 & ~n6705;
  assign n6707 = n6694 & n6706;
  assign n6708 = n6689 & n6707;
  assign n6709 = n6630 & ~n6708;
  assign n6710 = ~n6614 & n6709;
  assign n6711 = ~n6630 & ~n6708;
  assign n6712 = n6614 & n6711;
  assign n6713 = ~n6630 & n6708;
  assign n6714 = ~n6614 & n6713;
  assign n6715 = ~n6712 & ~n6714;
  assign n6716 = ~n6710 & n6715;
  assign n6717 = ~n6251 & ~n6318;
  assign n6718 = ~n6623 & ~n6691;
  assign n6719 = n6628 & n6718;
  assign n6720 = n6621 & n6719;
  assign n6721 = ~n6677 & ~n6681;
  assign n6722 = ~n6687 & n6721;
  assign n6723 = ~n6693 & ~n6700;
  assign n6724 = ~n6674 & ~n6705;
  assign n6725 = n6723 & n6724;
  assign n6726 = n6722 & n6725;
  assign n6727 = n6720 & n6726;
  assign n6728 = n6614 & n6727;
  assign n6729 = ~n6256 & ~n6728;
  assign n6730 = ~n6717 & n6729;
  assign n6731 = n6716 & n6730;
  assign n6732 = ~n6559 & n6731;
  assign n6733 = ~n6712 & ~n6728;
  assign n6734 = ~n6710 & ~n6714;
  assign n6735 = n6733 & n6734;
  assign n6736 = ~n6556 & n6735;
  assign n6737 = ~n6256 & ~n6717;
  assign n6738 = ~n6558 & ~n6737;
  assign n6739 = n6736 & n6738;
  assign n6740 = ~n6732 & ~n6739;
  assign n6741 = ~n6735 & ~n6737;
  assign n6742 = ~n6559 & n6741;
  assign n6743 = ~n6556 & n6737;
  assign n6744 = ~n6558 & ~n6735;
  assign n6745 = n6743 & n6744;
  assign n6746 = ~n6742 & ~n6745;
  assign n6747 = n6740 & n6746;
  assign n6748 = ~n6492 & n6747;
  assign n6749 = ~n6490 & n6748;
  assign n6750 = ~n6490 & ~n6492;
  assign n6751 = ~n6747 & ~n6750;
  assign n6752 = ~n6749 & ~n6751;
  assign n6753 = ~n6397 & ~n6404;
  assign n6754 = ~n6193 & ~n6753;
  assign n6755 = n6070 & ~n6181;
  assign n6756 = ~n6182 & n6755;
  assign n6757 = ~n6191 & ~n6756;
  assign n6758 = ~n6754 & ~n6757;
  assign n6759 = ~n6193 & n6757;
  assign n6760 = ~n6753 & n6759;
  assign n6761 = ~n6758 & ~n6760;
  assign n6762 = ~n6752 & n6761;
  assign n6763 = n6752 & ~n6761;
  assign n6764 = ~n6762 & ~n6763;
  assign n6765 = n6436 & n6764;
  assign n6766 = ~n6436 & ~n6764;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n6435 & n6767;
  assign n6769 = ~n6420 & ~n6767;
  assign n6770 = ~n6433 & n6769;
  assign n6771 = ~n6432 & n6770;
  assign po35 = ~n6768 & ~n6771;
  assign n6773 = n5166 & n6428;
  assign n6774 = n6427 & n6773;
  assign n6775 = ~n4864 & n6774;
  assign n6776 = ~n4863 & n6775;
  assign n6777 = n5480 & ~n5795;
  assign n6778 = n6124 & n6777;
  assign n6779 = ~n6134 & ~n6420;
  assign n6780 = ~n6778 & n6779;
  assign n6781 = ~n6419 & ~n6780;
  assign n6782 = n5173 & n6428;
  assign n6783 = n6427 & n6782;
  assign n6784 = ~n6781 & ~n6783;
  assign n6785 = ~n6776 & n6784;
  assign n6786 = ~n6765 & ~n6785;
  assign n6787 = ~n6766 & ~n6786;
  assign n6788 = n6752 & ~n6760;
  assign n6789 = ~n6758 & ~n6788;
  assign n6790 = n6181 & ~n6476;
  assign n6791 = ~n6477 & n6790;
  assign n6792 = ~n6486 & ~n6791;
  assign n6793 = ~n6732 & n6792;
  assign n6794 = ~n6739 & ~n6742;
  assign n6795 = ~n6745 & n6794;
  assign n6796 = n6793 & n6795;
  assign n6797 = ~n6489 & n6796;
  assign n6798 = ~n6559 & n6737;
  assign n6799 = n6559 & ~n6737;
  assign n6800 = n6735 & ~n6799;
  assign n6801 = ~n6798 & ~n6800;
  assign n6802 = ~n6550 & ~n6555;
  assign n6803 = ~n6449 & ~n6458;
  assign n6804 = ~n6456 & n6803;
  assign n6805 = ~n6447 & n6804;
  assign n6806 = ~n6472 & ~n6805;
  assign n6807 = pi05 & ~n5091;
  assign n6808 = ~n5092 & n6807;
  assign n6809 = ~n5178 & n6808;
  assign n6810 = pi06 & ~n5093;
  assign n6811 = ~n6809 & ~n6810;
  assign n6812 = pi63 & ~n6811;
  assign n6813 = ~pi63 & ~n6810;
  assign n6814 = ~n6809 & n6813;
  assign n6815 = ~n6812 & ~n6814;
  assign n6816 = pi07 & ~n4513;
  assign n6817 = ~n4514 & n6816;
  assign n6818 = ~n4577 & n6817;
  assign n6819 = pi08 & ~n4515;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = pi61 & ~n6820;
  assign n6822 = ~pi61 & ~n6819;
  assign n6823 = ~n6818 & n6822;
  assign n6824 = ~n6821 & ~n6823;
  assign n6825 = ~n6815 & n6824;
  assign n6826 = n6815 & ~n6824;
  assign n6827 = ~n6825 & ~n6826;
  assign n6828 = pi09 & ~n3959;
  assign n6829 = ~n3960 & n6828;
  assign n6830 = ~n4233 & n6829;
  assign n6831 = pi10 & ~n3961;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833 = pi59 & ~n6832;
  assign n6834 = ~pi59 & ~n6831;
  assign n6835 = ~n6830 & n6834;
  assign n6836 = ~n6833 & ~n6835;
  assign n6837 = ~n6827 & n6836;
  assign n6838 = ~n6825 & ~n6836;
  assign n6839 = ~n6826 & n6838;
  assign n6840 = ~n6837 & ~n6839;
  assign n6841 = ~n6806 & n6840;
  assign n6842 = n6806 & ~n6840;
  assign n6843 = ~n6841 & ~n6842;
  assign n6844 = n6476 & ~n6843;
  assign n6845 = ~n6476 & ~n6841;
  assign n6846 = ~n6842 & n6845;
  assign n6847 = ~n6844 & ~n6846;
  assign n6848 = ~n6549 & n6847;
  assign n6849 = ~n6802 & n6848;
  assign n6850 = ~n6549 & ~n6802;
  assign n6851 = ~n6847 & ~n6850;
  assign n6852 = ~n6849 & ~n6851;
  assign n6853 = ~n6801 & n6852;
  assign n6854 = ~n6798 & ~n6852;
  assign n6855 = ~n6800 & n6854;
  assign n6856 = ~n6505 & ~n6545;
  assign n6857 = pi11 & ~n3205;
  assign n6858 = ~n3206 & n6857;
  assign n6859 = ~n3463 & n6858;
  assign n6860 = pi12 & ~n3207;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = pi57 & ~n6861;
  assign n6863 = ~pi57 & ~n6860;
  assign n6864 = ~n6859 & n6863;
  assign n6865 = ~n6862 & ~n6864;
  assign n6866 = ~n6527 & n6537;
  assign n6867 = ~n6524 & ~n6866;
  assign n6868 = n6865 & ~n6867;
  assign n6869 = pi13 & ~n2876;
  assign n6870 = ~n2877 & n6869;
  assign n6871 = ~n2960 & n6870;
  assign n6872 = pi14 & ~n2878;
  assign n6873 = ~n6871 & ~n6872;
  assign n6874 = pi55 & ~n6873;
  assign n6875 = pi15 & ~n2288;
  assign n6876 = ~n2289 & n6875;
  assign n6877 = ~n2647 & n6876;
  assign n6878 = pi16 & ~n2290;
  assign n6879 = ~n6877 & ~n6878;
  assign n6880 = pi53 & ~n6879;
  assign n6881 = ~pi53 & ~n6878;
  assign n6882 = ~n6877 & n6881;
  assign n6883 = ~pi55 & ~n6872;
  assign n6884 = ~n6871 & n6883;
  assign n6885 = ~n6882 & ~n6884;
  assign n6886 = ~n6880 & n6885;
  assign n6887 = ~n6874 & n6886;
  assign n6888 = ~n6880 & ~n6882;
  assign n6889 = ~n6874 & ~n6884;
  assign n6890 = ~n6888 & ~n6889;
  assign n6891 = ~n6887 & ~n6890;
  assign n6892 = pi17 & ~n2023;
  assign n6893 = ~n2024 & n6892;
  assign n6894 = ~n2079 & n6893;
  assign n6895 = pi18 & ~n2025;
  assign n6896 = ~n6894 & ~n6895;
  assign n6897 = pi51 & ~n6896;
  assign n6898 = ~pi51 & ~n6895;
  assign n6899 = ~n6894 & n6898;
  assign n6900 = ~n6897 & ~n6899;
  assign n6901 = ~n6891 & n6900;
  assign n6902 = ~n6887 & ~n6900;
  assign n6903 = ~n6890 & n6902;
  assign n6904 = ~n6901 & ~n6903;
  assign n6905 = ~n6524 & ~n6865;
  assign n6906 = ~n6866 & n6905;
  assign n6907 = ~n6904 & ~n6906;
  assign n6908 = ~n6868 & n6907;
  assign n6909 = ~n6868 & ~n6906;
  assign n6910 = n6904 & ~n6909;
  assign n6911 = ~n6908 & ~n6910;
  assign n6912 = ~n6856 & n6911;
  assign n6913 = n6856 & ~n6911;
  assign n6914 = ~n6912 & ~n6913;
  assign n6915 = ~n6594 & ~n6606;
  assign n6916 = n6595 & ~n6597;
  assign n6917 = ~n6599 & ~n6916;
  assign n6918 = ~n6915 & ~n6917;
  assign n6919 = ~n6914 & n6918;
  assign n6920 = ~n6912 & ~n6918;
  assign n6921 = ~n6913 & n6920;
  assign n6922 = ~n6919 & ~n6921;
  assign n6923 = ~n6614 & ~n6630;
  assign n6924 = pi19 & ~n1607;
  assign n6925 = ~n1608 & n6924;
  assign n6926 = ~n1782 & n6925;
  assign n6927 = pi20 & ~n1609;
  assign n6928 = ~n6926 & ~n6927;
  assign n6929 = pi49 & ~n6928;
  assign n6930 = pi21 & ~n1212;
  assign n6931 = ~n1213 & n6930;
  assign n6932 = ~n1425 & n6931;
  assign n6933 = pi22 & ~n1214;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = pi47 & ~n6934;
  assign n6936 = ~pi47 & ~n6933;
  assign n6937 = ~n6932 & n6936;
  assign n6938 = ~pi49 & ~n6927;
  assign n6939 = ~n6926 & n6938;
  assign n6940 = ~n6937 & ~n6939;
  assign n6941 = ~n6935 & n6940;
  assign n6942 = ~n6929 & n6941;
  assign n6943 = ~n6935 & ~n6937;
  assign n6944 = ~n6929 & ~n6939;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = ~n6942 & ~n6945;
  assign n6947 = pi23 & ~n1006;
  assign n6948 = ~n1007 & n6947;
  assign n6949 = ~n1068 & n6948;
  assign n6950 = pi24 & ~n1008;
  assign n6951 = ~n6949 & ~n6950;
  assign n6952 = pi45 & ~n6951;
  assign n6953 = ~pi45 & ~n6950;
  assign n6954 = ~n6949 & n6953;
  assign n6955 = ~n6952 & ~n6954;
  assign n6956 = ~n6946 & n6955;
  assign n6957 = ~n6581 & n6591;
  assign n6958 = ~n6578 & ~n6957;
  assign n6959 = ~n6956 & n6958;
  assign n6960 = ~n6942 & ~n6955;
  assign n6961 = ~n6945 & n6960;
  assign n6962 = ~n6652 & n6671;
  assign n6963 = ~n6649 & ~n6962;
  assign n6964 = ~n6961 & ~n6963;
  assign n6965 = n6959 & n6964;
  assign n6966 = ~n6956 & n6963;
  assign n6967 = ~n6958 & ~n6961;
  assign n6968 = n6966 & n6967;
  assign n6969 = ~n6965 & ~n6968;
  assign n6970 = ~n6956 & ~n6961;
  assign n6971 = ~n6958 & ~n6963;
  assign n6972 = ~n6970 & n6971;
  assign n6973 = ~n6578 & ~n6649;
  assign n6974 = ~n6962 & n6973;
  assign n6975 = ~n6957 & n6974;
  assign n6976 = ~n6970 & n6975;
  assign n6977 = ~n6972 & ~n6976;
  assign n6978 = n6969 & n6977;
  assign n6979 = pi25 & ~n683;
  assign n6980 = ~n684 & n6979;
  assign n6981 = ~n1231 & n6980;
  assign n6982 = pi26 & ~n685;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = pi43 & ~n6983;
  assign n6985 = pi27 & ~n489;
  assign n6986 = ~n490 & n6985;
  assign n6987 = ~n572 & n6986;
  assign n6988 = pi28 & ~n491;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = pi41 & ~n6989;
  assign n6991 = ~pi41 & ~n6988;
  assign n6992 = ~n6987 & n6991;
  assign n6993 = ~pi43 & ~n6982;
  assign n6994 = ~n6981 & n6993;
  assign n6995 = ~n6992 & ~n6994;
  assign n6996 = ~n6990 & n6995;
  assign n6997 = ~n6984 & n6996;
  assign n6998 = ~n6990 & ~n6992;
  assign n6999 = ~n6984 & ~n6994;
  assign n7000 = ~n6998 & ~n6999;
  assign n7001 = ~n6997 & ~n7000;
  assign n7002 = pi29 & ~n304;
  assign n7003 = ~n305 & n7002;
  assign n7004 = ~n394 & n7003;
  assign n7005 = pi30 & ~n306;
  assign n7006 = ~n7004 & ~n7005;
  assign n7007 = pi39 & ~n7006;
  assign n7008 = ~pi39 & ~n7005;
  assign n7009 = ~n7004 & n7008;
  assign n7010 = ~n7007 & ~n7009;
  assign n7011 = n195 & n729;
  assign n7012 = pi31 & pi37;
  assign n7013 = ~n7011 & n7012;
  assign n7014 = pi31 & ~n7011;
  assign n7015 = ~pi37 & ~n7014;
  assign n7016 = ~n7013 & ~n7015;
  assign n7017 = n6662 & ~n7016;
  assign n7018 = ~n7010 & n7017;
  assign n7019 = ~n7001 & n7018;
  assign n7020 = n7010 & ~n7016;
  assign n7021 = ~n6662 & n7020;
  assign n7022 = ~n7001 & n7021;
  assign n7023 = ~n7019 & ~n7022;
  assign n7024 = ~n6662 & ~n7016;
  assign n7025 = ~n7010 & n7024;
  assign n7026 = n7001 & n7025;
  assign n7027 = ~n6661 & ~n7009;
  assign n7028 = ~n6659 & n7027;
  assign n7029 = ~n7007 & ~n7016;
  assign n7030 = n7028 & n7029;
  assign n7031 = ~n6997 & n7030;
  assign n7032 = ~n7000 & n7031;
  assign n7033 = ~n7026 & ~n7032;
  assign n7034 = n7023 & n7033;
  assign n7035 = ~n6662 & n7016;
  assign n7036 = ~n7010 & n7035;
  assign n7037 = ~n7001 & n7036;
  assign n7038 = n7016 & n7027;
  assign n7039 = ~n6659 & ~n7007;
  assign n7040 = n7038 & n7039;
  assign n7041 = ~n7001 & n7040;
  assign n7042 = ~n7037 & ~n7041;
  assign n7043 = n6662 & n7016;
  assign n7044 = ~n7010 & n7043;
  assign n7045 = n7001 & n7044;
  assign n7046 = n7010 & n7035;
  assign n7047 = n7001 & n7046;
  assign n7048 = ~n7045 & ~n7047;
  assign n7049 = n7042 & n7048;
  assign n7050 = n7034 & n7049;
  assign n7051 = ~n6649 & n6672;
  assign n7052 = ~n6652 & n7051;
  assign n7053 = n6311 & ~n6671;
  assign n7054 = n6653 & n7053;
  assign n7055 = ~n6653 & n6698;
  assign n7056 = ~n7054 & ~n7055;
  assign n7057 = ~n7052 & n7056;
  assign n7058 = n6311 & ~n6662;
  assign n7059 = ~n6653 & n6679;
  assign n7060 = ~n7058 & ~n7059;
  assign n7061 = n7057 & n7060;
  assign n7062 = ~n7050 & ~n7061;
  assign n7063 = n6978 & n7062;
  assign n7064 = n7050 & ~n7061;
  assign n7065 = ~n6978 & n7064;
  assign n7066 = ~n7063 & ~n7065;
  assign n7067 = ~n6923 & n7066;
  assign n7068 = n6614 & n6630;
  assign n7069 = n6708 & ~n7068;
  assign n7070 = ~n7037 & ~n7058;
  assign n7071 = ~n7041 & ~n7045;
  assign n7072 = ~n7019 & ~n7047;
  assign n7073 = n7071 & n7072;
  assign n7074 = n7070 & n7073;
  assign n7075 = ~n7022 & ~n7026;
  assign n7076 = ~n7032 & ~n7059;
  assign n7077 = n7075 & n7076;
  assign n7078 = n7057 & n7077;
  assign n7079 = n7074 & n7078;
  assign n7080 = n6978 & n7079;
  assign n7081 = ~n7050 & n7061;
  assign n7082 = ~n6978 & n7081;
  assign n7083 = ~n7080 & ~n7082;
  assign n7084 = ~n7069 & n7083;
  assign n7085 = n7067 & n7084;
  assign n7086 = ~n6922 & n7085;
  assign n7087 = n7066 & n7083;
  assign n7088 = ~n6923 & ~n7069;
  assign n7089 = ~n7087 & ~n7088;
  assign n7090 = ~n6922 & n7089;
  assign n7091 = ~n7086 & ~n7090;
  assign n7092 = ~n6919 & n7087;
  assign n7093 = ~n6921 & ~n7088;
  assign n7094 = n7092 & n7093;
  assign n7095 = ~n6919 & n7088;
  assign n7096 = ~n6921 & ~n7087;
  assign n7097 = n7095 & n7096;
  assign n7098 = ~n7094 & ~n7097;
  assign n7099 = n7091 & n7098;
  assign n7100 = ~n6855 & ~n7099;
  assign n7101 = ~n6853 & n7100;
  assign n7102 = ~n6487 & ~n6792;
  assign n7103 = ~n6747 & n7102;
  assign n7104 = n6491 & ~n6792;
  assign n7105 = ~n6488 & n7104;
  assign n7106 = ~n7103 & ~n7105;
  assign n7107 = ~n7101 & n7106;
  assign n7108 = ~n6797 & n7107;
  assign n7109 = ~n6853 & ~n6855;
  assign n7110 = n7099 & ~n7109;
  assign n7111 = ~n6484 & ~n6791;
  assign n7112 = ~n6486 & n7111;
  assign n7113 = ~n6732 & n7112;
  assign n7114 = n6795 & n7113;
  assign n7115 = ~n6489 & n7112;
  assign n7116 = ~n6392 & ~n6792;
  assign n7117 = ~n6488 & n7116;
  assign n7118 = ~n6747 & n7117;
  assign n7119 = ~n7115 & ~n7118;
  assign n7120 = ~n7114 & n7119;
  assign n7121 = ~n7110 & n7120;
  assign n7122 = n7108 & n7121;
  assign n7123 = ~n7101 & ~n7110;
  assign n7124 = ~n6797 & n7106;
  assign n7125 = n7120 & n7124;
  assign n7126 = ~n7123 & ~n7125;
  assign n7127 = ~n7122 & ~n7126;
  assign n7128 = ~n6789 & ~n7127;
  assign n7129 = n6789 & n7127;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~n6787 & n7130;
  assign n7132 = ~n6766 & ~n7130;
  assign n7133 = ~n6786 & n7132;
  assign po36 = ~n7131 & ~n7133;
  assign n7135 = n3434 & ~n3705;
  assign n7136 = ~n4549 & n7135;
  assign n7137 = ~n4550 & n7136;
  assign n7138 = ~n4854 & n6127;
  assign n7139 = n4557 & n6107;
  assign n7140 = n7138 & n7139;
  assign n7141 = n7137 & n7140;
  assign n7142 = ~n4854 & ~n7141;
  assign n7143 = n2710 & n3181;
  assign n7144 = n2051 & ~n2256;
  assign n7145 = ~n2259 & n7144;
  assign n7146 = ~n2474 & n7145;
  assign n7147 = n2947 & n7146;
  assign n7148 = n7143 & n7147;
  assign n7149 = ~n3179 & ~n4854;
  assign n7150 = ~n7148 & n7149;
  assign n7151 = ~n3198 & n7150;
  assign n7152 = ~n7142 & ~n7151;
  assign n7153 = n3447 & n4551;
  assign n7154 = ~n2944 & ~n3705;
  assign n7155 = n3188 & n7154;
  assign n7156 = n7139 & n7155;
  assign n7157 = n7138 & n7156;
  assign n7158 = n7153 & n7157;
  assign n7159 = ~n2062 & n7158;
  assign n7160 = ~n4550 & n4855;
  assign n7161 = ~n4561 & n7160;
  assign n7162 = n3431 & ~n3705;
  assign n7163 = ~n4549 & n7162;
  assign n7164 = ~n4550 & n7163;
  assign n7165 = n7140 & n7164;
  assign n7166 = ~n5159 & ~n7165;
  assign n7167 = ~n7161 & n7166;
  assign n7168 = ~n7159 & n7167;
  assign n7169 = ~n7152 & n7168;
  assign n7170 = n6421 & n6767;
  assign n7171 = n5797 & n6102;
  assign n7172 = ~n5160 & ~n7128;
  assign n7173 = ~n7129 & n7172;
  assign n7174 = n5481 & n7173;
  assign n7175 = n7171 & n7174;
  assign n7176 = n7170 & n7175;
  assign n7177 = ~n7169 & n7176;
  assign n7178 = ~n6766 & ~n7128;
  assign n7179 = ~n7129 & ~n7178;
  assign n7180 = ~n6419 & n7130;
  assign n7181 = n6767 & n7180;
  assign n7182 = ~n6780 & n7181;
  assign n7183 = ~n7179 & ~n7182;
  assign n7184 = ~n7177 & n7183;
  assign n7185 = ~n6490 & ~n6749;
  assign n7186 = ~n6792 & ~n7185;
  assign n7187 = n7123 & ~n7125;
  assign n7188 = ~n7186 & ~n7187;
  assign n7189 = n6922 & ~n7088;
  assign n7190 = ~n7090 & ~n7097;
  assign n7191 = ~n7189 & n7190;
  assign n7192 = ~n6913 & ~n6918;
  assign n7193 = ~n6814 & ~n6823;
  assign n7194 = ~n6821 & n7193;
  assign n7195 = ~n6812 & n7194;
  assign n7196 = ~n6837 & ~n7195;
  assign n7197 = pi06 & ~n5091;
  assign n7198 = ~n5092 & n7197;
  assign n7199 = ~n5178 & n7198;
  assign n7200 = pi07 & ~n5093;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = pi63 & ~n7201;
  assign n7203 = ~pi63 & ~n7200;
  assign n7204 = ~n7199 & n7203;
  assign n7205 = ~n7202 & ~n7204;
  assign n7206 = pi08 & ~n4513;
  assign n7207 = ~n4514 & n7206;
  assign n7208 = ~n4577 & n7207;
  assign n7209 = pi09 & ~n4515;
  assign n7210 = ~n7208 & ~n7209;
  assign n7211 = pi61 & ~n7210;
  assign n7212 = ~pi61 & ~n7209;
  assign n7213 = ~n7208 & n7212;
  assign n7214 = ~n7211 & ~n7213;
  assign n7215 = ~n7205 & n7214;
  assign n7216 = n7205 & ~n7214;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = pi10 & ~n3959;
  assign n7219 = ~n3960 & n7218;
  assign n7220 = ~n4233 & n7219;
  assign n7221 = pi11 & ~n3961;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = pi59 & ~n7222;
  assign n7224 = ~pi59 & ~n7221;
  assign n7225 = ~n7220 & n7224;
  assign n7226 = ~n7223 & ~n7225;
  assign n7227 = ~n7217 & n7226;
  assign n7228 = ~n7215 & ~n7226;
  assign n7229 = ~n7216 & n7228;
  assign n7230 = ~n7227 & ~n7229;
  assign n7231 = ~n7196 & n7230;
  assign n7232 = n7196 & ~n7230;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = n6841 & ~n7233;
  assign n7235 = ~n6841 & ~n7231;
  assign n7236 = ~n7232 & n7235;
  assign n7237 = ~n7234 & ~n7236;
  assign n7238 = ~n6912 & n7237;
  assign n7239 = ~n7192 & n7238;
  assign n7240 = ~n6912 & ~n7192;
  assign n7241 = ~n7237 & ~n7240;
  assign n7242 = ~n7239 & ~n7241;
  assign n7243 = ~n7191 & n7242;
  assign n7244 = ~n7189 & ~n7242;
  assign n7245 = n7190 & n7244;
  assign n7246 = ~n6868 & ~n6908;
  assign n7247 = pi12 & ~n3205;
  assign n7248 = ~n3206 & n7247;
  assign n7249 = ~n3463 & n7248;
  assign n7250 = pi13 & ~n3207;
  assign n7251 = ~n7249 & ~n7250;
  assign n7252 = pi57 & ~n7251;
  assign n7253 = ~pi57 & ~n7250;
  assign n7254 = ~n7249 & n7253;
  assign n7255 = ~n7252 & ~n7254;
  assign n7256 = ~n6890 & n6900;
  assign n7257 = ~n6887 & ~n7256;
  assign n7258 = n7255 & ~n7257;
  assign n7259 = pi14 & ~n2876;
  assign n7260 = ~n2877 & n7259;
  assign n7261 = ~n2960 & n7260;
  assign n7262 = pi15 & ~n2878;
  assign n7263 = ~n7261 & ~n7262;
  assign n7264 = pi55 & ~n7263;
  assign n7265 = pi16 & ~n2288;
  assign n7266 = ~n2289 & n7265;
  assign n7267 = ~n2647 & n7266;
  assign n7268 = pi17 & ~n2290;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = pi53 & ~n7269;
  assign n7271 = ~pi53 & ~n7268;
  assign n7272 = ~n7267 & n7271;
  assign n7273 = ~pi55 & ~n7262;
  assign n7274 = ~n7261 & n7273;
  assign n7275 = ~n7272 & ~n7274;
  assign n7276 = ~n7270 & n7275;
  assign n7277 = ~n7264 & n7276;
  assign n7278 = ~n7270 & ~n7272;
  assign n7279 = ~n7264 & ~n7274;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = ~n7277 & ~n7280;
  assign n7282 = pi18 & ~n2023;
  assign n7283 = ~n2024 & n7282;
  assign n7284 = ~n2079 & n7283;
  assign n7285 = pi19 & ~n2025;
  assign n7286 = ~n7284 & ~n7285;
  assign n7287 = pi51 & ~n7286;
  assign n7288 = ~pi51 & ~n7285;
  assign n7289 = ~n7284 & n7288;
  assign n7290 = ~n7287 & ~n7289;
  assign n7291 = ~n7281 & n7290;
  assign n7292 = ~n7277 & ~n7290;
  assign n7293 = ~n7280 & n7292;
  assign n7294 = ~n7291 & ~n7293;
  assign n7295 = ~n6887 & ~n7255;
  assign n7296 = ~n7256 & n7295;
  assign n7297 = ~n7294 & ~n7296;
  assign n7298 = ~n7258 & n7297;
  assign n7299 = ~n7258 & ~n7296;
  assign n7300 = n7294 & ~n7299;
  assign n7301 = ~n7298 & ~n7300;
  assign n7302 = ~n7246 & n7301;
  assign n7303 = n7246 & ~n7301;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = ~n6958 & ~n6970;
  assign n7306 = n6959 & ~n6961;
  assign n7307 = ~n6963 & ~n7306;
  assign n7308 = ~n7305 & ~n7307;
  assign n7309 = ~n7304 & n7308;
  assign n7310 = ~n7302 & ~n7308;
  assign n7311 = ~n7303 & n7310;
  assign n7312 = ~n7309 & ~n7311;
  assign n7313 = ~n6978 & ~n7061;
  assign n7314 = n6978 & n7061;
  assign n7315 = n7050 & ~n7314;
  assign n7316 = ~n7313 & ~n7315;
  assign n7317 = n6662 & ~n7010;
  assign n7318 = ~n6997 & n7317;
  assign n7319 = ~n7000 & n7318;
  assign n7320 = ~n7007 & n7028;
  assign n7321 = ~n7001 & n7320;
  assign n7322 = ~n7010 & ~n7016;
  assign n7323 = ~n6997 & n7322;
  assign n7324 = ~n7000 & n7323;
  assign n7325 = ~n7321 & ~n7324;
  assign n7326 = ~n7319 & n7325;
  assign n7327 = pi26 & ~n683;
  assign n7328 = ~n684 & n7327;
  assign n7329 = ~n1231 & n7328;
  assign n7330 = pi27 & ~n685;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = pi43 & ~n7331;
  assign n7333 = pi28 & ~n489;
  assign n7334 = ~n490 & n7333;
  assign n7335 = ~n572 & n7334;
  assign n7336 = pi29 & ~n491;
  assign n7337 = ~n7335 & ~n7336;
  assign n7338 = pi41 & ~n7337;
  assign n7339 = ~pi41 & ~n7336;
  assign n7340 = ~n7335 & n7339;
  assign n7341 = ~pi43 & ~n7330;
  assign n7342 = ~n7329 & n7341;
  assign n7343 = ~n7340 & ~n7342;
  assign n7344 = ~n7338 & n7343;
  assign n7345 = ~n7332 & n7344;
  assign n7346 = ~n7338 & ~n7340;
  assign n7347 = ~n7332 & ~n7342;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = ~n7345 & ~n7348;
  assign n7350 = pi30 & ~n304;
  assign n7351 = ~n305 & n7350;
  assign n7352 = ~n394 & n7351;
  assign n7353 = pi31 & ~n306;
  assign n7354 = ~n7352 & ~n7353;
  assign n7355 = pi39 & ~n7354;
  assign n7356 = ~pi39 & ~n7353;
  assign n7357 = ~n7352 & n7356;
  assign n7358 = ~n7355 & ~n7357;
  assign n7359 = ~n7349 & n7358;
  assign n7360 = ~n7017 & ~n7359;
  assign n7361 = ~n7345 & ~n7358;
  assign n7362 = ~n7348 & n7361;
  assign n7363 = ~n7001 & n7020;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = n7360 & n7364;
  assign n7366 = n7326 & n7365;
  assign n7367 = pi20 & ~n1607;
  assign n7368 = ~n1608 & n7367;
  assign n7369 = ~n1782 & n7368;
  assign n7370 = pi21 & ~n1609;
  assign n7371 = ~n7369 & ~n7370;
  assign n7372 = pi49 & ~n7371;
  assign n7373 = pi22 & ~n1212;
  assign n7374 = ~n1213 & n7373;
  assign n7375 = ~n1425 & n7374;
  assign n7376 = pi23 & ~n1214;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = pi47 & ~n7377;
  assign n7379 = ~pi47 & ~n7376;
  assign n7380 = ~n7375 & n7379;
  assign n7381 = ~pi49 & ~n7370;
  assign n7382 = ~n7369 & n7381;
  assign n7383 = ~n7380 & ~n7382;
  assign n7384 = ~n7378 & n7383;
  assign n7385 = ~n7372 & n7384;
  assign n7386 = ~n7378 & ~n7380;
  assign n7387 = ~n7372 & ~n7382;
  assign n7388 = ~n7386 & ~n7387;
  assign n7389 = ~n7385 & ~n7388;
  assign n7390 = pi24 & ~n1006;
  assign n7391 = ~n1007 & n7390;
  assign n7392 = ~n1068 & n7391;
  assign n7393 = pi25 & ~n1008;
  assign n7394 = ~n7392 & ~n7393;
  assign n7395 = pi45 & ~n7394;
  assign n7396 = ~pi45 & ~n7393;
  assign n7397 = ~n7392 & n7396;
  assign n7398 = ~n7395 & ~n7397;
  assign n7399 = ~n7389 & n7398;
  assign n7400 = ~n6945 & n6955;
  assign n7401 = ~n6942 & ~n7400;
  assign n7402 = ~n7399 & n7401;
  assign n7403 = ~n7385 & ~n7398;
  assign n7404 = ~n7388 & n7403;
  assign n7405 = ~n7000 & n7010;
  assign n7406 = ~n6997 & ~n7405;
  assign n7407 = ~n7404 & ~n7406;
  assign n7408 = n7402 & n7407;
  assign n7409 = ~n7399 & n7406;
  assign n7410 = ~n7401 & ~n7404;
  assign n7411 = n7409 & n7410;
  assign n7412 = ~n7408 & ~n7411;
  assign n7413 = ~n7399 & ~n7404;
  assign n7414 = ~n7401 & ~n7406;
  assign n7415 = ~n7413 & n7414;
  assign n7416 = ~n6942 & ~n6997;
  assign n7417 = ~n7405 & n7416;
  assign n7418 = ~n7400 & n7417;
  assign n7419 = ~n7413 & n7418;
  assign n7420 = ~n7415 & ~n7419;
  assign n7421 = n7412 & n7420;
  assign n7422 = n7366 & n7421;
  assign n7423 = ~n7411 & ~n7415;
  assign n7424 = ~n7419 & n7423;
  assign n7425 = ~n7017 & ~n7363;
  assign n7426 = n7326 & n7425;
  assign n7427 = ~n7359 & ~n7362;
  assign n7428 = ~n7408 & ~n7427;
  assign n7429 = ~n7426 & n7428;
  assign n7430 = n7424 & n7429;
  assign n7431 = ~n7422 & ~n7430;
  assign n7432 = ~n7426 & n7427;
  assign n7433 = ~n7421 & n7432;
  assign n7434 = n7425 & ~n7427;
  assign n7435 = n7326 & n7434;
  assign n7436 = ~n7421 & n7435;
  assign n7437 = ~n7433 & ~n7436;
  assign n7438 = n7431 & n7437;
  assign n7439 = ~n7316 & ~n7438;
  assign n7440 = ~n7312 & n7439;
  assign n7441 = ~n7309 & n7316;
  assign n7442 = ~n7311 & ~n7438;
  assign n7443 = n7441 & n7442;
  assign n7444 = ~n7440 & ~n7443;
  assign n7445 = ~n7430 & ~n7433;
  assign n7446 = ~n7436 & n7445;
  assign n7447 = ~n7313 & ~n7422;
  assign n7448 = ~n7315 & n7447;
  assign n7449 = n7446 & n7448;
  assign n7450 = ~n7312 & n7449;
  assign n7451 = ~n7309 & n7438;
  assign n7452 = ~n7311 & ~n7316;
  assign n7453 = n7451 & n7452;
  assign n7454 = ~n7450 & ~n7453;
  assign n7455 = n7444 & n7454;
  assign n7456 = ~n7245 & ~n7455;
  assign n7457 = ~n7243 & n7456;
  assign n7458 = ~n7243 & ~n7245;
  assign n7459 = n7455 & ~n7458;
  assign n7460 = ~n7457 & ~n7459;
  assign n7461 = n6476 & ~n6841;
  assign n7462 = ~n6842 & n7461;
  assign n7463 = ~n6851 & ~n7462;
  assign n7464 = ~n6798 & ~n7463;
  assign n7465 = n7098 & n7464;
  assign n7466 = ~n6800 & n7091;
  assign n7467 = n7465 & n7466;
  assign n7468 = ~n6852 & n7463;
  assign n7469 = ~n7099 & n7468;
  assign n7470 = ~n6801 & n7468;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = ~n7467 & n7471;
  assign n7473 = ~n6801 & n7463;
  assign n7474 = ~n7099 & n7473;
  assign n7475 = ~n6798 & n6852;
  assign n7476 = ~n7463 & n7475;
  assign n7477 = ~n6800 & n7476;
  assign n7478 = n6852 & ~n7086;
  assign n7479 = ~n7094 & ~n7463;
  assign n7480 = n7190 & n7479;
  assign n7481 = n7478 & n7480;
  assign n7482 = ~n7477 & ~n7481;
  assign n7483 = ~n7474 & n7482;
  assign n7484 = n7472 & n7483;
  assign n7485 = ~n7460 & ~n7484;
  assign n7486 = n7460 & n7484;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = n7188 & n7487;
  assign n7489 = ~n7188 & ~n7487;
  assign n7490 = ~n7488 & ~n7489;
  assign n7491 = ~n7184 & n7490;
  assign n7492 = ~n7179 & ~n7490;
  assign n7493 = ~n7182 & n7492;
  assign n7494 = ~n7177 & n7493;
  assign po37 = ~n7491 & ~n7494;
  assign n7496 = n5168 & ~n5489;
  assign n7497 = ~n5171 & n5501;
  assign n7498 = ~n7496 & n7497;
  assign n7499 = ~n6420 & ~n6765;
  assign n7500 = ~n6766 & n7499;
  assign n7501 = ~n6101 & ~n6419;
  assign n7502 = n6123 & n7501;
  assign n7503 = n7130 & n7490;
  assign n7504 = n6135 & n7503;
  assign n7505 = n7502 & n7504;
  assign n7506 = n7500 & n7505;
  assign n7507 = ~n7498 & n7506;
  assign n7508 = n7129 & ~n7489;
  assign n7509 = ~n7128 & ~n7489;
  assign n7510 = ~n6766 & n7509;
  assign n7511 = ~n7508 & ~n7510;
  assign n7512 = n6420 & n7130;
  assign n7513 = n6767 & n7512;
  assign n7514 = ~n7511 & ~n7513;
  assign n7515 = ~n7488 & ~n7514;
  assign n7516 = ~n6100 & ~n6419;
  assign n7517 = n7503 & n7516;
  assign n7518 = ~n6133 & n7517;
  assign n7519 = n7500 & n7518;
  assign n7520 = ~n7515 & ~n7519;
  assign n7521 = ~n7507 & n7520;
  assign n7522 = ~n6800 & n7475;
  assign n7523 = ~n7110 & ~n7522;
  assign n7524 = ~n7463 & ~n7523;
  assign n7525 = ~n7460 & n7484;
  assign n7526 = ~n7524 & ~n7525;
  assign n7527 = n7312 & ~n7316;
  assign n7528 = n7444 & ~n7527;
  assign n7529 = ~n7303 & ~n7308;
  assign n7530 = ~n7204 & ~n7213;
  assign n7531 = ~n7211 & n7530;
  assign n7532 = ~n7202 & n7531;
  assign n7533 = ~n7227 & ~n7532;
  assign n7534 = pi07 & ~n5091;
  assign n7535 = ~n5092 & n7534;
  assign n7536 = ~n5178 & n7535;
  assign n7537 = pi08 & ~n5093;
  assign n7538 = ~n7536 & ~n7537;
  assign n7539 = pi63 & ~n7538;
  assign n7540 = ~pi63 & ~n7537;
  assign n7541 = ~n7536 & n7540;
  assign n7542 = ~n7539 & ~n7541;
  assign n7543 = pi09 & ~n4513;
  assign n7544 = ~n4514 & n7543;
  assign n7545 = ~n4577 & n7544;
  assign n7546 = pi10 & ~n4515;
  assign n7547 = ~n7545 & ~n7546;
  assign n7548 = pi61 & ~n7547;
  assign n7549 = ~pi61 & ~n7546;
  assign n7550 = ~n7545 & n7549;
  assign n7551 = ~n7548 & ~n7550;
  assign n7552 = ~n7542 & n7551;
  assign n7553 = n7542 & ~n7551;
  assign n7554 = ~n7552 & ~n7553;
  assign n7555 = pi11 & ~n3959;
  assign n7556 = ~n3960 & n7555;
  assign n7557 = ~n4233 & n7556;
  assign n7558 = pi12 & ~n3961;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = pi59 & ~n7559;
  assign n7561 = ~pi59 & ~n7558;
  assign n7562 = ~n7557 & n7561;
  assign n7563 = ~n7560 & ~n7562;
  assign n7564 = ~n7554 & n7563;
  assign n7565 = ~n7552 & ~n7563;
  assign n7566 = ~n7553 & n7565;
  assign n7567 = ~n7564 & ~n7566;
  assign n7568 = ~n7533 & n7567;
  assign n7569 = n7533 & ~n7567;
  assign n7570 = ~n7568 & ~n7569;
  assign n7571 = n7231 & ~n7570;
  assign n7572 = ~n7231 & ~n7568;
  assign n7573 = ~n7569 & n7572;
  assign n7574 = ~n7571 & ~n7573;
  assign n7575 = ~n7302 & n7574;
  assign n7576 = ~n7529 & n7575;
  assign n7577 = ~n7302 & ~n7529;
  assign n7578 = ~n7574 & ~n7577;
  assign n7579 = ~n7576 & ~n7578;
  assign n7580 = ~n7528 & n7579;
  assign n7581 = ~n7527 & ~n7579;
  assign n7582 = n7444 & n7581;
  assign n7583 = ~n7580 & ~n7582;
  assign n7584 = ~n7258 & ~n7298;
  assign n7585 = ~n7280 & n7290;
  assign n7586 = pi13 & ~n3205;
  assign n7587 = ~n3206 & n7586;
  assign n7588 = ~n3463 & n7587;
  assign n7589 = pi14 & ~n3207;
  assign n7590 = ~n7588 & ~n7589;
  assign n7591 = pi57 & ~n7590;
  assign n7592 = ~pi57 & ~n7589;
  assign n7593 = ~n7588 & n7592;
  assign n7594 = ~n7591 & ~n7593;
  assign n7595 = ~n7277 & ~n7594;
  assign n7596 = ~n7585 & n7595;
  assign n7597 = ~n7277 & ~n7585;
  assign n7598 = n7594 & ~n7597;
  assign n7599 = ~n7596 & ~n7598;
  assign n7600 = pi15 & ~n2876;
  assign n7601 = ~n2877 & n7600;
  assign n7602 = ~n2960 & n7601;
  assign n7603 = pi16 & ~n2878;
  assign n7604 = ~n7602 & ~n7603;
  assign n7605 = pi55 & ~n7604;
  assign n7606 = pi17 & ~n2288;
  assign n7607 = ~n2289 & n7606;
  assign n7608 = ~n2647 & n7607;
  assign n7609 = pi18 & ~n2290;
  assign n7610 = ~n7608 & ~n7609;
  assign n7611 = pi53 & ~n7610;
  assign n7612 = ~pi53 & ~n7609;
  assign n7613 = ~n7608 & n7612;
  assign n7614 = ~pi55 & ~n7603;
  assign n7615 = ~n7602 & n7614;
  assign n7616 = ~n7613 & ~n7615;
  assign n7617 = ~n7611 & n7616;
  assign n7618 = ~n7605 & n7617;
  assign n7619 = ~n7611 & ~n7613;
  assign n7620 = ~n7605 & ~n7615;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = ~n7618 & ~n7621;
  assign n7623 = pi19 & ~n2023;
  assign n7624 = ~n2024 & n7623;
  assign n7625 = ~n2079 & n7624;
  assign n7626 = pi20 & ~n2025;
  assign n7627 = ~n7625 & ~n7626;
  assign n7628 = pi51 & ~n7627;
  assign n7629 = ~pi51 & ~n7626;
  assign n7630 = ~n7625 & n7629;
  assign n7631 = ~n7628 & ~n7630;
  assign n7632 = ~n7622 & n7631;
  assign n7633 = ~n7618 & ~n7631;
  assign n7634 = ~n7621 & n7633;
  assign n7635 = ~n7632 & ~n7634;
  assign n7636 = ~n7599 & n7635;
  assign n7637 = n7599 & ~n7635;
  assign n7638 = ~n7636 & ~n7637;
  assign n7639 = ~n7584 & n7638;
  assign n7640 = n7584 & ~n7638;
  assign n7641 = ~n7639 & ~n7640;
  assign n7642 = ~n7401 & ~n7413;
  assign n7643 = n7402 & ~n7404;
  assign n7644 = ~n7406 & ~n7643;
  assign n7645 = ~n7642 & ~n7644;
  assign n7646 = ~n7641 & n7645;
  assign n7647 = ~n7639 & ~n7645;
  assign n7648 = ~n7640 & n7647;
  assign n7649 = ~n7646 & ~n7648;
  assign n7650 = ~n7421 & ~n7426;
  assign n7651 = pi21 & ~n1607;
  assign n7652 = ~n1608 & n7651;
  assign n7653 = ~n1782 & n7652;
  assign n7654 = pi22 & ~n1609;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = pi49 & ~n7655;
  assign n7657 = pi23 & ~n1212;
  assign n7658 = ~n1213 & n7657;
  assign n7659 = ~n1425 & n7658;
  assign n7660 = pi24 & ~n1214;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = pi47 & ~n7661;
  assign n7663 = ~pi47 & ~n7660;
  assign n7664 = ~n7659 & n7663;
  assign n7665 = ~pi49 & ~n7654;
  assign n7666 = ~n7653 & n7665;
  assign n7667 = ~n7664 & ~n7666;
  assign n7668 = ~n7662 & n7667;
  assign n7669 = ~n7656 & n7668;
  assign n7670 = ~n7662 & ~n7664;
  assign n7671 = ~n7656 & ~n7666;
  assign n7672 = ~n7670 & ~n7671;
  assign n7673 = ~n7669 & ~n7672;
  assign n7674 = pi25 & ~n1006;
  assign n7675 = ~n1007 & n7674;
  assign n7676 = ~n1068 & n7675;
  assign n7677 = pi26 & ~n1008;
  assign n7678 = ~n7676 & ~n7677;
  assign n7679 = pi45 & ~n7678;
  assign n7680 = ~pi45 & ~n7677;
  assign n7681 = ~n7676 & n7680;
  assign n7682 = ~n7679 & ~n7681;
  assign n7683 = ~n7673 & n7682;
  assign n7684 = ~n7388 & n7398;
  assign n7685 = ~n7385 & ~n7684;
  assign n7686 = ~n7683 & n7685;
  assign n7687 = ~n7669 & ~n7682;
  assign n7688 = ~n7672 & n7687;
  assign n7689 = ~n7348 & n7358;
  assign n7690 = ~n7345 & ~n7689;
  assign n7691 = ~n7688 & ~n7690;
  assign n7692 = n7686 & n7691;
  assign n7693 = ~n7683 & n7690;
  assign n7694 = ~n7685 & ~n7688;
  assign n7695 = n7693 & n7694;
  assign n7696 = ~n7692 & ~n7695;
  assign n7697 = ~n7683 & ~n7688;
  assign n7698 = ~n7685 & ~n7690;
  assign n7699 = ~n7697 & n7698;
  assign n7700 = ~n7345 & ~n7385;
  assign n7701 = ~n7689 & n7700;
  assign n7702 = ~n7684 & n7701;
  assign n7703 = ~n7697 & n7702;
  assign n7704 = ~n7699 & ~n7703;
  assign n7705 = n7696 & n7704;
  assign n7706 = pi29 & ~n489;
  assign n7707 = ~n490 & n7706;
  assign n7708 = ~n572 & n7707;
  assign n7709 = pi30 & ~n491;
  assign n7710 = ~n7708 & ~n7709;
  assign n7711 = pi41 & ~n7710;
  assign n7712 = ~pi41 & ~n7709;
  assign n7713 = ~n7708 & n7712;
  assign n7714 = ~n7711 & ~n7713;
  assign n7715 = pi27 & ~n683;
  assign n7716 = ~n684 & n7715;
  assign n7717 = ~n1231 & n7716;
  assign n7718 = pi28 & ~n685;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = pi43 & ~n7719;
  assign n7721 = ~pi43 & ~n7718;
  assign n7722 = ~n7717 & n7721;
  assign n7723 = ~n7720 & ~n7722;
  assign n7724 = ~n7714 & ~n7723;
  assign n7725 = ~n7713 & ~n7722;
  assign n7726 = ~n7711 & n7725;
  assign n7727 = ~n7720 & n7726;
  assign n7728 = n306 & n394;
  assign n7729 = pi31 & pi39;
  assign n7730 = ~n7728 & n7729;
  assign n7731 = pi31 & ~n7728;
  assign n7732 = ~pi39 & ~n7731;
  assign n7733 = ~n7730 & ~n7732;
  assign n7734 = ~n7727 & ~n7733;
  assign n7735 = ~n7724 & n7734;
  assign n7736 = ~n7724 & ~n7727;
  assign n7737 = n7733 & ~n7736;
  assign n7738 = ~n7735 & ~n7737;
  assign n7739 = n7427 & ~n7738;
  assign n7740 = ~n7705 & n7739;
  assign n7741 = ~n7427 & n7738;
  assign n7742 = ~n7705 & n7741;
  assign n7743 = ~n7740 & ~n7742;
  assign n7744 = ~n7650 & n7743;
  assign n7745 = n7421 & n7426;
  assign n7746 = n7427 & ~n7745;
  assign n7747 = n7427 & n7738;
  assign n7748 = ~n7692 & n7747;
  assign n7749 = ~n7695 & ~n7699;
  assign n7750 = ~n7703 & n7749;
  assign n7751 = n7748 & n7750;
  assign n7752 = ~n7427 & ~n7738;
  assign n7753 = ~n7692 & n7752;
  assign n7754 = n7750 & n7753;
  assign n7755 = ~n7751 & ~n7754;
  assign n7756 = ~n7746 & n7755;
  assign n7757 = n7744 & n7756;
  assign n7758 = ~n7649 & n7757;
  assign n7759 = n7743 & n7755;
  assign n7760 = ~n7650 & ~n7746;
  assign n7761 = ~n7759 & ~n7760;
  assign n7762 = ~n7649 & n7761;
  assign n7763 = ~n7758 & ~n7762;
  assign n7764 = ~n7646 & n7759;
  assign n7765 = ~n7648 & ~n7760;
  assign n7766 = n7764 & n7765;
  assign n7767 = ~n7646 & n7760;
  assign n7768 = ~n7648 & ~n7759;
  assign n7769 = n7767 & n7768;
  assign n7770 = ~n7766 & ~n7769;
  assign n7771 = n7763 & n7770;
  assign n7772 = ~n7583 & n7771;
  assign n7773 = ~n7582 & ~n7771;
  assign n7774 = ~n7580 & n7773;
  assign n7775 = ~n7772 & ~n7774;
  assign n7776 = ~n7245 & n7455;
  assign n7777 = n6841 & ~n7231;
  assign n7778 = ~n7232 & n7777;
  assign n7779 = ~n7241 & ~n7778;
  assign n7780 = ~n7243 & ~n7779;
  assign n7781 = ~n7776 & n7780;
  assign n7782 = ~n7243 & ~n7776;
  assign n7783 = n7779 & ~n7782;
  assign n7784 = ~n7781 & ~n7783;
  assign n7785 = ~n7775 & ~n7784;
  assign n7786 = n7775 & n7784;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = ~n7526 & n7787;
  assign n7789 = n7526 & ~n7787;
  assign n7790 = ~n7788 & ~n7789;
  assign n7791 = ~n7521 & n7790;
  assign n7792 = ~n7515 & ~n7790;
  assign n7793 = ~n7519 & n7792;
  assign n7794 = ~n7507 & n7793;
  assign po38 = ~n7791 & ~n7794;
  assign n7796 = n7171 & n7503;
  assign n7797 = n7170 & n7796;
  assign n7798 = n5803 & n7797;
  assign n7799 = ~n3992 & n7798;
  assign n7800 = ~n5812 & n7797;
  assign n7801 = n7520 & ~n7800;
  assign n7802 = ~n7799 & n7801;
  assign n7803 = ~n7789 & ~n7802;
  assign n7804 = ~n7788 & ~n7803;
  assign n7805 = n7649 & ~n7760;
  assign n7806 = ~n7762 & ~n7769;
  assign n7807 = ~n7805 & n7806;
  assign n7808 = ~n7640 & ~n7645;
  assign n7809 = ~n7541 & ~n7550;
  assign n7810 = ~n7548 & n7809;
  assign n7811 = ~n7539 & n7810;
  assign n7812 = ~n7564 & ~n7811;
  assign n7813 = pi08 & ~n5091;
  assign n7814 = ~n5092 & n7813;
  assign n7815 = ~n5178 & n7814;
  assign n7816 = pi09 & ~n5093;
  assign n7817 = ~n7815 & ~n7816;
  assign n7818 = pi63 & ~n7817;
  assign n7819 = ~pi63 & ~n7816;
  assign n7820 = ~n7815 & n7819;
  assign n7821 = ~n7818 & ~n7820;
  assign n7822 = pi10 & ~n4513;
  assign n7823 = ~n4514 & n7822;
  assign n7824 = ~n4577 & n7823;
  assign n7825 = pi11 & ~n4515;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = pi61 & ~n7826;
  assign n7828 = ~pi61 & ~n7825;
  assign n7829 = ~n7824 & n7828;
  assign n7830 = ~n7827 & ~n7829;
  assign n7831 = ~n7821 & n7830;
  assign n7832 = n7821 & ~n7830;
  assign n7833 = ~n7831 & ~n7832;
  assign n7834 = pi12 & ~n3959;
  assign n7835 = ~n3960 & n7834;
  assign n7836 = ~n4233 & n7835;
  assign n7837 = pi13 & ~n3961;
  assign n7838 = ~n7836 & ~n7837;
  assign n7839 = pi59 & ~n7838;
  assign n7840 = ~pi59 & ~n7837;
  assign n7841 = ~n7836 & n7840;
  assign n7842 = ~n7839 & ~n7841;
  assign n7843 = ~n7833 & n7842;
  assign n7844 = ~n7831 & ~n7842;
  assign n7845 = ~n7832 & n7844;
  assign n7846 = ~n7843 & ~n7845;
  assign n7847 = ~n7812 & n7846;
  assign n7848 = n7812 & ~n7846;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = n7568 & ~n7849;
  assign n7851 = ~n7568 & ~n7847;
  assign n7852 = ~n7848 & n7851;
  assign n7853 = ~n7850 & ~n7852;
  assign n7854 = ~n7639 & n7853;
  assign n7855 = ~n7808 & n7854;
  assign n7856 = ~n7639 & ~n7808;
  assign n7857 = ~n7853 & ~n7856;
  assign n7858 = ~n7855 & ~n7857;
  assign n7859 = ~n7807 & n7858;
  assign n7860 = ~n7805 & ~n7858;
  assign n7861 = n7806 & n7860;
  assign n7862 = ~n7598 & ~n7637;
  assign n7863 = ~n7621 & n7631;
  assign n7864 = pi14 & ~n3205;
  assign n7865 = ~n3206 & n7864;
  assign n7866 = ~n3463 & n7865;
  assign n7867 = pi15 & ~n3207;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = pi57 & ~n7868;
  assign n7870 = ~pi57 & ~n7867;
  assign n7871 = ~n7866 & n7870;
  assign n7872 = ~n7869 & ~n7871;
  assign n7873 = ~n7618 & ~n7872;
  assign n7874 = ~n7863 & n7873;
  assign n7875 = ~n7618 & ~n7863;
  assign n7876 = n7872 & ~n7875;
  assign n7877 = ~n7874 & ~n7876;
  assign n7878 = pi16 & ~n2876;
  assign n7879 = ~n2877 & n7878;
  assign n7880 = ~n2960 & n7879;
  assign n7881 = pi17 & ~n2878;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = pi55 & ~n7882;
  assign n7884 = pi18 & ~n2288;
  assign n7885 = ~n2289 & n7884;
  assign n7886 = ~n2647 & n7885;
  assign n7887 = pi19 & ~n2290;
  assign n7888 = ~n7886 & ~n7887;
  assign n7889 = pi53 & ~n7888;
  assign n7890 = ~pi53 & ~n7887;
  assign n7891 = ~n7886 & n7890;
  assign n7892 = ~pi55 & ~n7881;
  assign n7893 = ~n7880 & n7892;
  assign n7894 = ~n7891 & ~n7893;
  assign n7895 = ~n7889 & n7894;
  assign n7896 = ~n7883 & n7895;
  assign n7897 = ~n7889 & ~n7891;
  assign n7898 = ~n7883 & ~n7893;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = ~n7896 & ~n7899;
  assign n7901 = pi20 & ~n2023;
  assign n7902 = ~n2024 & n7901;
  assign n7903 = ~n2079 & n7902;
  assign n7904 = pi21 & ~n2025;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = pi51 & ~n7905;
  assign n7907 = ~pi51 & ~n7904;
  assign n7908 = ~n7903 & n7907;
  assign n7909 = ~n7906 & ~n7908;
  assign n7910 = ~n7900 & n7909;
  assign n7911 = ~n7896 & ~n7909;
  assign n7912 = ~n7899 & n7911;
  assign n7913 = ~n7910 & ~n7912;
  assign n7914 = ~n7877 & n7913;
  assign n7915 = n7877 & ~n7913;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = ~n7862 & n7916;
  assign n7918 = n7862 & ~n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = ~n7685 & ~n7697;
  assign n7921 = n7686 & ~n7688;
  assign n7922 = ~n7690 & ~n7921;
  assign n7923 = ~n7920 & ~n7922;
  assign n7924 = ~n7919 & n7923;
  assign n7925 = ~n7917 & ~n7923;
  assign n7926 = ~n7918 & n7925;
  assign n7927 = ~n7924 & ~n7926;
  assign n7928 = n7427 & ~n7692;
  assign n7929 = n7750 & n7928;
  assign n7930 = n7738 & ~n7929;
  assign n7931 = pi22 & ~n1607;
  assign n7932 = ~n1608 & n7931;
  assign n7933 = ~n1782 & n7932;
  assign n7934 = pi23 & ~n1609;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = pi49 & ~n7935;
  assign n7937 = pi24 & ~n1212;
  assign n7938 = ~n1213 & n7937;
  assign n7939 = ~n1425 & n7938;
  assign n7940 = pi25 & ~n1214;
  assign n7941 = ~n7939 & ~n7940;
  assign n7942 = pi47 & ~n7941;
  assign n7943 = ~pi47 & ~n7940;
  assign n7944 = ~n7939 & n7943;
  assign n7945 = ~pi49 & ~n7934;
  assign n7946 = ~n7933 & n7945;
  assign n7947 = ~n7944 & ~n7946;
  assign n7948 = ~n7942 & n7947;
  assign n7949 = ~n7936 & n7948;
  assign n7950 = ~n7942 & ~n7944;
  assign n7951 = ~n7936 & ~n7946;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = ~n7949 & ~n7952;
  assign n7954 = pi26 & ~n1006;
  assign n7955 = ~n1007 & n7954;
  assign n7956 = ~n1068 & n7955;
  assign n7957 = pi27 & ~n1008;
  assign n7958 = ~n7956 & ~n7957;
  assign n7959 = pi45 & ~n7958;
  assign n7960 = ~pi45 & ~n7957;
  assign n7961 = ~n7956 & n7960;
  assign n7962 = ~n7959 & ~n7961;
  assign n7963 = ~n7953 & n7962;
  assign n7964 = ~n7672 & n7682;
  assign n7965 = ~n7669 & ~n7964;
  assign n7966 = ~n7963 & n7965;
  assign n7967 = ~n7949 & ~n7962;
  assign n7968 = ~n7952 & n7967;
  assign n7969 = ~n7724 & ~n7733;
  assign n7970 = ~n7727 & ~n7969;
  assign n7971 = ~n7968 & ~n7970;
  assign n7972 = n7966 & n7971;
  assign n7973 = ~n7963 & n7970;
  assign n7974 = ~n7965 & ~n7968;
  assign n7975 = n7973 & n7974;
  assign n7976 = ~n7972 & ~n7975;
  assign n7977 = ~n7963 & ~n7968;
  assign n7978 = ~n7965 & ~n7970;
  assign n7979 = ~n7977 & n7978;
  assign n7980 = ~n7669 & ~n7727;
  assign n7981 = ~n7969 & n7980;
  assign n7982 = ~n7964 & n7981;
  assign n7983 = ~n7977 & n7982;
  assign n7984 = ~n7979 & ~n7983;
  assign n7985 = n7976 & n7984;
  assign n7986 = pi30 & ~n489;
  assign n7987 = ~n490 & n7986;
  assign n7988 = ~n572 & n7987;
  assign n7989 = pi31 & ~n491;
  assign n7990 = ~n7988 & ~n7989;
  assign n7991 = pi41 & ~n7990;
  assign n7992 = pi28 & ~n683;
  assign n7993 = ~n684 & n7992;
  assign n7994 = ~n1231 & n7993;
  assign n7995 = pi29 & ~n685;
  assign n7996 = ~n7994 & ~n7995;
  assign n7997 = pi43 & ~n7996;
  assign n7998 = ~pi43 & ~n7995;
  assign n7999 = ~n7994 & n7998;
  assign n8000 = ~pi41 & ~n7989;
  assign n8001 = ~n7988 & n8000;
  assign n8002 = ~n7999 & ~n8001;
  assign n8003 = ~n7997 & n8002;
  assign n8004 = ~n7991 & n8003;
  assign n8005 = ~n7997 & ~n7999;
  assign n8006 = ~n7991 & ~n8001;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = ~n8004 & ~n8007;
  assign n8009 = ~n7985 & ~n8008;
  assign n8010 = ~n7972 & n8008;
  assign n8011 = ~n7975 & ~n7979;
  assign n8012 = ~n7983 & n8011;
  assign n8013 = n8010 & n8012;
  assign n8014 = ~n8009 & ~n8013;
  assign n8015 = ~n7427 & ~n7705;
  assign n8016 = ~n8014 & ~n8015;
  assign n8017 = ~n7930 & n8016;
  assign n8018 = ~n7927 & n8017;
  assign n8019 = ~n7930 & ~n8015;
  assign n8020 = n8014 & ~n8019;
  assign n8021 = ~n7927 & n8020;
  assign n8022 = ~n8018 & ~n8021;
  assign n8023 = ~n7924 & ~n8014;
  assign n8024 = ~n7926 & ~n8019;
  assign n8025 = n8023 & n8024;
  assign n8026 = n8014 & n8019;
  assign n8027 = n7927 & n8026;
  assign n8028 = ~n8025 & ~n8027;
  assign n8029 = n8022 & n8028;
  assign n8030 = ~n7861 & ~n8029;
  assign n8031 = ~n7859 & n8030;
  assign n8032 = ~n7859 & ~n7861;
  assign n8033 = n8029 & ~n8032;
  assign n8034 = ~n8031 & ~n8033;
  assign n8035 = ~n7582 & n7771;
  assign n8036 = n7231 & ~n7568;
  assign n8037 = ~n7569 & n8036;
  assign n8038 = ~n7578 & ~n8037;
  assign n8039 = ~n7580 & ~n8038;
  assign n8040 = ~n8035 & n8039;
  assign n8041 = ~n7580 & ~n8035;
  assign n8042 = n8038 & ~n8041;
  assign n8043 = ~n8040 & ~n8042;
  assign n8044 = ~n8034 & ~n8043;
  assign n8045 = n8034 & n8043;
  assign n8046 = ~n8044 & ~n8045;
  assign n8047 = ~n7779 & ~n7782;
  assign n8048 = ~n7785 & ~n8047;
  assign n8049 = ~n8046 & n8048;
  assign n8050 = n8046 & ~n8048;
  assign n8051 = ~n8049 & ~n8050;
  assign n8052 = ~n7804 & n8051;
  assign n8053 = ~n7788 & ~n8051;
  assign n8054 = ~n7803 & n8053;
  assign po39 = ~n8052 & ~n8054;
  assign n8056 = n4261 & ~n4853;
  assign n8057 = ~n4549 & n8056;
  assign n8058 = n5807 & n8057;
  assign n8059 = n5491 & n8058;
  assign n8060 = ~n5503 & ~n8059;
  assign n8061 = ~n5796 & ~n8060;
  assign n8062 = n6128 & n7139;
  assign n8063 = n5807 & n8062;
  assign n8064 = n3452 & ~n4550;
  assign n8065 = n6110 & n8064;
  assign n8066 = n6428 & n8065;
  assign n8067 = n8063 & n8066;
  assign n8068 = ~n2713 & n8067;
  assign n8069 = ~n3981 & ~n4261;
  assign n8070 = ~n4550 & n8069;
  assign n8071 = n6128 & n8070;
  assign n8072 = n5807 & n8071;
  assign n8073 = n6428 & n8072;
  assign n8074 = ~n6119 & n8073;
  assign n8075 = ~n5795 & ~n8074;
  assign n8076 = ~n8068 & n8075;
  assign n8077 = ~n8061 & n8076;
  assign n8078 = n7790 & n8051;
  assign n8079 = n6102 & n7503;
  assign n8080 = n8078 & n8079;
  assign n8081 = n7170 & n8080;
  assign n8082 = ~n8077 & n8081;
  assign n8083 = ~n7488 & ~n7788;
  assign n8084 = ~n7789 & ~n8049;
  assign n8085 = ~n8050 & n8084;
  assign n8086 = n8083 & n8085;
  assign n8087 = ~n7514 & n8086;
  assign n8088 = n6101 & ~n6419;
  assign n8089 = n7503 & n8088;
  assign n8090 = n8078 & n8089;
  assign n8091 = n7500 & n8090;
  assign n8092 = ~n7788 & ~n8050;
  assign n8093 = ~n8049 & ~n8092;
  assign n8094 = ~n8091 & ~n8093;
  assign n8095 = ~n8087 & n8094;
  assign n8096 = ~n8082 & n8095;
  assign n8097 = ~n8038 & ~n8041;
  assign n8098 = ~n8044 & ~n8097;
  assign n8099 = ~n7876 & ~n7915;
  assign n8100 = pi17 & ~n2876;
  assign n8101 = ~n2877 & n8100;
  assign n8102 = ~n2960 & n8101;
  assign n8103 = pi18 & ~n2878;
  assign n8104 = ~n8102 & ~n8103;
  assign n8105 = pi55 & ~n8104;
  assign n8106 = pi19 & ~n2288;
  assign n8107 = ~n2289 & n8106;
  assign n8108 = ~n2647 & n8107;
  assign n8109 = pi20 & ~n2290;
  assign n8110 = ~n8108 & ~n8109;
  assign n8111 = pi53 & ~n8110;
  assign n8112 = ~pi53 & ~n8109;
  assign n8113 = ~n8108 & n8112;
  assign n8114 = ~pi55 & ~n8103;
  assign n8115 = ~n8102 & n8114;
  assign n8116 = ~n8113 & ~n8115;
  assign n8117 = ~n8111 & n8116;
  assign n8118 = ~n8105 & n8117;
  assign n8119 = ~n8111 & ~n8113;
  assign n8120 = ~n8105 & ~n8115;
  assign n8121 = ~n8119 & ~n8120;
  assign n8122 = ~n8118 & ~n8121;
  assign n8123 = pi21 & ~n2023;
  assign n8124 = ~n2024 & n8123;
  assign n8125 = ~n2079 & n8124;
  assign n8126 = pi22 & ~n2025;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = pi51 & ~n8127;
  assign n8129 = ~pi51 & ~n8126;
  assign n8130 = ~n8125 & n8129;
  assign n8131 = ~n8128 & ~n8130;
  assign n8132 = ~n8122 & n8131;
  assign n8133 = ~n8118 & ~n8131;
  assign n8134 = ~n8121 & n8133;
  assign n8135 = ~n8132 & ~n8134;
  assign n8136 = ~n7899 & n7909;
  assign n8137 = ~n7896 & ~n8136;
  assign n8138 = pi15 & ~n3205;
  assign n8139 = ~n3206 & n8138;
  assign n8140 = ~n3463 & n8139;
  assign n8141 = pi16 & ~n3207;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = pi57 & ~n8142;
  assign n8144 = ~pi57 & ~n8141;
  assign n8145 = ~n8140 & n8144;
  assign n8146 = ~n8143 & ~n8145;
  assign n8147 = ~n8137 & n8146;
  assign n8148 = ~n7896 & ~n8146;
  assign n8149 = ~n8136 & n8148;
  assign n8150 = ~n8147 & ~n8149;
  assign n8151 = ~n8135 & ~n8150;
  assign n8152 = n8135 & n8150;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = ~n8099 & ~n8153;
  assign n8155 = n8099 & n8153;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = ~n7965 & ~n7977;
  assign n8158 = n7966 & ~n7968;
  assign n8159 = ~n7970 & ~n8158;
  assign n8160 = ~n8157 & ~n8159;
  assign n8161 = ~n8009 & n8160;
  assign n8162 = ~n8156 & n8161;
  assign n8163 = n8009 & ~n8160;
  assign n8164 = ~n8156 & n8163;
  assign n8165 = ~n8162 & ~n8164;
  assign n8166 = ~n8009 & ~n8160;
  assign n8167 = n8156 & n8166;
  assign n8168 = ~n8008 & ~n8157;
  assign n8169 = ~n8159 & n8168;
  assign n8170 = ~n7985 & n8169;
  assign n8171 = ~n8154 & n8170;
  assign n8172 = ~n8155 & n8171;
  assign n8173 = ~n8167 & ~n8172;
  assign n8174 = n8165 & n8173;
  assign n8175 = pi23 & ~n1607;
  assign n8176 = ~n1608 & n8175;
  assign n8177 = ~n1782 & n8176;
  assign n8178 = pi24 & ~n1609;
  assign n8179 = ~n8177 & ~n8178;
  assign n8180 = pi49 & ~n8179;
  assign n8181 = ~pi49 & ~n8178;
  assign n8182 = ~n8177 & n8181;
  assign n8183 = ~n8180 & ~n8182;
  assign n8184 = pi25 & ~n1212;
  assign n8185 = ~n1213 & n8184;
  assign n8186 = ~n1425 & n8185;
  assign n8187 = pi26 & ~n1214;
  assign n8188 = ~n8186 & ~n8187;
  assign n8189 = pi47 & ~n8188;
  assign n8190 = ~pi47 & ~n8187;
  assign n8191 = ~n8186 & n8190;
  assign n8192 = ~n8189 & ~n8191;
  assign n8193 = ~n8183 & n8192;
  assign n8194 = n8183 & ~n8192;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = pi27 & ~n1006;
  assign n8197 = ~n1007 & n8196;
  assign n8198 = ~n1068 & n8197;
  assign n8199 = pi28 & ~n1008;
  assign n8200 = ~n8198 & ~n8199;
  assign n8201 = pi45 & ~n8200;
  assign n8202 = ~pi45 & ~n8199;
  assign n8203 = ~n8198 & n8202;
  assign n8204 = ~n8201 & ~n8203;
  assign n8205 = ~n8195 & n8204;
  assign n8206 = ~n8193 & ~n8204;
  assign n8207 = ~n8194 & n8206;
  assign n8208 = ~n8205 & ~n8207;
  assign n8209 = ~n7952 & n7962;
  assign n8210 = ~n7949 & ~n8209;
  assign n8211 = n491 & n572;
  assign n8212 = pi31 & pi41;
  assign n8213 = ~n8211 & n8212;
  assign n8214 = pi31 & ~n8211;
  assign n8215 = ~pi41 & ~n8214;
  assign n8216 = ~n8213 & ~n8215;
  assign n8217 = pi29 & ~n683;
  assign n8218 = ~n684 & n8217;
  assign n8219 = ~n1231 & n8218;
  assign n8220 = pi30 & ~n685;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = pi43 & ~n8221;
  assign n8223 = ~pi43 & ~n8220;
  assign n8224 = ~n8219 & n8223;
  assign n8225 = ~n8222 & ~n8224;
  assign n8226 = ~n8216 & n8225;
  assign n8227 = n8216 & ~n8225;
  assign n8228 = ~n8226 & ~n8227;
  assign n8229 = ~n8007 & ~n8228;
  assign n8230 = ~n8210 & n8229;
  assign n8231 = ~n8208 & n8230;
  assign n8232 = ~n7949 & n8007;
  assign n8233 = ~n8209 & n8232;
  assign n8234 = ~n8228 & n8233;
  assign n8235 = ~n8208 & n8234;
  assign n8236 = ~n8231 & ~n8235;
  assign n8237 = ~n8207 & ~n8210;
  assign n8238 = n8007 & ~n8228;
  assign n8239 = ~n8205 & n8238;
  assign n8240 = n8237 & n8239;
  assign n8241 = ~n7949 & ~n8007;
  assign n8242 = ~n8209 & n8241;
  assign n8243 = ~n8228 & n8242;
  assign n8244 = n8208 & n8243;
  assign n8245 = ~n8240 & ~n8244;
  assign n8246 = n8236 & n8245;
  assign n8247 = n8007 & ~n8226;
  assign n8248 = ~n8227 & n8247;
  assign n8249 = ~n8210 & n8248;
  assign n8250 = ~n8208 & n8249;
  assign n8251 = n8228 & n8241;
  assign n8252 = ~n8209 & n8251;
  assign n8253 = ~n8208 & n8252;
  assign n8254 = ~n8250 & ~n8253;
  assign n8255 = ~n8007 & ~n8226;
  assign n8256 = ~n8227 & n8255;
  assign n8257 = ~n8205 & n8256;
  assign n8258 = n8237 & n8257;
  assign n8259 = ~n7949 & ~n8227;
  assign n8260 = n8247 & n8259;
  assign n8261 = ~n8209 & n8260;
  assign n8262 = n8208 & n8261;
  assign n8263 = ~n8258 & ~n8262;
  assign n8264 = n8254 & n8263;
  assign n8265 = n8246 & n8264;
  assign n8266 = ~n8174 & n8265;
  assign n8267 = ~n8162 & ~n8265;
  assign n8268 = ~n8164 & ~n8167;
  assign n8269 = ~n8172 & n8268;
  assign n8270 = n8267 & n8269;
  assign n8271 = ~n8266 & ~n8270;
  assign n8272 = n7927 & ~n8019;
  assign n8273 = ~n8021 & ~n8027;
  assign n8274 = ~n8272 & n8273;
  assign n8275 = ~n7918 & ~n7923;
  assign n8276 = ~n7820 & ~n7829;
  assign n8277 = ~n7827 & n8276;
  assign n8278 = ~n7818 & n8277;
  assign n8279 = ~n7843 & ~n8278;
  assign n8280 = pi09 & ~n5091;
  assign n8281 = ~n5092 & n8280;
  assign n8282 = ~n5178 & n8281;
  assign n8283 = pi10 & ~n5093;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = pi63 & ~n8284;
  assign n8286 = ~pi63 & ~n8283;
  assign n8287 = ~n8282 & n8286;
  assign n8288 = ~n8285 & ~n8287;
  assign n8289 = pi11 & ~n4513;
  assign n8290 = ~n4514 & n8289;
  assign n8291 = ~n4577 & n8290;
  assign n8292 = pi12 & ~n4515;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = pi61 & ~n8293;
  assign n8295 = ~pi61 & ~n8292;
  assign n8296 = ~n8291 & n8295;
  assign n8297 = ~n8294 & ~n8296;
  assign n8298 = ~n8288 & n8297;
  assign n8299 = n8288 & ~n8297;
  assign n8300 = ~n8298 & ~n8299;
  assign n8301 = pi13 & ~n3959;
  assign n8302 = ~n3960 & n8301;
  assign n8303 = ~n4233 & n8302;
  assign n8304 = pi14 & ~n3961;
  assign n8305 = ~n8303 & ~n8304;
  assign n8306 = pi59 & ~n8305;
  assign n8307 = ~pi59 & ~n8304;
  assign n8308 = ~n8303 & n8307;
  assign n8309 = ~n8306 & ~n8308;
  assign n8310 = ~n8300 & n8309;
  assign n8311 = ~n8298 & ~n8309;
  assign n8312 = ~n8299 & n8311;
  assign n8313 = ~n8310 & ~n8312;
  assign n8314 = ~n8279 & n8313;
  assign n8315 = n8279 & ~n8313;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = n7847 & ~n8316;
  assign n8318 = ~n7847 & ~n8314;
  assign n8319 = ~n8315 & n8318;
  assign n8320 = ~n8317 & ~n8319;
  assign n8321 = ~n7917 & n8320;
  assign n8322 = ~n8275 & n8321;
  assign n8323 = ~n7917 & ~n8275;
  assign n8324 = ~n8320 & ~n8323;
  assign n8325 = ~n8322 & ~n8324;
  assign n8326 = ~n8274 & n8325;
  assign n8327 = ~n8272 & ~n8325;
  assign n8328 = n8273 & n8327;
  assign n8329 = ~n8326 & ~n8328;
  assign n8330 = ~n8271 & ~n8329;
  assign n8331 = n8271 & ~n8328;
  assign n8332 = ~n8326 & n8331;
  assign n8333 = ~n8330 & ~n8332;
  assign n8334 = ~n7861 & n8029;
  assign n8335 = n7568 & ~n7847;
  assign n8336 = ~n7848 & n8335;
  assign n8337 = ~n7857 & ~n8336;
  assign n8338 = ~n7859 & ~n8337;
  assign n8339 = ~n8334 & n8338;
  assign n8340 = ~n7859 & ~n8334;
  assign n8341 = n8337 & ~n8340;
  assign n8342 = ~n8339 & ~n8341;
  assign n8343 = ~n8333 & ~n8342;
  assign n8344 = n8333 & n8342;
  assign n8345 = ~n8343 & ~n8344;
  assign n8346 = ~n8098 & n8345;
  assign n8347 = n8098 & ~n8345;
  assign n8348 = ~n8346 & ~n8347;
  assign n8349 = ~n8096 & n8348;
  assign n8350 = ~n8093 & ~n8348;
  assign n8351 = ~n8091 & n8350;
  assign n8352 = ~n8087 & n8351;
  assign n8353 = ~n8082 & n8352;
  assign po40 = ~n8349 & ~n8353;
  assign n8355 = n5166 & n7503;
  assign n8356 = n8078 & n8355;
  assign n8357 = n5497 & n7171;
  assign n8358 = n7170 & n8357;
  assign n8359 = n8356 & n8358;
  assign n8360 = ~n4273 & n8359;
  assign n8361 = n7503 & n8078;
  assign n8362 = n7170 & n8361;
  assign n8363 = ~n6138 & n8362;
  assign n8364 = ~n8087 & ~n8093;
  assign n8365 = ~n8363 & n8364;
  assign n8366 = ~n8360 & n8365;
  assign n8367 = ~n8347 & ~n8366;
  assign n8368 = ~n8346 & ~n8367;
  assign n8369 = ~n8337 & ~n8340;
  assign n8370 = ~n8343 & ~n8369;
  assign n8371 = ~n8155 & ~n8160;
  assign n8372 = ~n8287 & ~n8296;
  assign n8373 = ~n8294 & n8372;
  assign n8374 = ~n8285 & n8373;
  assign n8375 = ~n8310 & ~n8374;
  assign n8376 = pi10 & ~n5091;
  assign n8377 = ~n5092 & n8376;
  assign n8378 = ~n5178 & n8377;
  assign n8379 = pi11 & ~n5093;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = pi63 & ~n8380;
  assign n8382 = ~pi63 & ~n8379;
  assign n8383 = ~n8378 & n8382;
  assign n8384 = ~n8381 & ~n8383;
  assign n8385 = pi12 & ~n4513;
  assign n8386 = ~n4514 & n8385;
  assign n8387 = ~n4577 & n8386;
  assign n8388 = pi13 & ~n4515;
  assign n8389 = ~n8387 & ~n8388;
  assign n8390 = pi61 & ~n8389;
  assign n8391 = ~pi61 & ~n8388;
  assign n8392 = ~n8387 & n8391;
  assign n8393 = ~n8390 & ~n8392;
  assign n8394 = ~n8384 & n8393;
  assign n8395 = n8384 & ~n8393;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = pi14 & ~n3959;
  assign n8398 = ~n3960 & n8397;
  assign n8399 = ~n4233 & n8398;
  assign n8400 = pi15 & ~n3961;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = pi59 & ~n8401;
  assign n8403 = ~pi59 & ~n8400;
  assign n8404 = ~n8399 & n8403;
  assign n8405 = ~n8402 & ~n8404;
  assign n8406 = ~n8396 & n8405;
  assign n8407 = ~n8394 & ~n8405;
  assign n8408 = ~n8395 & n8407;
  assign n8409 = ~n8406 & ~n8408;
  assign n8410 = ~n8375 & n8409;
  assign n8411 = n8375 & ~n8409;
  assign n8412 = ~n8410 & ~n8411;
  assign n8413 = n8314 & ~n8412;
  assign n8414 = ~n8314 & ~n8410;
  assign n8415 = ~n8411 & n8414;
  assign n8416 = ~n8413 & ~n8415;
  assign n8417 = ~n8154 & n8416;
  assign n8418 = ~n8371 & n8417;
  assign n8419 = ~n8154 & ~n8371;
  assign n8420 = ~n8416 & ~n8419;
  assign n8421 = ~n8418 & ~n8420;
  assign n8422 = ~n8008 & ~n8250;
  assign n8423 = ~n8253 & ~n8258;
  assign n8424 = ~n8231 & ~n8262;
  assign n8425 = n8423 & n8424;
  assign n8426 = n8422 & n8425;
  assign n8427 = ~n8235 & ~n8240;
  assign n8428 = ~n8244 & n8427;
  assign n8429 = ~n7985 & n8428;
  assign n8430 = n8426 & n8429;
  assign n8431 = ~n8164 & ~n8430;
  assign n8432 = ~n8160 & n8265;
  assign n8433 = ~n8156 & n8432;
  assign n8434 = n8160 & n8265;
  assign n8435 = n8156 & n8434;
  assign n8436 = ~n8172 & ~n8435;
  assign n8437 = ~n8433 & n8436;
  assign n8438 = n8431 & n8437;
  assign n8439 = n8421 & ~n8438;
  assign n8440 = ~n8421 & n8438;
  assign n8441 = pi16 & ~n3205;
  assign n8442 = ~n3206 & n8441;
  assign n8443 = ~n3463 & n8442;
  assign n8444 = pi17 & ~n3207;
  assign n8445 = ~n8443 & ~n8444;
  assign n8446 = pi57 & ~n8445;
  assign n8447 = ~pi57 & ~n8444;
  assign n8448 = ~n8443 & n8447;
  assign n8449 = ~n8446 & ~n8448;
  assign n8450 = ~n8121 & n8131;
  assign n8451 = ~n8118 & ~n8450;
  assign n8452 = n8449 & ~n8451;
  assign n8453 = pi18 & ~n2876;
  assign n8454 = ~n2877 & n8453;
  assign n8455 = ~n2960 & n8454;
  assign n8456 = pi19 & ~n2878;
  assign n8457 = ~n8455 & ~n8456;
  assign n8458 = pi55 & ~n8457;
  assign n8459 = pi20 & ~n2288;
  assign n8460 = ~n2289 & n8459;
  assign n8461 = ~n2647 & n8460;
  assign n8462 = pi21 & ~n2290;
  assign n8463 = ~n8461 & ~n8462;
  assign n8464 = pi53 & ~n8463;
  assign n8465 = ~pi53 & ~n8462;
  assign n8466 = ~n8461 & n8465;
  assign n8467 = ~pi55 & ~n8456;
  assign n8468 = ~n8455 & n8467;
  assign n8469 = ~n8466 & ~n8468;
  assign n8470 = ~n8464 & n8469;
  assign n8471 = ~n8458 & n8470;
  assign n8472 = ~n8464 & ~n8466;
  assign n8473 = ~n8458 & ~n8468;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = ~n8471 & ~n8474;
  assign n8476 = pi22 & ~n2023;
  assign n8477 = ~n2024 & n8476;
  assign n8478 = ~n2079 & n8477;
  assign n8479 = pi23 & ~n2025;
  assign n8480 = ~n8478 & ~n8479;
  assign n8481 = pi51 & ~n8480;
  assign n8482 = ~pi51 & ~n8479;
  assign n8483 = ~n8478 & n8482;
  assign n8484 = ~n8481 & ~n8483;
  assign n8485 = ~n8475 & n8484;
  assign n8486 = ~n8471 & ~n8484;
  assign n8487 = ~n8474 & n8486;
  assign n8488 = ~n8485 & ~n8487;
  assign n8489 = ~n8118 & ~n8449;
  assign n8490 = ~n8450 & n8489;
  assign n8491 = ~n8488 & ~n8490;
  assign n8492 = ~n8452 & n8491;
  assign n8493 = ~n8135 & ~n8149;
  assign n8494 = ~n8147 & ~n8493;
  assign n8495 = ~n8492 & n8494;
  assign n8496 = ~n8452 & ~n8490;
  assign n8497 = n8488 & ~n8496;
  assign n8498 = ~n8005 & n8204;
  assign n8499 = ~n8006 & n8498;
  assign n8500 = ~n8195 & n8499;
  assign n8501 = n8007 & ~n8194;
  assign n8502 = n8206 & n8501;
  assign n8503 = ~n8233 & ~n8502;
  assign n8504 = ~n8500 & n8503;
  assign n8505 = ~n7949 & ~n8194;
  assign n8506 = n8206 & n8505;
  assign n8507 = ~n8209 & n8506;
  assign n8508 = ~n7949 & n8204;
  assign n8509 = ~n8195 & n8508;
  assign n8510 = ~n8209 & n8509;
  assign n8511 = ~n8507 & ~n8510;
  assign n8512 = n8504 & n8511;
  assign n8513 = ~n8497 & ~n8512;
  assign n8514 = n8495 & n8513;
  assign n8515 = ~n8492 & ~n8497;
  assign n8516 = ~n8494 & ~n8512;
  assign n8517 = ~n8515 & n8516;
  assign n8518 = ~n8492 & n8512;
  assign n8519 = ~n8494 & ~n8497;
  assign n8520 = n8518 & n8519;
  assign n8521 = ~n8517 & ~n8520;
  assign n8522 = ~n8514 & n8521;
  assign n8523 = ~n8182 & ~n8191;
  assign n8524 = ~n8189 & n8523;
  assign n8525 = ~n8180 & n8524;
  assign n8526 = ~n8205 & ~n8525;
  assign n8527 = pi24 & ~n1607;
  assign n8528 = ~n1608 & n8527;
  assign n8529 = ~n1782 & n8528;
  assign n8530 = pi25 & ~n1609;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = pi49 & ~n8531;
  assign n8533 = ~pi49 & ~n8530;
  assign n8534 = ~n8529 & n8533;
  assign n8535 = ~n8532 & ~n8534;
  assign n8536 = pi26 & ~n1212;
  assign n8537 = ~n1213 & n8536;
  assign n8538 = ~n1425 & n8537;
  assign n8539 = pi27 & ~n1214;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = pi47 & ~n8540;
  assign n8542 = ~pi47 & ~n8539;
  assign n8543 = ~n8538 & n8542;
  assign n8544 = ~n8541 & ~n8543;
  assign n8545 = ~n8535 & n8544;
  assign n8546 = n8535 & ~n8544;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = pi28 & ~n1006;
  assign n8549 = ~n1007 & n8548;
  assign n8550 = ~n1068 & n8549;
  assign n8551 = pi29 & ~n1008;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = pi45 & ~n8552;
  assign n8554 = ~pi45 & ~n8551;
  assign n8555 = ~n8550 & n8554;
  assign n8556 = ~n8553 & ~n8555;
  assign n8557 = ~n8547 & n8556;
  assign n8558 = ~n8545 & ~n8556;
  assign n8559 = ~n8546 & n8558;
  assign n8560 = ~n8557 & ~n8559;
  assign n8561 = ~n8526 & n8560;
  assign n8562 = n8526 & ~n8560;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = pi30 & ~n683;
  assign n8565 = ~n684 & n8564;
  assign n8566 = ~n1231 & n8565;
  assign n8567 = pi31 & ~n685;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = pi43 & ~n8568;
  assign n8570 = ~pi43 & ~n8567;
  assign n8571 = ~n8566 & n8570;
  assign n8572 = ~n8569 & ~n8571;
  assign n8573 = ~n8226 & n8572;
  assign n8574 = ~n8563 & n8573;
  assign n8575 = n8226 & ~n8572;
  assign n8576 = ~n8563 & n8575;
  assign n8577 = ~n8574 & ~n8576;
  assign n8578 = ~n8226 & ~n8572;
  assign n8579 = ~n8561 & n8578;
  assign n8580 = ~n8562 & n8579;
  assign n8581 = ~n8224 & ~n8571;
  assign n8582 = ~n8222 & n8581;
  assign n8583 = ~n8216 & ~n8569;
  assign n8584 = n8582 & n8583;
  assign n8585 = ~n8561 & n8584;
  assign n8586 = ~n8562 & n8585;
  assign n8587 = ~n8580 & ~n8586;
  assign n8588 = n8577 & n8587;
  assign n8589 = ~n8147 & ~n8507;
  assign n8590 = ~n8510 & n8589;
  assign n8591 = ~n8493 & n8504;
  assign n8592 = n8590 & n8591;
  assign n8593 = ~n8515 & n8592;
  assign n8594 = ~n8264 & ~n8593;
  assign n8595 = ~n8588 & n8594;
  assign n8596 = n8522 & n8595;
  assign n8597 = ~n8517 & ~n8593;
  assign n8598 = ~n8514 & ~n8520;
  assign n8599 = n8597 & n8598;
  assign n8600 = n8264 & ~n8588;
  assign n8601 = ~n8599 & n8600;
  assign n8602 = ~n8596 & ~n8601;
  assign n8603 = ~n8576 & ~n8580;
  assign n8604 = ~n8586 & n8603;
  assign n8605 = n8264 & ~n8574;
  assign n8606 = ~n8593 & n8605;
  assign n8607 = n8604 & n8606;
  assign n8608 = n8522 & n8607;
  assign n8609 = ~n8264 & ~n8574;
  assign n8610 = n8604 & n8609;
  assign n8611 = ~n8599 & n8610;
  assign n8612 = ~n8608 & ~n8611;
  assign n8613 = n8602 & n8612;
  assign n8614 = ~n8440 & ~n8613;
  assign n8615 = ~n8439 & n8614;
  assign n8616 = ~n8439 & ~n8440;
  assign n8617 = n8613 & ~n8616;
  assign n8618 = ~n8615 & ~n8617;
  assign n8619 = ~n8271 & ~n8328;
  assign n8620 = ~n8326 & ~n8619;
  assign n8621 = n7847 & ~n8314;
  assign n8622 = ~n8315 & n8621;
  assign n8623 = ~n8324 & ~n8622;
  assign n8624 = ~n8620 & ~n8623;
  assign n8625 = ~n8326 & n8623;
  assign n8626 = ~n8619 & n8625;
  assign n8627 = ~n8624 & ~n8626;
  assign n8628 = ~n8618 & n8627;
  assign n8629 = n8618 & ~n8627;
  assign n8630 = ~n8628 & ~n8629;
  assign n8631 = n8370 & n8630;
  assign n8632 = ~n8370 & ~n8630;
  assign n8633 = ~n8631 & ~n8632;
  assign n8634 = ~n8368 & n8633;
  assign n8635 = ~n8346 & ~n8633;
  assign n8636 = ~n8367 & n8635;
  assign po41 = ~n8634 & ~n8636;
  assign n8638 = ~n6765 & n7130;
  assign n8639 = ~n6766 & n8638;
  assign n8640 = ~n6784 & n8639;
  assign n8641 = n5166 & n6125;
  assign n8642 = n7180 & n8641;
  assign n8643 = ~n5479 & ~n6101;
  assign n8644 = n6123 & n8643;
  assign n8645 = n7500 & n8644;
  assign n8646 = n8642 & n8645;
  assign n8647 = ~n4864 & n8646;
  assign n8648 = ~n4863 & n8647;
  assign n8649 = ~n8640 & ~n8648;
  assign n8650 = n8348 & n8633;
  assign n8651 = n7490 & n8078;
  assign n8652 = n8650 & n8651;
  assign n8653 = ~n8649 & n8652;
  assign n8654 = n7489 & ~n7788;
  assign n8655 = n8085 & n8654;
  assign n8656 = ~n8093 & ~n8346;
  assign n8657 = ~n8655 & n8656;
  assign n8658 = ~n8347 & ~n8657;
  assign n8659 = ~n7129 & ~n7488;
  assign n8660 = ~n7489 & ~n7788;
  assign n8661 = n8084 & n8660;
  assign n8662 = n8659 & n8661;
  assign n8663 = ~n8050 & ~n8346;
  assign n8664 = ~n8347 & n8663;
  assign n8665 = ~n7178 & n8664;
  assign n8666 = n8662 & n8665;
  assign n8667 = ~n8658 & ~n8666;
  assign n8668 = ~n8631 & ~n8667;
  assign n8669 = ~n8632 & ~n8668;
  assign n8670 = ~n8653 & n8669;
  assign n8671 = n8618 & ~n8626;
  assign n8672 = ~n8624 & ~n8671;
  assign n8673 = n8314 & ~n8410;
  assign n8674 = ~n8411 & n8673;
  assign n8675 = ~n8430 & ~n8674;
  assign n8676 = ~n8164 & n8675;
  assign n8677 = ~n8420 & n8676;
  assign n8678 = n8437 & n8677;
  assign n8679 = n8613 & n8678;
  assign n8680 = ~n8420 & ~n8674;
  assign n8681 = ~n8421 & n8680;
  assign n8682 = n8613 & n8681;
  assign n8683 = n8421 & ~n8680;
  assign n8684 = ~n8613 & n8683;
  assign n8685 = ~n8682 & ~n8684;
  assign n8686 = ~n8679 & n8685;
  assign n8687 = ~n8438 & ~n8680;
  assign n8688 = ~n8613 & n8687;
  assign n8689 = ~n8438 & n8683;
  assign n8690 = ~n8421 & n8678;
  assign n8691 = ~n8689 & ~n8690;
  assign n8692 = ~n8688 & n8691;
  assign n8693 = n8686 & n8692;
  assign n8694 = ~n8452 & ~n8492;
  assign n8695 = pi17 & ~n3205;
  assign n8696 = ~n3206 & n8695;
  assign n8697 = ~n3463 & n8696;
  assign n8698 = pi18 & ~n3207;
  assign n8699 = ~n8697 & ~n8698;
  assign n8700 = pi57 & ~n8699;
  assign n8701 = ~pi57 & ~n8698;
  assign n8702 = ~n8697 & n8701;
  assign n8703 = ~n8700 & ~n8702;
  assign n8704 = ~n8474 & n8484;
  assign n8705 = ~n8471 & ~n8704;
  assign n8706 = n8703 & ~n8705;
  assign n8707 = pi19 & ~n2876;
  assign n8708 = ~n2877 & n8707;
  assign n8709 = ~n2960 & n8708;
  assign n8710 = pi20 & ~n2878;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = pi55 & ~n8711;
  assign n8713 = pi21 & ~n2288;
  assign n8714 = ~n2289 & n8713;
  assign n8715 = ~n2647 & n8714;
  assign n8716 = pi22 & ~n2290;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = pi53 & ~n8717;
  assign n8719 = ~pi53 & ~n8716;
  assign n8720 = ~n8715 & n8719;
  assign n8721 = ~pi55 & ~n8710;
  assign n8722 = ~n8709 & n8721;
  assign n8723 = ~n8720 & ~n8722;
  assign n8724 = ~n8718 & n8723;
  assign n8725 = ~n8712 & n8724;
  assign n8726 = ~n8718 & ~n8720;
  assign n8727 = ~n8712 & ~n8722;
  assign n8728 = ~n8726 & ~n8727;
  assign n8729 = ~n8725 & ~n8728;
  assign n8730 = pi23 & ~n2023;
  assign n8731 = ~n2024 & n8730;
  assign n8732 = ~n2079 & n8731;
  assign n8733 = pi24 & ~n2025;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = pi51 & ~n8734;
  assign n8736 = ~pi51 & ~n8733;
  assign n8737 = ~n8732 & n8736;
  assign n8738 = ~n8735 & ~n8737;
  assign n8739 = ~n8729 & n8738;
  assign n8740 = ~n8725 & ~n8738;
  assign n8741 = ~n8728 & n8740;
  assign n8742 = ~n8739 & ~n8741;
  assign n8743 = ~n8471 & ~n8703;
  assign n8744 = ~n8704 & n8743;
  assign n8745 = ~n8742 & ~n8744;
  assign n8746 = ~n8706 & n8745;
  assign n8747 = ~n8706 & ~n8744;
  assign n8748 = n8742 & ~n8747;
  assign n8749 = ~n8746 & ~n8748;
  assign n8750 = ~n8694 & n8749;
  assign n8751 = n8694 & ~n8749;
  assign n8752 = ~n8750 & ~n8751;
  assign n8753 = n8226 & ~n8562;
  assign n8754 = ~n8561 & ~n8753;
  assign n8755 = ~n8752 & n8754;
  assign n8756 = ~n8750 & ~n8754;
  assign n8757 = ~n8751 & n8756;
  assign n8758 = ~n8755 & ~n8757;
  assign n8759 = ~n8534 & ~n8543;
  assign n8760 = ~n8541 & n8759;
  assign n8761 = ~n8532 & n8760;
  assign n8762 = ~n8557 & ~n8761;
  assign n8763 = pi25 & ~n1607;
  assign n8764 = ~n1608 & n8763;
  assign n8765 = ~n1782 & n8764;
  assign n8766 = pi26 & ~n1609;
  assign n8767 = ~n8765 & ~n8766;
  assign n8768 = pi49 & ~n8767;
  assign n8769 = ~pi49 & ~n8766;
  assign n8770 = ~n8765 & n8769;
  assign n8771 = ~n8768 & ~n8770;
  assign n8772 = pi27 & ~n1212;
  assign n8773 = ~n1213 & n8772;
  assign n8774 = ~n1425 & n8773;
  assign n8775 = pi28 & ~n1214;
  assign n8776 = ~n8774 & ~n8775;
  assign n8777 = pi47 & ~n8776;
  assign n8778 = ~pi47 & ~n8775;
  assign n8779 = ~n8774 & n8778;
  assign n8780 = ~n8777 & ~n8779;
  assign n8781 = ~n8771 & n8780;
  assign n8782 = n8771 & ~n8780;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = pi29 & ~n1006;
  assign n8785 = ~n1007 & n8784;
  assign n8786 = ~n1068 & n8785;
  assign n8787 = pi30 & ~n1008;
  assign n8788 = ~n8786 & ~n8787;
  assign n8789 = pi45 & ~n8788;
  assign n8790 = ~pi45 & ~n8787;
  assign n8791 = ~n8786 & n8790;
  assign n8792 = ~n8789 & ~n8791;
  assign n8793 = ~n8783 & n8792;
  assign n8794 = ~n8781 & ~n8792;
  assign n8795 = ~n8782 & n8794;
  assign n8796 = ~n8793 & ~n8795;
  assign n8797 = ~n8762 & n8796;
  assign n8798 = n8762 & ~n8796;
  assign n8799 = ~n8797 & ~n8798;
  assign n8800 = n8572 & ~n8799;
  assign n8801 = ~n8572 & ~n8797;
  assign n8802 = ~n8798 & n8801;
  assign n8803 = ~n8800 & ~n8802;
  assign n8804 = n685 & n1231;
  assign n8805 = pi31 & pi43;
  assign n8806 = ~n8804 & n8805;
  assign n8807 = pi31 & ~n8804;
  assign n8808 = ~pi43 & ~n8807;
  assign n8809 = ~n8806 & ~n8808;
  assign n8810 = ~n8803 & ~n8809;
  assign n8811 = ~n8800 & n8809;
  assign n8812 = ~n8802 & n8811;
  assign n8813 = ~n8810 & ~n8812;
  assign n8814 = n8226 & ~n8563;
  assign n8815 = ~n8226 & ~n8561;
  assign n8816 = ~n8562 & n8815;
  assign n8817 = ~n8814 & ~n8816;
  assign n8818 = ~n8572 & ~n8817;
  assign n8819 = ~n8813 & n8818;
  assign n8820 = ~n8758 & n8819;
  assign n8821 = ~n8755 & ~n8818;
  assign n8822 = ~n8757 & ~n8813;
  assign n8823 = n8821 & n8822;
  assign n8824 = ~n8820 & ~n8823;
  assign n8825 = n8813 & ~n8818;
  assign n8826 = ~n8758 & n8825;
  assign n8827 = ~n8810 & n8818;
  assign n8828 = ~n8812 & n8827;
  assign n8829 = n8758 & n8828;
  assign n8830 = ~n8826 & ~n8829;
  assign n8831 = n8824 & n8830;
  assign n8832 = ~n8264 & ~n8599;
  assign n8833 = n8264 & ~n8593;
  assign n8834 = n8522 & n8833;
  assign n8835 = n8588 & ~n8834;
  assign n8836 = ~n8832 & ~n8835;
  assign n8837 = n8494 & ~n8515;
  assign n8838 = n8512 & ~n8837;
  assign n8839 = ~n8494 & n8515;
  assign n8840 = ~n8383 & ~n8392;
  assign n8841 = ~n8390 & n8840;
  assign n8842 = ~n8381 & n8841;
  assign n8843 = ~n8406 & ~n8842;
  assign n8844 = pi11 & ~n5091;
  assign n8845 = ~n5092 & n8844;
  assign n8846 = ~n5178 & n8845;
  assign n8847 = pi12 & ~n5093;
  assign n8848 = ~n8846 & ~n8847;
  assign n8849 = pi63 & ~n8848;
  assign n8850 = ~pi63 & ~n8847;
  assign n8851 = ~n8846 & n8850;
  assign n8852 = ~n8849 & ~n8851;
  assign n8853 = pi13 & ~n4513;
  assign n8854 = ~n4514 & n8853;
  assign n8855 = ~n4577 & n8854;
  assign n8856 = pi14 & ~n4515;
  assign n8857 = ~n8855 & ~n8856;
  assign n8858 = pi61 & ~n8857;
  assign n8859 = ~pi61 & ~n8856;
  assign n8860 = ~n8855 & n8859;
  assign n8861 = ~n8858 & ~n8860;
  assign n8862 = ~n8852 & n8861;
  assign n8863 = n8852 & ~n8861;
  assign n8864 = ~n8862 & ~n8863;
  assign n8865 = pi15 & ~n3959;
  assign n8866 = ~n3960 & n8865;
  assign n8867 = ~n4233 & n8866;
  assign n8868 = pi16 & ~n3961;
  assign n8869 = ~n8867 & ~n8868;
  assign n8870 = pi59 & ~n8869;
  assign n8871 = ~pi59 & ~n8868;
  assign n8872 = ~n8867 & n8871;
  assign n8873 = ~n8870 & ~n8872;
  assign n8874 = ~n8864 & n8873;
  assign n8875 = ~n8862 & ~n8873;
  assign n8876 = ~n8863 & n8875;
  assign n8877 = ~n8874 & ~n8876;
  assign n8878 = ~n8843 & n8877;
  assign n8879 = n8843 & ~n8877;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = n8410 & ~n8880;
  assign n8882 = ~n8410 & ~n8878;
  assign n8883 = ~n8879 & n8882;
  assign n8884 = ~n8881 & ~n8883;
  assign n8885 = ~n8839 & n8884;
  assign n8886 = ~n8838 & n8885;
  assign n8887 = ~n8838 & ~n8839;
  assign n8888 = ~n8884 & ~n8887;
  assign n8889 = ~n8886 & ~n8888;
  assign n8890 = ~n8836 & n8889;
  assign n8891 = n8836 & ~n8889;
  assign n8892 = ~n8890 & ~n8891;
  assign n8893 = ~n8831 & n8892;
  assign n8894 = n8831 & ~n8892;
  assign n8895 = ~n8893 & ~n8894;
  assign n8896 = ~n8693 & n8895;
  assign n8897 = n8693 & ~n8895;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = n8672 & n8898;
  assign n8900 = ~n8672 & ~n8898;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = ~n8670 & n8901;
  assign n8903 = ~n8632 & ~n8901;
  assign n8904 = ~n8668 & n8903;
  assign n8905 = ~n8653 & n8904;
  assign po42 = ~n8902 & ~n8905;
  assign n8907 = ~n7161 & ~n7165;
  assign n8908 = ~n7159 & n8907;
  assign n8909 = ~n7152 & n8908;
  assign n8910 = n8361 & n8650;
  assign n8911 = n5161 & ~n5479;
  assign n8912 = n6125 & n8911;
  assign n8913 = n7502 & n8912;
  assign n8914 = n7500 & n8913;
  assign n8915 = n8910 & n8914;
  assign n8916 = ~n8909 & n8915;
  assign n8917 = ~n6420 & n7501;
  assign n8918 = n5159 & ~n5479;
  assign n8919 = n6123 & n6125;
  assign n8920 = n8918 & n8919;
  assign n8921 = n8917 & n8920;
  assign n8922 = ~n6766 & ~n8921;
  assign n8923 = ~n6781 & n8922;
  assign n8924 = ~n6765 & n7503;
  assign n8925 = n8078 & n8650;
  assign n8926 = n8924 & n8925;
  assign n8927 = ~n8923 & n8926;
  assign n8928 = ~n8347 & ~n8631;
  assign n8929 = ~n8632 & n8928;
  assign n8930 = ~n8657 & n8929;
  assign n8931 = n8084 & n8663;
  assign n8932 = n7128 & ~n7488;
  assign n8933 = n8660 & n8932;
  assign n8934 = n8931 & n8933;
  assign n8935 = n8929 & n8934;
  assign n8936 = ~n8632 & ~n8935;
  assign n8937 = ~n8930 & n8936;
  assign n8938 = ~n8927 & n8937;
  assign n8939 = ~n8916 & n8938;
  assign n8940 = ~n8899 & ~n8939;
  assign n8941 = ~n8900 & ~n8940;
  assign n8942 = ~n8755 & n8818;
  assign n8943 = ~n8757 & n8942;
  assign n8944 = ~n8758 & ~n8818;
  assign n8945 = n8813 & ~n8944;
  assign n8946 = ~n8943 & ~n8945;
  assign n8947 = ~n8751 & ~n8754;
  assign n8948 = ~n8851 & ~n8860;
  assign n8949 = ~n8858 & n8948;
  assign n8950 = ~n8849 & n8949;
  assign n8951 = ~n8874 & ~n8950;
  assign n8952 = pi12 & ~n5091;
  assign n8953 = ~n5092 & n8952;
  assign n8954 = ~n5178 & n8953;
  assign n8955 = pi13 & ~n5093;
  assign n8956 = ~n8954 & ~n8955;
  assign n8957 = pi63 & ~n8956;
  assign n8958 = ~pi63 & ~n8955;
  assign n8959 = ~n8954 & n8958;
  assign n8960 = ~n8957 & ~n8959;
  assign n8961 = pi14 & ~n4513;
  assign n8962 = ~n4514 & n8961;
  assign n8963 = ~n4577 & n8962;
  assign n8964 = pi15 & ~n4515;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = pi61 & ~n8965;
  assign n8967 = ~pi61 & ~n8964;
  assign n8968 = ~n8963 & n8967;
  assign n8969 = ~n8966 & ~n8968;
  assign n8970 = ~n8960 & n8969;
  assign n8971 = n8960 & ~n8969;
  assign n8972 = ~n8970 & ~n8971;
  assign n8973 = pi16 & ~n3959;
  assign n8974 = ~n3960 & n8973;
  assign n8975 = ~n4233 & n8974;
  assign n8976 = pi17 & ~n3961;
  assign n8977 = ~n8975 & ~n8976;
  assign n8978 = pi59 & ~n8977;
  assign n8979 = ~pi59 & ~n8976;
  assign n8980 = ~n8975 & n8979;
  assign n8981 = ~n8978 & ~n8980;
  assign n8982 = ~n8972 & n8981;
  assign n8983 = ~n8970 & ~n8981;
  assign n8984 = ~n8971 & n8983;
  assign n8985 = ~n8982 & ~n8984;
  assign n8986 = ~n8951 & n8985;
  assign n8987 = n8951 & ~n8985;
  assign n8988 = ~n8986 & ~n8987;
  assign n8989 = n8878 & ~n8988;
  assign n8990 = ~n8878 & ~n8986;
  assign n8991 = ~n8987 & n8990;
  assign n8992 = ~n8989 & ~n8991;
  assign n8993 = ~n8750 & n8992;
  assign n8994 = ~n8947 & n8993;
  assign n8995 = ~n8750 & ~n8947;
  assign n8996 = ~n8992 & ~n8995;
  assign n8997 = ~n8994 & ~n8996;
  assign n8998 = ~n8946 & n8997;
  assign n8999 = ~n8943 & ~n8997;
  assign n9000 = ~n8945 & n8999;
  assign n9001 = ~n8998 & ~n9000;
  assign n9002 = ~n8706 & ~n8746;
  assign n9003 = pi18 & ~n3205;
  assign n9004 = ~n3206 & n9003;
  assign n9005 = ~n3463 & n9004;
  assign n9006 = pi19 & ~n3207;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = pi57 & ~n9007;
  assign n9009 = ~pi57 & ~n9006;
  assign n9010 = ~n9005 & n9009;
  assign n9011 = ~n9008 & ~n9010;
  assign n9012 = ~n8728 & n8738;
  assign n9013 = ~n8725 & ~n9012;
  assign n9014 = n9011 & ~n9013;
  assign n9015 = pi20 & ~n2876;
  assign n9016 = ~n2877 & n9015;
  assign n9017 = ~n2960 & n9016;
  assign n9018 = pi21 & ~n2878;
  assign n9019 = ~n9017 & ~n9018;
  assign n9020 = pi55 & ~n9019;
  assign n9021 = pi22 & ~n2288;
  assign n9022 = ~n2289 & n9021;
  assign n9023 = ~n2647 & n9022;
  assign n9024 = pi23 & ~n2290;
  assign n9025 = ~n9023 & ~n9024;
  assign n9026 = pi53 & ~n9025;
  assign n9027 = ~pi53 & ~n9024;
  assign n9028 = ~n9023 & n9027;
  assign n9029 = ~pi55 & ~n9018;
  assign n9030 = ~n9017 & n9029;
  assign n9031 = ~n9028 & ~n9030;
  assign n9032 = ~n9026 & n9031;
  assign n9033 = ~n9020 & n9032;
  assign n9034 = ~n9026 & ~n9028;
  assign n9035 = ~n9020 & ~n9030;
  assign n9036 = ~n9034 & ~n9035;
  assign n9037 = ~n9033 & ~n9036;
  assign n9038 = pi24 & ~n2023;
  assign n9039 = ~n2024 & n9038;
  assign n9040 = ~n2079 & n9039;
  assign n9041 = pi25 & ~n2025;
  assign n9042 = ~n9040 & ~n9041;
  assign n9043 = pi51 & ~n9042;
  assign n9044 = ~pi51 & ~n9041;
  assign n9045 = ~n9040 & n9044;
  assign n9046 = ~n9043 & ~n9045;
  assign n9047 = ~n9037 & n9046;
  assign n9048 = ~n9033 & ~n9046;
  assign n9049 = ~n9036 & n9048;
  assign n9050 = ~n9047 & ~n9049;
  assign n9051 = ~n8725 & ~n9011;
  assign n9052 = ~n9012 & n9051;
  assign n9053 = ~n9050 & ~n9052;
  assign n9054 = ~n9014 & n9053;
  assign n9055 = ~n9014 & ~n9052;
  assign n9056 = n9050 & ~n9055;
  assign n9057 = ~n9054 & ~n9056;
  assign n9058 = ~n9002 & n9057;
  assign n9059 = n9002 & ~n9057;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = n8572 & ~n8798;
  assign n9062 = ~n8797 & ~n9061;
  assign n9063 = ~n9060 & n9062;
  assign n9064 = ~n9058 & ~n9062;
  assign n9065 = ~n9059 & n9064;
  assign n9066 = ~n9063 & ~n9065;
  assign n9067 = ~n8770 & ~n8779;
  assign n9068 = ~n8777 & n9067;
  assign n9069 = ~n8768 & n9068;
  assign n9070 = ~n8793 & ~n9069;
  assign n9071 = pi26 & ~n1607;
  assign n9072 = ~n1608 & n9071;
  assign n9073 = ~n1782 & n9072;
  assign n9074 = pi27 & ~n1609;
  assign n9075 = ~n9073 & ~n9074;
  assign n9076 = pi49 & ~n9075;
  assign n9077 = ~pi49 & ~n9074;
  assign n9078 = ~n9073 & n9077;
  assign n9079 = ~n9076 & ~n9078;
  assign n9080 = pi28 & ~n1212;
  assign n9081 = ~n1213 & n9080;
  assign n9082 = ~n1425 & n9081;
  assign n9083 = pi29 & ~n1214;
  assign n9084 = ~n9082 & ~n9083;
  assign n9085 = pi47 & ~n9084;
  assign n9086 = ~pi47 & ~n9083;
  assign n9087 = ~n9082 & n9086;
  assign n9088 = ~n9085 & ~n9087;
  assign n9089 = n9079 & ~n9088;
  assign n9090 = pi30 & ~n1006;
  assign n9091 = ~n1007 & n9090;
  assign n9092 = ~n1068 & n9091;
  assign n9093 = pi31 & ~n1008;
  assign n9094 = ~n9092 & ~n9093;
  assign n9095 = pi45 & ~n9094;
  assign n9096 = ~pi45 & ~n9093;
  assign n9097 = ~n9092 & n9096;
  assign n9098 = ~n9095 & ~n9097;
  assign n9099 = ~n9079 & n9088;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = ~n9089 & n9100;
  assign n9102 = ~n9089 & ~n9099;
  assign n9103 = n9098 & ~n9102;
  assign n9104 = ~n9101 & ~n9103;
  assign n9105 = ~n9070 & n9104;
  assign n9106 = n9070 & ~n9104;
  assign n9107 = ~n9105 & ~n9106;
  assign n9108 = ~n8809 & ~n9107;
  assign n9109 = ~n8803 & n9108;
  assign n9110 = ~n9066 & n9109;
  assign n9111 = ~n8810 & ~n9107;
  assign n9112 = ~n9063 & n9111;
  assign n9113 = ~n9065 & n9112;
  assign n9114 = ~n9110 & ~n9113;
  assign n9115 = ~n8810 & n9107;
  assign n9116 = ~n9066 & n9115;
  assign n9117 = ~n8809 & ~n9105;
  assign n9118 = ~n9106 & n9117;
  assign n9119 = ~n8803 & n9118;
  assign n9120 = ~n9063 & n9119;
  assign n9121 = ~n9065 & n9120;
  assign n9122 = ~n9116 & ~n9121;
  assign n9123 = n9114 & n9122;
  assign n9124 = ~n9001 & n9123;
  assign n9125 = ~n9000 & ~n9123;
  assign n9126 = ~n8998 & n9125;
  assign n9127 = ~n9124 & ~n9126;
  assign n9128 = n8410 & ~n8878;
  assign n9129 = ~n8879 & n9128;
  assign n9130 = ~n8888 & ~n9129;
  assign n9131 = ~n8890 & n9130;
  assign n9132 = ~n8892 & n9131;
  assign n9133 = n8889 & ~n9130;
  assign n9134 = ~n8836 & n9133;
  assign n9135 = ~n9132 & ~n9134;
  assign n9136 = ~n8890 & ~n9130;
  assign n9137 = ~n8831 & ~n8891;
  assign n9138 = n9136 & n9137;
  assign n9139 = ~n8820 & n9130;
  assign n9140 = ~n8823 & ~n8826;
  assign n9141 = ~n8829 & n9140;
  assign n9142 = n9139 & n9141;
  assign n9143 = ~n8890 & n9142;
  assign n9144 = ~n9138 & ~n9143;
  assign n9145 = n9135 & n9144;
  assign n9146 = ~n9127 & ~n9145;
  assign n9147 = ~n9126 & ~n9138;
  assign n9148 = ~n9143 & n9147;
  assign n9149 = ~n9124 & n9135;
  assign n9150 = n9148 & n9149;
  assign n9151 = ~n9146 & ~n9150;
  assign n9152 = ~n8439 & n8680;
  assign n9153 = ~n8615 & n9152;
  assign n9154 = ~n8897 & ~n9153;
  assign n9155 = ~n9151 & n9154;
  assign n9156 = n9151 & ~n9154;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = ~n8941 & n9157;
  assign n9159 = ~n8900 & ~n9157;
  assign n9160 = ~n8940 & n9159;
  assign po43 = ~n9158 & ~n9160;
  assign n9162 = ~n3454 & n5168;
  assign n9163 = n5485 & ~n9162;
  assign n9164 = n6125 & n7180;
  assign n9165 = n8644 & n9164;
  assign n9166 = n7500 & n9165;
  assign n9167 = ~n9163 & n9166;
  assign n9168 = n3708 & ~n5479;
  assign n9169 = n4271 & n7160;
  assign n9170 = n9168 & n9169;
  assign n9171 = n2716 & ~n4549;
  assign n9172 = n4563 & n9171;
  assign n9173 = n9164 & n9172;
  assign n9174 = n5161 & ~n6101;
  assign n9175 = n6123 & n9174;
  assign n9176 = n7500 & n9175;
  assign n9177 = n9173 & n9176;
  assign n9178 = n9170 & n9177;
  assign n9179 = ~n2270 & n9178;
  assign n9180 = ~n7179 & ~n7489;
  assign n9181 = ~n7182 & n9180;
  assign n9182 = ~n9179 & n9181;
  assign n9183 = ~n9167 & n9182;
  assign n9184 = n8633 & n9157;
  assign n9185 = ~n8049 & n8901;
  assign n9186 = n8348 & n9185;
  assign n9187 = ~n7488 & ~n8050;
  assign n9188 = n7790 & n9187;
  assign n9189 = n9186 & n9188;
  assign n9190 = n9184 & n9189;
  assign n9191 = ~n9183 & n9190;
  assign n9192 = n8346 & n8901;
  assign n9193 = n8633 & n9192;
  assign n9194 = n8632 & n8901;
  assign n9195 = ~n8900 & ~n9155;
  assign n9196 = ~n9194 & n9195;
  assign n9197 = ~n9193 & n9196;
  assign n9198 = ~n9156 & ~n9197;
  assign n9199 = ~n8092 & n9186;
  assign n9200 = n9184 & n9199;
  assign n9201 = ~n9198 & ~n9200;
  assign n9202 = ~n9191 & n9201;
  assign n9203 = ~n8890 & ~n8893;
  assign n9204 = ~n9130 & ~n9203;
  assign n9205 = ~n9127 & n9145;
  assign n9206 = ~n9204 & ~n9205;
  assign n9207 = n8878 & ~n8986;
  assign n9208 = ~n8987 & n9207;
  assign n9209 = ~n8996 & ~n9208;
  assign n9210 = ~n8943 & n9209;
  assign n9211 = ~n8945 & n9210;
  assign n9212 = ~n9123 & n9211;
  assign n9213 = ~n8997 & n9210;
  assign n9214 = ~n8945 & n9213;
  assign n9215 = ~n8997 & n9209;
  assign n9216 = ~n9123 & n9215;
  assign n9217 = ~n9214 & ~n9216;
  assign n9218 = ~n9212 & n9217;
  assign n9219 = n9122 & ~n9209;
  assign n9220 = n9114 & n9219;
  assign n9221 = ~n8946 & n9220;
  assign n9222 = n8997 & ~n9209;
  assign n9223 = ~n8946 & n9222;
  assign n9224 = n9123 & n9222;
  assign n9225 = ~n9223 & ~n9224;
  assign n9226 = ~n9221 & n9225;
  assign n9227 = n9218 & n9226;
  assign n9228 = n8810 & ~n9063;
  assign n9229 = ~n9065 & n9228;
  assign n9230 = ~n8810 & ~n9066;
  assign n9231 = ~n9107 & ~n9230;
  assign n9232 = ~n9229 & ~n9231;
  assign n9233 = ~n9059 & ~n9062;
  assign n9234 = ~n8959 & ~n8968;
  assign n9235 = ~n8966 & n9234;
  assign n9236 = ~n8957 & n9235;
  assign n9237 = ~n8982 & ~n9236;
  assign n9238 = pi13 & ~n5091;
  assign n9239 = ~n5092 & n9238;
  assign n9240 = ~n5178 & n9239;
  assign n9241 = pi14 & ~n5093;
  assign n9242 = ~n9240 & ~n9241;
  assign n9243 = pi63 & ~n9242;
  assign n9244 = ~pi63 & ~n9241;
  assign n9245 = ~n9240 & n9244;
  assign n9246 = ~n9243 & ~n9245;
  assign n9247 = pi15 & ~n4513;
  assign n9248 = ~n4514 & n9247;
  assign n9249 = ~n4577 & n9248;
  assign n9250 = pi16 & ~n4515;
  assign n9251 = ~n9249 & ~n9250;
  assign n9252 = pi61 & ~n9251;
  assign n9253 = ~pi61 & ~n9250;
  assign n9254 = ~n9249 & n9253;
  assign n9255 = ~n9252 & ~n9254;
  assign n9256 = ~n9246 & n9255;
  assign n9257 = n9246 & ~n9255;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = pi17 & ~n3959;
  assign n9260 = ~n3960 & n9259;
  assign n9261 = ~n4233 & n9260;
  assign n9262 = pi18 & ~n3961;
  assign n9263 = ~n9261 & ~n9262;
  assign n9264 = pi59 & ~n9263;
  assign n9265 = ~pi59 & ~n9262;
  assign n9266 = ~n9261 & n9265;
  assign n9267 = ~n9264 & ~n9266;
  assign n9268 = ~n9258 & n9267;
  assign n9269 = ~n9256 & ~n9267;
  assign n9270 = ~n9257 & n9269;
  assign n9271 = ~n9268 & ~n9270;
  assign n9272 = n9237 & ~n9271;
  assign n9273 = ~n9237 & n9271;
  assign n9274 = n8986 & ~n9273;
  assign n9275 = ~n9272 & n9274;
  assign n9276 = ~n9272 & ~n9273;
  assign n9277 = ~n8986 & ~n9276;
  assign n9278 = ~n9275 & ~n9277;
  assign n9279 = ~n9058 & ~n9278;
  assign n9280 = ~n9233 & n9279;
  assign n9281 = ~n9058 & ~n9233;
  assign n9282 = n9278 & ~n9281;
  assign n9283 = ~n9280 & ~n9282;
  assign n9284 = ~n9232 & n9283;
  assign n9285 = ~n9229 & ~n9283;
  assign n9286 = ~n9231 & n9285;
  assign n9287 = ~n9014 & ~n9054;
  assign n9288 = ~n9036 & n9046;
  assign n9289 = pi19 & ~n3205;
  assign n9290 = ~n3206 & n9289;
  assign n9291 = ~n3463 & n9290;
  assign n9292 = pi20 & ~n3207;
  assign n9293 = ~n9291 & ~n9292;
  assign n9294 = pi57 & ~n9293;
  assign n9295 = ~pi57 & ~n9292;
  assign n9296 = ~n9291 & n9295;
  assign n9297 = ~n9294 & ~n9296;
  assign n9298 = ~n9033 & ~n9297;
  assign n9299 = ~n9288 & n9298;
  assign n9300 = ~n9033 & ~n9288;
  assign n9301 = n9297 & ~n9300;
  assign n9302 = ~n9299 & ~n9301;
  assign n9303 = pi21 & ~n2876;
  assign n9304 = ~n2877 & n9303;
  assign n9305 = ~n2960 & n9304;
  assign n9306 = pi22 & ~n2878;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = pi55 & ~n9307;
  assign n9309 = pi23 & ~n2288;
  assign n9310 = ~n2289 & n9309;
  assign n9311 = ~n2647 & n9310;
  assign n9312 = pi24 & ~n2290;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = pi53 & ~n9313;
  assign n9315 = ~pi53 & ~n9312;
  assign n9316 = ~n9311 & n9315;
  assign n9317 = ~pi55 & ~n9306;
  assign n9318 = ~n9305 & n9317;
  assign n9319 = ~n9316 & ~n9318;
  assign n9320 = ~n9314 & n9319;
  assign n9321 = ~n9308 & n9320;
  assign n9322 = ~n9314 & ~n9316;
  assign n9323 = ~n9308 & ~n9318;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = ~n9321 & ~n9324;
  assign n9326 = pi25 & ~n2023;
  assign n9327 = ~n2024 & n9326;
  assign n9328 = ~n2079 & n9327;
  assign n9329 = pi26 & ~n2025;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = pi51 & ~n9330;
  assign n9332 = ~pi51 & ~n9329;
  assign n9333 = ~n9328 & n9332;
  assign n9334 = ~n9331 & ~n9333;
  assign n9335 = ~n9325 & n9334;
  assign n9336 = ~n9321 & ~n9334;
  assign n9337 = ~n9324 & n9336;
  assign n9338 = ~n9335 & ~n9337;
  assign n9339 = ~n9302 & n9338;
  assign n9340 = n9302 & ~n9338;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = ~n9287 & n9341;
  assign n9343 = n9287 & ~n9341;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = n9106 & ~n9344;
  assign n9346 = ~n9106 & ~n9342;
  assign n9347 = ~n9343 & n9346;
  assign n9348 = ~n9345 & ~n9347;
  assign n9349 = ~n9078 & ~n9087;
  assign n9350 = ~n9085 & n9349;
  assign n9351 = ~n9076 & n9350;
  assign n9352 = ~n9103 & ~n9351;
  assign n9353 = pi27 & ~n1607;
  assign n9354 = ~n1608 & n9353;
  assign n9355 = ~n1782 & n9354;
  assign n9356 = pi28 & ~n1609;
  assign n9357 = ~n9355 & ~n9356;
  assign n9358 = pi49 & ~n9357;
  assign n9359 = ~pi49 & ~n9356;
  assign n9360 = ~n9355 & n9359;
  assign n9361 = ~n9358 & ~n9360;
  assign n9362 = pi29 & ~n1212;
  assign n9363 = ~n1213 & n9362;
  assign n9364 = ~n1425 & n9363;
  assign n9365 = pi30 & ~n1214;
  assign n9366 = ~n9364 & ~n9365;
  assign n9367 = pi47 & ~n9366;
  assign n9368 = ~pi47 & ~n9365;
  assign n9369 = ~n9364 & n9368;
  assign n9370 = ~n9367 & ~n9369;
  assign n9371 = ~n9361 & n9370;
  assign n9372 = n9361 & ~n9370;
  assign n9373 = ~n9371 & ~n9372;
  assign n9374 = n1008 & n1068;
  assign n9375 = pi31 & pi45;
  assign n9376 = ~n9374 & n9375;
  assign n9377 = pi31 & ~n9374;
  assign n9378 = ~pi45 & ~n9377;
  assign n9379 = ~n9376 & ~n9378;
  assign n9380 = ~n9373 & ~n9379;
  assign n9381 = ~n9371 & n9379;
  assign n9382 = ~n9372 & n9381;
  assign n9383 = ~n9380 & ~n9382;
  assign n9384 = ~n9352 & n9383;
  assign n9385 = n9352 & ~n9383;
  assign n9386 = ~n9384 & ~n9385;
  assign n9387 = ~n9348 & n9386;
  assign n9388 = ~n9345 & ~n9386;
  assign n9389 = ~n9347 & n9388;
  assign n9390 = ~n9387 & ~n9389;
  assign n9391 = ~n9286 & ~n9390;
  assign n9392 = ~n9284 & n9391;
  assign n9393 = ~n9284 & ~n9286;
  assign n9394 = n9390 & ~n9393;
  assign n9395 = ~n9392 & ~n9394;
  assign n9396 = ~n9227 & n9395;
  assign n9397 = n9227 & ~n9395;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = n9206 & n9398;
  assign n9400 = ~n9206 & ~n9398;
  assign n9401 = ~n9399 & ~n9400;
  assign n9402 = ~n9202 & n9401;
  assign n9403 = ~n9198 & ~n9401;
  assign n9404 = ~n9200 & n9403;
  assign n9405 = ~n9191 & n9404;
  assign po44 = ~n9402 & ~n9405;
  assign n9407 = ~n8632 & ~n9155;
  assign n9408 = ~n9156 & n9407;
  assign n9409 = n8663 & n8928;
  assign n9410 = n7790 & n9185;
  assign n9411 = n9409 & n9410;
  assign n9412 = n9408 & n9411;
  assign n9413 = ~n7802 & n9412;
  assign n9414 = n9201 & ~n9413;
  assign n9415 = ~n9399 & ~n9414;
  assign n9416 = ~n9400 & ~n9415;
  assign n9417 = ~n9000 & n9123;
  assign n9418 = ~n8998 & ~n9417;
  assign n9419 = ~n9209 & ~n9418;
  assign n9420 = n9227 & n9395;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = n9107 & ~n9342;
  assign n9423 = ~n9343 & n9422;
  assign n9424 = ~n9345 & n9386;
  assign n9425 = ~n9347 & n9424;
  assign n9426 = ~n9423 & ~n9425;
  assign n9427 = ~n9105 & ~n9342;
  assign n9428 = ~n9343 & ~n9427;
  assign n9429 = ~n9245 & ~n9254;
  assign n9430 = ~n9252 & n9429;
  assign n9431 = ~n9243 & n9430;
  assign n9432 = ~n9268 & ~n9431;
  assign n9433 = pi14 & ~n5091;
  assign n9434 = ~n5092 & n9433;
  assign n9435 = ~n5178 & n9434;
  assign n9436 = pi15 & ~n5093;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = pi63 & ~n9437;
  assign n9439 = ~pi63 & ~n9436;
  assign n9440 = ~n9435 & n9439;
  assign n9441 = ~n9438 & ~n9440;
  assign n9442 = pi16 & ~n4513;
  assign n9443 = ~n4514 & n9442;
  assign n9444 = ~n4577 & n9443;
  assign n9445 = pi17 & ~n4515;
  assign n9446 = ~n9444 & ~n9445;
  assign n9447 = pi61 & ~n9446;
  assign n9448 = ~pi61 & ~n9445;
  assign n9449 = ~n9444 & n9448;
  assign n9450 = ~n9447 & ~n9449;
  assign n9451 = ~n9441 & n9450;
  assign n9452 = n9441 & ~n9450;
  assign n9453 = ~n9451 & ~n9452;
  assign n9454 = pi18 & ~n3959;
  assign n9455 = ~n3960 & n9454;
  assign n9456 = ~n4233 & n9455;
  assign n9457 = pi19 & ~n3961;
  assign n9458 = ~n9456 & ~n9457;
  assign n9459 = pi59 & ~n9458;
  assign n9460 = ~pi59 & ~n9457;
  assign n9461 = ~n9456 & n9460;
  assign n9462 = ~n9459 & ~n9461;
  assign n9463 = ~n9453 & n9462;
  assign n9464 = ~n9451 & ~n9462;
  assign n9465 = ~n9452 & n9464;
  assign n9466 = ~n9463 & ~n9465;
  assign n9467 = ~n9432 & n9466;
  assign n9468 = n9432 & ~n9466;
  assign n9469 = ~n9467 & ~n9468;
  assign n9470 = n9273 & ~n9469;
  assign n9471 = ~n9273 & ~n9467;
  assign n9472 = ~n9468 & n9471;
  assign n9473 = ~n9470 & ~n9472;
  assign n9474 = ~n9428 & n9473;
  assign n9475 = ~n9343 & ~n9473;
  assign n9476 = ~n9427 & n9475;
  assign n9477 = ~n9474 & ~n9476;
  assign n9478 = n9426 & ~n9477;
  assign n9479 = ~n9426 & n9477;
  assign n9480 = ~n9301 & ~n9340;
  assign n9481 = pi20 & ~n3205;
  assign n9482 = ~n3206 & n9481;
  assign n9483 = ~n3463 & n9482;
  assign n9484 = pi21 & ~n3207;
  assign n9485 = ~n9483 & ~n9484;
  assign n9486 = pi57 & ~n9485;
  assign n9487 = ~pi57 & ~n9484;
  assign n9488 = ~n9483 & n9487;
  assign n9489 = ~n9486 & ~n9488;
  assign n9490 = ~n9324 & n9334;
  assign n9491 = ~n9321 & ~n9490;
  assign n9492 = n9489 & ~n9491;
  assign n9493 = pi22 & ~n2876;
  assign n9494 = ~n2877 & n9493;
  assign n9495 = ~n2960 & n9494;
  assign n9496 = pi23 & ~n2878;
  assign n9497 = ~n9495 & ~n9496;
  assign n9498 = pi55 & ~n9497;
  assign n9499 = pi24 & ~n2288;
  assign n9500 = ~n2289 & n9499;
  assign n9501 = ~n2647 & n9500;
  assign n9502 = pi25 & ~n2290;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = pi53 & ~n9503;
  assign n9505 = ~pi53 & ~n9502;
  assign n9506 = ~n9501 & n9505;
  assign n9507 = ~pi55 & ~n9496;
  assign n9508 = ~n9495 & n9507;
  assign n9509 = ~n9506 & ~n9508;
  assign n9510 = ~n9504 & n9509;
  assign n9511 = ~n9498 & n9510;
  assign n9512 = ~n9504 & ~n9506;
  assign n9513 = ~n9498 & ~n9508;
  assign n9514 = ~n9512 & ~n9513;
  assign n9515 = ~n9511 & ~n9514;
  assign n9516 = pi26 & ~n2023;
  assign n9517 = ~n2024 & n9516;
  assign n9518 = ~n2079 & n9517;
  assign n9519 = pi27 & ~n2025;
  assign n9520 = ~n9518 & ~n9519;
  assign n9521 = pi51 & ~n9520;
  assign n9522 = ~pi51 & ~n9519;
  assign n9523 = ~n9518 & n9522;
  assign n9524 = ~n9521 & ~n9523;
  assign n9525 = ~n9515 & n9524;
  assign n9526 = ~n9511 & ~n9524;
  assign n9527 = ~n9514 & n9526;
  assign n9528 = ~n9525 & ~n9527;
  assign n9529 = ~n9321 & ~n9489;
  assign n9530 = ~n9490 & n9529;
  assign n9531 = ~n9528 & ~n9530;
  assign n9532 = ~n9492 & n9531;
  assign n9533 = ~n9492 & ~n9530;
  assign n9534 = n9528 & ~n9533;
  assign n9535 = ~n9532 & ~n9534;
  assign n9536 = ~n9480 & n9535;
  assign n9537 = n9480 & ~n9535;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = ~n9384 & ~n9538;
  assign n9540 = n9384 & ~n9536;
  assign n9541 = ~n9537 & n9540;
  assign n9542 = ~n9360 & ~n9369;
  assign n9543 = ~n9367 & n9542;
  assign n9544 = ~n9358 & n9543;
  assign n9545 = ~n9380 & ~n9544;
  assign n9546 = pi30 & ~n1212;
  assign n9547 = ~n1213 & n9546;
  assign n9548 = ~n1425 & n9547;
  assign n9549 = pi31 & ~n1214;
  assign n9550 = ~n9548 & ~n9549;
  assign n9551 = pi47 & ~n9550;
  assign n9552 = pi28 & ~n1607;
  assign n9553 = ~n1608 & n9552;
  assign n9554 = ~n1782 & n9553;
  assign n9555 = pi29 & ~n1609;
  assign n9556 = ~n9554 & ~n9555;
  assign n9557 = pi49 & ~n9556;
  assign n9558 = ~pi49 & ~n9555;
  assign n9559 = ~n9554 & n9558;
  assign n9560 = ~pi47 & ~n9549;
  assign n9561 = ~n9548 & n9560;
  assign n9562 = ~n9559 & ~n9561;
  assign n9563 = ~n9557 & n9562;
  assign n9564 = ~n9551 & n9563;
  assign n9565 = ~n9557 & ~n9559;
  assign n9566 = ~n9551 & ~n9561;
  assign n9567 = ~n9565 & ~n9566;
  assign n9568 = ~n9564 & ~n9567;
  assign n9569 = ~n9545 & ~n9568;
  assign n9570 = ~n9544 & ~n9564;
  assign n9571 = ~n9567 & n9570;
  assign n9572 = ~n9380 & n9571;
  assign n9573 = ~n9569 & ~n9572;
  assign n9574 = ~n9541 & n9573;
  assign n9575 = ~n9539 & n9574;
  assign n9576 = ~n9539 & ~n9541;
  assign n9577 = ~n9573 & ~n9576;
  assign n9578 = ~n9575 & ~n9577;
  assign n9579 = ~n9479 & ~n9578;
  assign n9580 = ~n9478 & n9579;
  assign n9581 = ~n9478 & ~n9479;
  assign n9582 = n9578 & ~n9581;
  assign n9583 = ~n9580 & ~n9582;
  assign n9584 = ~n9275 & ~n9282;
  assign n9585 = ~n9229 & n9584;
  assign n9586 = ~n9283 & n9585;
  assign n9587 = ~n9231 & n9586;
  assign n9588 = ~n9283 & n9584;
  assign n9589 = n9390 & n9588;
  assign n9590 = n9283 & ~n9584;
  assign n9591 = ~n9390 & n9590;
  assign n9592 = ~n9589 & ~n9591;
  assign n9593 = ~n9587 & n9592;
  assign n9594 = ~n9390 & ~n9584;
  assign n9595 = ~n9232 & n9594;
  assign n9596 = n9390 & n9585;
  assign n9597 = ~n9231 & n9596;
  assign n9598 = ~n9232 & n9590;
  assign n9599 = ~n9597 & ~n9598;
  assign n9600 = ~n9595 & n9599;
  assign n9601 = n9593 & n9600;
  assign n9602 = ~n9583 & ~n9601;
  assign n9603 = ~n9580 & n9593;
  assign n9604 = ~n9582 & n9603;
  assign n9605 = n9600 & n9604;
  assign n9606 = ~n9602 & ~n9605;
  assign n9607 = n9421 & n9606;
  assign n9608 = ~n9421 & ~n9606;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = ~n9416 & n9609;
  assign n9611 = ~n9400 & ~n9609;
  assign n9612 = ~n9415 & n9611;
  assign po45 = ~n9610 & ~n9612;
  assign n9614 = ~n9400 & ~n9608;
  assign n9615 = ~n9607 & n9614;
  assign n9616 = ~n9156 & ~n9399;
  assign n9617 = n9407 & n9616;
  assign n9618 = ~n8346 & n8901;
  assign n9619 = n8928 & n9618;
  assign n9620 = n9617 & n9619;
  assign n9621 = n9615 & n9620;
  assign n9622 = ~n8096 & n9621;
  assign n9623 = n9615 & n9616;
  assign n9624 = ~n9197 & n9623;
  assign n9625 = ~n9607 & ~n9614;
  assign n9626 = ~n9284 & ~n9392;
  assign n9627 = ~n9584 & ~n9626;
  assign n9628 = ~n9583 & n9601;
  assign n9629 = ~n9627 & ~n9628;
  assign n9630 = ~n9440 & ~n9449;
  assign n9631 = ~n9447 & n9630;
  assign n9632 = ~n9438 & n9631;
  assign n9633 = ~n9463 & ~n9632;
  assign n9634 = pi15 & ~n5091;
  assign n9635 = ~n5092 & n9634;
  assign n9636 = ~n5178 & n9635;
  assign n9637 = pi16 & ~n5093;
  assign n9638 = ~n9636 & ~n9637;
  assign n9639 = pi63 & ~n9638;
  assign n9640 = ~pi63 & ~n9637;
  assign n9641 = ~n9636 & n9640;
  assign n9642 = ~n9639 & ~n9641;
  assign n9643 = pi17 & ~n4513;
  assign n9644 = ~n4514 & n9643;
  assign n9645 = ~n4577 & n9644;
  assign n9646 = pi18 & ~n4515;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = pi61 & ~n9647;
  assign n9649 = ~pi61 & ~n9646;
  assign n9650 = ~n9645 & n9649;
  assign n9651 = ~n9648 & ~n9650;
  assign n9652 = ~n9642 & n9651;
  assign n9653 = n9642 & ~n9651;
  assign n9654 = ~n9652 & ~n9653;
  assign n9655 = pi19 & ~n3959;
  assign n9656 = ~n3960 & n9655;
  assign n9657 = ~n4233 & n9656;
  assign n9658 = pi20 & ~n3961;
  assign n9659 = ~n9657 & ~n9658;
  assign n9660 = pi59 & ~n9659;
  assign n9661 = ~pi59 & ~n9658;
  assign n9662 = ~n9657 & n9661;
  assign n9663 = ~n9660 & ~n9662;
  assign n9664 = ~n9654 & n9663;
  assign n9665 = ~n9652 & ~n9663;
  assign n9666 = ~n9653 & n9665;
  assign n9667 = ~n9664 & ~n9666;
  assign n9668 = n9633 & ~n9667;
  assign n9669 = ~n9633 & n9667;
  assign n9670 = n9467 & ~n9669;
  assign n9671 = ~n9668 & n9670;
  assign n9672 = ~n9668 & ~n9669;
  assign n9673 = ~n9467 & ~n9672;
  assign n9674 = ~n9671 & ~n9673;
  assign n9675 = ~n9536 & ~n9541;
  assign n9676 = n9674 & ~n9675;
  assign n9677 = ~n9536 & ~n9674;
  assign n9678 = ~n9541 & n9677;
  assign n9679 = n9575 & ~n9678;
  assign n9680 = ~n9676 & n9679;
  assign n9681 = ~n9676 & ~n9678;
  assign n9682 = ~n9575 & ~n9681;
  assign n9683 = ~n9680 & ~n9682;
  assign n9684 = ~n9492 & ~n9532;
  assign n9685 = pi21 & ~n3205;
  assign n9686 = ~n3206 & n9685;
  assign n9687 = ~n3463 & n9686;
  assign n9688 = pi22 & ~n3207;
  assign n9689 = ~n9687 & ~n9688;
  assign n9690 = pi57 & ~n9689;
  assign n9691 = ~pi57 & ~n9688;
  assign n9692 = ~n9687 & n9691;
  assign n9693 = ~n9690 & ~n9692;
  assign n9694 = ~n9514 & n9524;
  assign n9695 = ~n9511 & ~n9694;
  assign n9696 = n9693 & ~n9695;
  assign n9697 = pi23 & ~n2876;
  assign n9698 = ~n2877 & n9697;
  assign n9699 = ~n2960 & n9698;
  assign n9700 = pi24 & ~n2878;
  assign n9701 = ~n9699 & ~n9700;
  assign n9702 = pi55 & ~n9701;
  assign n9703 = pi25 & ~n2288;
  assign n9704 = ~n2289 & n9703;
  assign n9705 = ~n2647 & n9704;
  assign n9706 = pi26 & ~n2290;
  assign n9707 = ~n9705 & ~n9706;
  assign n9708 = pi53 & ~n9707;
  assign n9709 = ~pi53 & ~n9706;
  assign n9710 = ~n9705 & n9709;
  assign n9711 = ~pi55 & ~n9700;
  assign n9712 = ~n9699 & n9711;
  assign n9713 = ~n9710 & ~n9712;
  assign n9714 = ~n9708 & n9713;
  assign n9715 = ~n9702 & n9714;
  assign n9716 = ~n9708 & ~n9710;
  assign n9717 = ~n9702 & ~n9712;
  assign n9718 = ~n9716 & ~n9717;
  assign n9719 = ~n9715 & ~n9718;
  assign n9720 = pi27 & ~n2023;
  assign n9721 = ~n2024 & n9720;
  assign n9722 = ~n2079 & n9721;
  assign n9723 = pi28 & ~n2025;
  assign n9724 = ~n9722 & ~n9723;
  assign n9725 = pi51 & ~n9724;
  assign n9726 = ~pi51 & ~n9723;
  assign n9727 = ~n9722 & n9726;
  assign n9728 = ~n9725 & ~n9727;
  assign n9729 = ~n9719 & n9728;
  assign n9730 = ~n9715 & ~n9728;
  assign n9731 = ~n9718 & n9730;
  assign n9732 = ~n9729 & ~n9731;
  assign n9733 = ~n9511 & ~n9693;
  assign n9734 = ~n9694 & n9733;
  assign n9735 = ~n9732 & ~n9734;
  assign n9736 = ~n9696 & n9735;
  assign n9737 = ~n9696 & ~n9734;
  assign n9738 = n9732 & ~n9737;
  assign n9739 = ~n9736 & ~n9738;
  assign n9740 = ~n9684 & n9739;
  assign n9741 = n9684 & ~n9739;
  assign n9742 = ~n9740 & ~n9741;
  assign n9743 = ~n9569 & ~n9742;
  assign n9744 = n9569 & ~n9740;
  assign n9745 = ~n9741 & n9744;
  assign n9746 = n1214 & n1425;
  assign n9747 = pi31 & pi47;
  assign n9748 = ~n9746 & n9747;
  assign n9749 = pi31 & ~n9746;
  assign n9750 = ~pi47 & ~n9749;
  assign n9751 = ~n9748 & ~n9750;
  assign n9752 = pi29 & ~n1607;
  assign n9753 = ~n1608 & n9752;
  assign n9754 = ~n1782 & n9753;
  assign n9755 = pi30 & ~n1609;
  assign n9756 = ~n9754 & ~n9755;
  assign n9757 = pi49 & ~n9756;
  assign n9758 = ~pi49 & ~n9755;
  assign n9759 = ~n9754 & n9758;
  assign n9760 = ~n9757 & ~n9759;
  assign n9761 = ~n9751 & n9760;
  assign n9762 = n9751 & ~n9760;
  assign n9763 = ~n9761 & ~n9762;
  assign n9764 = n9567 & ~n9763;
  assign n9765 = ~n9567 & ~n9761;
  assign n9766 = ~n9762 & n9765;
  assign n9767 = ~n9764 & ~n9766;
  assign n9768 = ~n9745 & n9767;
  assign n9769 = ~n9743 & n9768;
  assign n9770 = ~n9743 & ~n9745;
  assign n9771 = ~n9767 & ~n9770;
  assign n9772 = ~n9769 & ~n9771;
  assign n9773 = ~n9683 & n9772;
  assign n9774 = ~n9680 & ~n9772;
  assign n9775 = ~n9682 & n9774;
  assign n9776 = ~n9773 & ~n9775;
  assign n9777 = ~n9478 & n9578;
  assign n9778 = n9273 & ~n9467;
  assign n9779 = ~n9468 & n9778;
  assign n9780 = ~n9476 & ~n9779;
  assign n9781 = ~n9479 & ~n9780;
  assign n9782 = ~n9777 & n9781;
  assign n9783 = ~n9479 & ~n9777;
  assign n9784 = n9780 & ~n9783;
  assign n9785 = ~n9782 & ~n9784;
  assign n9786 = ~n9776 & ~n9785;
  assign n9787 = n9776 & n9785;
  assign n9788 = ~n9786 & ~n9787;
  assign n9789 = ~n9629 & n9788;
  assign n9790 = n9629 & ~n9788;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = ~n9625 & ~n9791;
  assign n9793 = ~n9624 & n9792;
  assign n9794 = ~n9622 & n9793;
  assign n9795 = ~n9624 & ~n9625;
  assign n9796 = ~n9622 & n9795;
  assign n9797 = n9791 & ~n9796;
  assign po46 = ~n9794 & ~n9797;
  assign n9799 = ~n9621 & n9795;
  assign n9800 = ~n8093 & ~n9625;
  assign n9801 = ~n9624 & n9800;
  assign n9802 = ~n8087 & n9801;
  assign n9803 = ~n8363 & n9802;
  assign n9804 = ~n8360 & n9803;
  assign n9805 = ~n9799 & ~n9804;
  assign n9806 = ~n9641 & ~n9650;
  assign n9807 = ~n9648 & n9806;
  assign n9808 = ~n9639 & n9807;
  assign n9809 = ~n9664 & ~n9808;
  assign n9810 = pi16 & ~n5091;
  assign n9811 = ~n5092 & n9810;
  assign n9812 = ~n5178 & n9811;
  assign n9813 = pi17 & ~n5093;
  assign n9814 = ~n9812 & ~n9813;
  assign n9815 = pi63 & ~n9814;
  assign n9816 = ~pi63 & ~n9813;
  assign n9817 = ~n9812 & n9816;
  assign n9818 = ~n9815 & ~n9817;
  assign n9819 = pi18 & ~n4513;
  assign n9820 = ~n4514 & n9819;
  assign n9821 = ~n4577 & n9820;
  assign n9822 = pi19 & ~n4515;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = pi61 & ~n9823;
  assign n9825 = ~pi61 & ~n9822;
  assign n9826 = ~n9821 & n9825;
  assign n9827 = ~n9824 & ~n9826;
  assign n9828 = ~n9818 & n9827;
  assign n9829 = n9818 & ~n9827;
  assign n9830 = ~n9828 & ~n9829;
  assign n9831 = pi20 & ~n3959;
  assign n9832 = ~n3960 & n9831;
  assign n9833 = ~n4233 & n9832;
  assign n9834 = pi21 & ~n3961;
  assign n9835 = ~n9833 & ~n9834;
  assign n9836 = pi59 & ~n9835;
  assign n9837 = ~pi59 & ~n9834;
  assign n9838 = ~n9833 & n9837;
  assign n9839 = ~n9836 & ~n9838;
  assign n9840 = ~n9830 & n9839;
  assign n9841 = ~n9828 & ~n9839;
  assign n9842 = ~n9829 & n9841;
  assign n9843 = ~n9840 & ~n9842;
  assign n9844 = ~n9809 & n9843;
  assign n9845 = n9809 & ~n9843;
  assign n9846 = ~n9844 & ~n9845;
  assign n9847 = n9669 & ~n9846;
  assign n9848 = ~n9669 & ~n9844;
  assign n9849 = ~n9845 & n9848;
  assign n9850 = ~n9847 & ~n9849;
  assign n9851 = ~n9740 & n9850;
  assign n9852 = ~n9745 & n9851;
  assign n9853 = ~n9740 & ~n9745;
  assign n9854 = ~n9850 & ~n9853;
  assign n9855 = ~n9852 & ~n9854;
  assign n9856 = ~n9769 & ~n9855;
  assign n9857 = n9769 & ~n9852;
  assign n9858 = ~n9854 & n9857;
  assign n9859 = ~n9696 & ~n9736;
  assign n9860 = ~n9718 & n9728;
  assign n9861 = pi22 & ~n3205;
  assign n9862 = ~n3206 & n9861;
  assign n9863 = ~n3463 & n9862;
  assign n9864 = pi23 & ~n3207;
  assign n9865 = ~n9863 & ~n9864;
  assign n9866 = pi57 & ~n9865;
  assign n9867 = ~pi57 & ~n9864;
  assign n9868 = ~n9863 & n9867;
  assign n9869 = ~n9866 & ~n9868;
  assign n9870 = ~n9715 & ~n9869;
  assign n9871 = ~n9860 & n9870;
  assign n9872 = ~n9715 & ~n9860;
  assign n9873 = n9869 & ~n9872;
  assign n9874 = ~n9871 & ~n9873;
  assign n9875 = pi24 & ~n2876;
  assign n9876 = ~n2877 & n9875;
  assign n9877 = ~n2960 & n9876;
  assign n9878 = pi25 & ~n2878;
  assign n9879 = ~n9877 & ~n9878;
  assign n9880 = pi55 & ~n9879;
  assign n9881 = pi26 & ~n2288;
  assign n9882 = ~n2289 & n9881;
  assign n9883 = ~n2647 & n9882;
  assign n9884 = pi27 & ~n2290;
  assign n9885 = ~n9883 & ~n9884;
  assign n9886 = pi53 & ~n9885;
  assign n9887 = ~pi53 & ~n9884;
  assign n9888 = ~n9883 & n9887;
  assign n9889 = ~pi55 & ~n9878;
  assign n9890 = ~n9877 & n9889;
  assign n9891 = ~n9888 & ~n9890;
  assign n9892 = ~n9886 & n9891;
  assign n9893 = ~n9880 & n9892;
  assign n9894 = ~n9886 & ~n9888;
  assign n9895 = ~n9880 & ~n9890;
  assign n9896 = ~n9894 & ~n9895;
  assign n9897 = ~n9893 & ~n9896;
  assign n9898 = pi28 & ~n2023;
  assign n9899 = ~n2024 & n9898;
  assign n9900 = ~n2079 & n9899;
  assign n9901 = pi29 & ~n2025;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = pi51 & ~n9902;
  assign n9904 = ~pi51 & ~n9901;
  assign n9905 = ~n9900 & n9904;
  assign n9906 = ~n9903 & ~n9905;
  assign n9907 = ~n9897 & n9906;
  assign n9908 = ~n9893 & ~n9906;
  assign n9909 = ~n9896 & n9908;
  assign n9910 = ~n9907 & ~n9909;
  assign n9911 = ~n9874 & n9910;
  assign n9912 = n9874 & ~n9910;
  assign n9913 = ~n9911 & ~n9912;
  assign n9914 = ~n9859 & n9913;
  assign n9915 = n9859 & ~n9913;
  assign n9916 = ~n9914 & ~n9915;
  assign n9917 = ~n9766 & ~n9916;
  assign n9918 = n9766 & ~n9914;
  assign n9919 = ~n9915 & n9918;
  assign n9920 = pi30 & ~n1607;
  assign n9921 = ~n1608 & n9920;
  assign n9922 = ~n1782 & n9921;
  assign n9923 = pi31 & ~n1609;
  assign n9924 = ~n9922 & ~n9923;
  assign n9925 = pi49 & ~n9924;
  assign n9926 = ~pi49 & ~n9923;
  assign n9927 = ~n9922 & n9926;
  assign n9928 = ~n9925 & ~n9927;
  assign n9929 = n9761 & ~n9928;
  assign n9930 = ~n9761 & n9928;
  assign n9931 = ~n9929 & ~n9930;
  assign n9932 = ~n9919 & n9931;
  assign n9933 = ~n9917 & n9932;
  assign n9934 = ~n9917 & ~n9919;
  assign n9935 = ~n9931 & ~n9934;
  assign n9936 = ~n9933 & ~n9935;
  assign n9937 = ~n9858 & ~n9936;
  assign n9938 = ~n9856 & n9937;
  assign n9939 = ~n9856 & ~n9858;
  assign n9940 = n9936 & ~n9939;
  assign n9941 = ~n9938 & ~n9940;
  assign n9942 = ~n9682 & n9772;
  assign n9943 = ~n9671 & ~n9676;
  assign n9944 = ~n9680 & ~n9943;
  assign n9945 = ~n9942 & n9944;
  assign n9946 = ~n9680 & ~n9942;
  assign n9947 = n9943 & ~n9946;
  assign n9948 = ~n9945 & ~n9947;
  assign n9949 = ~n9941 & ~n9948;
  assign n9950 = n9941 & n9948;
  assign n9951 = ~n9949 & ~n9950;
  assign n9952 = ~n9780 & ~n9783;
  assign n9953 = ~n9786 & ~n9952;
  assign n9954 = ~n9951 & n9953;
  assign n9955 = n9951 & ~n9953;
  assign n9956 = ~n9954 & ~n9955;
  assign n9957 = ~n9789 & ~n9956;
  assign n9958 = ~n9805 & n9957;
  assign n9959 = ~n9790 & ~n9954;
  assign n9960 = ~n9955 & n9959;
  assign n9961 = ~n9799 & n9960;
  assign n9962 = ~n9804 & n9961;
  assign n9963 = ~n9789 & n9790;
  assign n9964 = ~n9956 & n9963;
  assign n9965 = n9789 & ~n9954;
  assign n9966 = ~n9955 & n9965;
  assign n9967 = ~n9964 & ~n9966;
  assign n9968 = ~n9962 & n9967;
  assign po47 = ~n9958 & n9968;
  assign n9970 = ~n7488 & ~n7789;
  assign n9971 = n8663 & n9970;
  assign n9972 = n8660 & n9185;
  assign n9973 = n9971 & n9972;
  assign n9974 = ~n9607 & ~n9789;
  assign n9975 = ~n9790 & n9974;
  assign n9976 = n9614 & n9616;
  assign n9977 = n8928 & n9407;
  assign n9978 = n9976 & n9977;
  assign n9979 = n9975 & n9978;
  assign n9980 = n9973 & n9979;
  assign n9981 = ~n8649 & n9980;
  assign n9982 = ~n8631 & n8901;
  assign n9983 = n9407 & n9982;
  assign n9984 = n9976 & n9983;
  assign n9985 = n9975 & n9984;
  assign n9986 = ~n8667 & n9985;
  assign n9987 = n9155 & ~n9399;
  assign n9988 = n9615 & n9987;
  assign n9989 = ~n9625 & ~n9789;
  assign n9990 = ~n9988 & n9989;
  assign n9991 = ~n9790 & ~n9990;
  assign n9992 = n9609 & n9791;
  assign n9993 = n9157 & n9401;
  assign n9994 = n9194 & n9993;
  assign n9995 = n9992 & n9994;
  assign n9996 = n8900 & ~n9155;
  assign n9997 = n9976 & n9996;
  assign n9998 = n9975 & n9997;
  assign n9999 = ~n9955 & ~n9998;
  assign n10000 = ~n9995 & n9999;
  assign n10001 = ~n9991 & n10000;
  assign n10002 = ~n9986 & n10001;
  assign n10003 = ~n9981 & n10002;
  assign n10004 = ~n9817 & ~n9826;
  assign n10005 = ~n9824 & n10004;
  assign n10006 = ~n9815 & n10005;
  assign n10007 = ~n9840 & ~n10006;
  assign n10008 = pi17 & ~n5091;
  assign n10009 = ~n5092 & n10008;
  assign n10010 = ~n5178 & n10009;
  assign n10011 = pi18 & ~n5093;
  assign n10012 = ~n10010 & ~n10011;
  assign n10013 = pi63 & ~n10012;
  assign n10014 = ~pi63 & ~n10011;
  assign n10015 = ~n10010 & n10014;
  assign n10016 = ~n10013 & ~n10015;
  assign n10017 = pi19 & ~n4513;
  assign n10018 = ~n4514 & n10017;
  assign n10019 = ~n4577 & n10018;
  assign n10020 = pi20 & ~n4515;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = pi61 & ~n10021;
  assign n10023 = ~pi61 & ~n10020;
  assign n10024 = ~n10019 & n10023;
  assign n10025 = ~n10022 & ~n10024;
  assign n10026 = ~n10016 & n10025;
  assign n10027 = n10016 & ~n10025;
  assign n10028 = ~n10026 & ~n10027;
  assign n10029 = pi21 & ~n3959;
  assign n10030 = ~n3960 & n10029;
  assign n10031 = ~n4233 & n10030;
  assign n10032 = pi22 & ~n3961;
  assign n10033 = ~n10031 & ~n10032;
  assign n10034 = pi59 & ~n10033;
  assign n10035 = ~pi59 & ~n10032;
  assign n10036 = ~n10031 & n10035;
  assign n10037 = ~n10034 & ~n10036;
  assign n10038 = ~n10028 & n10037;
  assign n10039 = ~n10026 & ~n10037;
  assign n10040 = ~n10027 & n10039;
  assign n10041 = ~n10038 & ~n10040;
  assign n10042 = ~n10007 & n10041;
  assign n10043 = n10007 & ~n10041;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = n9844 & ~n10044;
  assign n10046 = ~n9844 & ~n10042;
  assign n10047 = ~n10043 & n10046;
  assign n10048 = ~n10045 & ~n10047;
  assign n10049 = ~n9914 & n10048;
  assign n10050 = ~n9919 & n10049;
  assign n10051 = ~n9914 & ~n9919;
  assign n10052 = ~n10048 & ~n10051;
  assign n10053 = ~n10050 & ~n10052;
  assign n10054 = ~n9933 & ~n10053;
  assign n10055 = n9933 & ~n10050;
  assign n10056 = ~n10052 & n10055;
  assign n10057 = ~n9873 & ~n9912;
  assign n10058 = ~n9896 & n9906;
  assign n10059 = pi23 & ~n3205;
  assign n10060 = ~n3206 & n10059;
  assign n10061 = ~n3463 & n10060;
  assign n10062 = pi24 & ~n3207;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = pi57 & ~n10063;
  assign n10065 = ~pi57 & ~n10062;
  assign n10066 = ~n10061 & n10065;
  assign n10067 = ~n10064 & ~n10066;
  assign n10068 = ~n9893 & ~n10067;
  assign n10069 = ~n10058 & n10068;
  assign n10070 = ~n9893 & ~n10058;
  assign n10071 = n10067 & ~n10070;
  assign n10072 = ~n10069 & ~n10071;
  assign n10073 = pi25 & ~n2876;
  assign n10074 = ~n2877 & n10073;
  assign n10075 = ~n2960 & n10074;
  assign n10076 = pi26 & ~n2878;
  assign n10077 = ~n10075 & ~n10076;
  assign n10078 = pi55 & ~n10077;
  assign n10079 = pi27 & ~n2288;
  assign n10080 = ~n2289 & n10079;
  assign n10081 = ~n2647 & n10080;
  assign n10082 = pi28 & ~n2290;
  assign n10083 = ~n10081 & ~n10082;
  assign n10084 = pi53 & ~n10083;
  assign n10085 = ~pi53 & ~n10082;
  assign n10086 = ~n10081 & n10085;
  assign n10087 = ~pi55 & ~n10076;
  assign n10088 = ~n10075 & n10087;
  assign n10089 = ~n10086 & ~n10088;
  assign n10090 = ~n10084 & n10089;
  assign n10091 = ~n10078 & n10090;
  assign n10092 = ~n10084 & ~n10086;
  assign n10093 = ~n10078 & ~n10088;
  assign n10094 = ~n10092 & ~n10093;
  assign n10095 = ~n10091 & ~n10094;
  assign n10096 = pi29 & ~n2023;
  assign n10097 = ~n2024 & n10096;
  assign n10098 = ~n2079 & n10097;
  assign n10099 = pi30 & ~n2025;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = pi51 & ~n10100;
  assign n10102 = ~pi51 & ~n10099;
  assign n10103 = ~n10098 & n10102;
  assign n10104 = ~n10101 & ~n10103;
  assign n10105 = ~n10095 & n10104;
  assign n10106 = ~n10091 & ~n10104;
  assign n10107 = ~n10094 & n10106;
  assign n10108 = ~n10105 & ~n10107;
  assign n10109 = ~n10072 & n10108;
  assign n10110 = n10072 & ~n10108;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10057 & n10111;
  assign n10113 = n10057 & ~n10111;
  assign n10114 = ~n10112 & ~n10113;
  assign n10115 = n9929 & ~n10114;
  assign n10116 = ~n9929 & ~n10112;
  assign n10117 = ~n10113 & n10116;
  assign n10118 = ~n10115 & ~n10117;
  assign n10119 = n1609 & n1782;
  assign n10120 = pi31 & pi49;
  assign n10121 = ~n10119 & n10120;
  assign n10122 = pi31 & ~n10119;
  assign n10123 = ~pi49 & ~n10122;
  assign n10124 = ~n10121 & ~n10123;
  assign n10125 = n9928 & ~n10124;
  assign n10126 = ~n9928 & n10124;
  assign n10127 = ~n10125 & ~n10126;
  assign n10128 = ~n10118 & n10127;
  assign n10129 = ~n10115 & ~n10127;
  assign n10130 = ~n10117 & n10129;
  assign n10131 = ~n10128 & ~n10130;
  assign n10132 = ~n10056 & ~n10131;
  assign n10133 = ~n10054 & n10132;
  assign n10134 = ~n10054 & ~n10056;
  assign n10135 = n10131 & ~n10134;
  assign n10136 = ~n10133 & ~n10135;
  assign n10137 = ~n9856 & n9936;
  assign n10138 = n9669 & ~n9844;
  assign n10139 = ~n9845 & n10138;
  assign n10140 = ~n9854 & ~n10139;
  assign n10141 = ~n9858 & ~n10140;
  assign n10142 = ~n10137 & n10141;
  assign n10143 = ~n9858 & ~n10137;
  assign n10144 = n10140 & ~n10143;
  assign n10145 = ~n10142 & ~n10144;
  assign n10146 = ~n10136 & ~n10145;
  assign n10147 = n10136 & n10145;
  assign n10148 = ~n10146 & ~n10147;
  assign n10149 = ~n9943 & ~n9946;
  assign n10150 = ~n9949 & ~n10149;
  assign n10151 = n10148 & ~n10150;
  assign n10152 = ~n10148 & n10150;
  assign n10153 = ~n9954 & ~n10152;
  assign n10154 = ~n10151 & n10153;
  assign n10155 = ~n10003 & n10154;
  assign n10156 = ~n10151 & ~n10152;
  assign n10157 = ~n9954 & ~n10003;
  assign n10158 = ~n10156 & ~n10157;
  assign po48 = ~n10155 & ~n10158;
  assign n10160 = ~n9991 & n9999;
  assign n10161 = n10154 & ~n10160;
  assign n10162 = n8937 & ~n10161;
  assign n10163 = ~n8927 & n10162;
  assign n10164 = ~n8916 & n10163;
  assign n10165 = n8901 & ~n9155;
  assign n10166 = n9976 & n10165;
  assign n10167 = ~n9955 & ~n10152;
  assign n10168 = ~n10151 & n10167;
  assign n10169 = n9959 & n9974;
  assign n10170 = n10168 & n10169;
  assign n10171 = n10166 & n10170;
  assign n10172 = ~n10161 & ~n10171;
  assign n10173 = ~n10164 & ~n10172;
  assign n10174 = ~n10140 & ~n10143;
  assign n10175 = ~n10146 & ~n10174;
  assign n10176 = ~n10054 & n10131;
  assign n10177 = ~n10056 & ~n10176;
  assign n10178 = n9844 & ~n10042;
  assign n10179 = ~n10043 & n10178;
  assign n10180 = ~n10052 & ~n10179;
  assign n10181 = ~n10177 & ~n10180;
  assign n10182 = ~n10056 & n10180;
  assign n10183 = ~n10176 & n10182;
  assign n10184 = ~n10181 & ~n10183;
  assign n10185 = n9929 & ~n10113;
  assign n10186 = ~n10015 & ~n10024;
  assign n10187 = ~n10022 & n10186;
  assign n10188 = ~n10013 & n10187;
  assign n10189 = ~n10038 & ~n10188;
  assign n10190 = pi18 & ~n5091;
  assign n10191 = ~n5092 & n10190;
  assign n10192 = ~n5178 & n10191;
  assign n10193 = pi19 & ~n5093;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = pi63 & ~n10194;
  assign n10196 = ~pi63 & ~n10193;
  assign n10197 = ~n10192 & n10196;
  assign n10198 = ~n10195 & ~n10197;
  assign n10199 = pi20 & ~n4513;
  assign n10200 = ~n4514 & n10199;
  assign n10201 = ~n4577 & n10200;
  assign n10202 = pi21 & ~n4515;
  assign n10203 = ~n10201 & ~n10202;
  assign n10204 = pi61 & ~n10203;
  assign n10205 = ~pi61 & ~n10202;
  assign n10206 = ~n10201 & n10205;
  assign n10207 = ~n10204 & ~n10206;
  assign n10208 = ~n10198 & n10207;
  assign n10209 = n10198 & ~n10207;
  assign n10210 = ~n10208 & ~n10209;
  assign n10211 = pi22 & ~n3959;
  assign n10212 = ~n3960 & n10211;
  assign n10213 = ~n4233 & n10212;
  assign n10214 = pi23 & ~n3961;
  assign n10215 = ~n10213 & ~n10214;
  assign n10216 = pi59 & ~n10215;
  assign n10217 = ~pi59 & ~n10214;
  assign n10218 = ~n10213 & n10217;
  assign n10219 = ~n10216 & ~n10218;
  assign n10220 = ~n10210 & n10219;
  assign n10221 = ~n10208 & ~n10219;
  assign n10222 = ~n10209 & n10221;
  assign n10223 = ~n10220 & ~n10222;
  assign n10224 = ~n10189 & n10223;
  assign n10225 = n10189 & ~n10223;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = n10042 & ~n10226;
  assign n10228 = ~n10042 & ~n10224;
  assign n10229 = ~n10225 & n10228;
  assign n10230 = ~n10227 & ~n10229;
  assign n10231 = ~n10112 & n10230;
  assign n10232 = ~n10185 & n10231;
  assign n10233 = ~n10112 & ~n10185;
  assign n10234 = ~n10230 & ~n10233;
  assign n10235 = ~n10232 & ~n10234;
  assign n10236 = ~n10128 & ~n10235;
  assign n10237 = n10127 & ~n10232;
  assign n10238 = ~n10118 & n10237;
  assign n10239 = ~n10234 & n10238;
  assign n10240 = ~n10071 & ~n10110;
  assign n10241 = pi24 & ~n3205;
  assign n10242 = ~n3206 & n10241;
  assign n10243 = ~n3463 & n10242;
  assign n10244 = pi25 & ~n3207;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = pi57 & ~n10245;
  assign n10247 = ~pi57 & ~n10244;
  assign n10248 = ~n10243 & n10247;
  assign n10249 = ~n10246 & ~n10248;
  assign n10250 = ~n10094 & n10104;
  assign n10251 = ~n10091 & ~n10250;
  assign n10252 = n10249 & ~n10251;
  assign n10253 = ~n10091 & ~n10249;
  assign n10254 = ~n10250 & n10253;
  assign n10255 = pi26 & ~n2876;
  assign n10256 = ~n2877 & n10255;
  assign n10257 = ~n2960 & n10256;
  assign n10258 = pi27 & ~n2878;
  assign n10259 = ~n10257 & ~n10258;
  assign n10260 = pi55 & ~n10259;
  assign n10261 = ~pi55 & ~n10258;
  assign n10262 = ~n10257 & n10261;
  assign n10263 = ~n10260 & ~n10262;
  assign n10264 = pi28 & ~n2288;
  assign n10265 = ~n2289 & n10264;
  assign n10266 = ~n2647 & n10265;
  assign n10267 = pi29 & ~n2290;
  assign n10268 = ~n10266 & ~n10267;
  assign n10269 = pi53 & ~n10268;
  assign n10270 = ~pi53 & ~n10267;
  assign n10271 = ~n10266 & n10270;
  assign n10272 = ~n10269 & ~n10271;
  assign n10273 = ~n10263 & n10272;
  assign n10274 = n10263 & ~n10272;
  assign n10275 = ~n10273 & ~n10274;
  assign n10276 = pi30 & ~n2023;
  assign n10277 = ~n2024 & n10276;
  assign n10278 = ~n2079 & n10277;
  assign n10279 = pi31 & ~n2025;
  assign n10280 = ~n10278 & ~n10279;
  assign n10281 = pi51 & ~n10280;
  assign n10282 = ~pi51 & ~n10279;
  assign n10283 = ~n10278 & n10282;
  assign n10284 = ~n10281 & ~n10283;
  assign n10285 = ~n10275 & n10284;
  assign n10286 = ~n10273 & ~n10284;
  assign n10287 = ~n10274 & n10286;
  assign n10288 = ~n10285 & ~n10287;
  assign n10289 = ~n10254 & n10288;
  assign n10290 = ~n10252 & n10289;
  assign n10291 = ~n10252 & ~n10254;
  assign n10292 = ~n10288 & ~n10291;
  assign n10293 = ~n10290 & ~n10292;
  assign n10294 = ~n10240 & n10293;
  assign n10295 = n10240 & ~n10293;
  assign n10296 = ~n10294 & ~n10295;
  assign n10297 = n10125 & ~n10296;
  assign n10298 = ~n10125 & ~n10294;
  assign n10299 = ~n10295 & n10298;
  assign n10300 = ~n10297 & ~n10299;
  assign n10301 = ~n10239 & n10300;
  assign n10302 = ~n10236 & n10301;
  assign n10303 = ~n10236 & ~n10239;
  assign n10304 = ~n10300 & ~n10303;
  assign n10305 = ~n10302 & ~n10304;
  assign n10306 = ~n10184 & n10305;
  assign n10307 = ~n10183 & ~n10305;
  assign n10308 = ~n10181 & n10307;
  assign n10309 = ~n10306 & ~n10308;
  assign n10310 = ~n10175 & ~n10309;
  assign n10311 = ~n10174 & ~n10308;
  assign n10312 = ~n10146 & n10311;
  assign n10313 = ~n10306 & n10312;
  assign n10314 = ~n10310 & ~n10313;
  assign n10315 = ~n10151 & ~n10314;
  assign n10316 = ~n10173 & n10315;
  assign n10317 = ~n10151 & ~n10173;
  assign n10318 = n10314 & ~n10317;
  assign po49 = ~n10316 & ~n10318;
  assign n10320 = n7183 & ~n9179;
  assign n10321 = ~n9167 & n10320;
  assign n10322 = n8929 & n9973;
  assign n10323 = ~n10321 & n10322;
  assign n10324 = ~n8347 & ~n8632;
  assign n10325 = n9982 & n10324;
  assign n10326 = ~n8657 & n10325;
  assign n10327 = n9196 & ~n10326;
  assign n10328 = ~n10323 & n10327;
  assign n10329 = n9614 & n9974;
  assign n10330 = n9616 & n10329;
  assign n10331 = ~n10151 & ~n10310;
  assign n10332 = ~n10313 & n10331;
  assign n10333 = n9959 & n10167;
  assign n10334 = n10332 & n10333;
  assign n10335 = n10330 & n10334;
  assign n10336 = ~n10328 & n10335;
  assign n10337 = ~n9614 & n9974;
  assign n10338 = n10333 & n10337;
  assign n10339 = n10332 & n10338;
  assign n10340 = n9965 & n10168;
  assign n10341 = n9955 & ~n10152;
  assign n10342 = ~n10151 & n10341;
  assign n10343 = n10331 & ~n10342;
  assign n10344 = ~n10340 & n10343;
  assign n10345 = ~n10313 & ~n10344;
  assign n10346 = ~n10339 & ~n10345;
  assign n10347 = ~n10336 & n10346;
  assign n10348 = ~n10183 & n10305;
  assign n10349 = ~n10181 & ~n10348;
  assign n10350 = n10042 & ~n10224;
  assign n10351 = ~n10225 & n10350;
  assign n10352 = ~n10234 & ~n10351;
  assign n10353 = ~n10239 & n10352;
  assign n10354 = ~n10303 & n10353;
  assign n10355 = n10300 & ~n10352;
  assign n10356 = ~n10239 & n10355;
  assign n10357 = ~n10236 & n10356;
  assign n10358 = n10239 & ~n10352;
  assign n10359 = ~n10300 & n10352;
  assign n10360 = ~n10239 & n10359;
  assign n10361 = ~n10358 & ~n10360;
  assign n10362 = ~n10357 & n10361;
  assign n10363 = ~n10354 & n10362;
  assign n10364 = n10125 & ~n10295;
  assign n10365 = ~n10197 & ~n10206;
  assign n10366 = ~n10204 & n10365;
  assign n10367 = ~n10195 & n10366;
  assign n10368 = ~n10220 & ~n10367;
  assign n10369 = pi19 & ~n5091;
  assign n10370 = ~n5092 & n10369;
  assign n10371 = ~n5178 & n10370;
  assign n10372 = pi20 & ~n5093;
  assign n10373 = ~n10371 & ~n10372;
  assign n10374 = pi63 & ~n10373;
  assign n10375 = ~pi63 & ~n10372;
  assign n10376 = ~n10371 & n10375;
  assign n10377 = ~n10374 & ~n10376;
  assign n10378 = pi21 & ~n4513;
  assign n10379 = ~n4514 & n10378;
  assign n10380 = ~n4577 & n10379;
  assign n10381 = pi22 & ~n4515;
  assign n10382 = ~n10380 & ~n10381;
  assign n10383 = pi61 & ~n10382;
  assign n10384 = ~pi61 & ~n10381;
  assign n10385 = ~n10380 & n10384;
  assign n10386 = ~n10383 & ~n10385;
  assign n10387 = ~n10377 & n10386;
  assign n10388 = n10377 & ~n10386;
  assign n10389 = ~n10387 & ~n10388;
  assign n10390 = pi23 & ~n3959;
  assign n10391 = ~n3960 & n10390;
  assign n10392 = ~n4233 & n10391;
  assign n10393 = pi24 & ~n3961;
  assign n10394 = ~n10392 & ~n10393;
  assign n10395 = pi59 & ~n10394;
  assign n10396 = ~pi59 & ~n10393;
  assign n10397 = ~n10392 & n10396;
  assign n10398 = ~n10395 & ~n10397;
  assign n10399 = ~n10389 & n10398;
  assign n10400 = ~n10387 & ~n10398;
  assign n10401 = ~n10388 & n10400;
  assign n10402 = ~n10399 & ~n10401;
  assign n10403 = ~n10368 & n10402;
  assign n10404 = n10368 & ~n10402;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = n10224 & ~n10405;
  assign n10407 = ~n10224 & ~n10403;
  assign n10408 = ~n10404 & n10407;
  assign n10409 = ~n10406 & ~n10408;
  assign n10410 = ~n10294 & n10409;
  assign n10411 = ~n10364 & n10410;
  assign n10412 = ~n10294 & ~n10364;
  assign n10413 = ~n10409 & ~n10412;
  assign n10414 = ~n10411 & ~n10413;
  assign n10415 = n10300 & ~n10414;
  assign n10416 = ~n10300 & ~n10411;
  assign n10417 = ~n10413 & n10416;
  assign n10418 = pi27 & ~n2876;
  assign n10419 = ~n2877 & n10418;
  assign n10420 = ~n2960 & n10419;
  assign n10421 = pi28 & ~n2878;
  assign n10422 = ~n10420 & ~n10421;
  assign n10423 = pi55 & ~n10422;
  assign n10424 = ~pi55 & ~n10421;
  assign n10425 = ~n10420 & n10424;
  assign n10426 = ~n10423 & ~n10425;
  assign n10427 = pi29 & ~n2288;
  assign n10428 = ~n2289 & n10427;
  assign n10429 = ~n2647 & n10428;
  assign n10430 = pi30 & ~n2290;
  assign n10431 = ~n10429 & ~n10430;
  assign n10432 = pi53 & ~n10431;
  assign n10433 = ~pi53 & ~n10430;
  assign n10434 = ~n10429 & n10433;
  assign n10435 = ~n10432 & ~n10434;
  assign n10436 = ~n10426 & n10435;
  assign n10437 = n10426 & ~n10435;
  assign n10438 = ~n10436 & ~n10437;
  assign n10439 = n2025 & n2079;
  assign n10440 = pi31 & pi51;
  assign n10441 = ~n10439 & n10440;
  assign n10442 = pi31 & ~n10439;
  assign n10443 = ~pi51 & ~n10442;
  assign n10444 = ~n10441 & ~n10443;
  assign n10445 = ~n10438 & ~n10444;
  assign n10446 = ~n10436 & n10444;
  assign n10447 = ~n10437 & n10446;
  assign n10448 = ~n10445 & ~n10447;
  assign n10449 = ~n10262 & ~n10271;
  assign n10450 = ~n10269 & n10449;
  assign n10451 = ~n10260 & n10450;
  assign n10452 = pi25 & ~n3205;
  assign n10453 = ~n3206 & n10452;
  assign n10454 = ~n3463 & n10453;
  assign n10455 = pi26 & ~n3207;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = pi57 & ~n10456;
  assign n10458 = ~pi57 & ~n10455;
  assign n10459 = ~n10454 & n10458;
  assign n10460 = ~n10457 & ~n10459;
  assign n10461 = ~n10451 & ~n10460;
  assign n10462 = ~n10285 & n10461;
  assign n10463 = ~n10285 & ~n10451;
  assign n10464 = n10460 & ~n10463;
  assign n10465 = ~n10462 & ~n10464;
  assign n10466 = ~n10448 & ~n10465;
  assign n10467 = ~n10252 & ~n10290;
  assign n10468 = n10448 & ~n10462;
  assign n10469 = ~n10464 & n10468;
  assign n10470 = ~n10467 & ~n10469;
  assign n10471 = ~n10466 & n10470;
  assign n10472 = ~n10466 & ~n10469;
  assign n10473 = n10467 & ~n10472;
  assign n10474 = ~n10471 & ~n10473;
  assign n10475 = ~n10417 & n10474;
  assign n10476 = ~n10415 & n10475;
  assign n10477 = ~n10415 & ~n10417;
  assign n10478 = ~n10474 & ~n10477;
  assign n10479 = ~n10476 & ~n10478;
  assign n10480 = ~n10363 & n10479;
  assign n10481 = n10363 & ~n10479;
  assign n10482 = ~n10480 & ~n10481;
  assign n10483 = ~n10349 & ~n10482;
  assign n10484 = n10349 & ~n10480;
  assign n10485 = ~n10481 & n10484;
  assign n10486 = ~n10483 & ~n10485;
  assign n10487 = ~n10347 & n10486;
  assign n10488 = ~n10339 & ~n10486;
  assign n10489 = ~n10345 & n10488;
  assign n10490 = ~n10336 & n10489;
  assign po50 = ~n10487 & ~n10490;
  assign n10492 = n10156 & n10314;
  assign n10493 = n9791 & n9956;
  assign n10494 = n9401 & n9609;
  assign n10495 = n10493 & n10494;
  assign n10496 = n10492 & n10495;
  assign n10497 = ~n9201 & n10496;
  assign n10498 = n7520 & n10346;
  assign n10499 = ~n10497 & n10498;
  assign n10500 = ~n7799 & ~n7800;
  assign n10501 = n10499 & n10500;
  assign n10502 = n9617 & n10329;
  assign n10503 = n10334 & n10502;
  assign n10504 = n9411 & n10503;
  assign n10505 = n10346 & ~n10504;
  assign n10506 = ~n10497 & n10505;
  assign n10507 = ~n10485 & ~n10506;
  assign n10508 = ~n10501 & n10507;
  assign n10509 = ~n10483 & ~n10508;
  assign n10510 = n10363 & n10479;
  assign n10511 = ~n10239 & ~n10302;
  assign n10512 = ~n10352 & ~n10511;
  assign n10513 = ~n10376 & ~n10385;
  assign n10514 = ~n10383 & n10513;
  assign n10515 = ~n10374 & n10514;
  assign n10516 = ~n10399 & ~n10515;
  assign n10517 = pi20 & ~n5091;
  assign n10518 = ~n5092 & n10517;
  assign n10519 = ~n5178 & n10518;
  assign n10520 = pi21 & ~n5093;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = pi63 & ~n10521;
  assign n10523 = ~pi63 & ~n10520;
  assign n10524 = ~n10519 & n10523;
  assign n10525 = ~n10522 & ~n10524;
  assign n10526 = pi22 & ~n4513;
  assign n10527 = ~n4514 & n10526;
  assign n10528 = ~n4577 & n10527;
  assign n10529 = pi23 & ~n4515;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = pi61 & ~n10530;
  assign n10532 = ~pi61 & ~n10529;
  assign n10533 = ~n10528 & n10532;
  assign n10534 = ~n10531 & ~n10533;
  assign n10535 = ~n10525 & n10534;
  assign n10536 = n10525 & ~n10534;
  assign n10537 = ~n10535 & ~n10536;
  assign n10538 = pi24 & ~n3959;
  assign n10539 = ~n3960 & n10538;
  assign n10540 = ~n4233 & n10539;
  assign n10541 = pi25 & ~n3961;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = pi59 & ~n10542;
  assign n10544 = ~pi59 & ~n10541;
  assign n10545 = ~n10540 & n10544;
  assign n10546 = ~n10543 & ~n10545;
  assign n10547 = ~n10537 & n10546;
  assign n10548 = ~n10535 & ~n10546;
  assign n10549 = ~n10536 & n10548;
  assign n10550 = ~n10547 & ~n10549;
  assign n10551 = n10516 & ~n10550;
  assign n10552 = ~n10516 & n10550;
  assign n10553 = n10403 & ~n10552;
  assign n10554 = ~n10551 & n10553;
  assign n10555 = ~n10551 & ~n10552;
  assign n10556 = ~n10403 & ~n10555;
  assign n10557 = ~n10554 & ~n10556;
  assign n10558 = n10471 & ~n10557;
  assign n10559 = ~n10471 & n10557;
  assign n10560 = ~n10558 & ~n10559;
  assign n10561 = ~n10425 & ~n10434;
  assign n10562 = ~n10432 & n10561;
  assign n10563 = ~n10423 & n10562;
  assign n10564 = pi26 & ~n3205;
  assign n10565 = ~n3206 & n10564;
  assign n10566 = ~n3463 & n10565;
  assign n10567 = pi27 & ~n3207;
  assign n10568 = ~n10566 & ~n10567;
  assign n10569 = pi57 & ~n10568;
  assign n10570 = ~pi57 & ~n10567;
  assign n10571 = ~n10566 & n10570;
  assign n10572 = ~n10569 & ~n10571;
  assign n10573 = ~n10563 & ~n10572;
  assign n10574 = ~n10445 & n10573;
  assign n10575 = ~n10445 & ~n10563;
  assign n10576 = n10572 & ~n10575;
  assign n10577 = ~n10574 & ~n10576;
  assign n10578 = pi30 & ~n2288;
  assign n10579 = ~n2289 & n10578;
  assign n10580 = ~n2647 & n10579;
  assign n10581 = pi31 & ~n2290;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = pi53 & ~n10582;
  assign n10584 = pi28 & ~n2876;
  assign n10585 = ~n2877 & n10584;
  assign n10586 = ~n2960 & n10585;
  assign n10587 = pi29 & ~n2878;
  assign n10588 = ~n10586 & ~n10587;
  assign n10589 = pi55 & ~n10588;
  assign n10590 = ~pi55 & ~n10587;
  assign n10591 = ~n10586 & n10590;
  assign n10592 = ~pi53 & ~n10581;
  assign n10593 = ~n10580 & n10592;
  assign n10594 = ~n10591 & ~n10593;
  assign n10595 = ~n10589 & n10594;
  assign n10596 = ~n10583 & n10595;
  assign n10597 = ~n10589 & ~n10591;
  assign n10598 = ~n10583 & ~n10593;
  assign n10599 = ~n10597 & ~n10598;
  assign n10600 = ~n10596 & ~n10599;
  assign n10601 = ~n10577 & n10600;
  assign n10602 = ~n10464 & ~n10469;
  assign n10603 = ~n10574 & ~n10600;
  assign n10604 = ~n10576 & n10603;
  assign n10605 = ~n10602 & ~n10604;
  assign n10606 = ~n10601 & n10605;
  assign n10607 = ~n10601 & ~n10604;
  assign n10608 = n10602 & ~n10607;
  assign n10609 = ~n10606 & ~n10608;
  assign n10610 = ~n10560 & n10609;
  assign n10611 = n10560 & ~n10609;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = n10224 & ~n10403;
  assign n10614 = ~n10404 & n10613;
  assign n10615 = ~n10413 & ~n10614;
  assign n10616 = ~n10417 & ~n10615;
  assign n10617 = ~n10612 & n10616;
  assign n10618 = ~n10476 & n10617;
  assign n10619 = ~n10610 & n10615;
  assign n10620 = ~n10611 & n10619;
  assign n10621 = ~n10417 & n10620;
  assign n10622 = ~n10476 & n10621;
  assign n10623 = ~n10618 & ~n10622;
  assign n10624 = ~n10512 & n10623;
  assign n10625 = ~n10417 & ~n10476;
  assign n10626 = n10612 & ~n10615;
  assign n10627 = ~n10625 & n10626;
  assign n10628 = ~n10612 & n10615;
  assign n10629 = ~n10625 & n10628;
  assign n10630 = ~n10627 & ~n10629;
  assign n10631 = n10624 & n10630;
  assign n10632 = ~n10510 & n10631;
  assign n10633 = ~n10510 & ~n10512;
  assign n10634 = n10623 & ~n10627;
  assign n10635 = ~n10629 & n10634;
  assign n10636 = ~n10633 & ~n10635;
  assign n10637 = ~n10632 & ~n10636;
  assign n10638 = ~n10509 & n10637;
  assign n10639 = ~n10483 & ~n10637;
  assign n10640 = ~n10508 & n10639;
  assign po51 = ~n10638 & ~n10640;
  assign n10642 = n10486 & n10637;
  assign n10643 = n8050 & ~n8347;
  assign n10644 = n9618 & n10643;
  assign n10645 = n9184 & n10644;
  assign n10646 = ~n9400 & ~n10645;
  assign n10647 = ~n9198 & n10646;
  assign n10648 = ~n9399 & ~n10647;
  assign n10649 = ~n10313 & n10642;
  assign n10650 = ~n10344 & n10649;
  assign n10651 = ~n10483 & ~n10636;
  assign n10652 = ~n10632 & ~n10651;
  assign n10653 = ~n9608 & ~n10652;
  assign n10654 = ~n10650 & n10653;
  assign n10655 = ~n10648 & n10654;
  assign n10656 = n9974 & n10642;
  assign n10657 = n10333 & n10656;
  assign n10658 = n10332 & n10657;
  assign n10659 = ~n10652 & ~n10658;
  assign n10660 = ~n10650 & n10659;
  assign n10661 = ~n10655 & ~n10660;
  assign n10662 = ~n10642 & ~n10661;
  assign n10663 = n8659 & n9185;
  assign n10664 = n6102 & n10663;
  assign n10665 = ~n7128 & ~n7789;
  assign n10666 = n8660 & n10665;
  assign n10667 = n9409 & n10666;
  assign n10668 = n10664 & n10667;
  assign n10669 = n7170 & n10668;
  assign n10670 = n10503 & n10669;
  assign n10671 = ~n8077 & n10670;
  assign n10672 = n7500 & n8089;
  assign n10673 = ~n7788 & ~n10672;
  assign n10674 = ~n7515 & n10673;
  assign n10675 = ~n7789 & ~n8050;
  assign n10676 = n9186 & n10675;
  assign n10677 = n9184 & n10494;
  assign n10678 = n10492 & n10493;
  assign n10679 = n10677 & n10678;
  assign n10680 = n10676 & n10679;
  assign n10681 = ~n10674 & n10680;
  assign n10682 = ~n10661 & ~n10681;
  assign n10683 = ~n10671 & n10682;
  assign n10684 = ~n10662 & ~n10683;
  assign n10685 = ~n10615 & ~n10625;
  assign n10686 = ~n10417 & n10615;
  assign n10687 = ~n10476 & n10686;
  assign n10688 = n10612 & ~n10687;
  assign n10689 = ~n10685 & ~n10688;
  assign n10690 = n10554 & ~n10610;
  assign n10691 = ~n10466 & ~n10554;
  assign n10692 = ~n10556 & n10691;
  assign n10693 = n10470 & n10692;
  assign n10694 = ~n10554 & ~n10606;
  assign n10695 = ~n10608 & n10694;
  assign n10696 = ~n10560 & n10695;
  assign n10697 = ~n10693 & ~n10696;
  assign n10698 = ~n10690 & n10697;
  assign n10699 = ~n10524 & ~n10533;
  assign n10700 = ~n10531 & n10699;
  assign n10701 = ~n10522 & n10700;
  assign n10702 = ~n10547 & ~n10701;
  assign n10703 = pi21 & ~n5091;
  assign n10704 = ~n5092 & n10703;
  assign n10705 = ~n5178 & n10704;
  assign n10706 = pi22 & ~n5093;
  assign n10707 = ~n10705 & ~n10706;
  assign n10708 = pi63 & ~n10707;
  assign n10709 = ~pi63 & ~n10706;
  assign n10710 = ~n10705 & n10709;
  assign n10711 = ~n10708 & ~n10710;
  assign n10712 = pi23 & ~n4513;
  assign n10713 = ~n4514 & n10712;
  assign n10714 = ~n4577 & n10713;
  assign n10715 = pi24 & ~n4515;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = pi61 & ~n10716;
  assign n10718 = ~pi61 & ~n10715;
  assign n10719 = ~n10714 & n10718;
  assign n10720 = ~n10717 & ~n10719;
  assign n10721 = ~n10711 & n10720;
  assign n10722 = n10711 & ~n10720;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = pi25 & ~n3959;
  assign n10725 = ~n3960 & n10724;
  assign n10726 = ~n4233 & n10725;
  assign n10727 = pi26 & ~n3961;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = pi59 & ~n10728;
  assign n10730 = ~pi59 & ~n10727;
  assign n10731 = ~n10726 & n10730;
  assign n10732 = ~n10729 & ~n10731;
  assign n10733 = ~n10723 & n10732;
  assign n10734 = ~n10721 & ~n10732;
  assign n10735 = ~n10722 & n10734;
  assign n10736 = ~n10733 & ~n10735;
  assign n10737 = n10702 & ~n10736;
  assign n10738 = ~n10702 & n10736;
  assign n10739 = n10552 & ~n10738;
  assign n10740 = ~n10737 & n10739;
  assign n10741 = ~n10737 & ~n10738;
  assign n10742 = ~n10552 & ~n10741;
  assign n10743 = ~n10740 & ~n10742;
  assign n10744 = n10606 & ~n10743;
  assign n10745 = ~n10606 & n10743;
  assign n10746 = ~n10744 & ~n10745;
  assign n10747 = pi27 & ~n3205;
  assign n10748 = ~n3206 & n10747;
  assign n10749 = ~n3463 & n10748;
  assign n10750 = pi28 & ~n3207;
  assign n10751 = ~n10749 & ~n10750;
  assign n10752 = pi57 & ~n10751;
  assign n10753 = ~pi57 & ~n10750;
  assign n10754 = ~n10749 & n10753;
  assign n10755 = ~n10752 & ~n10754;
  assign n10756 = ~n10599 & n10755;
  assign n10757 = n10599 & ~n10755;
  assign n10758 = n2290 & n2647;
  assign n10759 = pi31 & pi53;
  assign n10760 = ~n10758 & n10759;
  assign n10761 = pi31 & ~n10758;
  assign n10762 = ~pi53 & ~n10761;
  assign n10763 = ~n10760 & ~n10762;
  assign n10764 = pi29 & ~n2876;
  assign n10765 = ~n2877 & n10764;
  assign n10766 = ~n2960 & n10765;
  assign n10767 = pi30 & ~n2878;
  assign n10768 = ~n10766 & ~n10767;
  assign n10769 = pi55 & ~n10768;
  assign n10770 = ~pi55 & ~n10767;
  assign n10771 = ~n10766 & n10770;
  assign n10772 = ~n10769 & ~n10771;
  assign n10773 = ~n10763 & n10772;
  assign n10774 = n10763 & ~n10772;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = ~n10757 & n10775;
  assign n10777 = ~n10756 & n10776;
  assign n10778 = ~n10756 & ~n10757;
  assign n10779 = ~n10775 & ~n10778;
  assign n10780 = ~n10777 & ~n10779;
  assign n10781 = ~n10576 & ~n10780;
  assign n10782 = ~n10604 & n10781;
  assign n10783 = ~n10576 & ~n10604;
  assign n10784 = n10780 & ~n10783;
  assign n10785 = ~n10782 & ~n10784;
  assign n10786 = ~n10746 & n10785;
  assign n10787 = ~n10744 & ~n10785;
  assign n10788 = ~n10745 & n10787;
  assign n10789 = ~n10786 & ~n10788;
  assign n10790 = ~n10698 & n10789;
  assign n10791 = n10698 & ~n10789;
  assign n10792 = ~n10790 & ~n10791;
  assign n10793 = ~n10689 & n10792;
  assign n10794 = ~n10685 & ~n10792;
  assign n10795 = ~n10688 & n10794;
  assign n10796 = ~n10793 & ~n10795;
  assign n10797 = ~n10684 & ~n10796;
  assign n10798 = ~n10662 & n10796;
  assign n10799 = ~n10683 & n10798;
  assign po52 = ~n10797 & ~n10799;
  assign n10801 = n5172 & n7172;
  assign n10802 = ~n4549 & n10642;
  assign n10803 = n10801 & n10802;
  assign n10804 = n6126 & n10803;
  assign n10805 = n7500 & n7502;
  assign n10806 = n10804 & n10805;
  assign n10807 = n10329 & n10333;
  assign n10808 = n10332 & n10807;
  assign n10809 = n8660 & n10675;
  assign n10810 = n10663 & n10809;
  assign n10811 = ~n4853 & ~n8346;
  assign n10812 = n8928 & n10811;
  assign n10813 = n9617 & n10812;
  assign n10814 = n10810 & n10813;
  assign n10815 = n10808 & n10814;
  assign n10816 = n10806 & n10815;
  assign n10817 = ~n4273 & n10816;
  assign n10818 = n9619 & n10642;
  assign n10819 = n10503 & n10818;
  assign n10820 = ~n8364 & n10819;
  assign n10821 = ~n6419 & n10642;
  assign n10822 = n10663 & n10821;
  assign n10823 = n10667 & n10822;
  assign n10824 = n7500 & n10823;
  assign n10825 = n10503 & n10824;
  assign n10826 = ~n6138 & n10825;
  assign n10827 = n10493 & n10642;
  assign n10828 = n10492 & n10827;
  assign n10829 = ~n9795 & n10828;
  assign n10830 = ~n10650 & ~n10652;
  assign n10831 = ~n10829 & n10830;
  assign n10832 = ~n10826 & n10831;
  assign n10833 = ~n10820 & n10832;
  assign n10834 = ~n10817 & n10833;
  assign n10835 = ~n10795 & ~n10834;
  assign n10836 = ~n10793 & ~n10835;
  assign n10837 = n10554 & ~n10606;
  assign n10838 = ~n10608 & n10837;
  assign n10839 = ~n10560 & n10838;
  assign n10840 = ~n10790 & ~n10839;
  assign n10841 = n10740 & ~n10786;
  assign n10842 = ~n10601 & ~n10740;
  assign n10843 = ~n10742 & n10842;
  assign n10844 = n10605 & n10843;
  assign n10845 = ~n10740 & ~n10782;
  assign n10846 = ~n10784 & n10845;
  assign n10847 = ~n10746 & n10846;
  assign n10848 = ~n10844 & ~n10847;
  assign n10849 = ~n10841 & n10848;
  assign n10850 = ~n10710 & ~n10719;
  assign n10851 = ~n10717 & n10850;
  assign n10852 = ~n10708 & n10851;
  assign n10853 = ~n10733 & ~n10852;
  assign n10854 = pi22 & ~n5091;
  assign n10855 = ~n5092 & n10854;
  assign n10856 = ~n5178 & n10855;
  assign n10857 = pi23 & ~n5093;
  assign n10858 = ~n10856 & ~n10857;
  assign n10859 = pi63 & ~n10858;
  assign n10860 = ~pi63 & ~n10857;
  assign n10861 = ~n10856 & n10860;
  assign n10862 = ~n10859 & ~n10861;
  assign n10863 = pi24 & ~n4513;
  assign n10864 = ~n4514 & n10863;
  assign n10865 = ~n4577 & n10864;
  assign n10866 = pi25 & ~n4515;
  assign n10867 = ~n10865 & ~n10866;
  assign n10868 = pi61 & ~n10867;
  assign n10869 = ~pi61 & ~n10866;
  assign n10870 = ~n10865 & n10869;
  assign n10871 = ~n10868 & ~n10870;
  assign n10872 = ~n10862 & n10871;
  assign n10873 = n10862 & ~n10871;
  assign n10874 = ~n10872 & ~n10873;
  assign n10875 = pi26 & ~n3959;
  assign n10876 = ~n3960 & n10875;
  assign n10877 = ~n4233 & n10876;
  assign n10878 = pi27 & ~n3961;
  assign n10879 = ~n10877 & ~n10878;
  assign n10880 = pi59 & ~n10879;
  assign n10881 = ~pi59 & ~n10878;
  assign n10882 = ~n10877 & n10881;
  assign n10883 = ~n10880 & ~n10882;
  assign n10884 = ~n10874 & n10883;
  assign n10885 = ~n10872 & ~n10883;
  assign n10886 = ~n10873 & n10885;
  assign n10887 = ~n10884 & ~n10886;
  assign n10888 = n10853 & ~n10887;
  assign n10889 = ~n10853 & n10887;
  assign n10890 = n10738 & ~n10889;
  assign n10891 = ~n10888 & n10890;
  assign n10892 = ~n10888 & ~n10889;
  assign n10893 = ~n10738 & ~n10892;
  assign n10894 = ~n10891 & ~n10893;
  assign n10895 = n10784 & ~n10894;
  assign n10896 = ~n10784 & n10894;
  assign n10897 = ~n10895 & ~n10896;
  assign n10898 = pi30 & ~n2876;
  assign n10899 = ~n2877 & n10898;
  assign n10900 = ~n2960 & n10899;
  assign n10901 = pi31 & ~n2878;
  assign n10902 = ~n10900 & ~n10901;
  assign n10903 = pi55 & ~n10902;
  assign n10904 = ~pi55 & ~n10901;
  assign n10905 = ~n10900 & n10904;
  assign n10906 = ~n10903 & ~n10905;
  assign n10907 = pi28 & ~n3205;
  assign n10908 = ~n3206 & n10907;
  assign n10909 = ~n3463 & n10908;
  assign n10910 = pi29 & ~n3207;
  assign n10911 = ~n10909 & ~n10910;
  assign n10912 = pi57 & ~n10911;
  assign n10913 = ~pi57 & ~n10910;
  assign n10914 = ~n10909 & n10913;
  assign n10915 = ~n10912 & ~n10914;
  assign n10916 = n10773 & ~n10915;
  assign n10917 = ~n10773 & n10915;
  assign n10918 = ~n10916 & ~n10917;
  assign n10919 = ~n10906 & ~n10918;
  assign n10920 = n10906 & ~n10916;
  assign n10921 = ~n10917 & n10920;
  assign n10922 = ~n10919 & ~n10921;
  assign n10923 = ~n10756 & ~n10777;
  assign n10924 = ~n10922 & n10923;
  assign n10925 = n10922 & ~n10923;
  assign n10926 = ~n10924 & ~n10925;
  assign n10927 = ~n10897 & n10926;
  assign n10928 = ~n10895 & ~n10926;
  assign n10929 = ~n10896 & n10928;
  assign n10930 = ~n10927 & ~n10929;
  assign n10931 = ~n10849 & n10930;
  assign n10932 = n10848 & ~n10930;
  assign n10933 = ~n10841 & n10932;
  assign n10934 = ~n10931 & ~n10933;
  assign n10935 = ~n10840 & n10934;
  assign n10936 = n10840 & ~n10934;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = ~n10836 & n10937;
  assign n10939 = ~n10793 & ~n10937;
  assign n10940 = ~n10835 & n10939;
  assign po53 = ~n10938 & ~n10940;
  assign n10942 = ~n10793 & n10937;
  assign n10943 = ~n10795 & n10942;
  assign n10944 = ~n10310 & n10943;
  assign n10945 = n10649 & n10944;
  assign n10946 = n10310 & n10642;
  assign n10947 = ~n10652 & ~n10946;
  assign n10948 = n10796 & ~n10947;
  assign n10949 = ~n10485 & ~n10632;
  assign n10950 = ~n10636 & n10949;
  assign n10951 = n10148 & n10796;
  assign n10952 = ~n10150 & ~n10483;
  assign n10953 = n10951 & n10952;
  assign n10954 = n10314 & n10953;
  assign n10955 = n10950 & n10954;
  assign n10956 = ~n10793 & ~n10935;
  assign n10957 = ~n10955 & n10956;
  assign n10958 = ~n10948 & n10957;
  assign n10959 = ~n10936 & ~n10958;
  assign n10960 = ~n10945 & ~n10959;
  assign n10961 = ~n9995 & ~n9998;
  assign n10962 = ~n9991 & n10961;
  assign n10963 = ~n9986 & n10962;
  assign n10964 = n9956 & n10156;
  assign n10965 = ~n10963 & n10964;
  assign n10966 = ~n10342 & ~n10959;
  assign n10967 = ~n10965 & n10966;
  assign n10968 = ~n10960 & ~n10967;
  assign n10969 = ~n8050 & ~n10313;
  assign n10970 = n10156 & n10969;
  assign n10971 = n10495 & n10970;
  assign n10972 = n7490 & n7790;
  assign n10973 = n10642 & n10944;
  assign n10974 = n10972 & n10973;
  assign n10975 = n9184 & n9186;
  assign n10976 = n10974 & n10975;
  assign n10977 = n10971 & n10976;
  assign n10978 = ~n8649 & n10977;
  assign n10979 = ~n10968 & ~n10978;
  assign n10980 = n10891 & ~n10927;
  assign n10981 = n10784 & n10894;
  assign n10982 = ~n10891 & n10926;
  assign n10983 = ~n10897 & n10982;
  assign n10984 = ~n10981 & ~n10983;
  assign n10985 = ~n10980 & n10984;
  assign n10986 = ~n10861 & ~n10870;
  assign n10987 = ~n10868 & n10986;
  assign n10988 = ~n10859 & n10987;
  assign n10989 = ~n10884 & ~n10988;
  assign n10990 = pi23 & ~n5091;
  assign n10991 = ~n5092 & n10990;
  assign n10992 = ~n5178 & n10991;
  assign n10993 = pi24 & ~n5093;
  assign n10994 = ~n10992 & ~n10993;
  assign n10995 = pi63 & ~n10994;
  assign n10996 = ~pi63 & ~n10993;
  assign n10997 = ~n10992 & n10996;
  assign n10998 = ~n10995 & ~n10997;
  assign n10999 = pi25 & ~n4513;
  assign n11000 = ~n4514 & n10999;
  assign n11001 = ~n4577 & n11000;
  assign n11002 = pi26 & ~n4515;
  assign n11003 = ~n11001 & ~n11002;
  assign n11004 = pi61 & ~n11003;
  assign n11005 = ~pi61 & ~n11002;
  assign n11006 = ~n11001 & n11005;
  assign n11007 = ~n11004 & ~n11006;
  assign n11008 = ~n10998 & n11007;
  assign n11009 = n10998 & ~n11007;
  assign n11010 = ~n11008 & ~n11009;
  assign n11011 = pi27 & ~n3959;
  assign n11012 = ~n3960 & n11011;
  assign n11013 = ~n4233 & n11012;
  assign n11014 = pi28 & ~n3961;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = pi59 & ~n11015;
  assign n11017 = ~pi59 & ~n11014;
  assign n11018 = ~n11013 & n11017;
  assign n11019 = ~n11016 & ~n11018;
  assign n11020 = ~n11010 & n11019;
  assign n11021 = ~n11008 & ~n11019;
  assign n11022 = ~n11009 & n11021;
  assign n11023 = ~n11020 & ~n11022;
  assign n11024 = n10989 & ~n11023;
  assign n11025 = ~n10989 & n11023;
  assign n11026 = n10889 & ~n11025;
  assign n11027 = ~n11024 & n11026;
  assign n11028 = ~n11024 & ~n11025;
  assign n11029 = ~n10889 & ~n11028;
  assign n11030 = ~n11027 & ~n11029;
  assign n11031 = n10925 & ~n11030;
  assign n11032 = ~n10925 & ~n11027;
  assign n11033 = ~n11029 & n11032;
  assign n11034 = ~n11031 & ~n11033;
  assign n11035 = ~n10771 & ~n10914;
  assign n11036 = ~n10769 & n11035;
  assign n11037 = ~n10763 & ~n10912;
  assign n11038 = n11036 & n11037;
  assign n11039 = ~n10919 & ~n11038;
  assign n11040 = pi29 & ~n3205;
  assign n11041 = ~n3206 & n11040;
  assign n11042 = ~n3463 & n11041;
  assign n11043 = pi30 & ~n3207;
  assign n11044 = ~n11042 & ~n11043;
  assign n11045 = pi57 & ~n11044;
  assign n11046 = ~pi57 & ~n11043;
  assign n11047 = ~n11042 & n11046;
  assign n11048 = ~n11045 & ~n11047;
  assign n11049 = ~n10906 & n11048;
  assign n11050 = n10906 & ~n11048;
  assign n11051 = n2878 & n2960;
  assign n11052 = pi31 & pi55;
  assign n11053 = ~n11051 & n11052;
  assign n11054 = pi31 & ~n11051;
  assign n11055 = ~pi55 & ~n11054;
  assign n11056 = ~n11053 & ~n11055;
  assign n11057 = ~n11050 & n11056;
  assign n11058 = ~n11049 & n11057;
  assign n11059 = ~n11049 & ~n11050;
  assign n11060 = ~n11056 & ~n11059;
  assign n11061 = ~n11058 & ~n11060;
  assign n11062 = ~n11039 & n11061;
  assign n11063 = n11039 & ~n11061;
  assign n11064 = ~n11062 & ~n11063;
  assign n11065 = ~n11034 & n11064;
  assign n11066 = ~n11031 & ~n11064;
  assign n11067 = ~n11033 & n11066;
  assign n11068 = ~n11065 & ~n11067;
  assign n11069 = ~n10985 & n11068;
  assign n11070 = n10985 & ~n11068;
  assign n11071 = ~n11069 & ~n11070;
  assign n11072 = n10740 & ~n10782;
  assign n11073 = ~n10784 & n11072;
  assign n11074 = ~n10746 & n11073;
  assign n11075 = ~n10931 & ~n11074;
  assign n11076 = ~n11071 & n11075;
  assign n11077 = n11071 & ~n11075;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = ~n10979 & n11078;
  assign n11080 = ~n10978 & ~n11078;
  assign n11081 = ~n10968 & n11080;
  assign po54 = ~n11079 & ~n11081;
  assign n11083 = ~n10936 & ~n11076;
  assign n11084 = ~n10958 & n11083;
  assign n11085 = n10891 & n10926;
  assign n11086 = ~n10897 & n11085;
  assign n11087 = ~n11069 & ~n11086;
  assign n11088 = n11027 & ~n11065;
  assign n11089 = n10925 & ~n11027;
  assign n11090 = ~n11029 & n11089;
  assign n11091 = ~n11027 & n11064;
  assign n11092 = ~n11034 & n11091;
  assign n11093 = ~n11090 & ~n11092;
  assign n11094 = ~n11088 & n11093;
  assign n11095 = ~n10997 & ~n11006;
  assign n11096 = ~n11004 & n11095;
  assign n11097 = ~n10995 & n11096;
  assign n11098 = ~n11020 & ~n11097;
  assign n11099 = pi24 & ~n5091;
  assign n11100 = ~n5092 & n11099;
  assign n11101 = ~n5178 & n11100;
  assign n11102 = pi25 & ~n5093;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = pi63 & ~n11103;
  assign n11105 = ~pi63 & ~n11102;
  assign n11106 = ~n11101 & n11105;
  assign n11107 = ~n11104 & ~n11106;
  assign n11108 = pi26 & ~n4513;
  assign n11109 = ~n4514 & n11108;
  assign n11110 = ~n4577 & n11109;
  assign n11111 = pi27 & ~n4515;
  assign n11112 = ~n11110 & ~n11111;
  assign n11113 = pi61 & ~n11112;
  assign n11114 = ~pi61 & ~n11111;
  assign n11115 = ~n11110 & n11114;
  assign n11116 = ~n11113 & ~n11115;
  assign n11117 = ~n11107 & n11116;
  assign n11118 = n11107 & ~n11116;
  assign n11119 = ~n11117 & ~n11118;
  assign n11120 = pi28 & ~n3959;
  assign n11121 = ~n3960 & n11120;
  assign n11122 = ~n4233 & n11121;
  assign n11123 = pi29 & ~n3961;
  assign n11124 = ~n11122 & ~n11123;
  assign n11125 = pi59 & ~n11124;
  assign n11126 = ~pi59 & ~n11123;
  assign n11127 = ~n11122 & n11126;
  assign n11128 = ~n11125 & ~n11127;
  assign n11129 = ~n11119 & n11128;
  assign n11130 = ~n11117 & ~n11128;
  assign n11131 = ~n11118 & n11130;
  assign n11132 = ~n11129 & ~n11131;
  assign n11133 = n11098 & ~n11132;
  assign n11134 = ~n11098 & n11132;
  assign n11135 = n11025 & ~n11134;
  assign n11136 = ~n11133 & n11135;
  assign n11137 = ~n11133 & ~n11134;
  assign n11138 = ~n11025 & ~n11137;
  assign n11139 = ~n11136 & ~n11138;
  assign n11140 = n11062 & ~n11139;
  assign n11141 = ~n11062 & ~n11136;
  assign n11142 = ~n11138 & n11141;
  assign n11143 = ~n11140 & ~n11142;
  assign n11144 = ~n10905 & ~n11047;
  assign n11145 = ~n10903 & n11144;
  assign n11146 = ~n11045 & n11145;
  assign n11147 = pi30 & ~n3205;
  assign n11148 = ~n3206 & n11147;
  assign n11149 = ~n3463 & n11148;
  assign n11150 = pi31 & ~n3207;
  assign n11151 = ~n11149 & ~n11150;
  assign n11152 = pi57 & ~n11151;
  assign n11153 = ~pi57 & ~n11150;
  assign n11154 = ~n11149 & n11153;
  assign n11155 = ~n11152 & ~n11154;
  assign n11156 = ~n11146 & n11155;
  assign n11157 = ~n11060 & n11156;
  assign n11158 = ~n11060 & ~n11146;
  assign n11159 = ~n11155 & ~n11158;
  assign n11160 = ~n11157 & ~n11159;
  assign n11161 = ~n11143 & n11160;
  assign n11162 = ~n11140 & ~n11160;
  assign n11163 = ~n11142 & n11162;
  assign n11164 = ~n11161 & ~n11163;
  assign n11165 = ~n11094 & n11164;
  assign n11166 = n11094 & ~n11164;
  assign n11167 = ~n11165 & ~n11166;
  assign n11168 = ~n11087 & n11167;
  assign n11169 = n11087 & ~n11167;
  assign n11170 = ~n11168 & ~n11169;
  assign n11171 = ~n11077 & ~n11170;
  assign n11172 = ~n11084 & n11171;
  assign n11173 = ~n10173 & n11172;
  assign n11174 = ~n10935 & n11170;
  assign n11175 = ~n11077 & n11083;
  assign n11176 = n11174 & n11175;
  assign n11177 = n10796 & n11176;
  assign n11178 = ~n10310 & n11177;
  assign n11179 = n10649 & n11178;
  assign n11180 = ~n10172 & n11179;
  assign n11181 = ~n10164 & n11180;
  assign n11182 = ~n11077 & ~n11084;
  assign n11183 = n11170 & ~n11182;
  assign n11184 = n10937 & n11078;
  assign n11185 = ~n10793 & n11184;
  assign n11186 = ~n10795 & n11185;
  assign n11187 = ~n10310 & n11186;
  assign n11188 = n10649 & n11187;
  assign n11189 = n11171 & ~n11188;
  assign n11190 = ~n11084 & n11189;
  assign n11191 = ~n11183 & ~n11190;
  assign n11192 = ~n11181 & n11191;
  assign po55 = ~n11173 & n11192;
  assign n11194 = ~n10947 & n11177;
  assign n11195 = n10792 & ~n10935;
  assign n11196 = ~n10689 & n11195;
  assign n11197 = n11175 & n11196;
  assign n11198 = n10935 & ~n11076;
  assign n11199 = ~n11077 & ~n11168;
  assign n11200 = ~n11198 & n11199;
  assign n11201 = ~n11197 & n11200;
  assign n11202 = ~n11169 & ~n11201;
  assign n11203 = ~n11179 & ~n11202;
  assign n11204 = ~n11194 & n11203;
  assign n11205 = n9978 & n10170;
  assign n11206 = n9973 & n11205;
  assign n11207 = ~n10321 & n11206;
  assign n11208 = ~n8900 & ~n9194;
  assign n11209 = ~n10326 & n11208;
  assign n11210 = n9992 & n9993;
  assign n11211 = n10964 & n11210;
  assign n11212 = ~n11209 & n11211;
  assign n11213 = n9959 & n10168;
  assign n11214 = ~n9990 & n11213;
  assign n11215 = ~n10151 & ~n11202;
  assign n11216 = ~n10342 & n11215;
  assign n11217 = ~n11194 & n11216;
  assign n11218 = ~n11214 & n11217;
  assign n11219 = ~n11212 & n11218;
  assign n11220 = ~n11207 & n11219;
  assign n11221 = ~n11204 & ~n11220;
  assign n11222 = n11136 & ~n11161;
  assign n11223 = n11062 & ~n11136;
  assign n11224 = ~n11138 & n11223;
  assign n11225 = ~n11136 & n11160;
  assign n11226 = ~n11143 & n11225;
  assign n11227 = ~n11224 & ~n11226;
  assign n11228 = ~n11222 & n11227;
  assign n11229 = ~n11106 & ~n11115;
  assign n11230 = ~n11113 & n11229;
  assign n11231 = ~n11104 & n11230;
  assign n11232 = ~n11129 & ~n11231;
  assign n11233 = pi25 & ~n5091;
  assign n11234 = ~n5092 & n11233;
  assign n11235 = ~n5178 & n11234;
  assign n11236 = pi26 & ~n5093;
  assign n11237 = ~n11235 & ~n11236;
  assign n11238 = pi63 & ~n11237;
  assign n11239 = ~pi63 & ~n11236;
  assign n11240 = ~n11235 & n11239;
  assign n11241 = ~n11238 & ~n11240;
  assign n11242 = pi27 & ~n4513;
  assign n11243 = ~n4514 & n11242;
  assign n11244 = ~n4577 & n11243;
  assign n11245 = pi28 & ~n4515;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = pi61 & ~n11246;
  assign n11248 = ~pi61 & ~n11245;
  assign n11249 = ~n11244 & n11248;
  assign n11250 = ~n11247 & ~n11249;
  assign n11251 = ~n11241 & n11250;
  assign n11252 = n11241 & ~n11250;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = pi29 & ~n3959;
  assign n11255 = ~n3960 & n11254;
  assign n11256 = ~n4233 & n11255;
  assign n11257 = pi30 & ~n3961;
  assign n11258 = ~n11256 & ~n11257;
  assign n11259 = pi59 & ~n11258;
  assign n11260 = ~pi59 & ~n11257;
  assign n11261 = ~n11256 & n11260;
  assign n11262 = ~n11259 & ~n11261;
  assign n11263 = ~n11253 & n11262;
  assign n11264 = ~n11251 & ~n11262;
  assign n11265 = ~n11252 & n11264;
  assign n11266 = ~n11263 & ~n11265;
  assign n11267 = n11232 & ~n11266;
  assign n11268 = ~n11232 & n11266;
  assign n11269 = n11134 & ~n11268;
  assign n11270 = ~n11267 & n11269;
  assign n11271 = ~n11267 & ~n11268;
  assign n11272 = ~n11134 & ~n11271;
  assign n11273 = ~n11270 & ~n11272;
  assign n11274 = n11159 & ~n11273;
  assign n11275 = ~n11159 & ~n11270;
  assign n11276 = ~n11272 & n11275;
  assign n11277 = ~n11274 & ~n11276;
  assign n11278 = n3207 & n3463;
  assign n11279 = pi31 & pi57;
  assign n11280 = ~n11278 & n11279;
  assign n11281 = pi31 & ~n11278;
  assign n11282 = ~pi57 & ~n11281;
  assign n11283 = ~n11280 & ~n11282;
  assign n11284 = n11155 & ~n11283;
  assign n11285 = ~n11155 & n11283;
  assign n11286 = ~n11284 & ~n11285;
  assign n11287 = ~n11277 & n11286;
  assign n11288 = ~n11274 & ~n11286;
  assign n11289 = ~n11276 & n11288;
  assign n11290 = ~n11287 & ~n11289;
  assign n11291 = ~n11228 & n11290;
  assign n11292 = n11228 & ~n11290;
  assign n11293 = ~n11291 & ~n11292;
  assign n11294 = n11027 & n11064;
  assign n11295 = ~n11034 & n11294;
  assign n11296 = ~n11165 & ~n11295;
  assign n11297 = ~n11293 & n11296;
  assign n11298 = n11293 & ~n11296;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = ~n11221 & ~n11299;
  assign n11301 = ~n11204 & n11299;
  assign n11302 = ~n11220 & n11301;
  assign po56 = ~n11300 & ~n11302;
  assign n11304 = n11170 & ~n11297;
  assign n11305 = n11184 & n11304;
  assign n11306 = n10796 & n11305;
  assign n11307 = n10642 & n11306;
  assign n11308 = ~n10506 & n11307;
  assign n11309 = ~n10501 & n11308;
  assign n11310 = n10652 & n11177;
  assign n11311 = ~n11202 & ~n11310;
  assign n11312 = ~n11297 & ~n11311;
  assign n11313 = ~n11298 & ~n11312;
  assign n11314 = ~n11309 & n11313;
  assign n11315 = n11136 & n11160;
  assign n11316 = ~n11143 & n11315;
  assign n11317 = ~n11291 & ~n11316;
  assign n11318 = n11270 & ~n11287;
  assign n11319 = ~n11270 & n11286;
  assign n11320 = ~n11277 & n11319;
  assign n11321 = n11159 & ~n11270;
  assign n11322 = ~n11272 & n11321;
  assign n11323 = ~n11240 & ~n11249;
  assign n11324 = ~n11247 & n11323;
  assign n11325 = ~n11238 & n11324;
  assign n11326 = ~n11263 & ~n11325;
  assign n11327 = pi26 & ~n5091;
  assign n11328 = ~n5092 & n11327;
  assign n11329 = ~n5178 & n11328;
  assign n11330 = pi27 & ~n5093;
  assign n11331 = ~n11329 & ~n11330;
  assign n11332 = pi63 & ~n11331;
  assign n11333 = ~pi63 & ~n11330;
  assign n11334 = ~n11329 & n11333;
  assign n11335 = ~n11332 & ~n11334;
  assign n11336 = pi28 & ~n4513;
  assign n11337 = ~n4514 & n11336;
  assign n11338 = ~n4577 & n11337;
  assign n11339 = pi29 & ~n4515;
  assign n11340 = ~n11338 & ~n11339;
  assign n11341 = pi61 & ~n11340;
  assign n11342 = ~pi61 & ~n11339;
  assign n11343 = ~n11338 & n11342;
  assign n11344 = ~n11341 & ~n11343;
  assign n11345 = ~n11335 & n11344;
  assign n11346 = n11335 & ~n11344;
  assign n11347 = ~n11345 & ~n11346;
  assign n11348 = pi30 & ~n3959;
  assign n11349 = ~n3960 & n11348;
  assign n11350 = ~n4233 & n11349;
  assign n11351 = pi31 & ~n3961;
  assign n11352 = ~n11350 & ~n11351;
  assign n11353 = pi59 & ~n11352;
  assign n11354 = ~pi59 & ~n11351;
  assign n11355 = ~n11350 & n11354;
  assign n11356 = ~n11353 & ~n11355;
  assign n11357 = ~n11347 & n11356;
  assign n11358 = ~n11345 & ~n11356;
  assign n11359 = ~n11346 & n11358;
  assign n11360 = ~n11357 & ~n11359;
  assign n11361 = n11326 & ~n11360;
  assign n11362 = ~n11326 & n11360;
  assign n11363 = n11268 & ~n11362;
  assign n11364 = ~n11361 & n11363;
  assign n11365 = ~n11361 & ~n11362;
  assign n11366 = ~n11268 & ~n11365;
  assign n11367 = ~n11364 & ~n11366;
  assign n11368 = n11284 & ~n11367;
  assign n11369 = ~n11284 & ~n11364;
  assign n11370 = ~n11366 & n11369;
  assign n11371 = ~n11368 & ~n11370;
  assign n11372 = ~n11322 & ~n11371;
  assign n11373 = ~n11320 & n11372;
  assign n11374 = ~n11318 & n11373;
  assign n11375 = ~n11320 & ~n11322;
  assign n11376 = ~n11318 & n11375;
  assign n11377 = n11371 & ~n11376;
  assign n11378 = ~n11374 & ~n11377;
  assign n11379 = ~n11317 & n11378;
  assign n11380 = n11317 & ~n11378;
  assign n11381 = ~n11379 & ~n11380;
  assign n11382 = ~n11314 & n11381;
  assign n11383 = ~n11298 & ~n11381;
  assign n11384 = ~n11312 & n11383;
  assign n11385 = ~n11309 & n11384;
  assign po57 = ~n11382 & ~n11385;
  assign n11387 = ~n11169 & ~n11297;
  assign n11388 = ~n11298 & ~n11379;
  assign n11389 = ~n11380 & n11388;
  assign n11390 = n11387 & n11389;
  assign n11391 = ~n11201 & n11390;
  assign n11392 = n11299 & n11381;
  assign n11393 = ~n11380 & ~n11388;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = ~n11391 & n11394;
  assign n11396 = n7180 & n10972;
  assign n11397 = n10975 & n11396;
  assign n11398 = ~n6100 & n10642;
  assign n11399 = ~n6101 & n11178;
  assign n11400 = n11398 & n11399;
  assign n11401 = n7500 & n11400;
  assign n11402 = n11397 & n11401;
  assign n11403 = n10971 & n11402;
  assign n11404 = ~n8077 & n11403;
  assign n11405 = ~n10660 & n11177;
  assign n11406 = ~n10655 & n11405;
  assign n11407 = n10649 & n10807;
  assign n11408 = ~n8346 & ~n10151;
  assign n11409 = n9185 & n10675;
  assign n11410 = n11408 & n11409;
  assign n11411 = n8928 & n11178;
  assign n11412 = n9617 & n11411;
  assign n11413 = n11410 & n11412;
  assign n11414 = n11407 & n11413;
  assign n11415 = ~n10674 & n11414;
  assign n11416 = ~n11391 & ~n11393;
  assign n11417 = ~n11415 & n11416;
  assign n11418 = ~n11406 & n11417;
  assign n11419 = ~n11404 & n11418;
  assign n11420 = ~n11395 & ~n11419;
  assign n11421 = ~n11129 & n11286;
  assign n11422 = ~n11131 & n11421;
  assign n11423 = ~n11098 & n11422;
  assign n11424 = n11271 & n11423;
  assign n11425 = ~n11277 & n11424;
  assign n11426 = ~n11377 & ~n11425;
  assign n11427 = ~n11263 & n11284;
  assign n11428 = ~n11265 & n11427;
  assign n11429 = ~n11232 & n11428;
  assign n11430 = n11365 & n11429;
  assign n11431 = ~n11268 & ~n11284;
  assign n11432 = ~n11365 & n11431;
  assign n11433 = ~n11430 & ~n11432;
  assign n11434 = ~n11334 & ~n11343;
  assign n11435 = ~n11341 & n11434;
  assign n11436 = ~n11332 & n11435;
  assign n11437 = ~n11357 & ~n11436;
  assign n11438 = pi27 & ~n5091;
  assign n11439 = ~n5092 & n11438;
  assign n11440 = ~n5178 & n11439;
  assign n11441 = pi28 & ~n5093;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 = pi63 & ~n11442;
  assign n11444 = ~pi63 & ~n11441;
  assign n11445 = ~n11440 & n11444;
  assign n11446 = ~n11443 & ~n11445;
  assign n11447 = pi29 & ~n4513;
  assign n11448 = ~n4514 & n11447;
  assign n11449 = ~n4577 & n11448;
  assign n11450 = pi30 & ~n4515;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = pi61 & ~n11451;
  assign n11453 = ~pi61 & ~n11450;
  assign n11454 = ~n11449 & n11453;
  assign n11455 = ~n11452 & ~n11454;
  assign n11456 = ~n11446 & n11455;
  assign n11457 = n11446 & ~n11455;
  assign n11458 = ~n11456 & ~n11457;
  assign n11459 = n3961 & n4233;
  assign n11460 = pi31 & pi59;
  assign n11461 = ~n11459 & n11460;
  assign n11462 = pi31 & ~n11459;
  assign n11463 = ~pi59 & ~n11462;
  assign n11464 = ~n11461 & ~n11463;
  assign n11465 = ~n11458 & ~n11464;
  assign n11466 = ~n11456 & n11464;
  assign n11467 = ~n11457 & n11466;
  assign n11468 = ~n11465 & ~n11467;
  assign n11469 = n11437 & ~n11468;
  assign n11470 = ~n11437 & n11468;
  assign n11471 = n11362 & ~n11470;
  assign n11472 = ~n11469 & n11471;
  assign n11473 = ~n11469 & ~n11470;
  assign n11474 = ~n11362 & ~n11473;
  assign n11475 = ~n11472 & ~n11474;
  assign n11476 = ~n11433 & n11475;
  assign n11477 = n11433 & ~n11475;
  assign n11478 = ~n11476 & ~n11477;
  assign n11479 = ~n11426 & ~n11478;
  assign n11480 = ~n11425 & n11478;
  assign n11481 = ~n11377 & n11480;
  assign n11482 = ~n11479 & ~n11481;
  assign n11483 = ~n11420 & ~n11482;
  assign n11484 = ~n11395 & n11482;
  assign n11485 = ~n11419 & n11484;
  assign po58 = ~n11483 & ~n11485;
  assign n11487 = n11174 & n11392;
  assign n11488 = n11175 & n11487;
  assign n11489 = n10796 & n11488;
  assign n11490 = ~n11393 & ~n11489;
  assign n11491 = ~n11391 & n11490;
  assign n11492 = ~n10652 & n11416;
  assign n11493 = ~n10650 & n11492;
  assign n11494 = ~n10829 & n11493;
  assign n11495 = ~n10826 & n11494;
  assign n11496 = ~n10820 & n11495;
  assign n11497 = ~n10817 & n11496;
  assign n11498 = ~n11491 & ~n11497;
  assign n11499 = ~n11470 & ~n11472;
  assign n11500 = ~n11445 & ~n11454;
  assign n11501 = ~n11452 & n11500;
  assign n11502 = ~n11443 & n11501;
  assign n11503 = ~n11465 & ~n11502;
  assign n11504 = pi30 & ~n4513;
  assign n11505 = ~n4514 & n11504;
  assign n11506 = ~n4577 & n11505;
  assign n11507 = pi31 & ~n4515;
  assign n11508 = ~n11506 & ~n11507;
  assign n11509 = pi61 & ~n11508;
  assign n11510 = pi28 & ~n5091;
  assign n11511 = ~n5092 & n11510;
  assign n11512 = ~n5178 & n11511;
  assign n11513 = pi29 & ~n5093;
  assign n11514 = ~n11512 & ~n11513;
  assign n11515 = pi63 & ~n11514;
  assign n11516 = ~pi63 & ~n11513;
  assign n11517 = ~n11512 & n11516;
  assign n11518 = ~pi61 & ~n11507;
  assign n11519 = ~n11506 & n11518;
  assign n11520 = ~n11517 & ~n11519;
  assign n11521 = ~n11515 & n11520;
  assign n11522 = ~n11509 & n11521;
  assign n11523 = ~n11515 & ~n11517;
  assign n11524 = ~n11509 & ~n11519;
  assign n11525 = ~n11523 & ~n11524;
  assign n11526 = ~n11522 & ~n11525;
  assign n11527 = ~n11503 & ~n11526;
  assign n11528 = ~n11502 & ~n11522;
  assign n11529 = ~n11525 & n11528;
  assign n11530 = ~n11465 & n11529;
  assign n11531 = ~n11527 & ~n11530;
  assign n11532 = ~n11499 & n11531;
  assign n11533 = ~n11470 & ~n11531;
  assign n11534 = ~n11472 & n11533;
  assign n11535 = ~n11532 & ~n11534;
  assign n11536 = n11433 & n11475;
  assign n11537 = ~n11430 & ~n11536;
  assign n11538 = ~n11535 & n11537;
  assign n11539 = n11535 & ~n11537;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = ~n11479 & ~n11540;
  assign n11542 = ~n11498 & n11541;
  assign n11543 = ~n11481 & n11540;
  assign n11544 = ~n11491 & n11543;
  assign n11545 = ~n11497 & n11544;
  assign n11546 = n11480 & ~n11540;
  assign n11547 = ~n11377 & n11546;
  assign n11548 = ~n11479 & n11547;
  assign n11549 = ~n11478 & ~n11538;
  assign n11550 = ~n11539 & n11549;
  assign n11551 = ~n11426 & n11550;
  assign n11552 = ~n11548 & ~n11551;
  assign n11553 = ~n11545 & n11552;
  assign po59 = ~n11542 & n11553;
  assign n11555 = ~n11380 & ~n11479;
  assign n11556 = n11388 & n11555;
  assign n11557 = n11470 & n11531;
  assign n11558 = ~n11527 & ~n11557;
  assign n11559 = n4515 & n4577;
  assign n11560 = pi31 & pi61;
  assign n11561 = ~n11559 & n11560;
  assign n11562 = pi31 & ~n11559;
  assign n11563 = ~pi61 & ~n11562;
  assign n11564 = ~n11561 & ~n11563;
  assign n11565 = pi29 & ~n5091;
  assign n11566 = ~n5092 & n11565;
  assign n11567 = ~n5178 & n11566;
  assign n11568 = pi30 & ~n5093;
  assign n11569 = ~n11567 & ~n11568;
  assign n11570 = pi63 & ~n11569;
  assign n11571 = ~pi63 & ~n11568;
  assign n11572 = ~n11567 & n11571;
  assign n11573 = ~n11570 & ~n11572;
  assign n11574 = ~n11564 & n11573;
  assign n11575 = n11564 & ~n11573;
  assign n11576 = ~n11574 & ~n11575;
  assign n11577 = n11525 & ~n11576;
  assign n11578 = ~n11525 & ~n11574;
  assign n11579 = ~n11575 & n11578;
  assign n11580 = ~n11577 & ~n11579;
  assign n11581 = ~n11558 & n11580;
  assign n11582 = ~n11527 & ~n11580;
  assign n11583 = ~n11557 & n11582;
  assign n11584 = n11362 & n11473;
  assign n11585 = n11531 & n11584;
  assign n11586 = ~n11583 & n11585;
  assign n11587 = ~n11581 & n11586;
  assign n11588 = ~n11581 & ~n11583;
  assign n11589 = ~n11585 & ~n11588;
  assign n11590 = ~n11587 & ~n11589;
  assign n11591 = n11540 & n11590;
  assign n11592 = ~n11481 & n11591;
  assign n11593 = ~n11168 & n11592;
  assign n11594 = n11387 & n11593;
  assign n11595 = n11078 & n11594;
  assign n11596 = n11556 & n11595;
  assign n11597 = ~n10979 & n11596;
  assign n11598 = n11381 & ~n11479;
  assign n11599 = ~n11169 & n11543;
  assign n11600 = n11299 & n11599;
  assign n11601 = n11598 & n11600;
  assign n11602 = ~n11199 & n11601;
  assign n11603 = ~n11393 & ~n11479;
  assign n11604 = n11543 & ~n11603;
  assign n11605 = ~n11539 & ~n11590;
  assign n11606 = ~n11604 & n11605;
  assign n11607 = ~n11602 & n11606;
  assign n11608 = ~n10978 & n11607;
  assign n11609 = ~n10968 & n11608;
  assign n11610 = ~n11539 & ~n11604;
  assign n11611 = ~n11602 & n11610;
  assign n11612 = n11590 & ~n11611;
  assign n11613 = ~n11168 & ~n11297;
  assign n11614 = n11599 & n11613;
  assign n11615 = n11078 & n11614;
  assign n11616 = n11556 & n11615;
  assign n11617 = ~n11602 & ~n11616;
  assign n11618 = n11606 & n11617;
  assign n11619 = ~n11612 & ~n11618;
  assign n11620 = ~n11609 & n11619;
  assign po60 = ~n11597 & n11620;
  assign n11622 = n11556 & n11614;
  assign n11623 = n11184 & n11622;
  assign n11624 = n10796 & n11623;
  assign n11625 = ~n9156 & n11624;
  assign n11626 = n10165 & n11625;
  assign n11627 = n10494 & n11626;
  assign n11628 = n10828 & n11627;
  assign n11629 = n11610 & n11617;
  assign n11630 = ~n9954 & ~n10313;
  assign n11631 = n10156 & n11630;
  assign n11632 = n10973 & n11631;
  assign n11633 = ~n10160 & n11632;
  assign n11634 = ~n10959 & n11611;
  assign n11635 = ~n11633 & n11634;
  assign n11636 = ~n11629 & ~n11635;
  assign n11637 = ~n11628 & ~n11636;
  assign n11638 = n8939 & ~n11636;
  assign n11639 = ~n11637 & ~n11638;
  assign n11640 = ~n11574 & ~n11579;
  assign n11641 = pi30 & ~n5091;
  assign n11642 = ~n5092 & n11641;
  assign n11643 = ~n5178 & n11642;
  assign n11644 = pi31 & ~n5093;
  assign n11645 = ~n11643 & ~n11644;
  assign n11646 = pi63 & ~n11645;
  assign n11647 = ~pi63 & ~n11644;
  assign n11648 = ~n11643 & n11647;
  assign n11649 = ~n11646 & ~n11648;
  assign n11650 = ~n11640 & n11649;
  assign n11651 = ~n11526 & ~n11577;
  assign n11652 = ~n11579 & n11651;
  assign n11653 = ~n11574 & ~n11649;
  assign n11654 = ~n11579 & n11653;
  assign n11655 = ~n11503 & ~n11654;
  assign n11656 = n11652 & n11655;
  assign n11657 = ~n11650 & n11656;
  assign n11658 = ~n11503 & n11652;
  assign n11659 = ~n11650 & ~n11654;
  assign n11660 = ~n11658 & ~n11659;
  assign n11661 = ~n11657 & ~n11660;
  assign n11662 = n11468 & n11580;
  assign n11663 = ~n11437 & ~n11530;
  assign n11664 = n11662 & n11663;
  assign n11665 = ~n11527 & n11664;
  assign n11666 = ~n11661 & ~n11665;
  assign n11667 = ~n11657 & n11665;
  assign n11668 = ~n11660 & n11667;
  assign n11669 = ~n11666 & ~n11668;
  assign n11670 = ~n11587 & n11669;
  assign n11671 = ~n11639 & n11670;
  assign n11672 = ~n11589 & ~n11669;
  assign n11673 = ~n11637 & n11672;
  assign n11674 = ~n11638 & n11673;
  assign n11675 = ~n11585 & ~n11666;
  assign n11676 = ~n11668 & n11675;
  assign n11677 = ~n11587 & ~n11588;
  assign n11678 = n11676 & n11677;
  assign n11679 = n11587 & ~n11669;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = ~n11674 & n11680;
  assign po61 = ~n11671 & n11681;
  assign n11683 = ~n11539 & ~n11587;
  assign n11684 = ~n11604 & n11683;
  assign n11685 = n11672 & ~n11684;
  assign n11686 = ~n11661 & n11665;
  assign n11687 = ~n11525 & ~n11575;
  assign n11688 = n11653 & n11687;
  assign n11689 = n11658 & ~n11659;
  assign n11690 = ~n11688 & ~n11689;
  assign n11691 = n5093 & n5178;
  assign n11692 = pi31 & pi63;
  assign n11693 = ~n11691 & n11692;
  assign n11694 = pi31 & ~n11691;
  assign n11695 = ~pi63 & ~n11694;
  assign n11696 = ~n11693 & ~n11695;
  assign n11697 = ~n11653 & ~n11696;
  assign n11698 = ~n11649 & n11696;
  assign n11699 = ~n11574 & n11698;
  assign n11700 = ~n11697 & ~n11699;
  assign n11701 = ~n11690 & n11700;
  assign n11702 = ~n11688 & ~n11700;
  assign n11703 = ~n11689 & n11702;
  assign n11704 = ~n11701 & ~n11703;
  assign n11705 = ~n11686 & ~n11704;
  assign n11706 = ~n11685 & n11705;
  assign n11707 = ~n11221 & n11706;
  assign n11708 = ~n11587 & n11704;
  assign n11709 = n11540 & n11708;
  assign n11710 = n11672 & n11709;
  assign n11711 = ~n11481 & n11710;
  assign n11712 = ~n11297 & n11711;
  assign n11713 = n11556 & n11712;
  assign n11714 = ~n11204 & n11713;
  assign n11715 = ~n11220 & n11714;
  assign n11716 = ~n11685 & ~n11686;
  assign n11717 = n11704 & ~n11716;
  assign n11718 = ~n11587 & ~n11669;
  assign n11719 = ~n11538 & n11718;
  assign n11720 = ~n11539 & ~n11589;
  assign n11721 = n11719 & n11720;
  assign n11722 = ~n11481 & n11721;
  assign n11723 = ~n11297 & n11722;
  assign n11724 = n11556 & n11723;
  assign n11725 = n11705 & ~n11724;
  assign n11726 = ~n11685 & n11725;
  assign n11727 = ~n11717 & ~n11726;
  assign n11728 = ~n11715 & n11727;
  assign po62 = ~n11707 & n11728;
  assign n11730 = ~n11690 & ~n11699;
  assign n11731 = ~n11697 & ~n11730;
  assign n11732 = ~n11704 & n11731;
  assign n11733 = n10642 & n11177;
  assign n11734 = ~n10506 & n11733;
  assign n11735 = ~n10501 & n11734;
  assign n11736 = n11311 & ~n11735;
  assign n11737 = n11724 & ~n11736;
  assign n11738 = ~n11686 & n11731;
  assign n11739 = ~n11685 & n11738;
  assign n11740 = ~n11737 & n11739;
  assign po63 = n11732 | n11740;
endmodule


