module tv80 ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319,
    pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329,
    pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339,
    pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369,
    pi370, pi371, pi372,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318,
    pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328,
    pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338,
    pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348,
    pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278, po279,
    po280, po281, po282, po283, po284, po285, po286, po287, po288, po289,
    po290, po291, po292, po293, po294, po295, po296, po297, po298, po299,
    po300, po301, po302, po303, po304, po305, po306, po307, po308, po309,
    po310, po311, po312, po313, po314, po315, po316, po317, po318, po319,
    po320, po321, po322, po323, po324, po325, po326, po327, po328, po329,
    po330, po331, po332, po333, po334, po335, po336, po337, po338, po339,
    po340, po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368, po369,
    po370, po371, po372, po373, po374, po375, po376, po377, po378, po379,
    po380, po381, po382, po383, po384, po385, po386, po387, po388, po389,
    po390, po391, po392, po393, po394, po395, po396, po397, po398, po399,
    po400, po401, po402, po403;
  wire n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
    n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
    n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
    n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
    n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
    n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
    n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
    n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
    n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
    n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
    n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
    n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
    n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
    n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
    n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
    n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367, n3369, n3370, n3371, n3372,
    n3373, n3374, n3376, n3377, n3378, n3379, n3380, n3381, n3383, n3384,
    n3385, n3386, n3387, n3389, n3390, n3391, n3392, n3393, n3394, n3396,
    n3397, n3398, n3399, n3400, n3402, n3403, n3404, n3405, n3406, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3459,
    n3460, n3461, n3462, n3463, n3465, n3466, n3467, n3468, n3469, n3471,
    n3472, n3473, n3474, n3475, n3477, n3478, n3479, n3480, n3481, n3483,
    n3484, n3485, n3486, n3487, n3489, n3490, n3491, n3492, n3493, n3495,
    n3496, n3497, n3498, n3499, n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
    n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3551, n3552, n3553, n3554, n3555, n3557, n3558,
    n3559, n3560, n3561, n3563, n3564, n3565, n3566, n3567, n3569, n3570,
    n3571, n3572, n3573, n3575, n3576, n3577, n3578, n3579, n3581, n3582,
    n3583, n3584, n3585, n3587, n3588, n3589, n3590, n3591, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
    n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
    n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3665,
    n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
    n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
    n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
    n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
    n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
    n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
    n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4315,
    n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
    n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
    n4376, n4377, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4426, n4427,
    n4429, n4430, n4432, n4433, n4435, n4436, n4438, n4439, n4441, n4442,
    n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4513, n4514, n4515, n4516,
    n4517, n4519, n4520, n4521, n4522, n4523, n4524, n4526, n4527, n4528,
    n4529, n4530, n4532, n4533, n4534, n4535, n4536, n4538, n4539, n4540,
    n4541, n4542, n4543, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
    n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
    n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4603,
    n4604, n4605, n4606, n4607, n4609, n4610, n4611, n4612, n4613, n4615,
    n4616, n4617, n4618, n4619, n4621, n4622, n4623, n4624, n4625, n4627,
    n4628, n4629, n4630, n4631, n4633, n4634, n4635, n4636, n4637, n4639,
    n4640, n4641, n4642, n4643, n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
    n4691, n4692, n4693, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4728, n4729, n4730, n4731, n4732,
    n4734, n4735, n4736, n4737, n4738, n4740, n4741, n4742, n4743, n4744,
    n4746, n4747, n4748, n4749, n4750, n4752, n4753, n4754, n4755, n4756,
    n4758, n4759, n4760, n4761, n4762, n4764, n4765, n4766, n4767, n4768,
    n4770, n4771, n4772, n4773, n4774, n4776, n4777, n4778, n4779, n4780,
    n4782, n4783, n4784, n4785, n4786, n4788, n4789, n4790, n4791, n4792,
    n4794, n4795, n4796, n4797, n4798, n4800, n4801, n4802, n4803, n4804,
    n4806, n4807, n4808, n4809, n4810, n4812, n4813, n4814, n4815, n4816,
    n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4890, n4891, n4892, n4893, n4894, n4896, n4897, n4898, n4899,
    n4900, n4902, n4903, n4904, n4905, n4906, n4908, n4909, n4910, n4911,
    n4912, n4914, n4915, n4916, n4917, n4918, n4920, n4921, n4922, n4923,
    n4924, n4926, n4927, n4928, n4929, n4930, n4932, n4933, n4934, n4935,
    n4936, n4937, n4939, n4940, n4941, n4942, n4943, n4945, n4946, n4947,
    n4948, n4949, n4951, n4952, n4953, n4954, n4955, n4957, n4958, n4959,
    n4960, n4961, n4963, n4964, n4965, n4966, n4967, n4969, n4970, n4971,
    n4972, n4973, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
    n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
    n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
    n5087, n5088, n5089, n5090, n5091, n5092, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
    n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
    n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
    n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
    n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
    n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
    n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
    n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
    n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
    n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5308,
    n5309, n5310, n5311, n5312, n5314, n5315, n5316, n5317, n5318, n5320,
    n5321, n5322, n5323, n5324, n5326, n5327, n5328, n5329, n5330, n5332,
    n5333, n5334, n5335, n5336, n5338, n5339, n5340, n5341, n5342, n5344,
    n5345, n5346, n5347, n5348, n5350, n5351, n5352, n5353, n5354, n5356,
    n5357, n5358, n5359, n5360, n5362, n5363, n5364, n5365, n5366, n5368,
    n5369, n5370, n5371, n5372, n5374, n5375, n5376, n5377, n5378, n5380,
    n5381, n5382, n5383, n5384, n5386, n5387, n5388, n5389, n5390, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
    n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
    n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
    n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5582, n5583, n5584,
    n5585, n5586, n5588, n5589, n5590, n5591, n5592, n5594, n5595, n5596,
    n5597, n5598, n5600, n5601, n5602, n5603, n5604, n5606, n5607, n5608,
    n5609, n5610, n5612, n5613, n5614, n5615, n5616, n5618, n5619, n5620,
    n5621, n5622, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
    n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5715, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
    n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
    n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
    n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
    n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
    n6252, n6253, n6254, n6255, n6256, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6286, n6287, n6288, n6289, n6290, n6292, n6293, n6294,
    n6295, n6296, n6298, n6299, n6300, n6301, n6302, n6304, n6305, n6306,
    n6307, n6308, n6310, n6311, n6312, n6313, n6314, n6316, n6317, n6318,
    n6319, n6320, n6322, n6323, n6324, n6325, n6326, n6328, n6329, n6330,
    n6331, n6332, n6334, n6335, n6336, n6337, n6338, n6340, n6341, n6342,
    n6343, n6344, n6346, n6347, n6348, n6349, n6350, n6352, n6353, n6354,
    n6355, n6356, n6358, n6359, n6360, n6361, n6362, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6380, n6381, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
    n6419, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
    n6461, n6462, n6463, n6464, n6465, n6466, n6468, n6469, n6470, n6471,
    n6472, n6474, n6475, n6476, n6477, n6478, n6480, n6481, n6482, n6483,
    n6484, n6486, n6487, n6488, n6489, n6490, n6492, n6493, n6494, n6495,
    n6496, n6498, n6499, n6500, n6501, n6502, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
    n6528, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
    n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
    n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
    n6581, n6582, n6583, n6584, n6585, n6587, n6588, n6589, n6590, n6591,
    n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
    n6623, n6624, n6625, n6626, n6627, n6628, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
    n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
    n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
    n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
    n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6766,
    n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
    n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
    n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
    n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6837, n6838,
    n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
    n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6950, n6951,
    n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
    n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
    n6972, n6973, n6974, n6975, n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
    n7003, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7036, n7037, n7038, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
    n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
    n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
    n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
    n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
    n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
    n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
    n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
    n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826, n7828, n7829, n7830, n7831,
    n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
    n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7863, n7864, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
    n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
    n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
    n7934, n7935, n7936, n7937, n7938, n7939, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
    n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8056, n8057,
    n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
    n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
    n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
    n8088, n8089, n8090, n8091, n8092, n8093, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
    n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
    n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
    n8422, n8423, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8441, n8442, n8443,
    n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8543, n8544, n8545, n8546, n8547,
    n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
    n8558, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8594, n8595, n8596, n8597, n8598, n8600,
    n8601, n8603, n8604, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
    n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8623, n8624,
    n8625, n8626, n8627, n8629, n8630, n8631, n8632, n8633, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
    n8790, n8791, n8792, n8793, n8795, n8796, n8798, n8799, n8800, n8801,
    n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
    n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8820, n8821, n8822,
    n8823, n8824, n8826, n8827, n8829, n8830, n8832, n8833, n8835, n8836,
    n8837, n8838, n8840, n8842, n8843, n8845, n8846, n8848, n8849, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
    n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
    n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
    n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
    n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
    n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
    n8932, n8933, n8934, n8935, n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
    n9024, n9025, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9049, n9050, n9052, n9053, n9055, n9056, n9058,
    n9059, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
    n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
    n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
    n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
    n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
    n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
    n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
    n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
    n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
    n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
    n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
    n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
    n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
    n9250, n9251, n9252, n9253, n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9277, n9278, n9280, n9281, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9341, n9342, n9343, n9344, n9345, n9346,
    n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9383, n9384, n9385, n9386, n9387, n9388,
    n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9479, n9480, n9481, n9482, n9483, n9484,
    n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
    n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
    n9545, n9546, n9547, n9548, n9549, n9551, n9552, n9553, n9554, n9555,
    n9556, n9557, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9585, n9586, n9587, n9588,
    n9590, n9591, n9592, n9594, n9595, n9596, n9597, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
    n9622, n9623, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
    n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659, n9661, n9662, n9663, n9664,
    n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
    n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
    n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
    n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9737, n9738,
    n9739, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
    n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9760,
    n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9780, n9781,
    n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
    n9803, n9804, n9805, n9806, n9807, n9808, n9810, n9811, n9812, n9813,
    n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
    n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9840, n9841, n9842, n9843, n9844, n9845,
    n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9855, n9856,
    n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
    n9878, n9879, n9880, n9881, n9882, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9899,
    n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
    n9910, n9911, n9912, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
    n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
    n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
    n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10043, n10044, n10045, n10046, n10047, n10049,
    n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
    n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100, n10102, n10103, n10104,
    n10105, n10106, n10108, n10109, n10111, n10112, n10113, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121, n10123, n10124, n10125,
    n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10134, n10135,
    n10136, n10137, n10138, n10139, n10141, n10142, n10143, n10144, n10145,
    n10146, n10148, n10149, n10150, n10151, n10152, n10153, n10155, n10156,
    n10157, n10158, n10159, n10160, n10162, n10163, n10164, n10165, n10166,
    n10167, n10169, n10170, n10171, n10172, n10173, n10174, n10176, n10177,
    n10178, n10179, n10180, n10181, n10183, n10184, n10185, n10186, n10187,
    n10188, n10190, n10191, n10192, n10193, n10194, n10195, n10197, n10198,
    n10199, n10200, n10201, n10202, n10204, n10205, n10206, n10207, n10208,
    n10209, n10211, n10212, n10213, n10214, n10215, n10216, n10218, n10219,
    n10220, n10221, n10222, n10223, n10225, n10226, n10227, n10228, n10229,
    n10230, n10232, n10233, n10234, n10235, n10236, n10237, n10239, n10240,
    n10241, n10242, n10243, n10244, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10269,
    n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
    n10280, n10281, n10282, n10283, n10284, n10285, n10287, n10289, n10290,
    n10291, n10292, n10293, n10294, n10296, n10297, n10298, n10299, n10300,
    n10301, n10302, n10303, n10304, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10346, n10347, n10348, n10349, n10350,
    n10351, n10352, n10353, n10354, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10376, n10377, n10378, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387, n10389, n10390, n10391,
    n10392, n10393, n10395, n10396, n10398, n10399, n10401, n10402, n10404,
    n10405, n10407, n10408, n10410, n10411, n10413, n10414, n10416, n10417,
    n10419, n10420, n10421;
  assign n779 = ~pi189 & pi190;
  assign n780 = ~pi188 & n779;
  assign n781 = pi097 & pi098;
  assign n782 = ~pi099 & n781;
  assign n783 = n780 & n782;
  assign n784 = ~pi097 & pi098;
  assign n785 = ~pi099 & n784;
  assign n786 = ~n783 & ~n785;
  assign n787 = ~pi294 & ~pi301;
  assign n788 = pi188 & ~pi189;
  assign n789 = pi296 & ~pi297;
  assign n790 = pi300 & ~pi302;
  assign n791 = n789 & n790;
  assign n792 = ~pi298 & pi299;
  assign n793 = ~pi291 & pi303;
  assign n794 = n792 & n793;
  assign n795 = n791 & n794;
  assign n796 = ~pi297 & pi299;
  assign n797 = ~pi296 & pi300;
  assign n798 = ~pi291 & n797;
  assign n799 = n796 & n798;
  assign n800 = ~n795 & ~n799;
  assign n801 = n788 & ~n800;
  assign n802 = ~pi188 & pi189;
  assign n803 = ~pi190 & n802;
  assign n804 = pi190 & n788;
  assign n805 = ~n803 & ~n804;
  assign n806 = pi299 & n791;
  assign n807 = ~pi298 & pi303;
  assign n808 = pi291 & n807;
  assign n809 = n806 & n808;
  assign n810 = ~n805 & n809;
  assign n811 = ~pi190 & n788;
  assign n812 = ~n780 & ~n811;
  assign n813 = pi291 & pi299;
  assign n814 = ~pi297 & n813;
  assign n815 = pi296 & pi300;
  assign n816 = ~pi303 & n815;
  assign n817 = n814 & n816;
  assign n818 = ~n812 & n817;
  assign n819 = ~n810 & ~n818;
  assign n820 = ~pi300 & ~pi302;
  assign n821 = ~pi296 & ~pi297;
  assign n822 = ~pi298 & ~pi299;
  assign n823 = ~pi291 & ~pi303;
  assign n824 = n822 & n823;
  assign n825 = n821 & n824;
  assign n826 = n820 & n825;
  assign n827 = ~pi195 & ~pi196;
  assign n828 = ~n812 & ~n827;
  assign n829 = n826 & n828;
  assign n830 = pi297 & pi299;
  assign n831 = pi296 & n830;
  assign n832 = pi291 & pi300;
  assign n833 = n831 & n832;
  assign n834 = ~n812 & n833;
  assign n835 = ~n829 & ~n834;
  assign n836 = n819 & n835;
  assign n837 = pi291 & n797;
  assign n838 = n796 & n837;
  assign n839 = ~pi302 & pi303;
  assign n840 = ~pi298 & n839;
  assign n841 = pi131 & n840;
  assign n842 = pi298 & n839;
  assign n843 = pi102 & n842;
  assign n844 = pi302 & pi303;
  assign n845 = ~pi298 & n844;
  assign n846 = pi132 & n845;
  assign n847 = ~n843 & ~n846;
  assign n848 = ~n841 & n847;
  assign n849 = pi298 & pi302;
  assign n850 = ~pi303 & n849;
  assign n851 = ~pi178 & n850;
  assign n852 = ~pi302 & ~pi303;
  assign n853 = pi298 & n852;
  assign n854 = ~pi102 & n853;
  assign n855 = ~n851 & ~n854;
  assign n856 = n848 & n855;
  assign n857 = ~pi298 & n852;
  assign n858 = ~pi131 & n857;
  assign n859 = pi303 & n849;
  assign n860 = pi178 & n859;
  assign n861 = ~n858 & ~n860;
  assign n862 = pi302 & ~pi303;
  assign n863 = ~pi298 & n862;
  assign n864 = ~pi132 & n863;
  assign n865 = n861 & ~n864;
  assign n866 = n856 & n865;
  assign n867 = n804 & ~n866;
  assign n868 = ~n803 & ~n867;
  assign n869 = n838 & ~n868;
  assign n870 = ~pi291 & ~pi297;
  assign n871 = pi299 & ~pi303;
  assign n872 = n870 & n871;
  assign n873 = n815 & n872;
  assign n874 = n788 & n873;
  assign n875 = ~pi291 & ~pi299;
  assign n876 = pi297 & n875;
  assign n877 = pi296 & ~pi300;
  assign n878 = pi303 & n877;
  assign n879 = n876 & n878;
  assign n880 = n876 & n877;
  assign n881 = ~pi303 & n880;
  assign n882 = ~n879 & ~n881;
  assign n883 = pi296 & pi297;
  assign n884 = n790 & n883;
  assign n885 = n823 & n884;
  assign n886 = pi298 & pi299;
  assign n887 = n885 & n886;
  assign n888 = ~n788 & ~n802;
  assign n889 = pi190 & ~n888;
  assign n890 = n887 & n889;
  assign n891 = n882 & ~n890;
  assign n892 = ~n874 & n891;
  assign n893 = ~n869 & n892;
  assign n894 = n836 & n893;
  assign n895 = ~n801 & n894;
  assign n896 = n787 & ~n895;
  assign n897 = pi298 & pi300;
  assign n898 = ~pi296 & n897;
  assign n899 = ~pi299 & n898;
  assign n900 = ~pi297 & n899;
  assign n901 = ~pi291 & n900;
  assign n902 = ~pi291 & n897;
  assign n903 = pi296 & n902;
  assign n904 = ~pi297 & ~pi299;
  assign n905 = n903 & n904;
  assign n906 = ~n901 & ~n905;
  assign n907 = ~n812 & ~n906;
  assign n908 = ~pi297 & n877;
  assign n909 = n813 & n908;
  assign n910 = n788 & n909;
  assign n911 = ~n907 & ~n910;
  assign n912 = n804 & n901;
  assign n913 = n911 & ~n912;
  assign n914 = pi301 & ~n913;
  assign n915 = ~n896 & ~n914;
  assign n916 = pi302 & ~n882;
  assign n917 = ~n869 & ~n874;
  assign n918 = ~n890 & n917;
  assign n919 = n835 & n918;
  assign n920 = ~n916 & n919;
  assign n921 = ~n801 & n819;
  assign n922 = n920 & n921;
  assign n923 = n787 & ~n922;
  assign n924 = ~n910 & ~n912;
  assign n925 = pi301 & ~n924;
  assign n926 = ~n923 & ~n925;
  assign n927 = pi297 & ~pi299;
  assign n928 = pi296 & n927;
  assign n929 = n902 & n928;
  assign n930 = n804 & n929;
  assign n931 = ~pi296 & n927;
  assign n932 = n902 & n931;
  assign n933 = n804 & n932;
  assign n934 = ~n930 & ~n933;
  assign n935 = n811 & n905;
  assign n936 = n811 & n901;
  assign n937 = ~n935 & ~n936;
  assign n938 = ~n910 & n937;
  assign n939 = n934 & n938;
  assign n940 = pi301 & ~n939;
  assign n941 = pi298 & ~n882;
  assign n942 = ~n801 & ~n941;
  assign n943 = n819 & n942;
  assign n944 = n919 & n943;
  assign n945 = n787 & ~n944;
  assign n946 = ~n940 & ~n945;
  assign n947 = n926 & n946;
  assign n948 = ~n915 & n947;
  assign n949 = ~n786 & n948;
  assign n950 = ~pi257 & pi271;
  assign n951 = pi257 & pi273;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~pi257 & pi272;
  assign n954 = pi257 & pi275;
  assign n955 = ~n953 & ~n954;
  assign n956 = ~pi241 & pi257;
  assign n957 = pi241 & ~pi257;
  assign n958 = ~n956 & ~n957;
  assign n959 = pi256 & ~n958;
  assign n960 = pi243 & n959;
  assign n961 = ~pi198 & ~pi216;
  assign n962 = ~pi257 & pi274;
  assign n963 = pi257 & pi269;
  assign n964 = ~n962 & ~n963;
  assign n965 = n961 & n964;
  assign n966 = ~pi217 & n965;
  assign n967 = ~pi223 & n966;
  assign n968 = n960 & n967;
  assign n969 = ~pi257 & pi264;
  assign n970 = pi257 & pi270;
  assign n971 = ~n969 & ~n970;
  assign n972 = n968 & n971;
  assign n973 = n955 & n972;
  assign n974 = n952 & n973;
  assign n975 = ~pi241 & ~pi256;
  assign n976 = pi243 & ~pi257;
  assign n977 = n975 & n976;
  assign n978 = pi216 & n853;
  assign n979 = pi217 & n840;
  assign n980 = ~n978 & ~n979;
  assign n981 = pi298 & n862;
  assign n982 = pi216 & n981;
  assign n983 = pi217 & n842;
  assign n984 = ~n982 & ~n983;
  assign n985 = pi298 & n844;
  assign n986 = ~n845 & ~n985;
  assign n987 = pi217 & ~n986;
  assign n988 = ~n857 & ~n863;
  assign n989 = pi216 & ~n988;
  assign n990 = ~n987 & ~n989;
  assign n991 = n984 & n990;
  assign n992 = n980 & n991;
  assign n993 = ~n787 & n992;
  assign n994 = pi202 & n853;
  assign n995 = pi198 & n840;
  assign n996 = ~n994 & ~n995;
  assign n997 = pi202 & n981;
  assign n998 = pi198 & n842;
  assign n999 = ~n997 & ~n998;
  assign n1000 = pi198 & ~n986;
  assign n1001 = pi202 & ~n988;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = n999 & n1002;
  assign n1004 = n996 & n1003;
  assign n1005 = pi225 & n845;
  assign n1006 = pi223 & n857;
  assign n1007 = ~n840 & ~n842;
  assign n1008 = pi225 & ~n1007;
  assign n1009 = ~n1006 & ~n1008;
  assign n1010 = pi225 & n985;
  assign n1011 = pi132 & n863;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~n981 & n1012;
  assign n1014 = n1009 & n1013;
  assign n1015 = ~n1005 & n1014;
  assign n1016 = pi223 & n985;
  assign n1017 = pi198 & n857;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = pi223 & n845;
  assign n1020 = n1018 & ~n1019;
  assign n1021 = pi223 & n842;
  assign n1022 = pi198 & n863;
  assign n1023 = pi223 & n840;
  assign n1024 = ~n1022 & ~n1023;
  assign n1025 = ~n853 & ~n981;
  assign n1026 = pi198 & ~n1025;
  assign n1027 = n1024 & ~n1026;
  assign n1028 = ~n1021 & n1027;
  assign n1029 = n1020 & n1028;
  assign n1030 = n1015 & n1029;
  assign n1031 = pi217 & n981;
  assign n1032 = ~n1021 & ~n1031;
  assign n1033 = pi197 & n840;
  assign n1034 = pi217 & n857;
  assign n1035 = ~n846 & ~n1034;
  assign n1036 = ~n853 & ~n863;
  assign n1037 = pi217 & ~n1036;
  assign n1038 = n1035 & ~n1037;
  assign n1039 = ~n1033 & n1038;
  assign n1040 = n1032 & n1039;
  assign n1041 = n1030 & n1040;
  assign n1042 = n1004 & n1041;
  assign n1043 = n993 & n1042;
  assign n1044 = pi197 & n853;
  assign n1045 = pi215 & n840;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = pi197 & n981;
  assign n1048 = pi215 & n842;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = pi215 & ~n986;
  assign n1051 = pi197 & ~n988;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n1049 & n1052;
  assign n1054 = n1046 & n1053;
  assign n1055 = n1043 & n1054;
  assign n1056 = pi225 & n853;
  assign n1057 = pi202 & n840;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = pi225 & n981;
  assign n1060 = pi202 & n842;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = pi202 & ~n986;
  assign n1063 = pi225 & ~n988;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n1061 & n1064;
  assign n1066 = n1058 & n1065;
  assign n1067 = pi215 & n853;
  assign n1068 = pi216 & n840;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = pi215 & n981;
  assign n1071 = pi216 & n842;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = pi216 & ~n986;
  assign n1074 = pi215 & ~n988;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = n1072 & n1075;
  assign n1077 = n1069 & n1076;
  assign n1078 = n1066 & n1077;
  assign n1079 = n1055 & n1078;
  assign n1080 = pi131 & n787;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = n977 & ~n1081;
  assign n1083 = pi243 & n975;
  assign n1084 = pi257 & n1083;
  assign n1085 = ~n960 & ~n1084;
  assign n1086 = ~pi241 & pi256;
  assign n1087 = n976 & n1086;
  assign n1088 = ~n977 & ~n1087;
  assign n1089 = pi243 & n1088;
  assign n1090 = n1085 & n1089;
  assign n1091 = pi131 & n1090;
  assign n1092 = pi256 & ~pi257;
  assign n1093 = pi241 & ~n1092;
  assign n1094 = ~pi241 & pi270;
  assign n1095 = pi241 & ~pi270;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = pi216 & ~n1096;
  assign n1098 = ~pi241 & pi273;
  assign n1099 = pi241 & ~pi273;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~pi198 & n1100;
  assign n1102 = n1097 & ~n1101;
  assign n1103 = pi198 & ~n1100;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~pi241 & pi269;
  assign n1106 = pi241 & ~pi269;
  assign n1107 = ~n1105 & ~n1106;
  assign n1108 = pi217 & ~n1107;
  assign n1109 = ~pi217 & n1107;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1104 & ~n1110;
  assign n1112 = n1104 & n1110;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = ~n1101 & ~n1103;
  assign n1115 = n1097 & n1114;
  assign n1116 = ~n1097 & ~n1114;
  assign n1117 = ~n1115 & ~n1116;
  assign n1118 = ~pi216 & ~n1096;
  assign n1119 = pi216 & n1096;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~pi241 & pi274;
  assign n1122 = pi241 & ~pi274;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = pi215 & ~n1123;
  assign n1125 = ~pi241 & pi272;
  assign n1126 = pi241 & ~pi272;
  assign n1127 = ~n1125 & ~n1126;
  assign n1128 = pi202 & ~n1127;
  assign n1129 = ~n1124 & ~n1128;
  assign n1130 = ~pi202 & n1127;
  assign n1131 = n1127 & n1130;
  assign n1132 = ~n1129 & ~n1131;
  assign n1133 = ~pi202 & n1130;
  assign n1134 = n1132 & ~n1133;
  assign n1135 = ~pi241 & pi264;
  assign n1136 = pi241 & ~pi264;
  assign n1137 = ~n1135 & ~n1136;
  assign n1138 = pi197 & ~n1137;
  assign n1139 = ~pi241 & pi271;
  assign n1140 = pi241 & ~pi271;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = ~pi225 & n1141;
  assign n1143 = n1138 & ~n1142;
  assign n1144 = pi225 & ~n1141;
  assign n1145 = ~n1143 & ~n1144;
  assign n1146 = ~pi215 & n1123;
  assign n1147 = ~n1130 & ~n1146;
  assign n1148 = ~n1145 & n1147;
  assign n1149 = ~n1134 & ~n1148;
  assign n1150 = ~n1124 & ~n1146;
  assign n1151 = n1145 & ~n1150;
  assign n1152 = ~n1145 & n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1142 & ~n1144;
  assign n1155 = ~n1138 & n1154;
  assign n1156 = n1138 & ~n1154;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~pi197 & ~n1137;
  assign n1159 = pi197 & n1137;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = pi132 & ~pi256;
  assign n1162 = pi257 & n1161;
  assign n1163 = ~pi241 & n1162;
  assign n1164 = pi241 & ~n1162;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = ~n1160 & ~n1165;
  assign n1167 = ~n1157 & n1166;
  assign n1168 = n1153 & n1167;
  assign n1169 = ~n1128 & ~n1130;
  assign n1170 = ~n1145 & ~n1146;
  assign n1171 = ~n1124 & ~n1170;
  assign n1172 = n1169 & n1171;
  assign n1173 = ~n1169 & ~n1171;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = n1168 & ~n1174;
  assign n1176 = n1149 & n1175;
  assign n1177 = ~n1149 & ~n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1120 & ~n1178;
  assign n1180 = n1117 & n1179;
  assign n1181 = ~n1113 & ~n1180;
  assign n1182 = n1113 & n1180;
  assign n1183 = ~n1181 & ~n1182;
  assign n1184 = n1093 & ~n1183;
  assign n1185 = pi241 & n1092;
  assign n1186 = ~pi217 & ~pi269;
  assign n1187 = n1185 & ~n1186;
  assign n1188 = n975 & ~n1183;
  assign n1189 = pi257 & n1086;
  assign n1190 = ~pi217 & pi269;
  assign n1191 = pi217 & ~pi269;
  assign n1192 = ~n1190 & ~n1191;
  assign n1193 = n1189 & ~n1192;
  assign n1194 = ~n1188 & ~n1193;
  assign n1195 = ~pi241 & n1092;
  assign n1196 = pi269 & n1195;
  assign n1197 = pi217 & n1196;
  assign n1198 = n1194 & ~n1197;
  assign n1199 = ~n1187 & n1198;
  assign n1200 = ~n1184 & n1199;
  assign n1201 = ~n1117 & n1179;
  assign n1202 = n1117 & ~n1179;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = n1093 & ~n1203;
  assign n1205 = pi273 & n1195;
  assign n1206 = pi198 & n1205;
  assign n1207 = n975 & ~n1203;
  assign n1208 = ~pi198 & pi273;
  assign n1209 = pi198 & ~pi273;
  assign n1210 = ~n1208 & ~n1209;
  assign n1211 = n1189 & ~n1210;
  assign n1212 = ~n1207 & ~n1211;
  assign n1213 = ~pi198 & ~pi273;
  assign n1214 = n1185 & ~n1213;
  assign n1215 = n1212 & ~n1214;
  assign n1216 = ~n1206 & n1215;
  assign n1217 = ~n1204 & n1216;
  assign n1218 = n1200 & n1217;
  assign n1219 = ~pi223 & pi275;
  assign n1220 = pi223 & ~pi275;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = n1189 & ~n1221;
  assign n1223 = ~pi223 & ~pi275;
  assign n1224 = n1185 & ~n1223;
  assign n1225 = ~n1222 & ~n1224;
  assign n1226 = ~n1113 & n1180;
  assign n1227 = ~n975 & ~n1093;
  assign n1228 = ~n1108 & n1109;
  assign n1229 = ~n1103 & ~n1108;
  assign n1230 = ~n1228 & ~n1229;
  assign n1231 = ~n1101 & ~n1109;
  assign n1232 = n1097 & n1231;
  assign n1233 = ~n1230 & ~n1232;
  assign n1234 = ~pi241 & pi275;
  assign n1235 = pi241 & ~pi275;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = pi223 & ~n1236;
  assign n1238 = ~pi223 & n1236;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = n1233 & n1239;
  assign n1241 = ~n1227 & ~n1240;
  assign n1242 = ~n1233 & ~n1239;
  assign n1243 = n1241 & ~n1242;
  assign n1244 = n1226 & ~n1243;
  assign n1245 = ~n1233 & n1239;
  assign n1246 = ~n1227 & ~n1245;
  assign n1247 = n1233 & ~n1239;
  assign n1248 = n1246 & ~n1247;
  assign n1249 = ~n1226 & ~n1248;
  assign n1250 = ~n1244 & ~n1249;
  assign n1251 = pi223 & n1195;
  assign n1252 = pi275 & n1251;
  assign n1253 = ~n1250 & ~n1252;
  assign n1254 = n1225 & n1253;
  assign n1255 = n1218 & n1254;
  assign n1256 = ~pi225 & ~pi271;
  assign n1257 = n1185 & ~n1256;
  assign n1258 = n1157 & n1166;
  assign n1259 = ~n1157 & ~n1166;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = n975 & ~n1260;
  assign n1262 = ~n1257 & ~n1261;
  assign n1263 = n1093 & ~n1260;
  assign n1264 = pi225 & ~pi271;
  assign n1265 = ~pi225 & pi271;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n1189 & ~n1266;
  assign n1268 = ~n1263 & ~n1267;
  assign n1269 = pi271 & n1195;
  assign n1270 = pi225 & n1269;
  assign n1271 = n1268 & ~n1270;
  assign n1272 = n1262 & n1271;
  assign n1273 = n1160 & ~n1165;
  assign n1274 = ~n1160 & n1165;
  assign n1275 = ~n1273 & ~n1274;
  assign n1276 = n1093 & ~n1275;
  assign n1277 = ~pi197 & ~pi264;
  assign n1278 = n1185 & ~n1277;
  assign n1279 = n975 & ~n1275;
  assign n1280 = pi197 & ~pi264;
  assign n1281 = ~pi197 & pi264;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = n1189 & ~n1282;
  assign n1284 = ~n1279 & ~n1283;
  assign n1285 = pi264 & n1195;
  assign n1286 = pi197 & n1285;
  assign n1287 = n1284 & ~n1286;
  assign n1288 = ~n1278 & n1287;
  assign n1289 = ~n1276 & n1288;
  assign n1290 = n1272 & n1289;
  assign n1291 = ~n1120 & n1178;
  assign n1292 = n1120 & ~n1178;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n975 & ~n1293;
  assign n1295 = ~pi216 & ~pi270;
  assign n1296 = n1185 & ~n1295;
  assign n1297 = n1093 & ~n1293;
  assign n1298 = ~pi216 & pi270;
  assign n1299 = pi216 & ~pi270;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = n1189 & ~n1300;
  assign n1302 = ~n1297 & ~n1301;
  assign n1303 = pi270 & n1195;
  assign n1304 = pi216 & n1303;
  assign n1305 = n1302 & ~n1304;
  assign n1306 = ~n1296 & n1305;
  assign n1307 = ~n1294 & n1306;
  assign n1308 = n1290 & n1307;
  assign n1309 = ~pi202 & ~pi272;
  assign n1310 = n1185 & ~n1309;
  assign n1311 = n1168 & n1174;
  assign n1312 = ~n1168 & ~n1174;
  assign n1313 = ~n1311 & ~n1312;
  assign n1314 = n975 & ~n1313;
  assign n1315 = ~n1310 & ~n1314;
  assign n1316 = n1093 & ~n1313;
  assign n1317 = ~pi202 & pi272;
  assign n1318 = pi202 & ~pi272;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = n1189 & ~n1319;
  assign n1321 = ~n1316 & ~n1320;
  assign n1322 = pi272 & n1195;
  assign n1323 = pi202 & n1322;
  assign n1324 = n1321 & ~n1323;
  assign n1325 = n1315 & n1324;
  assign n1326 = ~n1153 & n1167;
  assign n1327 = n1153 & ~n1167;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = n975 & ~n1328;
  assign n1330 = pi274 & n1195;
  assign n1331 = pi215 & n1330;
  assign n1332 = n1093 & ~n1328;
  assign n1333 = pi215 & ~pi274;
  assign n1334 = ~pi215 & pi274;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = n1189 & ~n1335;
  assign n1337 = ~n1332 & ~n1336;
  assign n1338 = ~pi215 & ~pi274;
  assign n1339 = n1185 & ~n1338;
  assign n1340 = n1337 & ~n1339;
  assign n1341 = ~n1331 & n1340;
  assign n1342 = ~n1329 & n1341;
  assign n1343 = n1325 & n1342;
  assign n1344 = ~pi131 & pi278;
  assign n1345 = n1343 & ~n1344;
  assign n1346 = n1308 & n1345;
  assign n1347 = n1255 & n1346;
  assign n1348 = ~pi344 & n1347;
  assign n1349 = pi131 & pi344;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~pi243 & ~n1350;
  assign n1352 = ~n1091 & ~n1351;
  assign n1353 = ~pi298 & ~pi302;
  assign n1354 = ~pi303 & n1353;
  assign n1355 = pi264 & n1354;
  assign n1356 = pi269 & n850;
  assign n1357 = pi275 & n859;
  assign n1358 = pi298 & ~pi302;
  assign n1359 = ~pi303 & n1358;
  assign n1360 = pi270 & n1359;
  assign n1361 = pi303 & n1358;
  assign n1362 = pi273 & n1361;
  assign n1363 = ~n1360 & ~n1362;
  assign n1364 = ~n1357 & n1363;
  assign n1365 = ~n1356 & n1364;
  assign n1366 = pi303 & n1353;
  assign n1367 = pi271 & n1366;
  assign n1368 = n1084 & ~n1367;
  assign n1369 = n1365 & n1368;
  assign n1370 = ~n1355 & n1369;
  assign n1371 = ~pi298 & pi302;
  assign n1372 = ~pi303 & n1371;
  assign n1373 = pi274 & n1372;
  assign n1374 = pi303 & n1371;
  assign n1375 = pi272 & n1374;
  assign n1376 = ~n1373 & ~n1375;
  assign n1377 = n1370 & n1376;
  assign n1378 = n1352 & ~n1377;
  assign n1379 = ~pi215 & ~pi225;
  assign n1380 = pi202 & ~n1379;
  assign n1381 = ~pi184 & ~n1380;
  assign n1382 = pi202 & n1381;
  assign n1383 = ~pi202 & n1379;
  assign n1384 = ~n1380 & ~n1383;
  assign n1385 = ~n1381 & n1384;
  assign n1386 = ~n1382 & ~n1385;
  assign n1387 = ~pi129 & ~n1386;
  assign n1388 = pi215 & pi225;
  assign n1389 = ~pi202 & ~n1388;
  assign n1390 = pi202 & n1388;
  assign n1391 = ~n1389 & ~n1390;
  assign n1392 = ~n1381 & ~n1391;
  assign n1393 = ~n1382 & ~n1392;
  assign n1394 = pi129 & ~n1393;
  assign n1395 = ~n1387 & ~n1394;
  assign n1396 = pi225 & ~n1381;
  assign n1397 = ~pi225 & n1381;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = pi217 & n1381;
  assign n1400 = pi216 & n1380;
  assign n1401 = pi198 & n1400;
  assign n1402 = pi217 & n1401;
  assign n1403 = ~pi217 & ~n1401;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1381 & n1404;
  assign n1406 = ~n1399 & ~n1405;
  assign n1407 = pi198 & n1381;
  assign n1408 = ~pi198 & n1400;
  assign n1409 = pi198 & ~n1400;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1381 & ~n1410;
  assign n1412 = ~n1407 & ~n1411;
  assign n1413 = pi223 & n1401;
  assign n1414 = pi217 & n1413;
  assign n1415 = ~n1381 & n1414;
  assign n1416 = pi223 & n1381;
  assign n1417 = pi198 & pi217;
  assign n1418 = n1400 & n1417;
  assign n1419 = ~pi223 & ~n1418;
  assign n1420 = pi223 & n1418;
  assign n1421 = ~n1419 & ~n1420;
  assign n1422 = ~n1381 & n1421;
  assign n1423 = ~n1416 & ~n1422;
  assign n1424 = n1406 & n1412;
  assign n1425 = ~n1423 & ~n1424;
  assign n1426 = ~n1415 & ~n1425;
  assign n1427 = ~pi132 & n1426;
  assign n1428 = n1412 & ~n1427;
  assign n1429 = ~n1406 & ~n1428;
  assign n1430 = n1424 & ~n1427;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~pi129 & ~n1431;
  assign n1433 = ~pi198 & ~n1400;
  assign n1434 = ~pi217 & n1433;
  assign n1435 = pi223 & ~n1434;
  assign n1436 = ~pi132 & ~n1435;
  assign n1437 = ~pi202 & ~pi216;
  assign n1438 = ~n1388 & n1437;
  assign n1439 = ~pi198 & ~n1438;
  assign n1440 = pi198 & n1438;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~n1381 & n1441;
  assign n1443 = ~n1407 & ~n1442;
  assign n1444 = ~pi202 & n961;
  assign n1445 = ~n1388 & n1444;
  assign n1446 = pi217 & n1445;
  assign n1447 = ~pi217 & ~n1445;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1381 & n1448;
  assign n1450 = ~n1399 & ~n1449;
  assign n1451 = ~n1443 & n1450;
  assign n1452 = n1443 & ~n1450;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = ~n1436 & ~n1453;
  assign n1455 = n1436 & ~n1450;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = pi129 & ~n1456;
  assign n1458 = ~n1432 & ~n1457;
  assign n1459 = ~n1412 & n1427;
  assign n1460 = ~n1428 & ~n1459;
  assign n1461 = ~pi129 & n1460;
  assign n1462 = n1436 & n1443;
  assign n1463 = ~n1436 & ~n1443;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = pi129 & ~n1464;
  assign n1466 = ~n1461 & ~n1465;
  assign n1467 = pi216 & n1381;
  assign n1468 = ~pi216 & ~n1380;
  assign n1469 = ~n1400 & ~n1468;
  assign n1470 = ~n1381 & n1469;
  assign n1471 = ~n1467 & ~n1470;
  assign n1472 = ~pi129 & ~n1471;
  assign n1473 = ~pi216 & ~n1389;
  assign n1474 = pi216 & n1389;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = ~n1381 & n1475;
  assign n1477 = ~n1467 & ~n1476;
  assign n1478 = pi129 & ~n1477;
  assign n1479 = ~n1472 & ~n1478;
  assign n1480 = ~n1466 & n1479;
  assign n1481 = n1458 & n1480;
  assign n1482 = ~pi197 & n1087;
  assign n1483 = ~n1423 & n1427;
  assign n1484 = ~n1423 & n1424;
  assign n1485 = n1423 & ~n1424;
  assign n1486 = ~n1484 & ~n1485;
  assign n1487 = ~n1427 & ~n1486;
  assign n1488 = ~n1483 & ~n1487;
  assign n1489 = ~pi129 & ~n1488;
  assign n1490 = ~pi217 & n1445;
  assign n1491 = pi223 & n1490;
  assign n1492 = ~pi223 & ~n1490;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = ~n1381 & n1493;
  assign n1495 = ~n1416 & ~n1494;
  assign n1496 = ~n1443 & ~n1450;
  assign n1497 = ~n1495 & n1496;
  assign n1498 = n1495 & ~n1496;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1436 & ~n1499;
  assign n1501 = n1436 & ~n1495;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = pi129 & ~n1502;
  assign n1504 = ~n1489 & ~n1503;
  assign n1505 = n1482 & n1504;
  assign n1506 = n1481 & n1505;
  assign n1507 = pi215 & n1381;
  assign n1508 = pi215 & ~pi225;
  assign n1509 = ~pi215 & pi225;
  assign n1510 = ~n1508 & ~n1509;
  assign n1511 = ~n1381 & ~n1510;
  assign n1512 = ~n1507 & ~n1511;
  assign n1513 = pi129 & n1512;
  assign n1514 = ~n1379 & ~n1388;
  assign n1515 = ~n1381 & ~n1514;
  assign n1516 = ~n1507 & ~n1515;
  assign n1517 = ~pi129 & n1516;
  assign n1518 = ~n1513 & ~n1517;
  assign n1519 = n1506 & ~n1518;
  assign n1520 = ~n1398 & n1519;
  assign n1521 = n1395 & n1520;
  assign n1522 = n1378 & ~n1521;
  assign n1523 = ~n1082 & n1522;
  assign n1524 = ~n974 & n1523;
  assign n1525 = ~pi300 & pi302;
  assign n1526 = n821 & n1525;
  assign n1527 = n824 & n1526;
  assign n1528 = ~n812 & n1527;
  assign n1529 = n787 & n1528;
  assign n1530 = pi242 & n1529;
  assign n1531 = ~n1524 & n1530;
  assign n1532 = pi000 & ~n1530;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n949 & n1533;
  assign n1535 = pi303 & n804;
  assign n1536 = pi303 & n811;
  assign n1537 = ~n780 & ~n1536;
  assign n1538 = ~n1535 & n1537;
  assign n1539 = n901 & ~n1538;
  assign n1540 = n905 & ~n1537;
  assign n1541 = ~n929 & ~n932;
  assign n1542 = n1535 & ~n1541;
  assign n1543 = ~n1540 & ~n1542;
  assign n1544 = ~n1539 & n1543;
  assign n1545 = pi301 & ~n1544;
  assign n1546 = pi190 & n802;
  assign n1547 = n887 & n1546;
  assign n1548 = n835 & ~n879;
  assign n1549 = n838 & n867;
  assign n1550 = n803 & n838;
  assign n1551 = ~n1549 & ~n1550;
  assign n1552 = n819 & n1551;
  assign n1553 = n1548 & n1552;
  assign n1554 = ~n1547 & n1553;
  assign n1555 = n787 & ~n1554;
  assign n1556 = ~n1545 & ~n1555;
  assign n1557 = n787 & n883;
  assign n1558 = pi299 & pi300;
  assign n1559 = pi298 & n1558;
  assign n1560 = ~pi302 & n1559;
  assign n1561 = n1557 & n1560;
  assign n1562 = n793 & n1561;
  assign n1563 = n782 & n1562;
  assign n1564 = ~pi097 & ~pi098;
  assign n1565 = pi099 & n1564;
  assign n1566 = n1562 & n1565;
  assign n1567 = pi311 & ~n1566;
  assign n1568 = pi304 & n1566;
  assign n1569 = ~n1567 & ~n1568;
  assign n1570 = ~n1563 & ~n1569;
  assign n1571 = pi304 & n1563;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = n783 & ~n915;
  assign n1574 = ~n785 & ~n1573;
  assign n1575 = ~pi313 & ~pi314;
  assign n1576 = ~n1574 & n1575;
  assign n1577 = n926 & ~n1574;
  assign n1578 = ~n946 & n1577;
  assign n1579 = ~n1576 & ~n1578;
  assign n1580 = ~n1572 & n1579;
  assign n1581 = pi304 & n1576;
  assign n1582 = pi314 & n1578;
  assign n1583 = ~n1576 & n1582;
  assign n1584 = ~n1581 & ~n1583;
  assign n1585 = ~n1580 & n1584;
  assign n1586 = ~n1576 & n1578;
  assign n1587 = ~n926 & n1576;
  assign n1588 = ~pi312 & ~n1566;
  assign n1589 = ~n1576 & ~n1588;
  assign n1590 = ~n1563 & n1589;
  assign n1591 = ~n1587 & ~n1590;
  assign n1592 = ~n1586 & n1591;
  assign n1593 = pi309 & ~n1566;
  assign n1594 = ~n1563 & ~n1593;
  assign n1595 = ~n1576 & ~n1594;
  assign n1596 = ~n946 & n1576;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1586 & n1597;
  assign n1599 = ~n1592 & ~n1598;
  assign n1600 = ~n1585 & n1599;
  assign n1601 = pi080 & n1600;
  assign n1602 = n1592 & n1598;
  assign n1603 = ~n1585 & n1602;
  assign n1604 = pi078 & n1603;
  assign n1605 = n1585 & ~n1592;
  assign n1606 = n1598 & n1605;
  assign n1607 = pi075 & n1606;
  assign n1608 = n1585 & n1602;
  assign n1609 = pi074 & n1608;
  assign n1610 = ~n1607 & ~n1609;
  assign n1611 = ~n1604 & n1610;
  assign n1612 = ~n1601 & n1611;
  assign n1613 = n1585 & ~n1598;
  assign n1614 = n1592 & n1613;
  assign n1615 = pi076 & n1614;
  assign n1616 = ~n1598 & n1605;
  assign n1617 = pi077 & n1616;
  assign n1618 = n1592 & ~n1598;
  assign n1619 = ~n1585 & n1618;
  assign n1620 = pi079 & n1619;
  assign n1621 = ~n1585 & ~n1592;
  assign n1622 = n1598 & n1621;
  assign n1623 = pi065 & n1622;
  assign n1624 = ~n1620 & ~n1623;
  assign n1625 = ~n1617 & n1624;
  assign n1626 = ~n1615 & n1625;
  assign n1627 = n1612 & n1626;
  assign n1628 = n1556 & n1627;
  assign n1629 = pi023 & n1614;
  assign n1630 = pi022 & n1606;
  assign n1631 = pi021 & n1608;
  assign n1632 = pi024 & n1616;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n1630 & n1633;
  assign n1635 = ~n1629 & n1634;
  assign n1636 = pi028 & n1600;
  assign n1637 = pi025 & n1603;
  assign n1638 = pi026 & n1622;
  assign n1639 = pi027 & n1619;
  assign n1640 = ~n1638 & ~n1639;
  assign n1641 = ~n1637 & n1640;
  assign n1642 = ~n1636 & n1641;
  assign n1643 = n1635 & n1642;
  assign n1644 = n1556 & n1643;
  assign n1645 = ~n1628 & ~n1644;
  assign n1646 = pi093 & n1616;
  assign n1647 = pi092 & n1614;
  assign n1648 = ~n1646 & ~n1647;
  assign n1649 = pi091 & n1606;
  assign n1650 = pi090 & n1608;
  assign n1651 = ~n1649 & ~n1650;
  assign n1652 = pi095 & n1619;
  assign n1653 = pi094 & n1622;
  assign n1654 = ~n1652 & ~n1653;
  assign n1655 = pi081 & n1603;
  assign n1656 = pi096 & n1600;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = n1654 & n1657;
  assign n1659 = n1651 & n1658;
  assign n1660 = n1648 & n1659;
  assign n1661 = n1556 & n1660;
  assign n1662 = pi082 & n1600;
  assign n1663 = pi087 & n1603;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = pi083 & n1608;
  assign n1666 = pi084 & n1606;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = n1664 & n1667;
  assign n1669 = pi085 & n1614;
  assign n1670 = pi086 & n1616;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = pi088 & n1622;
  assign n1673 = pi089 & n1619;
  assign n1674 = ~n1672 & ~n1673;
  assign n1675 = n1671 & n1674;
  assign n1676 = n1668 & n1675;
  assign n1677 = n1556 & n1676;
  assign n1678 = ~n1661 & ~n1677;
  assign n1679 = pi069 & n1622;
  assign n1680 = pi072 & n1616;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = pi070 & n1619;
  assign n1683 = pi068 & n1614;
  assign n1684 = ~n1682 & ~n1683;
  assign n1685 = pi071 & n1600;
  assign n1686 = pi066 & n1608;
  assign n1687 = ~n1685 & ~n1686;
  assign n1688 = n1684 & n1687;
  assign n1689 = pi067 & n1606;
  assign n1690 = pi073 & n1603;
  assign n1691 = ~n1689 & ~n1690;
  assign n1692 = n1688 & n1691;
  assign n1693 = n1681 & n1692;
  assign n1694 = n1556 & n1693;
  assign n1695 = pi107 & n1622;
  assign n1696 = pi108 & n1619;
  assign n1697 = pi106 & n1603;
  assign n1698 = pi109 & n1600;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = ~n1696 & n1699;
  assign n1701 = ~n1695 & n1700;
  assign n1702 = pi101 & n1608;
  assign n1703 = pi103 & n1606;
  assign n1704 = pi104 & n1614;
  assign n1705 = pi105 & n1616;
  assign n1706 = ~n1704 & ~n1705;
  assign n1707 = ~n1703 & n1706;
  assign n1708 = ~n1702 & n1707;
  assign n1709 = n1701 & n1708;
  assign n1710 = n1556 & n1709;
  assign n1711 = ~n1694 & ~n1710;
  assign n1712 = n1678 & n1711;
  assign n1713 = pi112 & n1614;
  assign n1714 = pi113 & n1616;
  assign n1715 = pi115 & n1600;
  assign n1716 = pi100 & n1603;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = ~n1714 & n1717;
  assign n1719 = ~n1713 & n1718;
  assign n1720 = pi110 & n1608;
  assign n1721 = pi111 & n1606;
  assign n1722 = pi116 & n1622;
  assign n1723 = pi114 & n1619;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = ~n1721 & n1724;
  assign n1726 = ~n1720 & n1725;
  assign n1727 = n1719 & n1726;
  assign n1728 = ~n1556 & ~n1727;
  assign n1729 = n1556 & n1727;
  assign n1730 = pi121 & n1606;
  assign n1731 = pi120 & n1608;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = pi122 & n1616;
  assign n1734 = pi125 & n1614;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = pi119 & n1619;
  assign n1737 = pi118 & n1622;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = pi123 & n1603;
  assign n1740 = pi124 & n1600;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = n1738 & n1741;
  assign n1743 = n1735 & n1742;
  assign n1744 = n1732 & n1743;
  assign n1745 = ~n1556 & ~n1744;
  assign n1746 = ~n1729 & n1745;
  assign n1747 = ~n1728 & ~n1746;
  assign n1748 = n1556 & n1744;
  assign n1749 = ~n1729 & ~n1748;
  assign n1750 = pi147 & n1608;
  assign n1751 = pi152 & n1619;
  assign n1752 = pi151 & n1622;
  assign n1753 = pi148 & n1606;
  assign n1754 = ~n1752 & ~n1753;
  assign n1755 = ~n1751 & n1754;
  assign n1756 = ~n1750 & n1755;
  assign n1757 = pi149 & n1614;
  assign n1758 = pi175 & n1603;
  assign n1759 = pi153 & n1600;
  assign n1760 = pi150 & n1616;
  assign n1761 = ~n1759 & ~n1760;
  assign n1762 = ~n1758 & n1761;
  assign n1763 = ~n1757 & n1762;
  assign n1764 = n1756 & n1763;
  assign n1765 = n1556 & n1764;
  assign n1766 = pi165 & n1608;
  assign n1767 = pi167 & n1614;
  assign n1768 = pi166 & n1606;
  assign n1769 = pi168 & n1616;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~n1767 & n1770;
  assign n1772 = ~n1766 & n1771;
  assign n1773 = pi170 & n1622;
  assign n1774 = pi176 & n1619;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = pi171 & n1600;
  assign n1777 = pi169 & n1603;
  assign n1778 = ~n1776 & ~n1777;
  assign n1779 = n1775 & n1778;
  assign n1780 = n1772 & n1779;
  assign n1781 = ~n1765 & ~n1780;
  assign n1782 = pi154 & n1608;
  assign n1783 = pi156 & n1614;
  assign n1784 = pi155 & n1606;
  assign n1785 = pi157 & n1616;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = ~n1783 & n1786;
  assign n1788 = ~n1782 & n1787;
  assign n1789 = pi158 & n1622;
  assign n1790 = pi159 & n1619;
  assign n1791 = pi160 & n1600;
  assign n1792 = pi127 & n1603;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = ~n1790 & n1793;
  assign n1795 = ~n1789 & n1794;
  assign n1796 = n1788 & n1795;
  assign n1797 = n1556 & n1796;
  assign n1798 = n1781 & ~n1797;
  assign n1799 = n1749 & n1798;
  assign n1800 = ~n1556 & ~n1796;
  assign n1801 = ~n1765 & n1800;
  assign n1802 = ~n1556 & ~n1764;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = n1749 & ~n1803;
  assign n1805 = ~n1799 & ~n1804;
  assign n1806 = n1747 & n1805;
  assign n1807 = n1712 & ~n1806;
  assign n1808 = ~pi059 & n1614;
  assign n1809 = ~pi060 & n1616;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = ~pi063 & n1619;
  assign n1812 = ~pi062 & n1622;
  assign n1813 = ~n1811 & ~n1812;
  assign n1814 = ~pi064 & n1600;
  assign n1815 = ~pi061 & n1603;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = ~pi058 & n1606;
  assign n1818 = ~pi057 & n1608;
  assign n1819 = ~n1817 & ~n1818;
  assign n1820 = n1816 & n1819;
  assign n1821 = n1813 & n1820;
  assign n1822 = n1810 & n1821;
  assign n1823 = n1556 & n1822;
  assign n1824 = ~pi015 & n1614;
  assign n1825 = ~pi016 & n1616;
  assign n1826 = ~pi020 & n1600;
  assign n1827 = ~pi017 & n1603;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1825 & n1828;
  assign n1830 = ~n1824 & n1829;
  assign n1831 = ~pi018 & n1622;
  assign n1832 = ~pi014 & n1606;
  assign n1833 = ~pi019 & n1619;
  assign n1834 = ~n1832 & ~n1833;
  assign n1835 = ~pi013 & n1608;
  assign n1836 = n1834 & ~n1835;
  assign n1837 = ~n1831 & n1836;
  assign n1838 = n1830 & n1837;
  assign n1839 = n1556 & n1838;
  assign n1840 = ~n1823 & ~n1839;
  assign n1841 = n1807 & n1840;
  assign n1842 = n1645 & n1841;
  assign n1843 = ~pi052 & n1616;
  assign n1844 = ~pi056 & n1619;
  assign n1845 = ~n1843 & ~n1844;
  assign n1846 = ~pi051 & n1614;
  assign n1847 = ~pi055 & n1622;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~pi049 & n1608;
  assign n1850 = ~pi050 & n1606;
  assign n1851 = ~n1849 & ~n1850;
  assign n1852 = ~pi054 & n1600;
  assign n1853 = ~pi053 & n1603;
  assign n1854 = ~n1852 & ~n1853;
  assign n1855 = n1851 & n1854;
  assign n1856 = n1848 & n1855;
  assign n1857 = n1845 & n1856;
  assign n1858 = n1556 & n1857;
  assign n1859 = ~n1556 & ~n1857;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1842 & n1860;
  assign n1862 = ~n1556 & ~n1822;
  assign n1863 = ~n1839 & n1862;
  assign n1864 = ~n1556 & ~n1838;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1556 & ~n1643;
  assign n1867 = ~n1556 & ~n1627;
  assign n1868 = ~n1644 & n1867;
  assign n1869 = ~n1866 & ~n1868;
  assign n1870 = ~n1556 & ~n1709;
  assign n1871 = ~n1694 & n1870;
  assign n1872 = ~n1556 & ~n1693;
  assign n1873 = ~n1871 & ~n1872;
  assign n1874 = n1678 & ~n1873;
  assign n1875 = ~n1556 & ~n1660;
  assign n1876 = ~n1556 & ~n1676;
  assign n1877 = ~n1661 & n1876;
  assign n1878 = ~n1875 & ~n1877;
  assign n1879 = ~n1874 & n1878;
  assign n1880 = n1645 & ~n1879;
  assign n1881 = n1869 & ~n1880;
  assign n1882 = n1840 & ~n1881;
  assign n1883 = n1865 & ~n1882;
  assign n1884 = n1861 & n1883;
  assign n1885 = ~n1842 & n1883;
  assign n1886 = ~n1860 & ~n1885;
  assign n1887 = ~n1884 & ~n1886;
  assign n1888 = ~n1839 & ~n1864;
  assign n1889 = ~n1823 & n1866;
  assign n1890 = ~n1862 & ~n1889;
  assign n1891 = ~n1644 & ~n1823;
  assign n1892 = ~n1628 & n1875;
  assign n1893 = ~n1867 & ~n1892;
  assign n1894 = ~n1628 & ~n1661;
  assign n1895 = ~n1677 & n1872;
  assign n1896 = ~n1876 & ~n1895;
  assign n1897 = ~n1710 & n1728;
  assign n1898 = ~n1870 & ~n1897;
  assign n1899 = ~n1677 & ~n1694;
  assign n1900 = ~n1898 & n1899;
  assign n1901 = n1896 & ~n1900;
  assign n1902 = n1894 & ~n1901;
  assign n1903 = n1893 & ~n1902;
  assign n1904 = n1891 & ~n1903;
  assign n1905 = ~n1780 & ~n1797;
  assign n1906 = ~n1800 & ~n1905;
  assign n1907 = ~n1748 & ~n1765;
  assign n1908 = ~n1906 & n1907;
  assign n1909 = ~n1748 & n1802;
  assign n1910 = ~n1745 & ~n1909;
  assign n1911 = ~n1908 & n1910;
  assign n1912 = ~n1710 & ~n1729;
  assign n1913 = ~n1911 & n1912;
  assign n1914 = n1891 & n1913;
  assign n1915 = n1899 & n1914;
  assign n1916 = n1894 & n1915;
  assign n1917 = ~n1904 & ~n1916;
  assign n1918 = n1890 & n1917;
  assign n1919 = n1888 & n1918;
  assign n1920 = ~n1888 & ~n1918;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = n1887 & n1921;
  assign n1923 = ~n1628 & ~n1867;
  assign n1924 = ~n1807 & n1879;
  assign n1925 = n1923 & n1924;
  assign n1926 = ~n1923 & ~n1924;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1823 & ~n1862;
  assign n1929 = ~n1798 & n1803;
  assign n1930 = n1749 & ~n1929;
  assign n1931 = n1711 & n1930;
  assign n1932 = n1711 & ~n1729;
  assign n1933 = ~n1728 & ~n1745;
  assign n1934 = n1932 & ~n1933;
  assign n1935 = n1873 & ~n1934;
  assign n1936 = ~n1931 & n1935;
  assign n1937 = n1645 & n1678;
  assign n1938 = ~n1936 & n1937;
  assign n1939 = n1645 & ~n1878;
  assign n1940 = n1869 & ~n1939;
  assign n1941 = ~n1938 & n1940;
  assign n1942 = n1928 & n1941;
  assign n1943 = ~n1928 & ~n1941;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = n1927 & n1944;
  assign n1946 = ~n1644 & ~n1866;
  assign n1947 = n1898 & ~n1913;
  assign n1948 = n1894 & n1899;
  assign n1949 = ~n1947 & n1948;
  assign n1950 = n1894 & ~n1896;
  assign n1951 = n1893 & ~n1950;
  assign n1952 = ~n1949 & n1951;
  assign n1953 = n1946 & n1952;
  assign n1954 = ~n1946 & ~n1952;
  assign n1955 = ~n1953 & ~n1954;
  assign n1956 = ~n1661 & ~n1875;
  assign n1957 = n1899 & n1912;
  assign n1958 = ~n1911 & n1957;
  assign n1959 = n1901 & ~n1958;
  assign n1960 = n1956 & n1959;
  assign n1961 = ~n1956 & ~n1959;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = n1955 & n1962;
  assign n1964 = n1945 & n1963;
  assign n1965 = ~n1765 & ~n1802;
  assign n1966 = ~n1906 & ~n1965;
  assign n1967 = n1906 & n1965;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = ~n1797 & ~n1800;
  assign n1970 = ~n1780 & ~n1969;
  assign n1971 = n1780 & n1969;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = n1968 & n1972;
  assign n1974 = pi044 & n1616;
  assign n1975 = pi043 & n1614;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = pi045 & n1603;
  assign n1978 = pi048 & n1600;
  assign n1979 = ~n1977 & ~n1978;
  assign n1980 = pi042 & n1606;
  assign n1981 = pi041 & n1608;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = pi047 & n1619;
  assign n1984 = pi046 & n1622;
  assign n1985 = ~n1983 & ~n1984;
  assign n1986 = n1982 & n1985;
  assign n1987 = n1979 & n1986;
  assign n1988 = n1976 & n1987;
  assign n1989 = n1556 & n1988;
  assign n1990 = ~n1556 & ~n1988;
  assign n1991 = ~n1989 & ~n1990;
  assign n1992 = ~pi006 & n1606;
  assign n1993 = ~pi011 & n1619;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = ~pi010 & n1622;
  assign n1996 = ~pi005 & n1608;
  assign n1997 = ~n1995 & ~n1996;
  assign n1998 = n1994 & n1997;
  assign n1999 = ~pi007 & n1614;
  assign n2000 = ~pi008 & n1616;
  assign n2001 = ~pi012 & n1600;
  assign n2002 = ~pi009 & n1603;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = ~n2000 & n2003;
  assign n2005 = ~n1999 & n2004;
  assign n2006 = n1998 & n2005;
  assign n2007 = n1556 & n2006;
  assign n2008 = ~n1858 & ~n2007;
  assign n2009 = ~n1865 & n2008;
  assign n2010 = n1556 & n2007;
  assign n2011 = ~n1857 & ~n2007;
  assign n2012 = n2006 & ~n2011;
  assign n2013 = ~n2010 & ~n2012;
  assign n2014 = ~n1556 & n2013;
  assign n2015 = ~n2009 & ~n2014;
  assign n2016 = n1840 & n2008;
  assign n2017 = ~n1941 & n2016;
  assign n2018 = n2015 & ~n2017;
  assign n2019 = ~n1991 & ~n2018;
  assign n2020 = n1991 & n2018;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = ~n1745 & ~n1748;
  assign n2023 = n1929 & n2022;
  assign n2024 = ~n1929 & ~n2022;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = n2021 & n2025;
  assign n2027 = n1973 & n2026;
  assign n2028 = n1964 & n2027;
  assign n2029 = n1922 & n2028;
  assign n2030 = ~n1556 & ~n2006;
  assign n2031 = ~n2007 & ~n2030;
  assign n2032 = ~n1839 & ~n1858;
  assign n2033 = ~n1890 & n2032;
  assign n2034 = n1891 & n2032;
  assign n2035 = n1949 & n2034;
  assign n2036 = ~n2033 & ~n2035;
  assign n2037 = ~n1858 & n1864;
  assign n2038 = ~n1951 & n2034;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = n2036 & n2039;
  assign n2041 = ~n1859 & n2040;
  assign n2042 = n2031 & n2041;
  assign n2043 = ~n2031 & ~n2041;
  assign n2044 = ~n2042 & ~n2043;
  assign n2045 = ~n1677 & ~n1876;
  assign n2046 = ~n1936 & ~n2045;
  assign n2047 = n1936 & n2045;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~n1710 & ~n1870;
  assign n2050 = n1806 & n2049;
  assign n2051 = ~n1806 & ~n2049;
  assign n2052 = ~n2050 & ~n2051;
  assign n2053 = n2048 & n2052;
  assign n2054 = ~n1694 & ~n1872;
  assign n2055 = n1947 & n2054;
  assign n2056 = ~n1947 & ~n2054;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = ~n1728 & ~n1729;
  assign n2059 = n1911 & n2058;
  assign n2060 = ~n1911 & ~n2058;
  assign n2061 = ~n2059 & ~n2060;
  assign n2062 = n2057 & n2061;
  assign n2063 = n2053 & n2062;
  assign n2064 = ~n1780 & n2063;
  assign n2065 = n2044 & n2064;
  assign n2066 = n949 & n2065;
  assign n2067 = n2029 & n2066;
  assign po034 = ~n1534 & ~n2067;
  assign n2069 = pi001 & pi247;
  assign n2070 = ~pi099 & n780;
  assign n2071 = pi361 & n785;
  assign n2072 = pi295 & n2071;
  assign n2073 = pi001 & ~n2071;
  assign n2074 = ~n2072 & ~n2073;
  assign n2075 = n2070 & ~n2074;
  assign n2076 = pi189 & ~pi190;
  assign n2077 = pi188 & n2076;
  assign n2078 = ~n780 & ~n2077;
  assign n2079 = ~pi296 & pi297;
  assign n2080 = pi291 & n2079;
  assign n2081 = pi300 & ~n2080;
  assign n2082 = pi299 & n2081;
  assign n2083 = ~pi300 & ~n2080;
  assign n2084 = pi299 & n2083;
  assign n2085 = ~n2082 & ~n2084;
  assign n2086 = ~n780 & ~n2085;
  assign n2087 = pi291 & ~pi296;
  assign n2088 = ~pi300 & n2087;
  assign n2089 = n830 & n2088;
  assign n2090 = n812 & n2089;
  assign n2091 = ~pi299 & ~pi300;
  assign n2092 = ~n2080 & n2091;
  assign n2093 = ~n780 & n2092;
  assign n2094 = ~n2090 & ~n2093;
  assign n2095 = pi300 & n2087;
  assign n2096 = n927 & n2095;
  assign n2097 = pi297 & n2087;
  assign n2098 = n1558 & n2097;
  assign n2099 = ~n2096 & ~n2098;
  assign n2100 = n812 & ~n2099;
  assign n2101 = n2091 & n2097;
  assign n2102 = n812 & n2101;
  assign n2103 = ~pi299 & n2081;
  assign n2104 = ~n780 & n2103;
  assign n2105 = ~n2102 & ~n2104;
  assign n2106 = ~n2100 & n2105;
  assign n2107 = n2094 & n2106;
  assign n2108 = ~n2086 & n2107;
  assign n2109 = pi294 & ~pi301;
  assign n2110 = ~n2108 & n2109;
  assign n2111 = ~pi299 & ~n2097;
  assign n2112 = pi300 & n2111;
  assign n2113 = ~n780 & n2112;
  assign n2114 = pi291 & ~pi298;
  assign n2115 = n877 & n927;
  assign n2116 = n2114 & n2115;
  assign n2117 = pi300 & pi302;
  assign n2118 = n883 & n2117;
  assign n2119 = n794 & n2118;
  assign n2120 = ~n2116 & ~n2119;
  assign n2121 = ~n780 & ~n2120;
  assign n2122 = ~n780 & ~n804;
  assign n2123 = n809 & n2122;
  assign n2124 = ~n780 & n804;
  assign n2125 = n866 & n2124;
  assign n2126 = ~n2122 & ~n2125;
  assign n2127 = n838 & ~n2126;
  assign n2128 = ~n2123 & ~n2127;
  assign n2129 = ~n2121 & n2128;
  assign n2130 = pi298 & ~pi299;
  assign n2131 = n823 & n2130;
  assign n2132 = n1525 & n2079;
  assign n2133 = n2131 & n2132;
  assign n2134 = n793 & n2130;
  assign n2135 = n820 & n2079;
  assign n2136 = n2134 & n2135;
  assign n2137 = n793 & n886;
  assign n2138 = n884 & n2137;
  assign n2139 = ~n2136 & ~n2138;
  assign n2140 = n830 & n837;
  assign n2141 = n2139 & ~n2140;
  assign n2142 = ~n2133 & n2141;
  assign n2143 = ~n780 & ~n2142;
  assign n2144 = n2129 & ~n2143;
  assign n2145 = ~pi300 & ~n850;
  assign n2146 = ~n2097 & n2145;
  assign n2147 = pi299 & n2146;
  assign n2148 = n793 & n822;
  assign n2149 = n820 & n821;
  assign n2150 = n2148 & n2149;
  assign n2151 = pi291 & ~pi303;
  assign n2152 = n2130 & n2151;
  assign n2153 = n820 & n883;
  assign n2154 = n2152 & n2153;
  assign n2155 = n789 & n2117;
  assign n2156 = n794 & n2155;
  assign n2157 = ~n2154 & ~n2156;
  assign n2158 = ~n2150 & n2157;
  assign n2159 = ~n2147 & n2158;
  assign n2160 = n1525 & n2151;
  assign n2161 = n2130 & n2160;
  assign n2162 = n883 & n2161;
  assign n2163 = n2118 & n2137;
  assign n2164 = ~n2162 & ~n2163;
  assign n2165 = n2159 & n2164;
  assign n2166 = ~n780 & ~n2165;
  assign n2167 = n2144 & ~n2166;
  assign n2168 = ~n2113 & n2167;
  assign n2169 = n2137 & n2155;
  assign n2170 = n824 & n2132;
  assign n2171 = ~n780 & n2170;
  assign n2172 = n904 & n2145;
  assign n2173 = n2087 & n2172;
  assign n2174 = ~n780 & n2173;
  assign n2175 = ~n2171 & ~n2174;
  assign n2176 = n2135 & n2148;
  assign n2177 = ~n780 & n2176;
  assign n2178 = ~pi303 & n877;
  assign n2179 = n876 & n2178;
  assign n2180 = ~n2177 & ~n2179;
  assign n2181 = n2175 & n2180;
  assign n2182 = n792 & n885;
  assign n2183 = ~n780 & n2182;
  assign n2184 = n886 & n2118;
  assign n2185 = n823 & n2184;
  assign n2186 = ~n780 & n2185;
  assign n2187 = ~n2183 & ~n2186;
  assign n2188 = n2181 & n2187;
  assign n2189 = ~n2169 & n2188;
  assign n2190 = ~n780 & n873;
  assign n2191 = ~pi297 & n875;
  assign n2192 = n2178 & n2191;
  assign n2193 = n798 & n830;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = ~n780 & ~n2194;
  assign n2196 = n878 & n2191;
  assign n2197 = n789 & n2161;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = n812 & ~n2198;
  assign n2200 = ~n2195 & ~n2199;
  assign n2201 = ~n780 & n817;
  assign n2202 = n2131 & n2149;
  assign n2203 = n2122 & n2202;
  assign n2204 = ~n2201 & ~n2203;
  assign n2205 = ~n780 & ~n1546;
  assign n2206 = ~n804 & n2205;
  assign n2207 = n887 & n2206;
  assign n2208 = n2204 & ~n2207;
  assign n2209 = n2200 & n2208;
  assign n2210 = ~n2190 & n2209;
  assign n2211 = n2189 & n2210;
  assign n2212 = n794 & n884;
  assign n2213 = ~n780 & n2212;
  assign n2214 = n792 & n2118;
  assign n2215 = n823 & n2214;
  assign n2216 = ~n780 & n2215;
  assign n2217 = ~n2213 & ~n2216;
  assign n2218 = pi291 & pi303;
  assign n2219 = n791 & n2218;
  assign n2220 = n886 & n2219;
  assign n2221 = ~n780 & n2220;
  assign n2222 = n830 & n2087;
  assign n2223 = n2145 & n2222;
  assign n2224 = ~n780 & n2223;
  assign n2225 = n2087 & n2145;
  assign n2226 = n927 & n2225;
  assign n2227 = ~n780 & n2226;
  assign n2228 = ~n780 & n833;
  assign n2229 = ~n780 & n2122;
  assign n2230 = n1527 & n2229;
  assign n2231 = ~n879 & ~n2230;
  assign n2232 = ~n2228 & n2231;
  assign n2233 = ~n2227 & n2232;
  assign n2234 = ~n2224 & n2233;
  assign n2235 = ~n2221 & n2234;
  assign n2236 = n1526 & n2152;
  assign n2237 = n812 & n2236;
  assign n2238 = n2131 & n2135;
  assign n2239 = ~n780 & n2238;
  assign n2240 = ~n2237 & ~n2239;
  assign n2241 = n2132 & n2152;
  assign n2242 = ~n780 & n2241;
  assign n2243 = n1526 & n2134;
  assign n2244 = n2122 & n2243;
  assign n2245 = ~n2242 & ~n2244;
  assign n2246 = n2240 & n2245;
  assign n2247 = n2235 & n2246;
  assign n2248 = n2217 & n2247;
  assign n2249 = pi291 & n2172;
  assign n2250 = pi296 & n2249;
  assign n2251 = ~n780 & n2250;
  assign n2252 = n837 & n927;
  assign n2253 = ~n780 & n2252;
  assign n2254 = n824 & n2135;
  assign n2255 = ~n780 & n2254;
  assign n2256 = n2132 & n2148;
  assign n2257 = ~n780 & n2256;
  assign n2258 = ~n2255 & ~n2257;
  assign n2259 = ~n2253 & n2258;
  assign n2260 = ~n2251 & n2259;
  assign n2261 = n2248 & n2260;
  assign n2262 = n2130 & n2153;
  assign n2263 = n2218 & n2262;
  assign n2264 = n883 & n2218;
  assign n2265 = n2130 & n2264;
  assign n2266 = n1525 & n2265;
  assign n2267 = ~n2263 & ~n2266;
  assign n2268 = ~n780 & ~n2267;
  assign n2269 = n813 & n2155;
  assign n2270 = pi303 & n2269;
  assign n2271 = n791 & n2137;
  assign n2272 = ~n2270 & ~n2271;
  assign n2273 = ~n780 & ~n2272;
  assign n2274 = n1526 & n2131;
  assign n2275 = n2122 & n2274;
  assign n2276 = ~n2273 & ~n2275;
  assign n2277 = ~n2268 & n2276;
  assign n2278 = n2132 & n2151;
  assign n2279 = n886 & n2278;
  assign n2280 = n2132 & n2134;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = ~n780 & ~n2281;
  assign n2283 = pi298 & ~pi300;
  assign n2284 = pi302 & n2283;
  assign n2285 = n871 & n2284;
  assign n2286 = ~n2097 & n2285;
  assign n2287 = ~n780 & n2286;
  assign n2288 = n1526 & n2148;
  assign n2289 = n2134 & n2149;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = n2122 & ~n2290;
  assign n2292 = ~n780 & ~n800;
  assign n2293 = ~n2291 & ~n2292;
  assign n2294 = ~n780 & n827;
  assign n2295 = ~n804 & n812;
  assign n2296 = ~n780 & n2295;
  assign n2297 = ~n827 & n2296;
  assign n2298 = ~n2294 & ~n2297;
  assign n2299 = n826 & ~n2298;
  assign n2300 = n2293 & ~n2299;
  assign n2301 = ~n2287 & n2300;
  assign n2302 = ~n2282 & n2301;
  assign n2303 = n2277 & n2302;
  assign n2304 = n2261 & n2303;
  assign n2305 = n2211 & n2304;
  assign n2306 = n2168 & n2305;
  assign n2307 = n787 & ~n2306;
  assign n2308 = pi297 & ~pi302;
  assign n2309 = pi299 & pi303;
  assign n2310 = n2308 & n2309;
  assign n2311 = pi291 & n877;
  assign n2312 = pi298 & n2311;
  assign n2313 = n2310 & n2312;
  assign n2314 = n2122 & n2313;
  assign n2315 = pi291 & ~pi299;
  assign n2316 = ~n822 & ~n2315;
  assign n2317 = ~n1558 & n2316;
  assign n2318 = ~n2091 & n2317;
  assign n2319 = ~n780 & ~n2318;
  assign n2320 = pi302 & n830;
  assign n2321 = pi298 & ~pi303;
  assign n2322 = ~n807 & ~n2321;
  assign n2323 = pi296 & ~pi298;
  assign n2324 = ~pi296 & pi298;
  assign n2325 = ~n2323 & ~n2324;
  assign n2326 = pi291 & ~pi300;
  assign n2327 = n2325 & n2326;
  assign n2328 = ~n2322 & n2327;
  assign n2329 = n2320 & n2328;
  assign n2330 = ~n780 & n2329;
  assign n2331 = ~n780 & n909;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = ~n2319 & n2332;
  assign n2334 = ~n2314 & n2333;
  assign n2335 = ~pi291 & n877;
  assign n2336 = ~pi303 & n2335;
  assign n2337 = n830 & n2336;
  assign n2338 = ~n780 & n2337;
  assign n2339 = ~pi296 & ~pi300;
  assign n2340 = n814 & n2339;
  assign n2341 = ~n780 & n2340;
  assign n2342 = pi303 & n2335;
  assign n2343 = n830 & n2342;
  assign n2344 = ~n780 & n2343;
  assign n2345 = pi297 & pi302;
  assign n2346 = n2326 & n2345;
  assign n2347 = n886 & n2346;
  assign n2348 = pi303 & n2347;
  assign n2349 = ~n780 & n2348;
  assign n2350 = ~n2344 & ~n2349;
  assign n2351 = ~n2341 & n2350;
  assign n2352 = ~n2338 & n2351;
  assign n2353 = ~pi291 & n2339;
  assign n2354 = ~pi303 & n830;
  assign n2355 = n2353 & n2354;
  assign n2356 = n812 & n2355;
  assign n2357 = pi299 & n870;
  assign n2358 = n877 & n2357;
  assign n2359 = ~n780 & n2358;
  assign n2360 = n2339 & n2357;
  assign n2361 = ~n780 & n2360;
  assign n2362 = ~n2359 & ~n2361;
  assign n2363 = n871 & n2308;
  assign n2364 = n2312 & n2363;
  assign n2365 = n2122 & n2364;
  assign n2366 = n2362 & ~n2365;
  assign n2367 = ~pi188 & n2076;
  assign n2368 = ~n780 & ~n2367;
  assign n2369 = ~n804 & n2368;
  assign n2370 = ~n906 & n2369;
  assign n2371 = n2366 & ~n2370;
  assign n2372 = ~n2356 & n2371;
  assign n2373 = ~n780 & n929;
  assign n2374 = n2368 & n2373;
  assign n2375 = pi303 & n830;
  assign n2376 = n2353 & n2375;
  assign n2377 = n812 & n2376;
  assign n2378 = ~pi303 & n2346;
  assign n2379 = ~pi296 & n2378;
  assign n2380 = pi299 & n2379;
  assign n2381 = ~n780 & n2380;
  assign n2382 = ~pi302 & n2326;
  assign n2383 = ~pi296 & n2382;
  assign n2384 = n830 & n2383;
  assign n2385 = ~n780 & n2384;
  assign n2386 = n932 & n2369;
  assign n2387 = ~n2385 & ~n2386;
  assign n2388 = ~n2381 & n2387;
  assign n2389 = ~n2377 & n2388;
  assign n2390 = ~n2374 & n2389;
  assign n2391 = n2372 & n2390;
  assign n2392 = n2352 & n2391;
  assign n2393 = n2334 & n2392;
  assign n2394 = pi301 & ~n2393;
  assign n2395 = ~n2307 & ~n2394;
  assign n2396 = ~n2110 & n2395;
  assign n2397 = ~n2077 & ~n2396;
  assign n2398 = ~n2078 & ~n2397;
  assign n2399 = pi098 & ~n2398;
  assign n2400 = ~pi098 & n2398;
  assign n2401 = ~n2399 & ~n2400;
  assign n2402 = n2240 & ~n2251;
  assign n2403 = ~n2242 & n2402;
  assign n2404 = n780 & ~n804;
  assign n2405 = n2243 & ~n2404;
  assign n2406 = n2403 & ~n2405;
  assign n2407 = ~n2253 & n2406;
  assign n2408 = ~n2255 & n2407;
  assign n2409 = ~n2257 & n2408;
  assign n2410 = ~n1527 & n2409;
  assign n2411 = ~n2213 & ~n2221;
  assign n2412 = n2410 & n2411;
  assign n2413 = ~n2227 & n2412;
  assign n2414 = ~n2216 & n2413;
  assign n2415 = ~n833 & ~n2224;
  assign n2416 = n2414 & n2415;
  assign n2417 = n2175 & ~n2177;
  assign n2418 = n2416 & n2417;
  assign n2419 = n2144 & n2418;
  assign n2420 = n2200 & n2419;
  assign n2421 = ~n1546 & ~n2206;
  assign n2422 = n887 & ~n2421;
  assign n2423 = n2202 & ~n2404;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2166 & n2424;
  assign n2426 = ~n817 & n2425;
  assign n2427 = ~n2186 & ~n2190;
  assign n2428 = ~n2113 & ~n2183;
  assign n2429 = n2274 & ~n2404;
  assign n2430 = ~n2273 & ~n2429;
  assign n2431 = ~n2268 & n2430;
  assign n2432 = n2428 & n2431;
  assign n2433 = n2427 & n2432;
  assign n2434 = n2426 & n2433;
  assign n2435 = ~n780 & ~n2296;
  assign n2436 = ~n827 & ~n2435;
  assign n2437 = ~n2294 & ~n2436;
  assign n2438 = n826 & ~n2437;
  assign n2439 = n2289 & ~n2404;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = n2288 & ~n2404;
  assign n2442 = ~n799 & ~n2441;
  assign n2443 = n2440 & n2442;
  assign n2444 = ~n2282 & n2443;
  assign n2445 = n2434 & n2444;
  assign n2446 = ~n795 & n2445;
  assign n2447 = ~n2287 & n2446;
  assign n2448 = n2420 & n2447;
  assign n2449 = n787 & ~n2448;
  assign n2450 = n877 & n2114;
  assign n2451 = n2310 & n2450;
  assign n2452 = ~n2330 & ~n2451;
  assign n2453 = ~n2319 & n2452;
  assign n2454 = ~n2331 & n2453;
  assign n2455 = ~n2367 & ~n2369;
  assign n2456 = n932 & ~n2455;
  assign n2457 = n2454 & ~n2456;
  assign n2458 = ~n2344 & ~n2381;
  assign n2459 = n2457 & n2458;
  assign n2460 = ~n2377 & n2459;
  assign n2461 = ~n929 & n2460;
  assign n2462 = ~n2338 & ~n2349;
  assign n2463 = ~n2385 & n2462;
  assign n2464 = ~n2341 & n2463;
  assign n2465 = n2461 & n2464;
  assign n2466 = n2363 & n2450;
  assign n2467 = n2465 & ~n2466;
  assign n2468 = ~n2314 & n2467;
  assign n2469 = ~n804 & n2455;
  assign n2470 = ~n906 & ~n2469;
  assign n2471 = n2345 & n2450;
  assign n2472 = n871 & n2471;
  assign n2473 = n2309 & n2450;
  assign n2474 = n2345 & n2473;
  assign n2475 = ~n2472 & ~n2474;
  assign n2476 = ~n2470 & n2475;
  assign n2477 = n2362 & n2476;
  assign n2478 = ~n2365 & n2477;
  assign n2479 = ~n2356 & n2478;
  assign n2480 = n2468 & n2479;
  assign n2481 = pi301 & ~n2480;
  assign n2482 = ~n2110 & ~n2481;
  assign n2483 = ~n2449 & n2482;
  assign n2484 = ~n2077 & ~n2483;
  assign n2485 = ~n2078 & ~n2484;
  assign n2486 = pi097 & ~n2485;
  assign n2487 = ~pi097 & n2485;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n780 & n2103;
  assign n2490 = n780 & n2084;
  assign n2491 = ~n2096 & ~n2101;
  assign n2492 = ~n2098 & n2491;
  assign n2493 = ~n2089 & n2492;
  assign n2494 = ~n812 & ~n2493;
  assign n2495 = ~n2082 & ~n2092;
  assign n2496 = n780 & ~n2495;
  assign n2497 = ~n2494 & ~n2496;
  assign n2498 = ~n2490 & n2497;
  assign n2499 = ~n2489 & n2498;
  assign n2500 = n2109 & ~n2499;
  assign n2501 = ~n2122 & n2364;
  assign n2502 = ~n812 & n2355;
  assign n2503 = ~n2501 & ~n2502;
  assign n2504 = n780 & n2360;
  assign n2505 = n2503 & ~n2504;
  assign n2506 = n780 & n2358;
  assign n2507 = n780 & n2343;
  assign n2508 = n929 & ~n2368;
  assign n2509 = ~n2507 & ~n2508;
  assign n2510 = ~n909 & ~n2380;
  assign n2511 = n780 & ~n2510;
  assign n2512 = n2509 & ~n2511;
  assign n2513 = ~n812 & n2376;
  assign n2514 = n780 & ~n2318;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n780 & n2329;
  assign n2517 = n2515 & ~n2516;
  assign n2518 = ~n2451 & n2517;
  assign n2519 = n932 & ~n2369;
  assign n2520 = ~n2122 & n2313;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n2518 & n2521;
  assign n2523 = ~n2466 & n2522;
  assign n2524 = n2512 & n2523;
  assign n2525 = ~n2337 & ~n2348;
  assign n2526 = ~n2340 & ~n2384;
  assign n2527 = n2525 & n2526;
  assign n2528 = n780 & ~n2527;
  assign n2529 = n2524 & ~n2528;
  assign n2530 = ~n906 & ~n2369;
  assign n2531 = n2475 & ~n2530;
  assign n2532 = n2529 & n2531;
  assign n2533 = ~n2506 & n2532;
  assign n2534 = n2505 & n2533;
  assign n2535 = pi301 & ~n2534;
  assign n2536 = ~n2500 & ~n2535;
  assign n2537 = n780 & n2193;
  assign n2538 = ~n812 & n2197;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = n780 & n2173;
  assign n2541 = ~n812 & n2196;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = ~n833 & ~n2215;
  assign n2544 = ~n2212 & n2543;
  assign n2545 = n780 & ~n2544;
  assign n2546 = ~n879 & ~n2545;
  assign n2547 = ~n817 & ~n873;
  assign n2548 = ~n2185 & n2547;
  assign n2549 = n780 & ~n2548;
  assign n2550 = n2546 & ~n2549;
  assign n2551 = ~n2169 & n2550;
  assign n2552 = n887 & ~n2206;
  assign n2553 = ~n2122 & n2202;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = n1527 & ~n2229;
  assign n2556 = n780 & n2223;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = ~n2220 & ~n2226;
  assign n2559 = n780 & ~n2558;
  assign n2560 = n2557 & ~n2559;
  assign n2561 = ~n2112 & ~n2182;
  assign n2562 = n780 & ~n2561;
  assign n2563 = n2560 & ~n2562;
  assign n2564 = n2554 & n2563;
  assign n2565 = n2551 & n2564;
  assign n2566 = n780 & n2170;
  assign n2567 = ~n2176 & ~n2192;
  assign n2568 = n780 & ~n2567;
  assign n2569 = ~n2179 & ~n2568;
  assign n2570 = ~n2566 & n2569;
  assign n2571 = ~n2238 & ~n2241;
  assign n2572 = ~n2256 & n2571;
  assign n2573 = n780 & ~n2572;
  assign n2574 = n780 & n2254;
  assign n2575 = n780 & n2252;
  assign n2576 = ~n2122 & n2243;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = n780 & n2250;
  assign n2579 = ~n812 & n2236;
  assign n2580 = ~n2578 & ~n2579;
  assign n2581 = n2577 & n2580;
  assign n2582 = ~n2574 & n2581;
  assign n2583 = ~n2573 & n2582;
  assign n2584 = n2570 & n2583;
  assign n2585 = n2565 & n2584;
  assign n2586 = n2542 & n2585;
  assign n2587 = n2539 & n2586;
  assign n2588 = n780 & ~n2165;
  assign n2589 = n780 & ~n2272;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = n780 & ~n2267;
  assign n2592 = ~n2122 & n2274;
  assign n2593 = ~n2591 & ~n2592;
  assign n2594 = n780 & n2286;
  assign n2595 = ~n2122 & n2288;
  assign n2596 = ~n2594 & ~n2595;
  assign n2597 = n800 & n2281;
  assign n2598 = n780 & ~n2597;
  assign n2599 = n780 & n2295;
  assign n2600 = ~n804 & ~n2599;
  assign n2601 = n812 & n2600;
  assign n2602 = pi196 & ~n2601;
  assign n2603 = ~pi195 & n780;
  assign n2604 = pi195 & ~n2601;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = ~pi196 & ~n2605;
  assign n2607 = ~n2602 & ~n2606;
  assign n2608 = n826 & ~n2607;
  assign n2609 = ~n2122 & n2289;
  assign n2610 = ~n2608 & ~n2609;
  assign n2611 = ~n2598 & n2610;
  assign n2612 = n2596 & n2611;
  assign n2613 = n780 & ~n2142;
  assign n2614 = n2612 & ~n2613;
  assign n2615 = n809 & ~n2122;
  assign n2616 = ~n780 & ~n867;
  assign n2617 = n838 & ~n2616;
  assign n2618 = ~n2615 & ~n2617;
  assign n2619 = n780 & ~n2120;
  assign n2620 = n2618 & ~n2619;
  assign n2621 = n2614 & n2620;
  assign n2622 = n2593 & n2621;
  assign n2623 = n2590 & n2622;
  assign n2624 = n2587 & n2623;
  assign n2625 = n787 & ~n2624;
  assign n2626 = n2536 & ~n2625;
  assign n2627 = n780 & ~n2626;
  assign n2628 = ~n2077 & ~n2627;
  assign n2629 = ~pi099 & n2628;
  assign n2630 = pi099 & ~n2628;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = ~n2488 & ~n2631;
  assign n2633 = ~n2401 & n2632;
  assign n2634 = pi301 & n804;
  assign n2635 = n909 & n2634;
  assign n2636 = pi195 & ~pi196;
  assign n2637 = n1546 & n2636;
  assign n2638 = n826 & n2637;
  assign n2639 = n799 & n804;
  assign n2640 = ~n2638 & ~n2639;
  assign n2641 = n867 & n2193;
  assign n2642 = n2640 & ~n2641;
  assign n2643 = ~n795 & ~n2182;
  assign n2644 = n804 & ~n2643;
  assign n2645 = n2642 & ~n2644;
  assign n2646 = n787 & ~n2645;
  assign n2647 = ~n2635 & ~n2646;
  assign n2648 = n787 & n789;
  assign n2649 = n793 & n1560;
  assign n2650 = n2648 & n2649;
  assign n2651 = pi331 & ~pi333;
  assign n2652 = n804 & n2651;
  assign n2653 = pi195 & n2652;
  assign n2654 = ~pi277 & ~pi346;
  assign n2655 = pi285 & n2654;
  assign n2656 = pi155 & n2655;
  assign n2657 = pi277 & ~pi346;
  assign n2658 = ~pi285 & n2657;
  assign n2659 = pi156 & n2658;
  assign n2660 = ~n2656 & ~n2659;
  assign n2661 = ~pi285 & n2654;
  assign n2662 = pi154 & n2661;
  assign n2663 = pi277 & pi346;
  assign n2664 = pi285 & n2663;
  assign n2665 = pi160 & n2664;
  assign n2666 = ~n2662 & ~n2665;
  assign n2667 = ~pi277 & pi346;
  assign n2668 = pi285 & n2667;
  assign n2669 = pi158 & n2668;
  assign n2670 = ~pi285 & n2663;
  assign n2671 = pi159 & n2670;
  assign n2672 = ~n2669 & ~n2671;
  assign n2673 = pi285 & n2657;
  assign n2674 = pi157 & n2673;
  assign n2675 = ~pi285 & n2667;
  assign n2676 = pi127 & n2675;
  assign n2677 = ~n2674 & ~n2676;
  assign n2678 = n2672 & n2677;
  assign n2679 = n2666 & n2678;
  assign n2680 = n2660 & n2679;
  assign n2681 = pi188 & pi190;
  assign n2682 = ~pi189 & ~n2681;
  assign n2683 = ~pi188 & ~pi190;
  assign n2684 = n2682 & ~n2683;
  assign n2685 = n909 & ~n2684;
  assign n2686 = ~n811 & n929;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = ~n2329 & ~n2376;
  assign n2689 = ~n2313 & n2688;
  assign n2690 = ~n780 & n932;
  assign n2691 = n2318 & ~n2690;
  assign n2692 = n2689 & n2691;
  assign n2693 = n2687 & n2692;
  assign n2694 = ~n2380 & ~n2384;
  assign n2695 = ~n2348 & ~n2466;
  assign n2696 = n2694 & n2695;
  assign n2697 = n2693 & n2696;
  assign n2698 = ~n2343 & ~n2451;
  assign n2699 = ~n2337 & ~n2340;
  assign n2700 = n2698 & n2699;
  assign n2701 = ~n811 & n901;
  assign n2702 = n2475 & ~n2701;
  assign n2703 = n2700 & n2702;
  assign n2704 = n2697 & n2703;
  assign n2705 = ~n905 & ~n2364;
  assign n2706 = n2362 & n2705;
  assign n2707 = ~n2355 & n2706;
  assign n2708 = n2704 & n2707;
  assign n2709 = pi301 & ~n2708;
  assign n2710 = n805 & n809;
  assign n2711 = ~n2138 & ~n2140;
  assign n2712 = ~n2133 & ~n2136;
  assign n2713 = n2711 & n2712;
  assign n2714 = n804 & n866;
  assign n2715 = ~n805 & ~n2714;
  assign n2716 = n838 & ~n2715;
  assign n2717 = ~n811 & n2119;
  assign n2718 = ~n2716 & ~n2717;
  assign n2719 = ~n2116 & n2718;
  assign n2720 = n2713 & n2719;
  assign n2721 = ~n2710 & n2720;
  assign n2722 = ~n811 & n2215;
  assign n2723 = ~n879 & ~n2722;
  assign n2724 = n833 & ~n2684;
  assign n2725 = ~n2250 & ~n2724;
  assign n2726 = n2723 & n2725;
  assign n2727 = ~n2226 & n2258;
  assign n2728 = n2726 & n2727;
  assign n2729 = ~n2223 & n2728;
  assign n2730 = ~n2238 & ~n2252;
  assign n2731 = ~n2236 & ~n2241;
  assign n2732 = n2730 & n2731;
  assign n2733 = n2729 & n2732;
  assign n2734 = n2721 & n2733;
  assign n2735 = ~n2171 & ~n2177;
  assign n2736 = ~n2173 & ~n2192;
  assign n2737 = ~n2193 & n2736;
  assign n2738 = ~n2179 & n2737;
  assign n2739 = ~n1527 & n2738;
  assign n2740 = n2735 & n2739;
  assign n2741 = ~n2212 & ~n2220;
  assign n2742 = ~n2243 & n2741;
  assign n2743 = n2740 & n2742;
  assign n2744 = n2734 & n2743;
  assign n2745 = n2198 & n2744;
  assign n2746 = ~n2547 & ~n2684;
  assign n2747 = ~n2182 & ~n2746;
  assign n2748 = pi189 & ~n2683;
  assign n2749 = ~pi189 & ~pi190;
  assign n2750 = ~pi188 & n2749;
  assign n2751 = ~n2748 & ~n2750;
  assign n2752 = n887 & ~n2751;
  assign n2753 = n2159 & ~n2752;
  assign n2754 = ~n2169 & ~n2202;
  assign n2755 = ~n2112 & n2754;
  assign n2756 = n2753 & n2755;
  assign n2757 = n2747 & n2756;
  assign n2758 = ~n2185 & n2757;
  assign n2759 = n2267 & ~n2274;
  assign n2760 = n2164 & n2759;
  assign n2761 = ~n2271 & n2760;
  assign n2762 = ~n2270 & n2761;
  assign n2763 = n2758 & n2762;
  assign n2764 = ~n827 & n2684;
  assign n2765 = n826 & ~n2764;
  assign n2766 = n795 & ~n2684;
  assign n2767 = n780 & n866;
  assign n2768 = ~n812 & ~n2767;
  assign n2769 = n799 & ~n2768;
  assign n2770 = ~n2766 & ~n2769;
  assign n2771 = ~n2765 & n2770;
  assign n2772 = ~n2280 & n2290;
  assign n2773 = ~n2279 & n2772;
  assign n2774 = ~n2286 & n2773;
  assign n2775 = n2771 & n2774;
  assign n2776 = n2763 & n2775;
  assign n2777 = n2745 & n2776;
  assign n2778 = n787 & ~n2777;
  assign n2779 = ~n2709 & ~n2778;
  assign n2780 = ~n2109 & n2779;
  assign n2781 = ~n2109 & n2681;
  assign n2782 = pi189 & n2781;
  assign n2783 = ~n2077 & ~n2782;
  assign n2784 = n2780 & n2783;
  assign n2785 = pi189 & n2681;
  assign n2786 = ~n2109 & n2785;
  assign n2787 = ~pi291 & pi297;
  assign n2788 = pi296 & n2787;
  assign n2789 = n1353 & n2788;
  assign n2790 = n1558 & n2789;
  assign n2791 = pi303 & n2790;
  assign n2792 = pi291 & pi297;
  assign n2793 = ~pi296 & n2792;
  assign n2794 = n849 & n2793;
  assign n2795 = n2091 & n2794;
  assign n2796 = ~pi303 & n2795;
  assign n2797 = ~n2791 & ~n2796;
  assign n2798 = n2077 & ~n2797;
  assign n2799 = pi190 & n888;
  assign n2800 = n2089 & ~n2799;
  assign n2801 = ~pi190 & ~n788;
  assign n2802 = ~n802 & ~n2801;
  assign n2803 = ~n804 & n2802;
  assign n2804 = n2096 & ~n2803;
  assign n2805 = ~n2800 & ~n2804;
  assign n2806 = ~n2082 & ~n2103;
  assign n2807 = ~n2084 & ~n2092;
  assign n2808 = n2806 & n2807;
  assign n2809 = n2805 & n2808;
  assign n2810 = ~n2098 & ~n2101;
  assign n2811 = ~n2803 & ~n2810;
  assign n2812 = n2809 & ~n2811;
  assign n2813 = n2109 & ~n2812;
  assign n2814 = ~n879 & ~n2224;
  assign n2815 = ~n2226 & n2741;
  assign n2816 = ~n1527 & n2543;
  assign n2817 = n2815 & n2816;
  assign n2818 = n2814 & n2817;
  assign n2819 = ~n811 & n2241;
  assign n2820 = n2236 & ~n2684;
  assign n2821 = n2258 & ~n2820;
  assign n2822 = ~n2819 & n2821;
  assign n2823 = n2159 & n2762;
  assign n2824 = ~n2238 & ~n2243;
  assign n2825 = ~n2250 & n2824;
  assign n2826 = ~n2253 & n2825;
  assign n2827 = ~n809 & ~n838;
  assign n2828 = n2197 & ~n2684;
  assign n2829 = ~n2171 & ~n2828;
  assign n2830 = ~n2173 & n2829;
  assign n2831 = ~n2140 & n2830;
  assign n2832 = ~n2177 & n2831;
  assign n2833 = n2827 & n2832;
  assign n2834 = ~n2119 & n2833;
  assign n2835 = ~n2116 & ~n2193;
  assign n2836 = ~n2196 & n2835;
  assign n2837 = ~n2179 & n2836;
  assign n2838 = n2834 & n2837;
  assign n2839 = ~n2133 & ~n2192;
  assign n2840 = n2838 & n2839;
  assign n2841 = n2139 & n2840;
  assign n2842 = n2826 & n2841;
  assign n2843 = n2823 & n2842;
  assign n2844 = n2822 & n2843;
  assign n2845 = n2818 & n2844;
  assign n2846 = ~n2185 & ~n2279;
  assign n2847 = ~n2112 & ~n2287;
  assign n2848 = ~n799 & n2847;
  assign n2849 = ~n887 & n2848;
  assign n2850 = n2290 & n2849;
  assign n2851 = ~n2202 & n2850;
  assign n2852 = ~n795 & n2851;
  assign n2853 = ~n2280 & n2547;
  assign n2854 = ~n2169 & n2853;
  assign n2855 = n2852 & n2854;
  assign n2856 = ~n826 & ~n2182;
  assign n2857 = n2855 & n2856;
  assign n2858 = n2846 & n2857;
  assign n2859 = n2845 & n2858;
  assign n2860 = n787 & ~n2859;
  assign n2861 = n932 & ~n2684;
  assign n2862 = ~n909 & n2698;
  assign n2863 = ~n788 & n2313;
  assign n2864 = n929 & ~n2684;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = n2318 & n2865;
  assign n2867 = n2694 & n2866;
  assign n2868 = n2688 & n2867;
  assign n2869 = n2862 & n2868;
  assign n2870 = ~n2861 & n2869;
  assign n2871 = n2695 & n2870;
  assign n2872 = n2699 & n2871;
  assign n2873 = ~n788 & n2364;
  assign n2874 = ~n780 & n905;
  assign n2875 = ~n2873 & ~n2874;
  assign n2876 = n901 & ~n2684;
  assign n2877 = n2875 & ~n2876;
  assign n2878 = ~n2355 & ~n2361;
  assign n2879 = ~n2359 & n2878;
  assign n2880 = ~n2474 & n2879;
  assign n2881 = ~n2472 & n2880;
  assign n2882 = n2877 & n2881;
  assign n2883 = n2872 & n2882;
  assign n2884 = pi301 & ~n2883;
  assign n2885 = ~n2860 & ~n2884;
  assign n2886 = ~n2813 & n2885;
  assign n2887 = ~n2077 & ~n2886;
  assign n2888 = ~n2798 & ~n2887;
  assign n2889 = ~n2786 & ~n2888;
  assign n2890 = n2784 & ~n2889;
  assign n2891 = ~n2680 & n2890;
  assign n2892 = ~n780 & n901;
  assign n2893 = n2318 & ~n2861;
  assign n2894 = ~n2451 & n2893;
  assign n2895 = ~n2892 & n2894;
  assign n2896 = n805 & n2337;
  assign n2897 = n2475 & n2875;
  assign n2898 = ~n2896 & n2897;
  assign n2899 = ~n2359 & n2898;
  assign n2900 = n2895 & n2899;
  assign n2901 = n805 & n2343;
  assign n2902 = n2865 & ~n2901;
  assign n2903 = ~n909 & n2902;
  assign n2904 = n2688 & n2696;
  assign n2905 = ~n2340 & n2904;
  assign n2906 = n2878 & n2905;
  assign n2907 = n2903 & n2906;
  assign n2908 = n2900 & n2907;
  assign n2909 = pi301 & ~n2908;
  assign n2910 = ~n2813 & ~n2909;
  assign n2911 = ~n2202 & ~n2289;
  assign n2912 = ~n826 & ~n2112;
  assign n2913 = ~n804 & n2280;
  assign n2914 = n2912 & ~n2913;
  assign n2915 = ~n2287 & n2914;
  assign n2916 = ~n817 & ~n2169;
  assign n2917 = ~n2182 & ~n2288;
  assign n2918 = n2846 & n2917;
  assign n2919 = ~n873 & ~n887;
  assign n2920 = n2918 & n2919;
  assign n2921 = n2916 & n2920;
  assign n2922 = n2915 & n2921;
  assign n2923 = n2823 & n2922;
  assign n2924 = n800 & n2923;
  assign n2925 = n2911 & n2924;
  assign n2926 = ~n1527 & n2180;
  assign n2927 = ~n2212 & n2926;
  assign n2928 = n2814 & n2927;
  assign n2929 = ~n2250 & ~n2256;
  assign n2930 = ~n2243 & n2929;
  assign n2931 = ~n2253 & n2930;
  assign n2932 = n805 & n2238;
  assign n2933 = n2931 & ~n2932;
  assign n2934 = ~n2255 & n2933;
  assign n2935 = ~n2819 & n2934;
  assign n2936 = ~n2820 & n2935;
  assign n2937 = ~n2722 & n2936;
  assign n2938 = ~n833 & n2558;
  assign n2939 = n2827 & ~n2828;
  assign n2940 = n2938 & n2939;
  assign n2941 = ~n2170 & ~n2196;
  assign n2942 = n2737 & n2941;
  assign n2943 = n2940 & n2942;
  assign n2944 = n805 & n2136;
  assign n2945 = ~n804 & n2133;
  assign n2946 = ~n2944 & ~n2945;
  assign n2947 = n2711 & n2946;
  assign n2948 = ~n2717 & n2947;
  assign n2949 = ~n2116 & n2948;
  assign n2950 = n2943 & n2949;
  assign n2951 = n2937 & n2950;
  assign n2952 = n2928 & n2951;
  assign n2953 = n2925 & n2952;
  assign n2954 = n787 & ~n2953;
  assign n2955 = n2910 & ~n2954;
  assign n2956 = ~n2077 & ~n2955;
  assign n2957 = ~n2798 & ~n2956;
  assign n2958 = ~n2786 & ~n2957;
  assign n2959 = n2784 & n2889;
  assign n2960 = ~n2958 & n2959;
  assign n2961 = pi349 & n2960;
  assign n2962 = n2958 & n2959;
  assign n2963 = pi130 & n2962;
  assign n2964 = ~n2961 & ~n2963;
  assign n2965 = ~n2784 & ~n2958;
  assign n2966 = ~n2889 & n2965;
  assign n2967 = n849 & n2151;
  assign n2968 = n2079 & n2967;
  assign n2969 = n780 & n2968;
  assign n2970 = n2091 & n2969;
  assign n2971 = n883 & n1558;
  assign n2972 = n780 & n1353;
  assign n2973 = n793 & n2972;
  assign n2974 = n2971 & n2973;
  assign n2975 = ~n2966 & ~n2974;
  assign n2976 = ~n2970 & n2975;
  assign n2977 = ~pi305 & ~n1575;
  assign n2978 = ~n2976 & n2977;
  assign n2979 = pi206 & n2978;
  assign n2980 = pi276 & ~n2978;
  assign n2981 = ~n2979 & ~n2980;
  assign n2982 = ~n1575 & ~n2981;
  assign n2983 = n1575 & ~n2680;
  assign n2984 = ~n2982 & ~n2983;
  assign n2985 = n2966 & ~n2984;
  assign n2986 = n2889 & n2965;
  assign n2987 = pi276 & ~pi282;
  assign n2988 = ~pi276 & pi282;
  assign n2989 = ~n2987 & ~n2988;
  assign n2990 = n803 & n2238;
  assign n2991 = n803 & n2136;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = n787 & ~n2992;
  assign n2994 = ~n2337 & ~n2343;
  assign n2995 = pi301 & n803;
  assign n2996 = ~n2994 & n2995;
  assign n2997 = ~n2993 & ~n2996;
  assign n2998 = ~n2989 & ~n2997;
  assign n2999 = pi276 & n2997;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = n2986 & ~n3000;
  assign n3002 = ~n2784 & n2958;
  assign n3003 = pi206 & n3002;
  assign n3004 = ~n3001 & ~n3003;
  assign n3005 = ~n2985 & n3004;
  assign n3006 = n2964 & n3005;
  assign n3007 = ~n2891 & n3006;
  assign n3008 = n787 & n833;
  assign n3009 = n804 & n3008;
  assign n3010 = n787 & ~n2827;
  assign n3011 = n1546 & n3010;
  assign n3012 = ~n3009 & ~n3011;
  assign n3013 = ~n3007 & n3012;
  assign n3014 = ~n2653 & n3013;
  assign n3015 = pi276 & n2653;
  assign n3016 = ~pi190 & pi307;
  assign n3017 = pi190 & ~pi307;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~pi188 & pi310;
  assign n3020 = pi188 & ~pi310;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = n3018 & n3021;
  assign n3023 = ~pi189 & pi308;
  assign n3024 = pi189 & ~pi308;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = n3022 & n3025;
  assign n3027 = pi196 & n3026;
  assign n3028 = ~n3015 & ~n3027;
  assign n3029 = n3012 & ~n3028;
  assign n3030 = pi276 & ~n3012;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n3014 & n3031;
  assign n3033 = ~n2650 & ~n3032;
  assign n3034 = n2650 & ~n2680;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = n2647 & ~n3035;
  assign n3037 = pi276 & ~n2647;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = n2633 & ~n3038;
  assign n3040 = pi001 & ~n2633;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n2070 & ~n3041;
  assign n3043 = ~n2075 & ~n3042;
  assign n3044 = ~pi247 & ~n3043;
  assign n3045 = ~n2069 & ~n3044;
  assign po037 = pi359 & ~n3045;
  assign n3047 = pi002 & pi247;
  assign n3048 = pi289 & n2071;
  assign n3049 = pi002 & ~n2071;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = n2070 & ~n3050;
  assign n3052 = pi148 & n2655;
  assign n3053 = pi149 & n2658;
  assign n3054 = ~n3052 & ~n3053;
  assign n3055 = pi147 & n2661;
  assign n3056 = pi153 & n2664;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = pi151 & n2668;
  assign n3059 = pi152 & n2670;
  assign n3060 = ~n3058 & ~n3059;
  assign n3061 = pi150 & n2673;
  assign n3062 = pi175 & n2675;
  assign n3063 = ~n3061 & ~n3062;
  assign n3064 = n3060 & n3063;
  assign n3065 = n3057 & n3064;
  assign n3066 = n3054 & n3065;
  assign n3067 = n2890 & ~n3066;
  assign n3068 = pi351 & n2960;
  assign n3069 = pi172 & n2962;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = pi207 & n2978;
  assign n3072 = pi268 & ~n2978;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = ~n1575 & ~n3073;
  assign n3075 = n1575 & ~n3066;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = n2966 & ~n3076;
  assign n3078 = pi276 & pi282;
  assign n3079 = ~pi268 & n3078;
  assign n3080 = pi268 & ~n3078;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = ~n2997 & ~n3081;
  assign n3083 = pi268 & n2997;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = n2986 & ~n3084;
  assign n3086 = pi207 & n3002;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = ~n3077 & n3087;
  assign n3089 = n3070 & n3088;
  assign n3090 = ~n3067 & n3089;
  assign n3091 = n3012 & ~n3090;
  assign n3092 = ~n2653 & n3091;
  assign n3093 = pi268 & n2653;
  assign n3094 = ~n3027 & ~n3093;
  assign n3095 = n3012 & ~n3094;
  assign n3096 = pi268 & ~n3012;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = ~n3092 & n3097;
  assign n3099 = ~n2650 & ~n3098;
  assign n3100 = n2650 & ~n3066;
  assign n3101 = ~n3099 & ~n3100;
  assign n3102 = n2647 & ~n3101;
  assign n3103 = pi268 & ~n2647;
  assign n3104 = ~n3102 & ~n3103;
  assign n3105 = n2633 & ~n3104;
  assign n3106 = pi002 & ~n2633;
  assign n3107 = ~n3105 & ~n3106;
  assign n3108 = ~n2070 & ~n3107;
  assign n3109 = ~n3051 & ~n3108;
  assign n3110 = ~pi247 & ~n3109;
  assign n3111 = ~n3047 & ~n3110;
  assign po038 = pi359 & ~n3111;
  assign n3113 = pi003 & pi247;
  assign n3114 = pi287 & n2071;
  assign n3115 = pi003 & ~n2071;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = n2070 & ~n3116;
  assign n3118 = pi103 & n2655;
  assign n3119 = pi104 & n2658;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = pi101 & n2661;
  assign n3122 = pi109 & n2664;
  assign n3123 = ~n3121 & ~n3122;
  assign n3124 = pi107 & n2668;
  assign n3125 = pi108 & n2670;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = pi105 & n2673;
  assign n3128 = pi106 & n2675;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = n3126 & n3129;
  assign n3131 = n3123 & n3130;
  assign n3132 = n3120 & n3131;
  assign n3133 = n2890 & ~n3132;
  assign n3134 = pi353 & n2960;
  assign n3135 = pi144 & n2962;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = pi210 & n2978;
  assign n3138 = pi246 & ~n2978;
  assign n3139 = ~n3137 & ~n3138;
  assign n3140 = ~n1575 & ~n3139;
  assign n3141 = n1575 & ~n3132;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = n2966 & ~n3142;
  assign n3144 = pi246 & n2997;
  assign n3145 = pi259 & pi265;
  assign n3146 = n3078 & n3145;
  assign n3147 = pi268 & n3146;
  assign n3148 = pi246 & n3147;
  assign n3149 = ~pi246 & ~n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = ~n2997 & n3150;
  assign n3152 = ~n3144 & ~n3151;
  assign n3153 = n2986 & ~n3152;
  assign n3154 = pi210 & n3002;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n3143 & n3155;
  assign n3157 = n3136 & n3156;
  assign n3158 = ~n3133 & n3157;
  assign n3159 = n3012 & ~n3158;
  assign n3160 = ~n2653 & n3159;
  assign n3161 = pi246 & n2653;
  assign n3162 = ~n3027 & ~n3161;
  assign n3163 = n3012 & ~n3162;
  assign n3164 = pi246 & ~n3012;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = ~n3160 & n3165;
  assign n3167 = ~n2650 & ~n3166;
  assign n3168 = n2650 & ~n3132;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = n2647 & ~n3169;
  assign n3171 = pi246 & ~n2647;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = n2633 & ~n3172;
  assign n3174 = pi003 & ~n2633;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = ~n2070 & ~n3175;
  assign n3177 = ~n3117 & ~n3176;
  assign n3178 = ~pi247 & ~n3177;
  assign n3179 = ~n3113 & ~n3178;
  assign po039 = pi359 & ~n3179;
  assign n3181 = pi004 & pi247;
  assign n3182 = pi286 & n2071;
  assign n3183 = pi004 & ~n2071;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = n2070 & ~n3184;
  assign n3186 = pi067 & n2655;
  assign n3187 = pi068 & n2658;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = pi066 & n2661;
  assign n3190 = pi071 & n2664;
  assign n3191 = ~n3189 & ~n3190;
  assign n3192 = pi072 & n2673;
  assign n3193 = pi073 & n2675;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = pi069 & n2668;
  assign n3196 = pi070 & n2670;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = n3194 & n3197;
  assign n3199 = n3191 & n3198;
  assign n3200 = n3188 & n3199;
  assign n3201 = n2890 & ~n3200;
  assign n3202 = pi347 & n2960;
  assign n3203 = pi137 & n2962;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = pi211 & n2978;
  assign n3206 = pi233 & ~n2978;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n1575 & ~n3207;
  assign n3209 = n1575 & ~n3200;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n2966 & ~n3210;
  assign n3212 = pi233 & n2997;
  assign n3213 = pi268 & n3078;
  assign n3214 = pi265 & n3213;
  assign n3215 = pi246 & n3214;
  assign n3216 = pi259 & n3215;
  assign n3217 = pi233 & n3216;
  assign n3218 = ~pi233 & ~n3216;
  assign n3219 = ~n3217 & ~n3218;
  assign n3220 = ~n2997 & n3219;
  assign n3221 = ~n3212 & ~n3220;
  assign n3222 = n2986 & ~n3221;
  assign n3223 = pi211 & n3002;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = ~n3211 & n3224;
  assign n3226 = n3204 & n3225;
  assign n3227 = ~n3201 & n3226;
  assign n3228 = n3012 & ~n3227;
  assign n3229 = ~n2653 & n3228;
  assign n3230 = pi233 & n2653;
  assign n3231 = ~n3027 & ~n3230;
  assign n3232 = n3012 & ~n3231;
  assign n3233 = pi233 & ~n3012;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = ~n3229 & n3234;
  assign n3236 = ~n2650 & ~n3235;
  assign n3237 = n2650 & ~n3200;
  assign n3238 = ~n3236 & ~n3237;
  assign n3239 = n2647 & ~n3238;
  assign n3240 = pi233 & ~n2647;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = n2633 & ~n3241;
  assign n3243 = pi004 & ~n2633;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = ~n2070 & ~n3244;
  assign n3246 = ~n3185 & ~n3245;
  assign n3247 = ~pi247 & ~n3246;
  assign n3248 = ~n3181 & ~n3247;
  assign po040 = pi359 & ~n3248;
  assign n3250 = ~pi234 & ~pi240;
  assign n3251 = ~pi231 & ~n3250;
  assign n3252 = pi251 & n3251;
  assign n3253 = pi239 & n3252;
  assign n3254 = pi097 & ~pi098;
  assign n3255 = ~pi099 & n3254;
  assign n3256 = ~pi252 & n3255;
  assign n3257 = ~pi242 & ~n3256;
  assign n3258 = pi241 & pi257;
  assign n3259 = pi256 & n3258;
  assign n3260 = ~pi243 & n3259;
  assign n3261 = pi242 & n3260;
  assign n3262 = ~n3257 & ~n3261;
  assign n3263 = n3253 & n3262;
  assign n3264 = ~n926 & ~n946;
  assign n3265 = ~n780 & n2071;
  assign n3266 = ~n915 & n3265;
  assign n3267 = ~n1573 & ~n3266;
  assign n3268 = ~n3264 & ~n3267;
  assign n3269 = ~n3263 & ~n3268;
  assign n3270 = ~n1563 & ~n1566;
  assign n3271 = n3269 & n3270;
  assign po078 = ~pi247 & ~n3271;
  assign n3273 = ~pi005 & ~po078;
  assign n3274 = pi005 & ~n1608;
  assign n3275 = pi280 & ~n1563;
  assign n3276 = ~n1571 & ~n3275;
  assign n3277 = pi284 & ~n1563;
  assign n3278 = ~pi283 & ~n1563;
  assign n3279 = ~n3277 & ~n3278;
  assign n3280 = ~n3276 & n3279;
  assign n3281 = ~pi010 & n3280;
  assign n3282 = ~n3277 & n3278;
  assign n3283 = ~n3276 & n3282;
  assign n3284 = ~pi009 & n3283;
  assign n3285 = ~n3281 & ~n3284;
  assign n3286 = n3277 & n3278;
  assign n3287 = n3276 & n3286;
  assign n3288 = ~pi007 & n3287;
  assign n3289 = n3277 & ~n3278;
  assign n3290 = n3276 & n3289;
  assign n3291 = ~pi008 & n3290;
  assign n3292 = ~n3288 & ~n3291;
  assign n3293 = ~n3276 & n3286;
  assign n3294 = ~pi011 & n3293;
  assign n3295 = ~n3276 & n3289;
  assign n3296 = ~pi012 & n3295;
  assign n3297 = ~n3294 & ~n3296;
  assign n3298 = n3276 & n3282;
  assign n3299 = ~pi005 & n3298;
  assign n3300 = n3276 & n3279;
  assign n3301 = ~pi006 & n3300;
  assign n3302 = ~n3299 & ~n3301;
  assign n3303 = n3297 & n3302;
  assign n3304 = n3292 & n3303;
  assign n3305 = n3285 & n3304;
  assign n3306 = n1563 & ~n3305;
  assign n3307 = ~n780 & n785;
  assign n3308 = ~n915 & n3307;
  assign n3309 = ~n1573 & ~n3308;
  assign n3310 = ~n1566 & ~n3309;
  assign n3311 = ~n2033 & n2039;
  assign n3312 = ~n1859 & ~n2035;
  assign n3313 = n3311 & n3312;
  assign n3314 = n2031 & ~n3313;
  assign n3315 = ~n1859 & ~n2031;
  assign n3316 = n2039 & n3315;
  assign n3317 = n2036 & n3316;
  assign n3318 = ~n3314 & ~n3317;
  assign n3319 = n3310 & n3318;
  assign n3320 = ~n1563 & n3319;
  assign n3321 = ~n1566 & n3309;
  assign n3322 = pi299 & ~pi300;
  assign n3323 = ~n850 & n3322;
  assign n3324 = n787 & n3323;
  assign n3325 = ~n2793 & n3324;
  assign n3326 = pi269 & n3325;
  assign n3327 = ~pi242 & pi347;
  assign n3328 = pi243 & ~pi256;
  assign n3329 = n3258 & n3328;
  assign n3330 = pi269 & n3329;
  assign n3331 = ~n850 & n3330;
  assign n3332 = ~pi269 & ~n850;
  assign n3333 = pi241 & n976;
  assign n3334 = ~pi256 & n3333;
  assign n3335 = ~n3332 & n3334;
  assign n3336 = ~pi243 & ~n1200;
  assign n3337 = ~n3335 & ~n3336;
  assign n3338 = n1087 & ~n1458;
  assign n3339 = n977 & ~n1029;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = n1084 & n1356;
  assign n3342 = pi217 & n960;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = n3340 & n3343;
  assign n3345 = n3337 & n3344;
  assign n3346 = ~n3331 & n3345;
  assign n3347 = pi242 & ~n3346;
  assign n3348 = ~n3327 & ~n3347;
  assign n3349 = ~n3325 & ~n3348;
  assign n3350 = ~n3326 & ~n3349;
  assign n3351 = n3321 & ~n3350;
  assign n3352 = ~pi250 & n1566;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~n1563 & ~n3353;
  assign n3355 = ~n3320 & ~n3354;
  assign n3356 = ~n3306 & n3355;
  assign n3357 = n1608 & n3356;
  assign n3358 = ~n3274 & ~n3357;
  assign n3359 = po078 & n3358;
  assign po041 = n3273 | n3359;
  assign n3361 = ~pi006 & ~po078;
  assign n3362 = ~n1592 & n1598;
  assign n3363 = n1585 & n3362;
  assign n3364 = n3356 & n3363;
  assign n3365 = pi006 & ~n3363;
  assign n3366 = po078 & ~n3365;
  assign n3367 = ~n3364 & n3366;
  assign po042 = n3361 | n3367;
  assign n3369 = ~pi007 & ~po078;
  assign n3370 = n1585 & n1618;
  assign n3371 = n3356 & n3370;
  assign n3372 = pi007 & ~n3370;
  assign n3373 = po078 & ~n3372;
  assign n3374 = ~n3371 & n3373;
  assign po043 = n3369 | n3374;
  assign n3376 = ~pi008 & ~po078;
  assign n3377 = n1585 & n1599;
  assign n3378 = pi008 & ~n3377;
  assign n3379 = n3356 & n3377;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = po078 & n3380;
  assign po044 = n3376 | n3381;
  assign n3383 = ~pi009 & ~po078;
  assign n3384 = pi009 & ~n1603;
  assign n3385 = n1603 & n3356;
  assign n3386 = ~n3384 & ~n3385;
  assign n3387 = po078 & n3386;
  assign po045 = n3383 | n3387;
  assign n3389 = ~pi010 & ~po078;
  assign n3390 = ~n1585 & n3362;
  assign n3391 = n3356 & n3390;
  assign n3392 = pi010 & ~n3390;
  assign n3393 = po078 & ~n3392;
  assign n3394 = ~n3391 & n3393;
  assign po046 = n3389 | n3394;
  assign n3396 = ~pi011 & ~po078;
  assign n3397 = n1619 & n3356;
  assign n3398 = pi011 & ~n1619;
  assign n3399 = po078 & ~n3398;
  assign n3400 = ~n3397 & n3399;
  assign po047 = n3396 | n3400;
  assign n3402 = ~pi012 & ~po078;
  assign n3403 = pi012 & ~n1600;
  assign n3404 = n1600 & n3356;
  assign n3405 = ~n3403 & ~n3404;
  assign n3406 = po078 & n3405;
  assign po048 = n3402 | n3406;
  assign n3408 = ~pi013 & ~po078;
  assign n3409 = ~pi018 & n3280;
  assign n3410 = ~pi017 & n3283;
  assign n3411 = ~n3409 & ~n3410;
  assign n3412 = ~pi019 & n3293;
  assign n3413 = ~pi020 & n3295;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~pi013 & n3298;
  assign n3416 = ~pi014 & n3300;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = ~pi015 & n3287;
  assign n3419 = ~pi016 & n3290;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = n3417 & n3420;
  assign n3422 = n3414 & n3421;
  assign n3423 = n3411 & n3422;
  assign n3424 = n1563 & ~n3423;
  assign n3425 = ~n1563 & n3310;
  assign n3426 = ~n1921 & n3425;
  assign n3427 = pi270 & n3325;
  assign n3428 = ~pi242 & pi352;
  assign n3429 = pi270 & ~n1359;
  assign n3430 = n3329 & n3429;
  assign n3431 = ~pi270 & ~n1359;
  assign n3432 = n3334 & ~n3431;
  assign n3433 = ~pi243 & ~n1307;
  assign n3434 = ~n3432 & ~n3433;
  assign n3435 = n1087 & ~n1479;
  assign n3436 = n977 & ~n1004;
  assign n3437 = ~n3435 & ~n3436;
  assign n3438 = n1084 & n1360;
  assign n3439 = pi216 & n960;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = n3437 & n3440;
  assign n3442 = n3434 & n3441;
  assign n3443 = ~n3430 & n3442;
  assign n3444 = pi242 & ~n3443;
  assign n3445 = ~n3428 & ~n3444;
  assign n3446 = ~n3325 & ~n3445;
  assign n3447 = ~n3427 & ~n3446;
  assign n3448 = n3321 & ~n3447;
  assign n3449 = ~pi249 & n1566;
  assign n3450 = ~n3448 & ~n3449;
  assign n3451 = ~n1563 & ~n3450;
  assign n3452 = ~n3426 & ~n3451;
  assign n3453 = ~n3424 & n3452;
  assign n3454 = n1608 & n3453;
  assign n3455 = pi013 & ~n1608;
  assign n3456 = po078 & ~n3455;
  assign n3457 = ~n3454 & n3456;
  assign po049 = n3408 | n3457;
  assign n3459 = ~pi014 & ~po078;
  assign n3460 = pi014 & ~n3363;
  assign n3461 = n3363 & n3453;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = po078 & n3462;
  assign po050 = n3459 | n3463;
  assign n3465 = ~pi015 & ~po078;
  assign n3466 = n3370 & n3453;
  assign n3467 = pi015 & ~n3370;
  assign n3468 = po078 & ~n3467;
  assign n3469 = ~n3466 & n3468;
  assign po051 = n3465 | n3469;
  assign n3471 = ~pi016 & ~po078;
  assign n3472 = pi016 & ~n3377;
  assign n3473 = n3377 & n3453;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = po078 & n3474;
  assign po052 = n3471 | n3475;
  assign n3477 = ~pi017 & ~po078;
  assign n3478 = pi017 & ~n1603;
  assign n3479 = n1603 & n3453;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = po078 & n3480;
  assign po053 = n3477 | n3481;
  assign n3483 = ~pi018 & ~po078;
  assign n3484 = n3390 & n3453;
  assign n3485 = pi018 & ~n3390;
  assign n3486 = po078 & ~n3485;
  assign n3487 = ~n3484 & n3486;
  assign po054 = n3483 | n3487;
  assign n3489 = ~pi019 & ~po078;
  assign n3490 = n1619 & n3453;
  assign n3491 = pi019 & ~n1619;
  assign n3492 = po078 & ~n3491;
  assign n3493 = ~n3490 & n3492;
  assign po055 = n3489 | n3493;
  assign n3495 = ~pi020 & ~po078;
  assign n3496 = pi020 & ~n1600;
  assign n3497 = n1600 & n3453;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = po078 & n3498;
  assign po056 = n3495 | n3499;
  assign n3501 = pi021 & ~po078;
  assign n3502 = ~pi021 & ~n1608;
  assign n3503 = ~n1955 & n3425;
  assign n3504 = pi026 & n3280;
  assign n3505 = pi025 & n3283;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = pi027 & n3293;
  assign n3508 = pi028 & n3295;
  assign n3509 = ~n3507 & ~n3508;
  assign n3510 = pi021 & n3298;
  assign n3511 = pi022 & n3300;
  assign n3512 = ~n3510 & ~n3511;
  assign n3513 = pi023 & n3287;
  assign n3514 = pi024 & n3290;
  assign n3515 = ~n3513 & ~n3514;
  assign n3516 = n3512 & n3515;
  assign n3517 = n3509 & n3516;
  assign n3518 = n3506 & n3517;
  assign n3519 = n1563 & ~n3518;
  assign n3520 = ~pi248 & n1566;
  assign n3521 = pi274 & n3325;
  assign n3522 = ~pi242 & pi351;
  assign n3523 = pi274 & ~n1372;
  assign n3524 = n3329 & n3523;
  assign n3525 = ~pi274 & ~n1372;
  assign n3526 = n3334 & ~n3525;
  assign n3527 = ~pi243 & ~n1342;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = n1087 & n1518;
  assign n3530 = n977 & ~n1066;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = n1084 & n1373;
  assign n3533 = n960 & ~n964;
  assign n3534 = ~n3532 & ~n3533;
  assign n3535 = n3531 & n3534;
  assign n3536 = n3528 & n3535;
  assign n3537 = ~n3524 & n3536;
  assign n3538 = pi242 & ~n3537;
  assign n3539 = ~n3522 & ~n3538;
  assign n3540 = ~n3325 & ~n3539;
  assign n3541 = ~n3521 & ~n3540;
  assign n3542 = n3321 & ~n3541;
  assign n3543 = ~n3520 & ~n3542;
  assign n3544 = ~n1563 & ~n3543;
  assign n3545 = ~n3519 & ~n3544;
  assign n3546 = ~n3503 & n3545;
  assign n3547 = n1608 & n3546;
  assign n3548 = ~n3502 & ~n3547;
  assign n3549 = po078 & n3548;
  assign po057 = n3501 | n3549;
  assign n3551 = pi022 & ~po078;
  assign n3552 = n3363 & n3546;
  assign n3553 = ~pi022 & ~n3363;
  assign n3554 = po078 & ~n3553;
  assign n3555 = ~n3552 & n3554;
  assign po058 = n3551 | n3555;
  assign n3557 = pi023 & ~po078;
  assign n3558 = n3370 & n3546;
  assign n3559 = ~pi023 & ~n3370;
  assign n3560 = po078 & ~n3559;
  assign n3561 = ~n3558 & n3560;
  assign po059 = n3557 | n3561;
  assign n3563 = pi024 & ~po078;
  assign n3564 = ~pi024 & ~n3377;
  assign n3565 = n3377 & n3546;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = po078 & n3566;
  assign po060 = n3563 | n3567;
  assign n3569 = pi025 & ~po078;
  assign n3570 = ~pi025 & ~n1603;
  assign n3571 = n1603 & n3546;
  assign n3572 = ~n3570 & ~n3571;
  assign n3573 = po078 & n3572;
  assign po061 = n3569 | n3573;
  assign n3575 = pi026 & ~po078;
  assign n3576 = n3390 & n3546;
  assign n3577 = ~pi026 & ~n3390;
  assign n3578 = po078 & ~n3577;
  assign n3579 = ~n3576 & n3578;
  assign po062 = n3575 | n3579;
  assign n3581 = pi027 & ~po078;
  assign n3582 = n1619 & n3546;
  assign n3583 = ~pi027 & ~n1619;
  assign n3584 = po078 & ~n3583;
  assign n3585 = ~n3582 & n3584;
  assign po063 = n3581 | n3585;
  assign n3587 = pi028 & ~po078;
  assign n3588 = ~pi028 & ~n1600;
  assign n3589 = n1600 & n3546;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = po078 & n3590;
  assign po064 = n3587 | n3591;
  assign n3593 = pi343 & n2071;
  assign n3594 = pi029 & ~n2071;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = n2070 & ~n3595;
  assign n3597 = pi343 & n2653;
  assign n3598 = ~pi062 & n2668;
  assign n3599 = ~pi063 & n2670;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = ~pi057 & n2661;
  assign n3602 = ~pi064 & n2664;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = ~pi058 & n2655;
  assign n3605 = ~pi059 & n2658;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = ~pi060 & n2673;
  assign n3608 = ~pi061 & n2675;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = n3606 & n3609;
  assign n3611 = n3603 & n3610;
  assign n3612 = n3600 & n3611;
  assign n3613 = n2890 & ~n3612;
  assign n3614 = pi138 & n2960;
  assign n3615 = pi186 & n2962;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617 = pi203 & n2978;
  assign n3618 = pi229 & ~n2978;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = ~n1575 & ~n3619;
  assign n3621 = n1575 & ~n3612;
  assign n3622 = ~n3620 & ~n3621;
  assign n3623 = n2966 & ~n3622;
  assign n3624 = pi348 & n2997;
  assign n3625 = pi232 & pi238;
  assign n3626 = pi244 & n3625;
  assign n3627 = pi222 & n3626;
  assign n3628 = pi233 & pi246;
  assign n3629 = n3213 & n3628;
  assign n3630 = n3145 & n3629;
  assign n3631 = n3627 & n3630;
  assign n3632 = pi229 & n3631;
  assign n3633 = ~pi229 & ~n3631;
  assign n3634 = ~n3632 & ~n3633;
  assign n3635 = ~n2997 & n3634;
  assign n3636 = ~n3624 & ~n3635;
  assign n3637 = n2986 & ~n3636;
  assign n3638 = pi203 & n3002;
  assign n3639 = ~n3637 & ~n3638;
  assign n3640 = ~n3623 & n3639;
  assign n3641 = n3616 & n3640;
  assign n3642 = ~n3613 & n3641;
  assign n3643 = ~n2653 & ~n3642;
  assign n3644 = ~n3597 & ~n3643;
  assign n3645 = ~n3009 & ~n3027;
  assign n3646 = ~n3011 & n3645;
  assign n3647 = ~n3644 & n3646;
  assign n3648 = pi229 & ~n3012;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = ~n2650 & ~n3649;
  assign n3651 = n2650 & ~n3612;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = n2647 & ~n3652;
  assign n3654 = pi348 & ~n2647;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = n2633 & ~n3655;
  assign n3657 = pi029 & ~n2633;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = ~n2070 & ~n3658;
  assign n3660 = ~n3596 & ~n3659;
  assign n3661 = ~pi247 & ~n3660;
  assign n3662 = pi029 & pi247;
  assign n3663 = ~n3661 & ~n3662;
  assign po065 = pi359 & ~n3663;
  assign n3665 = pi338 & n2071;
  assign n3666 = pi030 & ~n2071;
  assign n3667 = ~n3665 & ~n3666;
  assign n3668 = n2070 & ~n3667;
  assign n3669 = pi338 & n2653;
  assign n3670 = ~pi014 & n2655;
  assign n3671 = ~pi015 & n2658;
  assign n3672 = ~n3670 & ~n3671;
  assign n3673 = ~pi013 & n2661;
  assign n3674 = ~pi020 & n2664;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = ~pi018 & n2668;
  assign n3677 = ~pi019 & n2670;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = ~pi016 & n2673;
  assign n3680 = ~pi017 & n2675;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = n3678 & n3681;
  assign n3683 = n3675 & n3682;
  assign n3684 = n3672 & n3683;
  assign n3685 = n2890 & ~n3684;
  assign n3686 = pi143 & n2960;
  assign n3687 = pi177 & n2962;
  assign n3688 = ~n3686 & ~n3687;
  assign n3689 = pi204 & n2978;
  assign n3690 = pi226 & ~n2978;
  assign n3691 = ~n3689 & ~n3690;
  assign n3692 = ~n1575 & ~n3691;
  assign n3693 = n1575 & ~n3684;
  assign n3694 = ~n3692 & ~n3693;
  assign n3695 = n2966 & ~n3694;
  assign n3696 = pi352 & n2997;
  assign n3697 = pi259 & n3214;
  assign n3698 = pi246 & n3697;
  assign n3699 = pi244 & n3698;
  assign n3700 = pi233 & n3699;
  assign n3701 = n3625 & n3700;
  assign n3702 = pi229 & n3701;
  assign n3703 = pi222 & n3702;
  assign n3704 = pi226 & n3703;
  assign n3705 = ~pi226 & ~n3703;
  assign n3706 = ~n3704 & ~n3705;
  assign n3707 = ~n2997 & n3706;
  assign n3708 = ~n3696 & ~n3707;
  assign n3709 = n2986 & ~n3708;
  assign n3710 = pi204 & n3002;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = ~n3695 & n3711;
  assign n3713 = n3688 & n3712;
  assign n3714 = ~n3685 & n3713;
  assign n3715 = ~n2653 & ~n3714;
  assign n3716 = ~n3669 & ~n3715;
  assign n3717 = n3646 & ~n3716;
  assign n3718 = pi226 & ~n3012;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = ~n2650 & ~n3719;
  assign n3721 = n2650 & ~n3684;
  assign n3722 = ~n3720 & ~n3721;
  assign n3723 = n2647 & ~n3722;
  assign n3724 = pi352 & ~n2647;
  assign n3725 = ~n3723 & ~n3724;
  assign n3726 = n2633 & ~n3725;
  assign n3727 = pi030 & ~n2633;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~n2070 & ~n3728;
  assign n3730 = ~n3668 & ~n3729;
  assign n3731 = ~pi247 & ~n3730;
  assign n3732 = pi030 & pi247;
  assign n3733 = ~n3731 & ~n3732;
  assign po066 = pi359 & ~n3733;
  assign n3735 = pi336 & n2071;
  assign n3736 = pi031 & ~n2071;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = n2070 & ~n3737;
  assign n3739 = pi336 & n2653;
  assign n3740 = ~pi055 & n2668;
  assign n3741 = ~pi056 & n2670;
  assign n3742 = ~n3740 & ~n3741;
  assign n3743 = ~pi049 & n2661;
  assign n3744 = ~pi054 & n2664;
  assign n3745 = ~n3743 & ~n3744;
  assign n3746 = ~pi050 & n2655;
  assign n3747 = ~pi051 & n2658;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = ~pi052 & n2673;
  assign n3750 = ~pi053 & n2675;
  assign n3751 = ~n3749 & ~n3750;
  assign n3752 = n3748 & n3751;
  assign n3753 = n3745 & n3752;
  assign n3754 = n3742 & n3753;
  assign n3755 = n2890 & ~n3754;
  assign n3756 = pi139 & n2960;
  assign n3757 = pi183 & n2962;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = pi205 & n2978;
  assign n3760 = pi227 & ~n2978;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = ~n1575 & ~n3761;
  assign n3763 = n1575 & ~n3754;
  assign n3764 = ~n3762 & ~n3763;
  assign n3765 = n2966 & ~n3764;
  assign n3766 = pi353 & n2997;
  assign n3767 = pi244 & n3628;
  assign n3768 = pi238 & n3767;
  assign n3769 = pi222 & n3768;
  assign n3770 = n3147 & n3769;
  assign n3771 = pi229 & n3770;
  assign n3772 = pi232 & n3771;
  assign n3773 = pi226 & n3772;
  assign n3774 = pi227 & n3773;
  assign n3775 = ~pi227 & ~n3773;
  assign n3776 = ~n3774 & ~n3775;
  assign n3777 = ~n2997 & n3776;
  assign n3778 = ~n3766 & ~n3777;
  assign n3779 = n2986 & ~n3778;
  assign n3780 = pi205 & n3002;
  assign n3781 = ~n3779 & ~n3780;
  assign n3782 = ~n3765 & n3781;
  assign n3783 = n3758 & n3782;
  assign n3784 = ~n3755 & n3783;
  assign n3785 = ~n2653 & ~n3784;
  assign n3786 = ~n3739 & ~n3785;
  assign n3787 = n3646 & ~n3786;
  assign n3788 = pi227 & ~n3012;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = ~n2650 & ~n3789;
  assign n3791 = n2650 & ~n3754;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = n2647 & ~n3792;
  assign n3794 = pi353 & ~n2647;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = n2633 & ~n3795;
  assign n3797 = pi031 & ~n2633;
  assign n3798 = ~n3796 & ~n3797;
  assign n3799 = ~n2070 & ~n3798;
  assign n3800 = ~n3738 & ~n3799;
  assign n3801 = ~pi247 & ~n3800;
  assign n3802 = pi031 & pi247;
  assign n3803 = ~n3801 & ~n3802;
  assign po067 = pi359 & ~n3803;
  assign n3805 = pi340 & n2071;
  assign n3806 = pi032 & ~n2071;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = n2070 & ~n3807;
  assign n3809 = pi340 & n2653;
  assign n3810 = ~pi010 & n2668;
  assign n3811 = ~pi011 & n2670;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = ~pi005 & n2661;
  assign n3814 = ~pi012 & n2664;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = ~pi006 & n2655;
  assign n3817 = ~pi007 & n2658;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = ~pi008 & n2673;
  assign n3820 = ~pi009 & n2675;
  assign n3821 = ~n3819 & ~n3820;
  assign n3822 = n3818 & n3821;
  assign n3823 = n3815 & n3822;
  assign n3824 = n3812 & n3823;
  assign n3825 = n2890 & ~n3824;
  assign n3826 = pi140 & n2960;
  assign n3827 = pi117 & n2962;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = pi347 & n2997;
  assign n3830 = pi226 & pi227;
  assign n3831 = pi233 & n3626;
  assign n3832 = n3216 & n3831;
  assign n3833 = pi222 & n3832;
  assign n3834 = pi229 & n3833;
  assign n3835 = n3830 & n3834;
  assign n3836 = pi191 & n3835;
  assign n3837 = ~pi191 & ~n3835;
  assign n3838 = ~n3836 & ~n3837;
  assign n3839 = ~n2997 & n3838;
  assign n3840 = ~n3829 & ~n3839;
  assign n3841 = n2986 & ~n3840;
  assign n3842 = pi219 & n3002;
  assign n3843 = ~n3841 & ~n3842;
  assign n3844 = pi219 & n2978;
  assign n3845 = pi191 & ~n2978;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = ~n1575 & ~n3846;
  assign n3848 = n1575 & ~n3824;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n2966 & ~n3849;
  assign n3851 = n3843 & ~n3850;
  assign n3852 = n3828 & n3851;
  assign n3853 = ~n3825 & n3852;
  assign n3854 = ~n2653 & ~n3853;
  assign n3855 = ~n3809 & ~n3854;
  assign n3856 = n3646 & ~n3855;
  assign n3857 = pi191 & ~n3012;
  assign n3858 = ~n3856 & ~n3857;
  assign n3859 = ~n2650 & ~n3858;
  assign n3860 = n2650 & ~n3824;
  assign n3861 = ~n3859 & ~n3860;
  assign n3862 = n2647 & ~n3861;
  assign n3863 = pi347 & ~n2647;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = n2633 & ~n3864;
  assign n3866 = pi032 & ~n2633;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = ~n2070 & ~n3867;
  assign n3869 = ~n3808 & ~n3868;
  assign n3870 = ~pi247 & ~n3869;
  assign n3871 = pi032 & pi247;
  assign n3872 = ~n3870 & ~n3871;
  assign po068 = pi359 & ~n3872;
  assign n3874 = pi337 & n2071;
  assign n3875 = pi033 & ~n2071;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = n2070 & ~n3876;
  assign n3878 = pi337 & n2653;
  assign n3879 = pi026 & n2668;
  assign n3880 = pi027 & n2670;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = pi021 & n2661;
  assign n3883 = pi028 & n2664;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = pi022 & n2655;
  assign n3886 = pi023 & n2658;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = pi024 & n2673;
  assign n3889 = pi025 & n2675;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = n3887 & n3890;
  assign n3892 = n3884 & n3891;
  assign n3893 = n3881 & n3892;
  assign n3894 = n2890 & ~n3893;
  assign n3895 = pi141 & n2960;
  assign n3896 = pi182 & n2962;
  assign n3897 = ~n3895 & ~n3896;
  assign n3898 = pi221 & n2978;
  assign n3899 = pi222 & ~n2978;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = ~n1575 & ~n3900;
  assign n3902 = n1575 & ~n3893;
  assign n3903 = ~n3901 & ~n3902;
  assign n3904 = n2966 & ~n3903;
  assign n3905 = pi222 & ~n3832;
  assign n3906 = ~pi222 & n3832;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = ~n2997 & ~n3907;
  assign n3909 = pi351 & n2997;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = n2986 & ~n3910;
  assign n3912 = pi221 & n3002;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = ~n3904 & n3913;
  assign n3915 = n3897 & n3914;
  assign n3916 = ~n3894 & n3915;
  assign n3917 = ~n2653 & ~n3916;
  assign n3918 = ~n3878 & ~n3917;
  assign n3919 = n3646 & ~n3918;
  assign n3920 = pi222 & ~n3012;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = ~n2650 & ~n3921;
  assign n3923 = n2650 & ~n3893;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = n2647 & ~n3924;
  assign n3926 = pi351 & ~n2647;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = n2633 & ~n3927;
  assign n3929 = pi033 & ~n2633;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = ~n2070 & ~n3930;
  assign n3932 = ~n3877 & ~n3931;
  assign n3933 = ~pi247 & ~n3932;
  assign n3934 = pi033 & pi247;
  assign n3935 = ~n3933 & ~n3934;
  assign po069 = pi359 & ~n3935;
  assign n3937 = pi290 & n2071;
  assign n3938 = pi034 & ~n2071;
  assign n3939 = ~n3937 & ~n3938;
  assign n3940 = n2070 & ~n3939;
  assign n3941 = pi259 & n2653;
  assign n3942 = pi111 & n2655;
  assign n3943 = pi112 & n2658;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = pi110 & n2661;
  assign n3946 = pi115 & n2664;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = pi116 & n2668;
  assign n3949 = pi114 & n2670;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = pi113 & n2673;
  assign n3952 = pi100 & n2675;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = n3950 & n3953;
  assign n3955 = n3947 & n3954;
  assign n3956 = n3944 & n3955;
  assign n3957 = n2890 & ~n3956;
  assign n3958 = pi352 & n2960;
  assign n3959 = pi146 & n2962;
  assign n3960 = ~n3958 & ~n3959;
  assign n3961 = pi209 & n2978;
  assign n3962 = pi259 & ~n2978;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = ~n1575 & ~n3963;
  assign n3965 = n1575 & ~n3956;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = n2966 & ~n3966;
  assign n3968 = pi259 & n2997;
  assign n3969 = ~pi259 & ~n3214;
  assign n3970 = ~n3697 & ~n3969;
  assign n3971 = ~n2997 & n3970;
  assign n3972 = ~n3968 & ~n3971;
  assign n3973 = n2986 & ~n3972;
  assign n3974 = pi209 & n3002;
  assign n3975 = ~n3973 & ~n3974;
  assign n3976 = ~n3967 & n3975;
  assign n3977 = n3960 & n3976;
  assign n3978 = ~n3957 & n3977;
  assign n3979 = ~n2653 & ~n3978;
  assign n3980 = ~n3941 & ~n3979;
  assign n3981 = n3646 & ~n3980;
  assign n3982 = pi259 & ~n3012;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n2650 & ~n3983;
  assign n3985 = n2650 & ~n3956;
  assign n3986 = ~n3984 & ~n3985;
  assign n3987 = n2647 & ~n3986;
  assign n3988 = pi259 & ~n2647;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = n2633 & ~n3989;
  assign n3991 = pi034 & ~n2633;
  assign n3992 = ~n3990 & ~n3991;
  assign n3993 = ~n2070 & ~n3992;
  assign n3994 = ~n3940 & ~n3993;
  assign n3995 = ~pi247 & ~n3994;
  assign n3996 = pi034 & pi247;
  assign n3997 = ~n3995 & ~n3996;
  assign po070 = pi359 & ~n3997;
  assign n3999 = pi292 & n2071;
  assign n4000 = pi035 & ~n2071;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = n2070 & ~n4001;
  assign n4003 = pi166 & n2655;
  assign n4004 = pi167 & n2658;
  assign n4005 = ~n4003 & ~n4004;
  assign n4006 = pi165 & n2661;
  assign n4007 = pi171 & n2664;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = pi170 & n2668;
  assign n4010 = pi176 & n2670;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = pi168 & n2673;
  assign n4013 = pi169 & n2675;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = n4011 & n4014;
  assign n4016 = n4008 & n4015;
  assign n4017 = n4005 & n4016;
  assign n4018 = n2890 & ~n4017;
  assign n4019 = pi354 & n2960;
  assign n4020 = pi174 & n2962;
  assign n4021 = ~n4019 & ~n4020;
  assign n4022 = pi282 & n2997;
  assign n4023 = ~pi282 & ~n2997;
  assign n4024 = ~n4022 & ~n4023;
  assign n4025 = n2986 & ~n4024;
  assign n4026 = pi220 & n3002;
  assign n4027 = ~n4025 & ~n4026;
  assign n4028 = pi220 & n2978;
  assign n4029 = pi282 & ~n2978;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = ~n1575 & ~n4030;
  assign n4032 = n1575 & ~n4017;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = n2966 & ~n4033;
  assign n4035 = n4027 & ~n4034;
  assign n4036 = n4021 & n4035;
  assign n4037 = ~n4018 & n4036;
  assign n4038 = n3646 & ~n4037;
  assign n4039 = ~n2653 & n4038;
  assign n4040 = pi282 & ~n3012;
  assign n4041 = pi282 & n2653;
  assign n4042 = n3646 & n4041;
  assign n4043 = ~n4040 & ~n4042;
  assign n4044 = ~n4039 & n4043;
  assign n4045 = ~n2650 & ~n4044;
  assign n4046 = n2650 & ~n4017;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = n2647 & ~n4047;
  assign n4049 = pi282 & ~n2647;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = n2633 & ~n4050;
  assign n4052 = pi035 & ~n2633;
  assign n4053 = ~n4051 & ~n4052;
  assign n4054 = ~n2070 & ~n4053;
  assign n4055 = ~n4002 & ~n4054;
  assign n4056 = ~pi247 & ~n4055;
  assign n4057 = pi035 & pi247;
  assign n4058 = ~n4056 & ~n4057;
  assign po071 = pi359 & ~n4058;
  assign n4060 = pi288 & n2071;
  assign n4061 = pi036 & ~n2071;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n2070 & ~n4062;
  assign n4064 = pi265 & n2653;
  assign n4065 = pi118 & n2668;
  assign n4066 = pi119 & n2670;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = pi121 & n2655;
  assign n4069 = pi125 & n2658;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = pi122 & n2673;
  assign n4072 = pi123 & n2675;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = pi120 & n2661;
  assign n4075 = pi124 & n2664;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = n4073 & n4076;
  assign n4078 = n4070 & n4077;
  assign n4079 = n4067 & n4078;
  assign n4080 = n2890 & ~n4079;
  assign n4081 = pi348 & n2960;
  assign n4082 = pi173 & n2962;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = pi208 & n2978;
  assign n4085 = pi265 & ~n2978;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = ~n1575 & ~n4086;
  assign n4088 = n1575 & ~n4079;
  assign n4089 = ~n4087 & ~n4088;
  assign n4090 = n2966 & ~n4089;
  assign n4091 = pi265 & ~n3213;
  assign n4092 = ~pi265 & n3213;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = ~n2997 & ~n4093;
  assign n4095 = pi265 & n2997;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = n2986 & ~n4096;
  assign n4098 = pi208 & n3002;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = ~n4090 & n4099;
  assign n4101 = n4083 & n4100;
  assign n4102 = ~n4080 & n4101;
  assign n4103 = ~n2653 & ~n4102;
  assign n4104 = ~n4064 & ~n4103;
  assign n4105 = n3646 & ~n4104;
  assign n4106 = pi265 & ~n3012;
  assign n4107 = ~n4105 & ~n4106;
  assign n4108 = ~n2650 & ~n4107;
  assign n4109 = n2650 & ~n4079;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = n2647 & ~n4110;
  assign n4112 = pi265 & ~n2647;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = n2633 & ~n4113;
  assign n4115 = pi036 & ~n2633;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = ~n2070 & ~n4116;
  assign n4118 = ~n4063 & ~n4117;
  assign n4119 = ~pi247 & ~n4118;
  assign n4120 = pi036 & pi247;
  assign n4121 = ~n4119 & ~n4120;
  assign po072 = pi359 & ~n4121;
  assign n4123 = pi339 & n2071;
  assign n4124 = pi037 & ~n2071;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = n2070 & ~n4125;
  assign n4127 = pi339 & n2653;
  assign n4128 = pi046 & n2668;
  assign n4129 = pi047 & n2670;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = pi042 & n2655;
  assign n4132 = pi043 & n2658;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = pi041 & n2661;
  assign n4135 = pi048 & n2664;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = pi044 & n2673;
  assign n4138 = pi045 & n2675;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = n4136 & n4139;
  assign n4141 = n4133 & n4140;
  assign n4142 = n4130 & n4141;
  assign n4143 = n2890 & ~n4142;
  assign n4144 = pi133 & n2960;
  assign n4145 = pi179 & n2962;
  assign n4146 = ~n4144 & ~n4145;
  assign n4147 = pi350 & n2997;
  assign n4148 = pi191 & pi227;
  assign n4149 = pi226 & n3632;
  assign n4150 = n4148 & n4149;
  assign n4151 = ~pi224 & n4150;
  assign n4152 = pi224 & ~n4150;
  assign n4153 = ~n4151 & ~n4152;
  assign n4154 = ~n2997 & n4153;
  assign n4155 = ~n4147 & ~n4154;
  assign n4156 = n2986 & ~n4155;
  assign n4157 = pi218 & n3002;
  assign n4158 = ~n4156 & ~n4157;
  assign n4159 = pi218 & n2978;
  assign n4160 = ~pi224 & ~n2978;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = ~n1575 & ~n4161;
  assign n4163 = n1575 & ~n4142;
  assign n4164 = ~n4162 & ~n4163;
  assign n4165 = n2966 & ~n4164;
  assign n4166 = n4158 & ~n4165;
  assign n4167 = n4146 & n4166;
  assign n4168 = ~n4143 & n4167;
  assign n4169 = ~n2653 & ~n4168;
  assign n4170 = ~n4127 & ~n4169;
  assign n4171 = n3646 & ~n4170;
  assign n4172 = ~pi224 & ~n3012;
  assign n4173 = ~n4171 & ~n4172;
  assign n4174 = ~n2650 & ~n4173;
  assign n4175 = n2650 & ~n4142;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = n2647 & ~n4176;
  assign n4178 = pi350 & ~n2647;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = n2633 & ~n4179;
  assign n4181 = pi037 & ~n2633;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n2070 & ~n4182;
  assign n4184 = ~n4126 & ~n4183;
  assign n4185 = ~pi247 & ~n4184;
  assign n4186 = pi037 & pi247;
  assign n4187 = ~n4185 & ~n4186;
  assign po073 = pi359 & ~n4187;
  assign n4189 = pi341 & n2071;
  assign n4190 = pi038 & ~n2071;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = n2070 & ~n4191;
  assign n4193 = pi341 & n2653;
  assign n4194 = pi091 & n2655;
  assign n4195 = pi092 & n2658;
  assign n4196 = ~n4194 & ~n4195;
  assign n4197 = pi090 & n2661;
  assign n4198 = pi096 & n2664;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = pi094 & n2668;
  assign n4201 = pi095 & n2670;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = pi093 & n2673;
  assign n4204 = pi081 & n2675;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = n4202 & n4205;
  assign n4207 = n4199 & n4206;
  assign n4208 = n4196 & n4207;
  assign n4209 = n2890 & ~n4208;
  assign n4210 = pi126 & n2960;
  assign n4211 = pi187 & n2962;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = pi354 & n2997;
  assign n4214 = pi238 & n3700;
  assign n4215 = ~pi238 & ~n3700;
  assign n4216 = ~n4214 & ~n4215;
  assign n4217 = ~n2997 & n4216;
  assign n4218 = ~n4213 & ~n4217;
  assign n4219 = n2986 & ~n4218;
  assign n4220 = pi212 & n3002;
  assign n4221 = ~n4219 & ~n4220;
  assign n4222 = pi212 & n2978;
  assign n4223 = pi238 & ~n2978;
  assign n4224 = ~n4222 & ~n4223;
  assign n4225 = ~n1575 & ~n4224;
  assign n4226 = n1575 & ~n4208;
  assign n4227 = ~n4225 & ~n4226;
  assign n4228 = n2966 & ~n4227;
  assign n4229 = n4221 & ~n4228;
  assign n4230 = n4212 & n4229;
  assign n4231 = ~n4209 & n4230;
  assign n4232 = ~n2653 & ~n4231;
  assign n4233 = ~n4193 & ~n4232;
  assign n4234 = n3646 & ~n4233;
  assign n4235 = pi238 & ~n3012;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = ~n2650 & ~n4236;
  assign n4238 = n2650 & ~n4208;
  assign n4239 = ~n4237 & ~n4238;
  assign n4240 = n2647 & ~n4239;
  assign n4241 = pi354 & ~n2647;
  assign n4242 = ~n4240 & ~n4241;
  assign n4243 = n2633 & ~n4242;
  assign n4244 = pi038 & ~n2633;
  assign n4245 = ~n4243 & ~n4244;
  assign n4246 = ~n2070 & ~n4245;
  assign n4247 = ~n4192 & ~n4246;
  assign n4248 = ~pi247 & ~n4247;
  assign n4249 = pi038 & pi247;
  assign n4250 = ~n4248 & ~n4249;
  assign po074 = pi359 & ~n4250;
  assign n4252 = pi332 & n2071;
  assign n4253 = pi039 & ~n2071;
  assign n4254 = ~n4252 & ~n4253;
  assign n4255 = n2070 & ~n4254;
  assign n4256 = pi244 & n2653;
  assign n4257 = pi084 & n2655;
  assign n4258 = pi085 & n2658;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260 = pi083 & n2661;
  assign n4261 = pi082 & n2664;
  assign n4262 = ~n4260 & ~n4261;
  assign n4263 = pi088 & n2668;
  assign n4264 = pi089 & n2670;
  assign n4265 = ~n4263 & ~n4264;
  assign n4266 = pi086 & n2673;
  assign n4267 = pi087 & n2675;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = n4265 & n4268;
  assign n4270 = n4262 & n4269;
  assign n4271 = n4259 & n4270;
  assign n4272 = n2890 & ~n4271;
  assign n4273 = pi350 & n2960;
  assign n4274 = pi135 & n2962;
  assign n4275 = ~n4273 & ~n4274;
  assign n4276 = pi244 & ~n3630;
  assign n4277 = ~pi244 & n3630;
  assign n4278 = ~n4276 & ~n4277;
  assign n4279 = ~n2997 & ~n4278;
  assign n4280 = pi244 & n2997;
  assign n4281 = ~n4279 & ~n4280;
  assign n4282 = n2986 & ~n4281;
  assign n4283 = pi200 & n3002;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = pi200 & n2978;
  assign n4286 = pi244 & ~n2978;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = ~n1575 & ~n4287;
  assign n4289 = n1575 & ~n4271;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = n2966 & ~n4290;
  assign n4292 = n4284 & ~n4291;
  assign n4293 = n4275 & n4292;
  assign n4294 = ~n4272 & n4293;
  assign n4295 = ~n2653 & ~n4294;
  assign n4296 = ~n4256 & ~n4295;
  assign n4297 = n3646 & ~n4296;
  assign n4298 = pi244 & ~n3012;
  assign n4299 = ~n4297 & ~n4298;
  assign n4300 = ~n2650 & ~n4299;
  assign n4301 = n2650 & ~n4271;
  assign n4302 = ~n4300 & ~n4301;
  assign n4303 = n2647 & ~n4302;
  assign n4304 = pi244 & ~n2647;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = n2633 & ~n4305;
  assign n4307 = pi039 & ~n2633;
  assign n4308 = ~n4306 & ~n4307;
  assign n4309 = ~n2070 & ~n4308;
  assign n4310 = ~n4255 & ~n4309;
  assign n4311 = ~pi247 & ~n4310;
  assign n4312 = pi039 & pi247;
  assign n4313 = ~n4311 & ~n4312;
  assign po075 = pi359 & ~n4313;
  assign n4315 = pi342 & n2071;
  assign n4316 = pi040 & ~n2071;
  assign n4317 = ~n4315 & ~n4316;
  assign n4318 = n2070 & ~n4317;
  assign n4319 = pi342 & n2653;
  assign n4320 = pi075 & n2655;
  assign n4321 = pi076 & n2658;
  assign n4322 = ~n4320 & ~n4321;
  assign n4323 = pi074 & n2661;
  assign n4324 = pi080 & n2664;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = pi065 & n2668;
  assign n4327 = pi079 & n2670;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = pi077 & n2673;
  assign n4330 = pi078 & n2675;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = n4328 & n4331;
  assign n4333 = n4325 & n4332;
  assign n4334 = n4322 & n4333;
  assign n4335 = n2890 & ~n4334;
  assign n4336 = pi142 & n2960;
  assign n4337 = pi185 & n2962;
  assign n4338 = ~n4336 & ~n4337;
  assign n4339 = pi199 & n2978;
  assign n4340 = pi232 & ~n2978;
  assign n4341 = ~n4339 & ~n4340;
  assign n4342 = ~n1575 & ~n4341;
  assign n4343 = n1575 & ~n4334;
  assign n4344 = ~n4342 & ~n4343;
  assign n4345 = n2966 & ~n4344;
  assign n4346 = n3147 & n3768;
  assign n4347 = pi232 & ~n4346;
  assign n4348 = ~pi232 & n4346;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = ~n2997 & ~n4349;
  assign n4351 = pi349 & n2997;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = n2986 & ~n4352;
  assign n4354 = pi199 & n3002;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = ~n4345 & n4355;
  assign n4357 = n4338 & n4356;
  assign n4358 = ~n4335 & n4357;
  assign n4359 = ~n2653 & ~n4358;
  assign n4360 = ~n4319 & ~n4359;
  assign n4361 = n3646 & ~n4360;
  assign n4362 = pi232 & ~n3012;
  assign n4363 = ~n4361 & ~n4362;
  assign n4364 = ~n2650 & ~n4363;
  assign n4365 = n2650 & ~n4334;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = n2647 & ~n4366;
  assign n4368 = pi349 & ~n2647;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = n2633 & ~n4369;
  assign n4371 = pi040 & ~n2633;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = ~n2070 & ~n4372;
  assign n4374 = ~n4318 & ~n4373;
  assign n4375 = ~pi247 & ~n4374;
  assign n4376 = pi040 & pi247;
  assign n4377 = ~n4375 & ~n4376;
  assign po076 = pi359 & ~n4377;
  assign n4379 = ~n2021 & n3310;
  assign n4380 = pi275 & n3325;
  assign n4381 = ~pi242 & pi350;
  assign n4382 = ~n859 & n3329;
  assign n4383 = pi275 & n4382;
  assign n4384 = ~pi275 & ~n859;
  assign n4385 = n3334 & ~n4384;
  assign n4386 = n1087 & ~n1504;
  assign n4387 = ~n4385 & ~n4386;
  assign n4388 = ~pi243 & ~n1254;
  assign n4389 = n977 & ~n1040;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = n1084 & n1357;
  assign n4392 = pi223 & n960;
  assign n4393 = ~n4391 & ~n4392;
  assign n4394 = n4390 & n4393;
  assign n4395 = n4387 & n4394;
  assign n4396 = ~n4383 & n4395;
  assign n4397 = pi242 & ~n4396;
  assign n4398 = ~n4381 & ~n4397;
  assign n4399 = ~n3325 & ~n4398;
  assign n4400 = ~n4380 & ~n4399;
  assign n4401 = n3321 & ~n4400;
  assign n4402 = ~pi253 & n1566;
  assign n4403 = ~n4401 & ~n4402;
  assign n4404 = ~n1563 & n4403;
  assign n4405 = ~n4379 & n4404;
  assign n4406 = pi044 & n3290;
  assign n4407 = pi043 & n3287;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = pi042 & n3300;
  assign n4410 = pi041 & n3298;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = n4408 & n4411;
  assign n4413 = pi045 & n3283;
  assign n4414 = pi046 & n3280;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = pi047 & n3293;
  assign n4417 = pi048 & n3295;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = n4415 & n4418;
  assign n4420 = n4412 & n4419;
  assign n4421 = n1563 & n4420;
  assign n4422 = ~n4405 & ~n4421;
  assign n4423 = n1608 & ~n4422;
  assign n4424 = ~pi041 & ~n1608;
  assign po079 = ~n4423 & ~n4424;
  assign n4426 = n3363 & ~n4422;
  assign n4427 = ~pi042 & ~n3363;
  assign po081 = ~n4426 & ~n4427;
  assign n4429 = n3370 & ~n4422;
  assign n4430 = ~pi043 & ~n3370;
  assign po083 = ~n4429 & ~n4430;
  assign n4432 = n3377 & ~n4422;
  assign n4433 = ~pi044 & ~n3377;
  assign po085 = ~n4432 & ~n4433;
  assign n4435 = n1603 & ~n4422;
  assign n4436 = ~pi045 & ~n1603;
  assign po087 = ~n4435 & ~n4436;
  assign n4438 = n3390 & ~n4422;
  assign n4439 = ~pi046 & ~n3390;
  assign po089 = ~n4438 & ~n4439;
  assign n4441 = n1619 & ~n4422;
  assign n4442 = ~pi047 & ~n1619;
  assign po091 = ~n4441 & ~n4442;
  assign n4444 = pi048 & ~n1600;
  assign n4445 = ~n4379 & n4403;
  assign n4446 = n1600 & ~n4445;
  assign n4447 = ~n1563 & n4446;
  assign n4448 = n1600 & ~n4420;
  assign n4449 = n1563 & n4448;
  assign n4450 = ~n4447 & ~n4449;
  assign po093 = n4444 | ~n4450;
  assign n4452 = ~pi049 & ~po078;
  assign n4453 = pi049 & ~n1608;
  assign n4454 = ~n1887 & ~n3309;
  assign n4455 = ~n1566 & n4454;
  assign n4456 = ~n1563 & n4455;
  assign n4457 = pi273 & n3325;
  assign n4458 = ~pi242 & pi353;
  assign n4459 = pi273 & ~n1361;
  assign n4460 = n3329 & n4459;
  assign n4461 = ~pi273 & ~n1361;
  assign n4462 = n3334 & ~n4461;
  assign n4463 = n1087 & n1466;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = n1084 & n1362;
  assign n4466 = ~pi243 & ~n1217;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = n977 & ~n992;
  assign n4469 = pi198 & n960;
  assign n4470 = ~n4468 & ~n4469;
  assign n4471 = n4467 & n4470;
  assign n4472 = n4464 & n4471;
  assign n4473 = ~n4460 & n4472;
  assign n4474 = pi242 & ~n4473;
  assign n4475 = ~n4458 & ~n4474;
  assign n4476 = ~n3325 & ~n4475;
  assign n4477 = ~n4457 & ~n4476;
  assign n4478 = n3321 & ~n4477;
  assign n4479 = ~pi236 & n1566;
  assign n4480 = ~n4478 & ~n4479;
  assign n4481 = ~n1563 & ~n4480;
  assign n4482 = ~pi055 & n3280;
  assign n4483 = ~pi053 & n3283;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~pi056 & n3293;
  assign n4486 = ~pi054 & n3295;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~pi049 & n3298;
  assign n4489 = ~pi050 & n3300;
  assign n4490 = ~n4488 & ~n4489;
  assign n4491 = ~pi051 & n3287;
  assign n4492 = ~pi052 & n3290;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = n4490 & n4493;
  assign n4495 = n4487 & n4494;
  assign n4496 = n4484 & n4495;
  assign n4497 = n1563 & ~n4496;
  assign n4498 = ~n4481 & ~n4497;
  assign n4499 = ~n4456 & n4498;
  assign n4500 = n1608 & n4499;
  assign n4501 = ~n4453 & ~n4500;
  assign n4502 = po078 & n4501;
  assign po094 = n4452 | n4502;
  assign n4504 = ~pi050 & ~po078;
  assign n4505 = n3363 & ~n4497;
  assign n4506 = ~n1887 & n3425;
  assign n4507 = ~n4481 & ~n4506;
  assign n4508 = n4505 & n4507;
  assign n4509 = pi050 & ~n3363;
  assign n4510 = po078 & ~n4509;
  assign n4511 = ~n4508 & n4510;
  assign po095 = n4504 | n4511;
  assign n4513 = n3370 & n4499;
  assign n4514 = pi051 & ~n3370;
  assign n4515 = ~n4513 & ~n4514;
  assign n4516 = po078 & n4515;
  assign n4517 = ~pi051 & ~po078;
  assign po096 = n4516 | n4517;
  assign n4519 = ~pi052 & ~po078;
  assign n4520 = pi052 & ~n3377;
  assign n4521 = ~n4497 & n4507;
  assign n4522 = n3377 & n4521;
  assign n4523 = ~n4520 & ~n4522;
  assign n4524 = po078 & n4523;
  assign po097 = n4519 | n4524;
  assign n4526 = ~pi053 & ~po078;
  assign n4527 = pi053 & ~n1603;
  assign n4528 = n1603 & n4499;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = po078 & n4529;
  assign po098 = n4526 | n4530;
  assign n4532 = ~pi054 & ~po078;
  assign n4533 = pi054 & ~n1600;
  assign n4534 = n1600 & n4499;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = po078 & n4535;
  assign po099 = n4532 | n4536;
  assign n4538 = n3390 & ~n4497;
  assign n4539 = n4507 & n4538;
  assign n4540 = pi055 & ~n3390;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = po078 & n4541;
  assign n4543 = ~pi055 & ~po078;
  assign po100 = n4542 | n4543;
  assign n4545 = n1619 & ~n4497;
  assign n4546 = ~n4481 & n4545;
  assign n4547 = ~n4456 & n4546;
  assign n4548 = pi056 & ~n1619;
  assign n4549 = po078 & ~n4548;
  assign n4550 = ~n4547 & n4549;
  assign n4551 = ~pi056 & ~po078;
  assign po101 = n4550 | n4551;
  assign n4553 = ~pi057 & ~po078;
  assign n4554 = pi057 & ~n1608;
  assign n4555 = ~pi059 & n3287;
  assign n4556 = ~pi060 & n3290;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = ~pi063 & n3293;
  assign n4559 = ~pi064 & n3295;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = ~pi062 & n3280;
  assign n4562 = ~pi061 & n3283;
  assign n4563 = ~n4561 & ~n4562;
  assign n4564 = ~pi057 & n3298;
  assign n4565 = ~pi058 & n3300;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = n4563 & n4566;
  assign n4568 = n4560 & n4567;
  assign n4569 = n4557 & n4568;
  assign n4570 = n1563 & ~n4569;
  assign n4571 = pi272 & n3325;
  assign n4572 = ~pi242 & pi348;
  assign n4573 = pi272 & ~n1374;
  assign n4574 = n3329 & n4573;
  assign n4575 = n1084 & n1375;
  assign n4576 = ~pi243 & ~n1325;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = ~n955 & n960;
  assign n4579 = n977 & ~n1077;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~pi272 & ~n1374;
  assign n4582 = n3334 & ~n4581;
  assign n4583 = n1087 & ~n1395;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = n4580 & n4584;
  assign n4586 = n4577 & n4585;
  assign n4587 = ~n4574 & n4586;
  assign n4588 = pi242 & ~n4587;
  assign n4589 = ~n4572 & ~n4588;
  assign n4590 = ~n3325 & ~n4589;
  assign n4591 = ~n4571 & ~n4590;
  assign n4592 = n3321 & ~n4591;
  assign n4593 = ~pi245 & n1566;
  assign n4594 = ~n4592 & ~n4593;
  assign n4595 = ~n1944 & n3310;
  assign n4596 = n4594 & ~n4595;
  assign n4597 = ~n1563 & ~n4596;
  assign n4598 = ~n4570 & ~n4597;
  assign n4599 = n1608 & n4598;
  assign n4600 = ~n4554 & ~n4599;
  assign n4601 = po078 & n4600;
  assign po102 = n4553 | n4601;
  assign n4603 = ~pi058 & ~po078;
  assign n4604 = pi058 & ~n3363;
  assign n4605 = n3363 & n4598;
  assign n4606 = ~n4604 & ~n4605;
  assign n4607 = po078 & n4606;
  assign po103 = n4603 | n4607;
  assign n4609 = ~pi059 & ~po078;
  assign n4610 = pi059 & ~n3370;
  assign n4611 = n3370 & n4598;
  assign n4612 = ~n4610 & ~n4611;
  assign n4613 = po078 & n4612;
  assign po104 = n4609 | n4613;
  assign n4615 = ~pi060 & ~po078;
  assign n4616 = pi060 & ~n3377;
  assign n4617 = n3377 & n4598;
  assign n4618 = ~n4616 & ~n4617;
  assign n4619 = po078 & n4618;
  assign po105 = n4615 | n4619;
  assign n4621 = ~pi061 & ~po078;
  assign n4622 = pi061 & ~n1603;
  assign n4623 = n1603 & n4598;
  assign n4624 = ~n4622 & ~n4623;
  assign n4625 = po078 & n4624;
  assign po106 = n4621 | n4625;
  assign n4627 = ~pi062 & ~po078;
  assign n4628 = pi062 & ~n3390;
  assign n4629 = n3390 & n4598;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = po078 & n4630;
  assign po107 = n4627 | n4631;
  assign n4633 = ~pi063 & ~po078;
  assign n4634 = pi063 & ~n1619;
  assign n4635 = n1619 & n4598;
  assign n4636 = ~n4634 & ~n4635;
  assign n4637 = po078 & n4636;
  assign po108 = n4633 | n4637;
  assign n4639 = ~pi064 & ~po078;
  assign n4640 = pi064 & ~n1600;
  assign n4641 = n1600 & n4598;
  assign n4642 = ~n4640 & ~n4641;
  assign n4643 = po078 & n4642;
  assign po109 = n4639 | n4643;
  assign n4645 = pi065 & ~po078;
  assign n4646 = ~pi065 & ~n3390;
  assign n4647 = pi271 & n3325;
  assign n4648 = ~pi242 & pi349;
  assign n4649 = pi271 & ~n1366;
  assign n4650 = n3329 & n4649;
  assign n4651 = ~pi271 & ~n1366;
  assign n4652 = n3334 & ~n4651;
  assign n4653 = ~pi243 & ~n1272;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = n1084 & n1367;
  assign n4656 = ~n952 & n960;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = n1087 & n1398;
  assign n4659 = n977 & ~n1054;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = n4657 & n4660;
  assign n4662 = n4654 & n4661;
  assign n4663 = ~n4650 & n4662;
  assign n4664 = pi242 & ~n4663;
  assign n4665 = ~n4648 & ~n4664;
  assign n4666 = ~n3325 & ~n4665;
  assign n4667 = ~n4647 & ~n4666;
  assign n4668 = n3321 & ~n4667;
  assign n4669 = ~pi255 & n1566;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = ~n1563 & ~n4670;
  assign n4672 = ~n1927 & n3425;
  assign n4673 = pi065 & n3280;
  assign n4674 = pi078 & n3283;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = pi079 & n3293;
  assign n4677 = pi080 & n3295;
  assign n4678 = ~n4676 & ~n4677;
  assign n4679 = pi074 & n3298;
  assign n4680 = pi075 & n3300;
  assign n4681 = ~n4679 & ~n4680;
  assign n4682 = pi076 & n3287;
  assign n4683 = pi077 & n3290;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = n4681 & n4684;
  assign n4686 = n4678 & n4685;
  assign n4687 = n4675 & n4686;
  assign n4688 = n1563 & ~n4687;
  assign n4689 = ~n4672 & ~n4688;
  assign n4690 = ~n4671 & n4689;
  assign n4691 = n3390 & n4690;
  assign n4692 = ~n4646 & ~n4691;
  assign n4693 = po078 & n4692;
  assign po110 = n4645 | n4693;
  assign n4695 = n3252 & n3262;
  assign n4696 = ~pi239 & n4695;
  assign n4697 = ~n3268 & ~n4696;
  assign n4698 = n3270 & n4697;
  assign n4699 = ~pi247 & ~n4698;
  assign n4700 = pi066 & ~n4699;
  assign n4701 = pi070 & n3293;
  assign n4702 = pi071 & n3295;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = pi066 & n3298;
  assign n4705 = pi067 & n3300;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = pi069 & n3280;
  assign n4708 = pi073 & n3283;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = pi068 & n3287;
  assign n4711 = pi072 & n3290;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = n4709 & n4712;
  assign n4714 = n4706 & n4713;
  assign n4715 = n4703 & n4714;
  assign n4716 = n1563 & ~n4715;
  assign n4717 = ~pi263 & n1566;
  assign n4718 = ~n3351 & ~n4717;
  assign n4719 = ~n2057 & n3310;
  assign n4720 = n4718 & ~n4719;
  assign n4721 = ~n1563 & ~n4720;
  assign n4722 = ~n4716 & ~n4721;
  assign n4723 = n1608 & n4722;
  assign n4724 = ~pi066 & ~n1608;
  assign n4725 = n4699 & ~n4724;
  assign n4726 = ~n4723 & n4725;
  assign po111 = n4700 | n4726;
  assign n4728 = pi067 & ~n4699;
  assign n4729 = n3363 & n4722;
  assign n4730 = ~pi067 & ~n3363;
  assign n4731 = n4699 & ~n4730;
  assign n4732 = ~n4729 & n4731;
  assign po112 = n4728 | n4732;
  assign n4734 = pi068 & ~n4699;
  assign n4735 = n3370 & n4722;
  assign n4736 = ~pi068 & ~n3370;
  assign n4737 = n4699 & ~n4736;
  assign n4738 = ~n4735 & n4737;
  assign po113 = n4734 | n4738;
  assign n4740 = pi069 & ~n4699;
  assign n4741 = n3390 & n4722;
  assign n4742 = ~pi069 & ~n3390;
  assign n4743 = n4699 & ~n4742;
  assign n4744 = ~n4741 & n4743;
  assign po114 = n4740 | n4744;
  assign n4746 = pi070 & ~n4699;
  assign n4747 = n1619 & n4722;
  assign n4748 = ~pi070 & ~n1619;
  assign n4749 = n4699 & ~n4748;
  assign n4750 = ~n4747 & n4749;
  assign po115 = n4746 | n4750;
  assign n4752 = pi071 & ~n4699;
  assign n4753 = n1600 & n4722;
  assign n4754 = ~pi071 & ~n1600;
  assign n4755 = n4699 & ~n4754;
  assign n4756 = ~n4753 & n4755;
  assign po116 = n4752 | n4756;
  assign n4758 = pi072 & ~n4699;
  assign n4759 = n3377 & n4722;
  assign n4760 = ~pi072 & ~n3377;
  assign n4761 = n4699 & ~n4760;
  assign n4762 = ~n4759 & n4761;
  assign po117 = n4758 | n4762;
  assign n4764 = pi073 & ~n4699;
  assign n4765 = n1603 & n4722;
  assign n4766 = ~pi073 & ~n1603;
  assign n4767 = n4699 & ~n4766;
  assign n4768 = ~n4765 & n4767;
  assign po118 = n4764 | n4768;
  assign n4770 = pi074 & ~po078;
  assign n4771 = n1608 & n4690;
  assign n4772 = ~pi074 & ~n1608;
  assign n4773 = po078 & ~n4772;
  assign n4774 = ~n4771 & n4773;
  assign po119 = n4770 | n4774;
  assign n4776 = pi075 & ~po078;
  assign n4777 = n3363 & n4690;
  assign n4778 = ~pi075 & ~n3363;
  assign n4779 = po078 & ~n4778;
  assign n4780 = ~n4777 & n4779;
  assign po120 = n4776 | n4780;
  assign n4782 = pi076 & ~po078;
  assign n4783 = ~pi076 & ~n3370;
  assign n4784 = n3370 & n4690;
  assign n4785 = ~n4783 & ~n4784;
  assign n4786 = po078 & n4785;
  assign po121 = n4782 | n4786;
  assign n4788 = pi077 & ~po078;
  assign n4789 = ~pi077 & ~n3377;
  assign n4790 = n3377 & n4690;
  assign n4791 = ~n4789 & ~n4790;
  assign n4792 = po078 & n4791;
  assign po122 = n4788 | n4792;
  assign n4794 = pi078 & ~po078;
  assign n4795 = ~pi078 & ~n1603;
  assign n4796 = n1603 & n4690;
  assign n4797 = ~n4795 & ~n4796;
  assign n4798 = po078 & n4797;
  assign po123 = n4794 | n4798;
  assign n4800 = pi079 & ~po078;
  assign n4801 = n1619 & n4690;
  assign n4802 = ~pi079 & ~n1619;
  assign n4803 = po078 & ~n4802;
  assign n4804 = ~n4801 & n4803;
  assign po124 = n4800 | n4804;
  assign n4806 = pi080 & ~po078;
  assign n4807 = ~pi080 & ~n1600;
  assign n4808 = n1600 & n4690;
  assign n4809 = ~n4807 & ~n4808;
  assign n4810 = po078 & n4809;
  assign po125 = n4806 | n4810;
  assign n4812 = pi081 & ~po078;
  assign n4813 = ~pi081 & ~n1603;
  assign n4814 = pi264 & n3325;
  assign n4815 = ~pi242 & pi354;
  assign n4816 = n1084 & n1355;
  assign n4817 = ~pi264 & ~n1354;
  assign n4818 = n3334 & ~n4817;
  assign n4819 = pi264 & n3329;
  assign n4820 = ~n1354 & n4819;
  assign n4821 = ~n4818 & ~n4820;
  assign n4822 = ~pi243 & ~n1289;
  assign n4823 = n977 & ~n1015;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = n960 & ~n971;
  assign n4826 = pi197 & n1087;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = n4824 & n4827;
  assign n4829 = n4821 & n4828;
  assign n4830 = ~n4816 & n4829;
  assign n4831 = pi242 & ~n4830;
  assign n4832 = ~n4815 & ~n4831;
  assign n4833 = ~n3325 & ~n4832;
  assign n4834 = ~n4814 & ~n4833;
  assign n4835 = n3321 & ~n4834;
  assign n4836 = ~pi258 & n1566;
  assign n4837 = ~n4835 & ~n4836;
  assign n4838 = ~n1962 & n3310;
  assign n4839 = n4837 & ~n4838;
  assign n4840 = ~n1563 & ~n4839;
  assign n4841 = pi095 & n3293;
  assign n4842 = pi096 & n3295;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = pi092 & n3287;
  assign n4845 = pi093 & n3290;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = pi090 & n3298;
  assign n4848 = pi091 & n3300;
  assign n4849 = ~n4847 & ~n4848;
  assign n4850 = pi094 & n3280;
  assign n4851 = pi081 & n3283;
  assign n4852 = ~n4850 & ~n4851;
  assign n4853 = n4849 & n4852;
  assign n4854 = n4846 & n4853;
  assign n4855 = n4843 & n4854;
  assign n4856 = n1563 & ~n4855;
  assign n4857 = ~n4840 & ~n4856;
  assign n4858 = n1603 & n4857;
  assign n4859 = ~n4813 & ~n4858;
  assign n4860 = po078 & n4859;
  assign po126 = n4812 | n4860;
  assign n4862 = pi082 & ~n4699;
  assign n4863 = pi087 & n3283;
  assign n4864 = pi088 & n3280;
  assign n4865 = ~n4863 & ~n4864;
  assign n4866 = pi082 & n3295;
  assign n4867 = pi089 & n3293;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = pi084 & n3300;
  assign n4870 = pi083 & n3298;
  assign n4871 = ~n4869 & ~n4870;
  assign n4872 = pi086 & n3290;
  assign n4873 = pi085 & n3287;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = n4871 & n4874;
  assign n4876 = n4868 & n4875;
  assign n4877 = n4865 & n4876;
  assign n4878 = n1563 & ~n4877;
  assign n4879 = ~pi254 & n1566;
  assign n4880 = ~n4401 & ~n4879;
  assign n4881 = ~n1563 & ~n4880;
  assign n4882 = ~n4878 & ~n4881;
  assign n4883 = ~n2048 & n3425;
  assign n4884 = n4882 & ~n4883;
  assign n4885 = n1600 & n4884;
  assign n4886 = ~pi082 & ~n1600;
  assign n4887 = n4699 & ~n4886;
  assign n4888 = ~n4885 & n4887;
  assign po127 = n4862 | n4888;
  assign n4890 = pi083 & ~n4699;
  assign n4891 = n1608 & n4884;
  assign n4892 = ~pi083 & ~n1608;
  assign n4893 = n4699 & ~n4892;
  assign n4894 = ~n4891 & n4893;
  assign po128 = n4890 | n4894;
  assign n4896 = pi084 & ~n4699;
  assign n4897 = n3363 & n4884;
  assign n4898 = ~pi084 & ~n3363;
  assign n4899 = n4699 & ~n4898;
  assign n4900 = ~n4897 & n4899;
  assign po129 = n4896 | n4900;
  assign n4902 = pi085 & ~n4699;
  assign n4903 = n3370 & n4884;
  assign n4904 = ~pi085 & ~n3370;
  assign n4905 = n4699 & ~n4904;
  assign n4906 = ~n4903 & n4905;
  assign po130 = n4902 | n4906;
  assign n4908 = pi086 & ~n4699;
  assign n4909 = n3377 & n4884;
  assign n4910 = ~pi086 & ~n3377;
  assign n4911 = n4699 & ~n4910;
  assign n4912 = ~n4909 & n4911;
  assign po131 = n4908 | n4912;
  assign n4914 = pi087 & ~n4699;
  assign n4915 = n1603 & n4884;
  assign n4916 = ~pi087 & ~n1603;
  assign n4917 = n4699 & ~n4916;
  assign n4918 = ~n4915 & n4917;
  assign po132 = n4914 | n4918;
  assign n4920 = pi088 & ~n4699;
  assign n4921 = n3390 & n4884;
  assign n4922 = ~pi088 & ~n3390;
  assign n4923 = n4699 & ~n4922;
  assign n4924 = ~n4921 & n4923;
  assign po133 = n4920 | n4924;
  assign n4926 = pi089 & ~n4699;
  assign n4927 = n1619 & n4884;
  assign n4928 = ~pi089 & ~n1619;
  assign n4929 = n4699 & ~n4928;
  assign n4930 = ~n4927 & n4929;
  assign po134 = n4926 | n4930;
  assign n4932 = ~pi090 & ~n1608;
  assign n4933 = n1608 & ~n4856;
  assign n4934 = ~n4840 & n4933;
  assign n4935 = po078 & ~n4934;
  assign n4936 = ~n4932 & n4935;
  assign n4937 = pi090 & ~po078;
  assign po135 = n4936 | n4937;
  assign n4939 = pi091 & ~po078;
  assign n4940 = ~pi091 & ~n3363;
  assign n4941 = n3363 & n4857;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = po078 & n4942;
  assign po136 = n4939 | n4943;
  assign n4945 = pi092 & ~po078;
  assign n4946 = ~pi092 & ~n3370;
  assign n4947 = n3370 & n4857;
  assign n4948 = ~n4946 & ~n4947;
  assign n4949 = po078 & n4948;
  assign po137 = n4945 | n4949;
  assign n4951 = pi093 & ~po078;
  assign n4952 = ~pi093 & ~n3377;
  assign n4953 = n3377 & n4857;
  assign n4954 = ~n4952 & ~n4953;
  assign n4955 = po078 & n4954;
  assign po138 = n4951 | n4955;
  assign n4957 = pi094 & ~po078;
  assign n4958 = ~pi094 & ~n3390;
  assign n4959 = n3390 & n4857;
  assign n4960 = ~n4958 & ~n4959;
  assign n4961 = po078 & n4960;
  assign po139 = n4957 | n4961;
  assign n4963 = pi095 & ~po078;
  assign n4964 = ~pi095 & ~n1619;
  assign n4965 = n1619 & n4857;
  assign n4966 = ~n4964 & ~n4965;
  assign n4967 = po078 & n4966;
  assign po140 = n4963 | n4967;
  assign n4969 = pi096 & ~po078;
  assign n4970 = ~pi096 & ~n1600;
  assign n4971 = n1600 & n4857;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = po078 & n4972;
  assign po141 = n4969 | n4973;
  assign n4975 = ~pi097 & pi356;
  assign n4976 = n2633 & ~n4975;
  assign n4977 = n811 & n2358;
  assign n4978 = n811 & n2360;
  assign n4979 = n811 & n932;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = ~n4977 & n4980;
  assign n4982 = ~n930 & n4981;
  assign n4983 = pi301 & ~n4982;
  assign n4984 = n804 & n2119;
  assign n4985 = n804 & n2215;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = n787 & ~n4986;
  assign n4988 = ~n4983 & ~n4987;
  assign n4989 = ~pi252 & ~n4988;
  assign n4990 = pi237 & ~n4989;
  assign n4991 = pi195 & n780;
  assign n4992 = pi196 & n780;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = pi252 & n4993;
  assign n4995 = ~n4990 & ~n4994;
  assign n4996 = n4988 & n4993;
  assign n4997 = n4995 & ~n4996;
  assign n4998 = pi097 & n4997;
  assign n4999 = ~pi097 & ~n4997;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = ~n2633 & ~n5000;
  assign n5002 = ~n4976 & ~n5001;
  assign n5003 = ~pi361 & n785;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = pi247 & pi356;
  assign n5006 = n5004 & ~n5005;
  assign n5007 = ~n5003 & ~n5005;
  assign n5008 = pi097 & ~n5007;
  assign n5009 = ~n5006 & ~n5008;
  assign po142 = pi359 & ~n5009;
  assign n5011 = pi098 & ~n5007;
  assign n5012 = ~n3254 & ~n4997;
  assign n5013 = ~n784 & n5012;
  assign n5014 = ~pi098 & n4997;
  assign n5015 = ~n2633 & ~n5014;
  assign n5016 = ~n5013 & n5015;
  assign n5017 = pi098 & pi356;
  assign n5018 = n2633 & n5017;
  assign n5019 = ~n5016 & ~n5018;
  assign n5020 = ~n5003 & ~n5019;
  assign n5021 = ~n5005 & n5020;
  assign n5022 = ~n5011 & ~n5021;
  assign po143 = pi359 & ~n5022;
  assign n5024 = pi099 & pi356;
  assign n5025 = n2633 & ~n5024;
  assign n5026 = pi099 & ~n781;
  assign n5027 = ~n782 & ~n5026;
  assign n5028 = ~n4997 & ~n5027;
  assign n5029 = pi099 & n4997;
  assign n5030 = ~n5028 & ~n5029;
  assign n5031 = ~n2633 & n5030;
  assign n5032 = ~n5025 & ~n5031;
  assign n5033 = ~n5005 & n5032;
  assign n5034 = ~n5003 & n5033;
  assign n5035 = pi099 & ~n5007;
  assign n5036 = ~n5034 & ~n5035;
  assign po144 = pi359 & ~n5036;
  assign n5038 = pi100 & ~n4699;
  assign n5039 = pi114 & n3293;
  assign n5040 = pi115 & n3295;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = pi116 & n3280;
  assign n5043 = pi100 & n3283;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = pi110 & n3298;
  assign n5046 = pi111 & n3300;
  assign n5047 = ~n5045 & ~n5046;
  assign n5048 = pi112 & n3287;
  assign n5049 = pi113 & n3290;
  assign n5050 = ~n5048 & ~n5049;
  assign n5051 = n5047 & n5050;
  assign n5052 = n5044 & n5051;
  assign n5053 = n5041 & n5052;
  assign n5054 = n1563 & ~n5053;
  assign n5055 = ~pi266 & n1566;
  assign n5056 = ~n3448 & ~n5055;
  assign n5057 = ~n2061 & n3310;
  assign n5058 = n5056 & ~n5057;
  assign n5059 = ~n1563 & ~n5058;
  assign n5060 = ~n5054 & ~n5059;
  assign n5061 = n1603 & n5060;
  assign n5062 = ~pi100 & ~n1603;
  assign n5063 = n4699 & ~n5062;
  assign n5064 = ~n5061 & n5063;
  assign po145 = n5038 | n5064;
  assign n5066 = pi101 & ~n4699;
  assign n5067 = pi101 & n3298;
  assign n5068 = pi103 & n3300;
  assign n5069 = ~n5067 & ~n5068;
  assign n5070 = pi104 & n3287;
  assign n5071 = pi105 & n3290;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = pi108 & n3293;
  assign n5074 = pi109 & n3295;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = pi107 & n3280;
  assign n5077 = pi106 & n3283;
  assign n5078 = ~n5076 & ~n5077;
  assign n5079 = n5075 & n5078;
  assign n5080 = n5072 & n5079;
  assign n5081 = n5069 & n5080;
  assign n5082 = n1563 & ~n5081;
  assign n5083 = ~pi262 & n1566;
  assign n5084 = ~n4478 & ~n5083;
  assign n5085 = ~n2052 & n3310;
  assign n5086 = n5084 & ~n5085;
  assign n5087 = ~n1563 & ~n5086;
  assign n5088 = ~n5082 & ~n5087;
  assign n5089 = n1608 & n5088;
  assign n5090 = ~pi101 & ~n1608;
  assign n5091 = ~n5089 & ~n5090;
  assign n5092 = n4699 & n5091;
  assign po146 = n5066 | n5092;
  assign n5094 = pi301 & n912;
  assign n5095 = n905 & n2634;
  assign n5096 = ~n5094 & ~n5095;
  assign n5097 = pi242 & ~n1529;
  assign n5098 = n956 & n3328;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = ~n1015 & n1040;
  assign n5101 = n1015 & ~n1040;
  assign n5102 = ~n5100 & ~n5101;
  assign n5103 = ~n1004 & n1066;
  assign n5104 = n1004 & ~n1066;
  assign n5105 = ~n5103 & ~n5104;
  assign n5106 = ~n5102 & n5105;
  assign n5107 = n5102 & ~n5105;
  assign n5108 = ~n5106 & ~n5107;
  assign n5109 = ~n1029 & n1054;
  assign n5110 = n1029 & ~n1054;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = ~n992 & n1077;
  assign n5113 = n992 & ~n1077;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = ~n5111 & n5114;
  assign n5116 = n5111 & ~n5114;
  assign n5117 = ~n5115 & ~n5116;
  assign n5118 = ~n5108 & n5117;
  assign n5119 = n5108 & ~n5117;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = ~n787 & n5120;
  assign n5122 = pi102 & n787;
  assign n5123 = ~n5121 & ~n5122;
  assign n5124 = n977 & ~n5123;
  assign n5125 = pi216 & n964;
  assign n5126 = ~pi216 & ~n964;
  assign n5127 = ~n5125 & ~n5126;
  assign n5128 = pi223 & n971;
  assign n5129 = ~pi223 & ~n971;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = ~n5127 & n5130;
  assign n5132 = n5127 & ~n5130;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = pi198 & n955;
  assign n5135 = ~pi198 & ~n955;
  assign n5136 = ~n5134 & ~n5135;
  assign n5137 = ~pi217 & ~n952;
  assign n5138 = pi217 & n952;
  assign n5139 = ~n5137 & ~n5138;
  assign n5140 = ~n5136 & n5139;
  assign n5141 = n5136 & ~n5139;
  assign n5142 = ~n5140 & ~n5141;
  assign n5143 = ~n5133 & n5142;
  assign n5144 = n5133 & ~n5142;
  assign n5145 = ~n5143 & ~n5144;
  assign n5146 = n960 & n5145;
  assign n5147 = ~n5124 & ~n5146;
  assign n5148 = n1466 & n1479;
  assign n5149 = ~n1466 & ~n1479;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~n1518 & n5150;
  assign n5152 = n1518 & ~n5150;
  assign n5153 = ~n5151 & ~n5152;
  assign n5154 = ~n1398 & n1504;
  assign n5155 = n1398 & ~n1504;
  assign n5156 = ~n5154 & ~n5155;
  assign n5157 = ~n1415 & n1425;
  assign n5158 = n1415 & ~n1425;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = ~n1427 & ~n5159;
  assign n5161 = n1415 & n1427;
  assign n5162 = ~n5160 & ~n5161;
  assign n5163 = ~pi129 & ~n5162;
  assign n5164 = ~n1443 & ~n1477;
  assign n5165 = ~n1450 & n5164;
  assign n5166 = n1495 & ~n5165;
  assign n5167 = ~n1496 & n5166;
  assign n5168 = ~n1436 & ~n5167;
  assign n5169 = pi129 & n5168;
  assign n5170 = ~n5163 & ~n5169;
  assign n5171 = pi197 & ~n5170;
  assign n5172 = ~pi197 & n5170;
  assign n5173 = ~n5171 & ~n5172;
  assign n5174 = n1395 & ~n1458;
  assign n5175 = ~n1395 & n1458;
  assign n5176 = ~n5174 & ~n5175;
  assign n5177 = ~n5173 & n5176;
  assign n5178 = n5173 & ~n5176;
  assign n5179 = ~n5177 & ~n5178;
  assign n5180 = ~n5156 & n5179;
  assign n5181 = n5156 & ~n5179;
  assign n5182 = ~n5180 & ~n5181;
  assign n5183 = ~n5153 & n5182;
  assign n5184 = n5153 & ~n5182;
  assign n5185 = ~n5183 & ~n5184;
  assign n5186 = n1087 & ~n5185;
  assign n5187 = n5147 & ~n5186;
  assign n5188 = pi102 & n1090;
  assign n5189 = pi256 & ~n3258;
  assign n5190 = ~n1185 & ~n1195;
  assign n5191 = pi102 & ~n5190;
  assign n5192 = ~n1226 & ~n1233;
  assign n5193 = n1226 & n1233;
  assign n5194 = ~n5192 & ~n5193;
  assign n5195 = n1239 & ~n5194;
  assign n5196 = ~n1237 & n5195;
  assign n5197 = n1237 & ~n5195;
  assign n5198 = ~n5196 & ~n5197;
  assign n5199 = ~n5194 & n5198;
  assign n5200 = n5194 & ~n5198;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = ~n1227 & ~n5201;
  assign n5203 = pi102 & n1189;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = ~n5191 & n5204;
  assign n5206 = ~n5189 & ~n5205;
  assign n5207 = n1307 & ~n1342;
  assign n5208 = ~n1307 & n1342;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = n1254 & ~n1289;
  assign n5211 = ~n1254 & n1289;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = ~n5209 & n5212;
  assign n5214 = n5209 & ~n5212;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = n1217 & ~n1325;
  assign n5217 = ~n1217 & n1325;
  assign n5218 = ~n5216 & ~n5217;
  assign n5219 = n1200 & ~n1272;
  assign n5220 = ~n1200 & n1272;
  assign n5221 = ~n5219 & ~n5220;
  assign n5222 = ~n5218 & n5221;
  assign n5223 = n5218 & ~n5221;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5215 & ~n5224;
  assign n5226 = n5215 & n5224;
  assign n5227 = ~n5225 & ~n5226;
  assign n5228 = n5189 & ~n5227;
  assign n5229 = ~n5206 & ~n5228;
  assign n5230 = ~pi344 & n5229;
  assign n5231 = ~pi102 & pi344;
  assign n5232 = ~n5230 & ~n5231;
  assign n5233 = ~pi243 & n5232;
  assign n5234 = ~n5188 & ~n5233;
  assign n5235 = ~n1377 & n5234;
  assign n5236 = n5187 & n5235;
  assign n5237 = ~n5099 & ~n5236;
  assign n5238 = pi291 & pi301;
  assign n5239 = ~pi302 & n5238;
  assign n5240 = n883 & n3322;
  assign n5241 = ~pi298 & n5240;
  assign n5242 = n5239 & n5241;
  assign n5243 = ~pi193 & ~n5242;
  assign n5244 = n870 & n1366;
  assign n5245 = n787 & n5244;
  assign n5246 = ~pi296 & n5245;
  assign n5247 = n2091 & n5246;
  assign n5248 = pi323 & n5247;
  assign n5249 = pi102 & ~n5247;
  assign n5250 = ~n5248 & ~n5249;
  assign n5251 = ~n2070 & ~n5250;
  assign n5252 = pi102 & n2070;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = n5242 & ~n5253;
  assign n5255 = ~n5243 & ~n5254;
  assign n5256 = n2114 & n3322;
  assign n5257 = pi301 & n5256;
  assign n5258 = n883 & n5257;
  assign n5259 = n782 & n5258;
  assign n5260 = ~n5255 & n5259;
  assign n5261 = ~n5253 & ~n5259;
  assign n5262 = ~n5260 & ~n5261;
  assign n5263 = n5099 & ~n5262;
  assign n5264 = ~n5237 & ~n5263;
  assign n5265 = pi301 & n4978;
  assign n5266 = n2633 & n5265;
  assign n5267 = n5264 & ~n5266;
  assign n5268 = ~pi348 & pi353;
  assign n5269 = pi348 & ~pi353;
  assign n5270 = ~n5268 & ~n5269;
  assign n5271 = pi347 & ~pi349;
  assign n5272 = ~pi347 & pi349;
  assign n5273 = ~n5271 & ~n5272;
  assign n5274 = ~n5270 & n5273;
  assign n5275 = n5270 & ~n5273;
  assign n5276 = ~n5274 & ~n5275;
  assign n5277 = ~pi351 & pi352;
  assign n5278 = pi351 & ~pi352;
  assign n5279 = ~n5277 & ~n5278;
  assign n5280 = ~pi350 & pi354;
  assign n5281 = pi350 & ~pi354;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = ~n5279 & n5282;
  assign n5284 = n5279 & ~n5282;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = ~n5276 & n5285;
  assign n5287 = n5276 & ~n5285;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = n5266 & ~n5288;
  assign n5290 = ~n5267 & ~n5289;
  assign n5291 = n5096 & n5290;
  assign n5292 = pi000 & ~n5096;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n3262 & ~n5293;
  assign n5295 = ~pi231 & ~pi251;
  assign n5296 = ~pi240 & n5295;
  assign n5297 = ~pi239 & n5296;
  assign n5298 = pi234 & n5297;
  assign n5299 = n3541 & n5298;
  assign n5300 = n5293 & ~n5298;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = n3262 & n5301;
  assign n5303 = ~n5294 & ~n5302;
  assign n5304 = ~pi247 & ~n5303;
  assign n5305 = pi102 & pi247;
  assign n5306 = ~n5304 & ~n5305;
  assign po147 = ~pi359 | ~n5306;
  assign n5308 = pi103 & ~n4699;
  assign n5309 = n3363 & n5088;
  assign n5310 = ~pi103 & ~n3363;
  assign n5311 = n4699 & ~n5310;
  assign n5312 = ~n5309 & n5311;
  assign po148 = n5308 | n5312;
  assign n5314 = pi104 & ~n4699;
  assign n5315 = n3370 & n5088;
  assign n5316 = ~pi104 & ~n3370;
  assign n5317 = ~n5315 & ~n5316;
  assign n5318 = n4699 & n5317;
  assign po149 = n5314 | n5318;
  assign n5320 = pi105 & ~n4699;
  assign n5321 = n3377 & n5088;
  assign n5322 = ~pi105 & ~n3377;
  assign n5323 = n4699 & ~n5322;
  assign n5324 = ~n5321 & n5323;
  assign po150 = n5320 | n5324;
  assign n5326 = pi106 & ~n4699;
  assign n5327 = n1603 & n5088;
  assign n5328 = ~pi106 & ~n1603;
  assign n5329 = n4699 & ~n5328;
  assign n5330 = ~n5327 & n5329;
  assign po151 = n5326 | n5330;
  assign n5332 = pi107 & ~n4699;
  assign n5333 = n3390 & n5088;
  assign n5334 = ~pi107 & ~n3390;
  assign n5335 = n4699 & ~n5334;
  assign n5336 = ~n5333 & n5335;
  assign po152 = n5332 | n5336;
  assign n5338 = pi108 & ~n4699;
  assign n5339 = n1619 & n5088;
  assign n5340 = ~pi108 & ~n1619;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = n4699 & n5341;
  assign po153 = n5338 | n5342;
  assign n5344 = pi109 & ~n4699;
  assign n5345 = n1600 & n5088;
  assign n5346 = ~pi109 & ~n1600;
  assign n5347 = n4699 & ~n5346;
  assign n5348 = ~n5345 & n5347;
  assign po154 = n5344 | n5348;
  assign n5350 = pi110 & ~n4699;
  assign n5351 = n1608 & n5060;
  assign n5352 = ~pi110 & ~n1608;
  assign n5353 = n4699 & ~n5352;
  assign n5354 = ~n5351 & n5353;
  assign po155 = n5350 | n5354;
  assign n5356 = pi111 & ~n4699;
  assign n5357 = n3363 & n5060;
  assign n5358 = ~pi111 & ~n3363;
  assign n5359 = n4699 & ~n5358;
  assign n5360 = ~n5357 & n5359;
  assign po156 = n5356 | n5360;
  assign n5362 = pi112 & ~n4699;
  assign n5363 = n3370 & n5060;
  assign n5364 = ~pi112 & ~n3370;
  assign n5365 = n4699 & ~n5364;
  assign n5366 = ~n5363 & n5365;
  assign po157 = n5362 | n5366;
  assign n5368 = pi113 & ~n4699;
  assign n5369 = n3377 & n5060;
  assign n5370 = ~pi113 & ~n3377;
  assign n5371 = n4699 & ~n5370;
  assign n5372 = ~n5369 & n5371;
  assign po158 = n5368 | n5372;
  assign n5374 = pi114 & ~n4699;
  assign n5375 = n1619 & n5060;
  assign n5376 = ~pi114 & ~n1619;
  assign n5377 = n4699 & ~n5376;
  assign n5378 = ~n5375 & n5377;
  assign po159 = n5374 | n5378;
  assign n5380 = pi115 & ~n4699;
  assign n5381 = n1600 & n5060;
  assign n5382 = ~pi115 & ~n1600;
  assign n5383 = n4699 & ~n5382;
  assign n5384 = ~n5381 & n5383;
  assign po160 = n5380 | n5384;
  assign n5386 = pi116 & ~n4699;
  assign n5387 = n3390 & n5060;
  assign n5388 = ~pi116 & ~n3390;
  assign n5389 = n4699 & ~n5388;
  assign n5390 = ~n5387 & n5389;
  assign po161 = n5386 | n5390;
  assign n5392 = n793 & n1559;
  assign n5393 = pi302 & n5392;
  assign n5394 = n2648 & n5393;
  assign n5395 = ~n3824 & n5394;
  assign n5396 = n780 & n1565;
  assign n5397 = ~pi117 & ~n2071;
  assign n5398 = ~n5396 & n5397;
  assign n5399 = ~n5394 & ~n5398;
  assign n5400 = ~n915 & n3264;
  assign n5401 = n782 & ~n3824;
  assign n5402 = pi117 & ~n782;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = ~n782 & ~n1556;
  assign n5405 = pi350 & n782;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = ~n5403 & ~n5406;
  assign n5408 = n5403 & n5406;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = n782 & ~n3754;
  assign n5411 = pi183 & ~n782;
  assign n5412 = ~n5410 & ~n5411;
  assign n5413 = n5406 & n5412;
  assign n5414 = n782 & ~n3684;
  assign n5415 = pi177 & ~n782;
  assign n5416 = ~n5414 & ~n5415;
  assign n5417 = n5406 & n5416;
  assign n5418 = n782 & ~n4334;
  assign n5419 = pi185 & ~n782;
  assign n5420 = ~n5418 & ~n5419;
  assign n5421 = ~n5406 & ~n5420;
  assign n5422 = n5406 & n5420;
  assign n5423 = n782 & ~n4208;
  assign n5424 = pi187 & ~n782;
  assign n5425 = ~n5423 & ~n5424;
  assign n5426 = ~n5406 & ~n5425;
  assign n5427 = ~n5422 & n5426;
  assign n5428 = ~n5421 & ~n5427;
  assign n5429 = n782 & ~n4271;
  assign n5430 = pi135 & ~n782;
  assign n5431 = ~n5429 & ~n5430;
  assign n5432 = ~n5406 & ~n5431;
  assign n5433 = n5406 & n5431;
  assign n5434 = n782 & ~n3200;
  assign n5435 = pi137 & ~n782;
  assign n5436 = ~n5434 & ~n5435;
  assign n5437 = pi347 & n782;
  assign n5438 = ~n5404 & ~n5437;
  assign n5439 = ~n5436 & ~n5438;
  assign n5440 = ~n5433 & n5439;
  assign n5441 = ~n5432 & ~n5440;
  assign n5442 = n782 & ~n3066;
  assign n5443 = pi172 & ~n782;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = pi351 & n782;
  assign n5446 = ~n5404 & ~n5445;
  assign n5447 = n5444 & n5446;
  assign n5448 = n782 & ~n4017;
  assign n5449 = pi174 & ~n782;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~pi354 & n782;
  assign n5452 = ~n5450 & ~n5451;
  assign n5453 = n782 & ~n2680;
  assign n5454 = pi130 & ~n782;
  assign n5455 = ~n5453 & ~n5454;
  assign n5456 = pi349 & n782;
  assign n5457 = ~n5404 & ~n5456;
  assign n5458 = n5455 & n5457;
  assign n5459 = n5452 & ~n5458;
  assign n5460 = ~n5455 & ~n5457;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = n782 & ~n4079;
  assign n5463 = pi173 & ~n782;
  assign n5464 = ~n5462 & ~n5463;
  assign n5465 = pi348 & n782;
  assign n5466 = ~n5404 & ~n5465;
  assign n5467 = n5464 & n5466;
  assign n5468 = ~n5461 & ~n5467;
  assign n5469 = ~n5447 & n5468;
  assign n5470 = ~n5464 & ~n5466;
  assign n5471 = ~n5444 & ~n5446;
  assign n5472 = ~n5467 & n5471;
  assign n5473 = ~n5470 & ~n5472;
  assign n5474 = ~n5469 & n5473;
  assign n5475 = n782 & ~n3956;
  assign n5476 = pi146 & ~n782;
  assign n5477 = ~n5475 & ~n5476;
  assign n5478 = pi352 & n782;
  assign n5479 = ~n5404 & ~n5478;
  assign n5480 = n5477 & n5479;
  assign n5481 = n782 & ~n3132;
  assign n5482 = pi144 & ~n782;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = pi353 & n782;
  assign n5485 = ~n5404 & ~n5484;
  assign n5486 = n5483 & n5485;
  assign n5487 = ~n5480 & ~n5486;
  assign n5488 = ~n5474 & n5487;
  assign n5489 = ~n5483 & ~n5485;
  assign n5490 = ~n5477 & ~n5479;
  assign n5491 = ~n5486 & n5490;
  assign n5492 = ~n5489 & ~n5491;
  assign n5493 = ~n5488 & n5492;
  assign n5494 = n5436 & n5438;
  assign n5495 = ~n5433 & ~n5494;
  assign n5496 = ~n5493 & n5495;
  assign n5497 = n5441 & ~n5496;
  assign n5498 = n5406 & n5425;
  assign n5499 = ~n5422 & ~n5498;
  assign n5500 = ~n5497 & n5499;
  assign n5501 = n5428 & ~n5500;
  assign n5502 = n782 & ~n3612;
  assign n5503 = pi186 & ~n782;
  assign n5504 = ~n5502 & ~n5503;
  assign n5505 = n5406 & n5504;
  assign n5506 = n782 & ~n3893;
  assign n5507 = pi182 & ~n782;
  assign n5508 = ~n5506 & ~n5507;
  assign n5509 = n5406 & n5508;
  assign n5510 = ~n5505 & ~n5509;
  assign n5511 = ~n5501 & n5510;
  assign n5512 = ~n5417 & n5511;
  assign n5513 = ~n5413 & n5512;
  assign n5514 = ~n5406 & ~n5412;
  assign n5515 = ~n5406 & ~n5504;
  assign n5516 = ~n5406 & ~n5508;
  assign n5517 = ~n5505 & n5516;
  assign n5518 = ~n5515 & ~n5517;
  assign n5519 = ~n5417 & ~n5518;
  assign n5520 = ~n5406 & ~n5416;
  assign n5521 = ~n5519 & ~n5520;
  assign n5522 = ~n5413 & ~n5521;
  assign n5523 = ~n5514 & ~n5522;
  assign n5524 = ~n5513 & n5523;
  assign n5525 = n5409 & n5524;
  assign n5526 = ~n5409 & ~n5524;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = n5400 & ~n5527;
  assign n5529 = ~n2071 & ~n5396;
  assign n5530 = n5400 & ~n5529;
  assign n5531 = pi117 & ~n5530;
  assign n5532 = ~n5528 & ~n5531;
  assign n5533 = n5399 & ~n5532;
  assign n5534 = ~n5395 & ~n5533;
  assign n5535 = ~n2070 & ~n5534;
  assign n5536 = pi117 & n2070;
  assign n5537 = ~n5535 & ~n5536;
  assign n5538 = ~n3262 & ~n5537;
  assign n5539 = pi234 & pi240;
  assign n5540 = n5295 & n5539;
  assign n5541 = pi239 & n5540;
  assign n5542 = ~pi239 & n5540;
  assign n5543 = ~n5541 & ~n5542;
  assign n5544 = ~n5541 & ~n5543;
  assign n5545 = ~n5537 & ~n5544;
  assign n5546 = ~n3350 & n5542;
  assign n5547 = ~n5545 & ~n5546;
  assign n5548 = n3262 & ~n5547;
  assign n5549 = ~n5538 & ~n5548;
  assign n5550 = ~pi247 & ~n5549;
  assign n5551 = pi117 & pi247;
  assign n5552 = ~n5550 & ~n5551;
  assign po162 = ~pi359 | ~n5552;
  assign n5554 = pi118 & ~n4699;
  assign n5555 = pi125 & n3287;
  assign n5556 = pi122 & n3290;
  assign n5557 = ~n5555 & ~n5556;
  assign n5558 = pi118 & n3280;
  assign n5559 = pi123 & n3283;
  assign n5560 = ~n5558 & ~n5559;
  assign n5561 = pi119 & n3293;
  assign n5562 = pi124 & n3295;
  assign n5563 = ~n5561 & ~n5562;
  assign n5564 = pi120 & n3298;
  assign n5565 = pi121 & n3300;
  assign n5566 = ~n5564 & ~n5565;
  assign n5567 = n5563 & n5566;
  assign n5568 = n5560 & n5567;
  assign n5569 = n5557 & n5568;
  assign n5570 = n1563 & ~n5569;
  assign n5571 = ~pi267 & n1566;
  assign n5572 = ~n4592 & ~n5571;
  assign n5573 = ~n2025 & n3310;
  assign n5574 = n5572 & ~n5573;
  assign n5575 = ~n1563 & ~n5574;
  assign n5576 = ~n5570 & ~n5575;
  assign n5577 = n3390 & n5576;
  assign n5578 = ~pi118 & ~n3390;
  assign n5579 = n4699 & ~n5578;
  assign n5580 = ~n5577 & n5579;
  assign po163 = n5554 | n5580;
  assign n5582 = pi119 & ~n4699;
  assign n5583 = n1619 & n5576;
  assign n5584 = ~pi119 & ~n1619;
  assign n5585 = n4699 & ~n5584;
  assign n5586 = ~n5583 & n5585;
  assign po164 = n5582 | n5586;
  assign n5588 = pi120 & ~n4699;
  assign n5589 = n1608 & n5576;
  assign n5590 = ~pi120 & ~n1608;
  assign n5591 = n4699 & ~n5590;
  assign n5592 = ~n5589 & n5591;
  assign po165 = n5588 | n5592;
  assign n5594 = pi121 & ~n4699;
  assign n5595 = n3363 & n5576;
  assign n5596 = ~pi121 & ~n3363;
  assign n5597 = n4699 & ~n5596;
  assign n5598 = ~n5595 & n5597;
  assign po166 = n5594 | n5598;
  assign n5600 = pi122 & ~n4699;
  assign n5601 = n3377 & n5576;
  assign n5602 = ~pi122 & ~n3377;
  assign n5603 = n4699 & ~n5602;
  assign n5604 = ~n5601 & n5603;
  assign po167 = n5600 | n5604;
  assign n5606 = pi123 & ~n4699;
  assign n5607 = n1603 & n5576;
  assign n5608 = ~pi123 & ~n1603;
  assign n5609 = n4699 & ~n5608;
  assign n5610 = ~n5607 & n5609;
  assign po168 = n5606 | n5610;
  assign n5612 = pi124 & ~n4699;
  assign n5613 = n1600 & n5576;
  assign n5614 = ~pi124 & ~n1600;
  assign n5615 = n4699 & ~n5614;
  assign n5616 = ~n5613 & n5615;
  assign po169 = n5612 | n5616;
  assign n5618 = pi125 & ~n4699;
  assign n5619 = n3370 & n5576;
  assign n5620 = ~pi125 & ~n3370;
  assign n5621 = n4699 & ~n5620;
  assign n5622 = ~n5619 & n5621;
  assign po170 = n5618 | n5622;
  assign n5624 = pi326 & n5247;
  assign n5625 = pi126 & ~n2633;
  assign n5626 = pi298 & n2091;
  assign n5627 = n787 & n5626;
  assign n5628 = n2218 & n5627;
  assign n5629 = ~pi302 & n5628;
  assign n5630 = n883 & n5629;
  assign n5631 = pi126 & n5630;
  assign n5632 = ~pi126 & ~n5630;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = n2633 & n5633;
  assign n5635 = ~n5625 & ~n5634;
  assign n5636 = ~n5247 & ~n5635;
  assign n5637 = ~n5624 & ~n5636;
  assign n5638 = ~n2070 & ~n5637;
  assign n5639 = pi126 & n2070;
  assign n5640 = ~n5638 & ~n5639;
  assign n5641 = ~n5259 & ~n5640;
  assign n5642 = n5238 & n5241;
  assign n5643 = pi303 & n5642;
  assign n5644 = ~n5242 & ~n5643;
  assign n5645 = pi341 & n5644;
  assign n5646 = n5242 & ~n5640;
  assign n5647 = ~n5242 & n5643;
  assign n5648 = pi292 & n5647;
  assign n5649 = ~n5646 & ~n5648;
  assign n5650 = ~n5645 & n5649;
  assign n5651 = n5258 & ~n5650;
  assign n5652 = n782 & n5651;
  assign n5653 = ~n5641 & ~n5652;
  assign n5654 = ~n3262 & ~n5653;
  assign n5655 = pi251 & n3250;
  assign n5656 = ~pi231 & n5655;
  assign n5657 = ~pi239 & n5656;
  assign n5658 = n5653 & ~n5657;
  assign n5659 = n4834 & n5657;
  assign n5660 = ~n5658 & ~n5659;
  assign n5661 = n3262 & n5660;
  assign n5662 = ~n5654 & ~n5661;
  assign n5663 = ~pi247 & ~n5662;
  assign n5664 = pi126 & pi247;
  assign n5665 = ~n5663 & ~n5664;
  assign po171 = ~pi359 | ~n5665;
  assign n5667 = pi127 & ~n4699;
  assign n5668 = ~pi127 & ~n1603;
  assign n5669 = ~pi260 & n1566;
  assign n5670 = ~n4668 & ~n5669;
  assign n5671 = ~n1972 & n3310;
  assign n5672 = n5670 & ~n5671;
  assign n5673 = ~n1563 & ~n5672;
  assign n5674 = pi158 & n3280;
  assign n5675 = pi127 & n3283;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = pi159 & n3293;
  assign n5678 = pi160 & n3295;
  assign n5679 = ~n5677 & ~n5678;
  assign n5680 = pi154 & n3298;
  assign n5681 = pi155 & n3300;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = pi156 & n3287;
  assign n5684 = pi157 & n3290;
  assign n5685 = ~n5683 & ~n5684;
  assign n5686 = n5682 & n5685;
  assign n5687 = n5679 & n5686;
  assign n5688 = n5676 & n5687;
  assign n5689 = n1563 & ~n5688;
  assign n5690 = ~n5673 & ~n5689;
  assign n5691 = n1603 & n5690;
  assign n5692 = ~n5668 & ~n5691;
  assign n5693 = n4699 & n5692;
  assign po172 = n5667 | n5693;
  assign n5695 = n2364 & n2995;
  assign n5696 = n2313 & n2995;
  assign n5697 = pi273 & ~n5696;
  assign n5698 = pi271 & n5696;
  assign n5699 = ~n5697 & ~n5698;
  assign n5700 = ~n5695 & ~n5699;
  assign n5701 = pi225 & n5695;
  assign n5702 = ~n5700 & ~n5701;
  assign n5703 = n3256 & ~n5702;
  assign n5704 = pi128 & ~n3256;
  assign n5705 = ~n5703 & ~n5704;
  assign n5706 = ~n3262 & ~n5705;
  assign n5707 = pi239 & n5656;
  assign n5708 = n5705 & ~n5707;
  assign n5709 = n4477 & n5707;
  assign n5710 = ~n5708 & ~n5709;
  assign n5711 = n3262 & n5710;
  assign n5712 = ~n5706 & ~n5711;
  assign n5713 = ~pi247 & ~n5712;
  assign n5714 = pi128 & pi247;
  assign n5715 = ~n5713 & ~n5714;
  assign po173 = pi359 & ~n5715;
  assign n5717 = n3255 & n5094;
  assign n5718 = ~n5266 & ~n5717;
  assign n5719 = pi320 & n5247;
  assign n5720 = pi129 & ~n2633;
  assign n5721 = pi302 & n5626;
  assign n5722 = n787 & n5721;
  assign n5723 = n2264 & n5722;
  assign n5724 = ~pi129 & ~n5630;
  assign n5725 = n2633 & ~n5724;
  assign n5726 = n2151 & n5722;
  assign n5727 = n883 & n5726;
  assign n5728 = n5725 & ~n5727;
  assign n5729 = ~n5723 & n5728;
  assign n5730 = ~n5720 & ~n5729;
  assign n5731 = ~n5247 & ~n5730;
  assign n5732 = ~n5719 & ~n5731;
  assign n5733 = ~n2070 & n5099;
  assign n5734 = ~n5732 & n5733;
  assign n5735 = pi129 & n2070;
  assign n5736 = n5099 & n5735;
  assign n5737 = ~n5734 & ~n5736;
  assign n5738 = pi129 & n1090;
  assign n5739 = ~pi243 & n1093;
  assign n5740 = ~n5738 & ~n5739;
  assign n5741 = ~n5099 & ~n5740;
  assign n5742 = n5737 & ~n5741;
  assign n5743 = pi129 & n1087;
  assign n5744 = ~n5099 & n5743;
  assign n5745 = n5742 & ~n5744;
  assign n5746 = n5718 & ~n5745;
  assign n5747 = ~n3262 & n5746;
  assign n5748 = n4667 & n5298;
  assign n5749 = ~n5298 & ~n5746;
  assign n5750 = ~n5748 & ~n5749;
  assign n5751 = n3262 & n5750;
  assign n5752 = ~n5747 & ~n5751;
  assign n5753 = ~pi247 & ~n5752;
  assign n5754 = pi129 & pi247;
  assign n5755 = ~n5753 & ~n5754;
  assign po174 = ~pi359 | ~n5755;
  assign n5757 = pi130 & n2070;
  assign n5758 = pi130 & ~n5400;
  assign n5759 = ~n5458 & ~n5460;
  assign n5760 = n5452 & ~n5759;
  assign n5761 = ~n5452 & n5759;
  assign n5762 = ~n5760 & ~n5761;
  assign n5763 = n5400 & ~n5762;
  assign n5764 = ~n5758 & ~n5763;
  assign n5765 = ~n5529 & ~n5764;
  assign n5766 = pi130 & n5529;
  assign n5767 = ~n5765 & ~n5766;
  assign n5768 = ~n5394 & ~n5767;
  assign n5769 = ~n2680 & n5394;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = ~n2070 & ~n5770;
  assign n5772 = ~n5757 & ~n5771;
  assign n5773 = ~n3262 & ~n5772;
  assign n5774 = ~n5542 & ~n5543;
  assign n5775 = ~n5772 & ~n5774;
  assign n5776 = ~n4667 & n5541;
  assign n5777 = ~n5775 & ~n5776;
  assign n5778 = n3262 & ~n5777;
  assign n5779 = ~n5773 & ~n5778;
  assign n5780 = ~pi247 & ~n5779;
  assign n5781 = pi130 & pi247;
  assign n5782 = ~n5780 & ~n5781;
  assign po175 = ~pi359 | ~n5782;
  assign n5784 = ~n1524 & ~n5099;
  assign n5785 = pi131 & n2070;
  assign n5786 = pi325 & n5247;
  assign n5787 = pi131 & ~n5247;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = ~n2070 & ~n5788;
  assign n5790 = ~n5785 & ~n5789;
  assign n5791 = n5099 & ~n5790;
  assign n5792 = ~n5784 & ~n5791;
  assign n5793 = ~n5266 & ~n5792;
  assign n5794 = ~pi347 & ~pi350;
  assign n5795 = ~pi352 & ~pi354;
  assign n5796 = n5266 & n5795;
  assign n5797 = ~pi353 & n5796;
  assign n5798 = n5794 & n5797;
  assign n5799 = ~pi349 & n5798;
  assign n5800 = ~pi348 & ~pi351;
  assign n5801 = n5799 & n5800;
  assign n5802 = ~n5793 & ~n5801;
  assign n5803 = ~n3262 & ~n5802;
  assign n5804 = n3350 & n5298;
  assign n5805 = ~n5298 & n5802;
  assign n5806 = ~n5804 & ~n5805;
  assign n5807 = n3262 & n5806;
  assign n5808 = ~n5803 & ~n5807;
  assign n5809 = ~pi247 & ~n5808;
  assign n5810 = pi131 & pi247;
  assign n5811 = ~n5809 & ~n5810;
  assign po176 = ~pi359 | ~n5811;
  assign n5813 = pi322 & n5247;
  assign n5814 = pi132 & n5723;
  assign n5815 = ~pi132 & ~n5723;
  assign n5816 = ~n5814 & ~n5815;
  assign n5817 = ~n5727 & ~n5816;
  assign n5818 = n2633 & ~n5817;
  assign n5819 = pi132 & ~n2633;
  assign n5820 = ~n5818 & ~n5819;
  assign n5821 = ~n5247 & ~n5820;
  assign n5822 = ~n5813 & ~n5821;
  assign n5823 = ~n2070 & ~n5822;
  assign n5824 = pi132 & n2070;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = pi335 & ~n5825;
  assign n5827 = ~pi132 & n5170;
  assign n5828 = n1087 & ~n5827;
  assign n5829 = pi223 & ~n1036;
  assign n5830 = pi197 & n842;
  assign n5831 = pi223 & n981;
  assign n5832 = ~n5830 & ~n5831;
  assign n5833 = pi197 & ~n986;
  assign n5834 = ~n1006 & ~n5833;
  assign n5835 = ~n1033 & n5834;
  assign n5836 = n5832 & n5835;
  assign n5837 = ~n5829 & n5836;
  assign n5838 = n977 & ~n5837;
  assign n5839 = ~n5828 & ~n5838;
  assign n5840 = n1093 & n5198;
  assign n5841 = n975 & ~n5198;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~pi243 & ~n5842;
  assign n5844 = n5839 & ~n5843;
  assign n5845 = n1085 & ~n1090;
  assign n5846 = pi132 & ~n5845;
  assign n5847 = n5844 & ~n5846;
  assign n5848 = ~pi335 & ~n5847;
  assign n5849 = ~n5826 & ~n5848;
  assign n5850 = ~n5099 & ~n5849;
  assign n5851 = n5099 & ~n5825;
  assign n5852 = ~n5850 & ~n5851;
  assign n5853 = ~n3262 & ~n5852;
  assign n5854 = n4834 & n5298;
  assign n5855 = ~n5298 & n5852;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = n3262 & n5856;
  assign n5858 = ~n5853 & ~n5857;
  assign n5859 = ~pi247 & ~n5858;
  assign n5860 = pi132 & pi247;
  assign n5861 = ~n5859 & ~n5860;
  assign po177 = ~pi359 | ~n5861;
  assign n5863 = pi330 & n5247;
  assign n5864 = pi133 & ~n2633;
  assign n5865 = pi133 & n5630;
  assign n5866 = ~pi133 & ~n5630;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = n2633 & n5867;
  assign n5869 = ~n5864 & ~n5868;
  assign n5870 = ~n5247 & ~n5869;
  assign n5871 = ~n5863 & ~n5870;
  assign n5872 = ~n2070 & ~n5871;
  assign n5873 = pi133 & n2070;
  assign n5874 = ~n5872 & ~n5873;
  assign n5875 = ~n5259 & ~n5874;
  assign n5876 = n5242 & ~n5874;
  assign n5877 = pi332 & n5647;
  assign n5878 = ~n5876 & ~n5877;
  assign n5879 = pi339 & n5644;
  assign n5880 = n5878 & ~n5879;
  assign n5881 = n5258 & ~n5880;
  assign n5882 = n782 & n5881;
  assign n5883 = ~n5875 & ~n5882;
  assign n5884 = ~n3262 & ~n5883;
  assign n5885 = ~n5657 & ~n5883;
  assign n5886 = ~n4400 & n5657;
  assign n5887 = ~n5885 & ~n5886;
  assign n5888 = n3262 & ~n5887;
  assign n5889 = ~n5884 & ~n5888;
  assign n5890 = ~pi247 & ~n5889;
  assign n5891 = pi133 & pi247;
  assign n5892 = ~n5890 & ~n5891;
  assign po178 = ~pi359 | ~n5892;
  assign n5894 = pi275 & ~n5696;
  assign n5895 = pi272 & n5696;
  assign n5896 = ~n5894 & ~n5895;
  assign n5897 = ~n5695 & ~n5896;
  assign n5898 = pi202 & n5695;
  assign n5899 = ~n5897 & ~n5898;
  assign n5900 = n3256 & ~n5899;
  assign n5901 = pi134 & ~n3256;
  assign n5902 = ~n5900 & ~n5901;
  assign n5903 = ~n3262 & ~n5902;
  assign n5904 = ~n5707 & ~n5902;
  assign n5905 = ~n4400 & n5707;
  assign n5906 = ~n5904 & ~n5905;
  assign n5907 = n3262 & ~n5906;
  assign n5908 = ~n5903 & ~n5907;
  assign n5909 = ~pi247 & ~n5908;
  assign n5910 = pi134 & pi247;
  assign n5911 = ~n5909 & ~n5910;
  assign po179 = pi359 & ~n5911;
  assign n5913 = pi135 & n2070;
  assign n5914 = pi135 & ~n5400;
  assign n5915 = ~n5432 & ~n5433;
  assign n5916 = n5489 & ~n5494;
  assign n5917 = ~n5439 & ~n5916;
  assign n5918 = ~n5486 & ~n5494;
  assign n5919 = n5470 & ~n5480;
  assign n5920 = ~n5490 & ~n5919;
  assign n5921 = n5918 & ~n5920;
  assign n5922 = n5917 & ~n5921;
  assign n5923 = ~n5447 & n5459;
  assign n5924 = ~n5447 & n5460;
  assign n5925 = ~n5471 & ~n5924;
  assign n5926 = ~n5923 & n5925;
  assign n5927 = ~n5467 & ~n5480;
  assign n5928 = n5918 & n5927;
  assign n5929 = ~n5926 & n5928;
  assign n5930 = n5922 & ~n5929;
  assign n5931 = ~n5915 & ~n5930;
  assign n5932 = n5915 & n5930;
  assign n5933 = ~n5931 & ~n5932;
  assign n5934 = n5400 & ~n5933;
  assign n5935 = ~n5914 & ~n5934;
  assign n5936 = ~n5529 & ~n5935;
  assign n5937 = pi135 & n5529;
  assign n5938 = ~n5936 & ~n5937;
  assign n5939 = ~n5394 & ~n5938;
  assign n5940 = ~n4271 & n5394;
  assign n5941 = ~n5939 & ~n5940;
  assign n5942 = ~n2070 & ~n5941;
  assign n5943 = ~n5913 & ~n5942;
  assign n5944 = ~n3262 & ~n5943;
  assign n5945 = ~n4400 & n5541;
  assign n5946 = ~n5774 & ~n5943;
  assign n5947 = ~n5945 & ~n5946;
  assign n5948 = n3262 & ~n5947;
  assign n5949 = ~n5944 & ~n5948;
  assign n5950 = ~pi247 & ~n5949;
  assign n5951 = pi135 & pi247;
  assign n5952 = ~n5950 & ~n5951;
  assign po180 = ~pi359 | ~n5952;
  assign n5954 = pi269 & ~n5696;
  assign n5955 = pi274 & n5696;
  assign n5956 = ~n5954 & ~n5955;
  assign n5957 = ~n5695 & ~n5956;
  assign n5958 = pi215 & n5695;
  assign n5959 = ~n5957 & ~n5958;
  assign n5960 = n3256 & ~n5959;
  assign n5961 = pi136 & ~n3256;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = ~n3262 & ~n5962;
  assign n5964 = ~n5707 & n5962;
  assign n5965 = n3350 & n5707;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = n3262 & n5966;
  assign n5968 = ~n5963 & ~n5967;
  assign n5969 = ~pi247 & ~n5968;
  assign n5970 = pi136 & pi247;
  assign n5971 = ~n5969 & ~n5970;
  assign po181 = pi359 & ~n5971;
  assign n5973 = pi137 & n2070;
  assign n5974 = pi137 & ~n5400;
  assign n5975 = ~n5439 & ~n5494;
  assign n5976 = n5493 & n5975;
  assign n5977 = ~n5493 & ~n5975;
  assign n5978 = ~n5976 & ~n5977;
  assign n5979 = n5400 & ~n5978;
  assign n5980 = ~n5974 & ~n5979;
  assign n5981 = ~n5529 & ~n5980;
  assign n5982 = pi137 & n5529;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = ~n5394 & ~n5983;
  assign n5985 = ~n3200 & n5394;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = ~n2070 & ~n5986;
  assign n5988 = ~n5973 & ~n5987;
  assign n5989 = ~n3262 & ~n5988;
  assign n5990 = ~n3350 & n5541;
  assign n5991 = ~n5774 & ~n5988;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = n3262 & ~n5992;
  assign n5994 = ~n5989 & ~n5993;
  assign n5995 = ~pi247 & ~n5994;
  assign n5996 = pi137 & pi247;
  assign n5997 = ~n5995 & ~n5996;
  assign po182 = ~pi359 | ~n5997;
  assign n5999 = pi316 & n5247;
  assign n6000 = n2633 & n5630;
  assign n6001 = pi138 & ~n6000;
  assign n6002 = ~pi138 & n5630;
  assign n6003 = n2633 & n6002;
  assign n6004 = ~n6001 & ~n6003;
  assign n6005 = ~n5247 & ~n6004;
  assign n6006 = ~n5999 & ~n6005;
  assign n6007 = ~n2070 & ~n6006;
  assign n6008 = pi138 & n2070;
  assign n6009 = ~n6007 & ~n6008;
  assign n6010 = ~n5259 & ~n6009;
  assign n6011 = pi343 & n5644;
  assign n6012 = n5242 & ~n6009;
  assign n6013 = pi288 & n5647;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = ~n6011 & n6014;
  assign n6016 = n5258 & ~n6015;
  assign n6017 = n782 & n6016;
  assign n6018 = ~n6010 & ~n6017;
  assign n6019 = ~n3262 & ~n6018;
  assign n6020 = ~n5657 & n6018;
  assign n6021 = n4591 & n5657;
  assign n6022 = ~n6020 & ~n6021;
  assign n6023 = n3262 & n6022;
  assign n6024 = ~n6019 & ~n6023;
  assign n6025 = ~pi247 & ~n6024;
  assign n6026 = pi138 & pi247;
  assign n6027 = ~n6025 & ~n6026;
  assign po183 = ~pi359 | ~n6027;
  assign n6029 = pi317 & n5247;
  assign n6030 = pi139 & ~n6000;
  assign n6031 = ~pi139 & n5630;
  assign n6032 = n2633 & n6031;
  assign n6033 = ~n6030 & ~n6032;
  assign n6034 = ~n5247 & ~n6033;
  assign n6035 = ~n6029 & ~n6034;
  assign n6036 = ~n2070 & ~n6035;
  assign n6037 = pi139 & n2070;
  assign n6038 = ~n6036 & ~n6037;
  assign n6039 = ~n5259 & ~n6038;
  assign n6040 = pi336 & n5644;
  assign n6041 = n5242 & ~n6038;
  assign n6042 = pi287 & n5647;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = ~n6040 & n6043;
  assign n6045 = n5258 & ~n6044;
  assign n6046 = n782 & n6045;
  assign n6047 = ~n6039 & ~n6046;
  assign n6048 = ~n3262 & ~n6047;
  assign n6049 = ~n5657 & n6047;
  assign n6050 = n4477 & n5657;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = n3262 & n6051;
  assign n6053 = ~n6048 & ~n6052;
  assign n6054 = ~pi247 & ~n6053;
  assign n6055 = pi139 & pi247;
  assign n6056 = ~n6054 & ~n6055;
  assign po184 = ~pi359 | ~n6056;
  assign n6058 = pi329 & n5247;
  assign n6059 = pi140 & ~n2633;
  assign n6060 = pi140 & n5630;
  assign n6061 = ~pi140 & ~n5630;
  assign n6062 = ~n6060 & ~n6061;
  assign n6063 = n2633 & n6062;
  assign n6064 = ~n6059 & ~n6063;
  assign n6065 = ~n5247 & ~n6064;
  assign n6066 = ~n6058 & ~n6065;
  assign n6067 = ~n2070 & ~n6066;
  assign n6068 = pi140 & n2070;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~n5259 & ~n6069;
  assign n6071 = n5242 & ~n6069;
  assign n6072 = pi286 & n5647;
  assign n6073 = ~n6071 & ~n6072;
  assign n6074 = pi340 & n5644;
  assign n6075 = n6073 & ~n6074;
  assign n6076 = n5258 & ~n6075;
  assign n6077 = n782 & n6076;
  assign n6078 = ~n6070 & ~n6077;
  assign n6079 = ~n3262 & ~n6078;
  assign n6080 = ~n5657 & n6078;
  assign n6081 = n3350 & n5657;
  assign n6082 = ~n6080 & ~n6081;
  assign n6083 = n3262 & n6082;
  assign n6084 = ~n6079 & ~n6083;
  assign n6085 = ~pi247 & ~n6084;
  assign n6086 = pi140 & pi247;
  assign n6087 = ~n6085 & ~n6086;
  assign po185 = ~pi359 | ~n6087;
  assign n6089 = pi327 & n5247;
  assign n6090 = pi141 & ~n2633;
  assign n6091 = pi141 & n5630;
  assign n6092 = ~pi141 & ~n5630;
  assign n6093 = ~n6091 & ~n6092;
  assign n6094 = n2633 & n6093;
  assign n6095 = ~n6090 & ~n6094;
  assign n6096 = ~n5247 & ~n6095;
  assign n6097 = ~n6089 & ~n6096;
  assign n6098 = ~n2070 & ~n6097;
  assign n6099 = pi141 & n2070;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = ~n5259 & ~n6100;
  assign n6102 = pi337 & n5644;
  assign n6103 = n5242 & ~n6100;
  assign n6104 = pi289 & n5647;
  assign n6105 = ~n6103 & ~n6104;
  assign n6106 = ~n6102 & n6105;
  assign n6107 = n5258 & ~n6106;
  assign n6108 = n782 & n6107;
  assign n6109 = ~n6101 & ~n6108;
  assign n6110 = ~n3262 & ~n6109;
  assign n6111 = ~n5657 & n6109;
  assign n6112 = n3541 & n5657;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = n3262 & n6113;
  assign n6115 = ~n6110 & ~n6114;
  assign n6116 = ~pi247 & ~n6115;
  assign n6117 = pi141 & pi247;
  assign n6118 = ~n6116 & ~n6117;
  assign po186 = ~pi359 | ~n6118;
  assign n6120 = pi319 & n5247;
  assign n6121 = pi142 & ~n2633;
  assign n6122 = pi142 & n5630;
  assign n6123 = ~pi142 & ~n5630;
  assign n6124 = ~n6122 & ~n6123;
  assign n6125 = n2633 & n6124;
  assign n6126 = ~n6121 & ~n6125;
  assign n6127 = ~n5247 & ~n6126;
  assign n6128 = ~n6120 & ~n6127;
  assign n6129 = ~n2070 & ~n6128;
  assign n6130 = pi142 & n2070;
  assign n6131 = ~n6129 & ~n6130;
  assign n6132 = ~n5259 & ~n6131;
  assign n6133 = n5242 & ~n6131;
  assign n6134 = pi295 & n5647;
  assign n6135 = ~n6133 & ~n6134;
  assign n6136 = pi342 & n5644;
  assign n6137 = n6135 & ~n6136;
  assign n6138 = n5258 & ~n6137;
  assign n6139 = n782 & n6138;
  assign n6140 = ~n6132 & ~n6139;
  assign n6141 = ~n3262 & ~n6140;
  assign n6142 = ~n5657 & n6140;
  assign n6143 = n4667 & n5657;
  assign n6144 = ~n6142 & ~n6143;
  assign n6145 = n3262 & n6144;
  assign n6146 = ~n6141 & ~n6145;
  assign n6147 = ~pi247 & ~n6146;
  assign n6148 = pi142 & pi247;
  assign n6149 = ~n6147 & ~n6148;
  assign po187 = ~pi359 | ~n6149;
  assign n6151 = pi328 & n5247;
  assign n6152 = pi143 & ~n2633;
  assign n6153 = pi143 & n5630;
  assign n6154 = ~pi143 & ~n5630;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = n2633 & n6155;
  assign n6157 = ~n6152 & ~n6156;
  assign n6158 = ~n5247 & ~n6157;
  assign n6159 = ~n6151 & ~n6158;
  assign n6160 = ~n2070 & ~n6159;
  assign n6161 = pi143 & n2070;
  assign n6162 = ~n6160 & ~n6161;
  assign n6163 = ~n5259 & ~n6162;
  assign n6164 = n5242 & ~n6162;
  assign n6165 = pi290 & n5647;
  assign n6166 = ~n6164 & ~n6165;
  assign n6167 = pi338 & n5644;
  assign n6168 = n6166 & ~n6167;
  assign n6169 = n5258 & ~n6168;
  assign n6170 = n782 & n6169;
  assign n6171 = ~n6163 & ~n6170;
  assign n6172 = ~n3262 & ~n6171;
  assign n6173 = ~n5657 & n6171;
  assign n6174 = n3447 & n5657;
  assign n6175 = ~n6173 & ~n6174;
  assign n6176 = n3262 & n6175;
  assign n6177 = ~n6172 & ~n6176;
  assign n6178 = ~pi247 & ~n6177;
  assign n6179 = pi143 & pi247;
  assign n6180 = ~n6178 & ~n6179;
  assign po188 = ~pi359 | ~n6180;
  assign n6182 = pi144 & n2070;
  assign n6183 = pi144 & ~n5400;
  assign n6184 = ~n5486 & ~n5489;
  assign n6185 = n5459 & n5927;
  assign n6186 = ~n5447 & n6185;
  assign n6187 = ~n5925 & n5927;
  assign n6188 = n5920 & ~n6187;
  assign n6189 = ~n6186 & n6188;
  assign n6190 = n6184 & n6189;
  assign n6191 = ~n6184 & ~n6189;
  assign n6192 = ~n6190 & ~n6191;
  assign n6193 = n5400 & ~n6192;
  assign n6194 = ~n6183 & ~n6193;
  assign n6195 = ~n5529 & ~n6194;
  assign n6196 = pi144 & n5529;
  assign n6197 = ~n6195 & ~n6196;
  assign n6198 = ~n5394 & ~n6197;
  assign n6199 = ~n3132 & n5394;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n2070 & ~n6200;
  assign n6202 = ~n6182 & ~n6201;
  assign n6203 = ~n3262 & ~n6202;
  assign n6204 = ~n4477 & n5541;
  assign n6205 = ~n5774 & ~n6202;
  assign n6206 = ~n6204 & ~n6205;
  assign n6207 = n3262 & ~n6206;
  assign n6208 = ~n6203 & ~n6207;
  assign n6209 = ~pi247 & ~n6208;
  assign n6210 = pi144 & pi247;
  assign n6211 = ~n6209 & ~n6210;
  assign po189 = ~pi359 | ~n6211;
  assign n6213 = pi270 & ~n5696;
  assign n6214 = pi264 & n5696;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = ~n5695 & ~n6215;
  assign n6217 = pi197 & n5695;
  assign n6218 = ~n6216 & ~n6217;
  assign n6219 = n3256 & ~n6218;
  assign n6220 = pi145 & ~n3256;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = ~n3262 & ~n6221;
  assign n6223 = ~n5707 & n6221;
  assign n6224 = n3447 & n5707;
  assign n6225 = ~n6223 & ~n6224;
  assign n6226 = n3262 & n6225;
  assign n6227 = ~n6222 & ~n6226;
  assign n6228 = ~pi247 & ~n6227;
  assign n6229 = pi145 & pi247;
  assign n6230 = ~n6228 & ~n6229;
  assign po190 = pi359 & ~n6230;
  assign n6232 = pi146 & n2070;
  assign n6233 = pi146 & ~n5400;
  assign n6234 = ~n5480 & ~n5490;
  assign n6235 = n5474 & n6234;
  assign n6236 = ~n5474 & ~n6234;
  assign n6237 = ~n6235 & ~n6236;
  assign n6238 = n5400 & ~n6237;
  assign n6239 = ~n6233 & ~n6238;
  assign n6240 = ~n5529 & ~n6239;
  assign n6241 = pi146 & n5529;
  assign n6242 = ~n6240 & ~n6241;
  assign n6243 = ~n5394 & ~n6242;
  assign n6244 = ~n3956 & n5394;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = ~n2070 & ~n6245;
  assign n6247 = ~n6232 & ~n6246;
  assign n6248 = ~n3262 & ~n6247;
  assign n6249 = ~n3447 & n5541;
  assign n6250 = ~n5774 & ~n6247;
  assign n6251 = ~n6249 & ~n6250;
  assign n6252 = n3262 & ~n6251;
  assign n6253 = ~n6248 & ~n6252;
  assign n6254 = ~pi247 & ~n6253;
  assign n6255 = pi146 & pi247;
  assign n6256 = ~n6254 & ~n6255;
  assign po191 = ~pi359 | ~n6256;
  assign n6258 = pi147 & ~n4699;
  assign n6259 = ~pi147 & ~n1608;
  assign n6260 = ~pi261 & n1566;
  assign n6261 = ~n3542 & ~n6260;
  assign n6262 = ~n1968 & n3310;
  assign n6263 = n6261 & ~n6262;
  assign n6264 = ~n1563 & ~n6263;
  assign n6265 = pi151 & n3280;
  assign n6266 = pi175 & n3283;
  assign n6267 = ~n6265 & ~n6266;
  assign n6268 = pi152 & n3293;
  assign n6269 = pi153 & n3295;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = pi147 & n3298;
  assign n6272 = pi148 & n3300;
  assign n6273 = ~n6271 & ~n6272;
  assign n6274 = pi149 & n3287;
  assign n6275 = pi150 & n3290;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = n6273 & n6276;
  assign n6278 = n6270 & n6277;
  assign n6279 = n6267 & n6278;
  assign n6280 = n1563 & ~n6279;
  assign n6281 = ~n6264 & ~n6280;
  assign n6282 = n1608 & n6281;
  assign n6283 = ~n6259 & ~n6282;
  assign n6284 = n4699 & n6283;
  assign po192 = n6258 | n6284;
  assign n6286 = pi148 & ~n4699;
  assign n6287 = ~pi148 & ~n3363;
  assign n6288 = n3363 & n6281;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = n4699 & n6289;
  assign po193 = n6286 | n6290;
  assign n6292 = pi149 & ~n4699;
  assign n6293 = ~pi149 & ~n3370;
  assign n6294 = n3370 & n6281;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = n4699 & n6295;
  assign po194 = n6292 | n6296;
  assign n6298 = pi150 & ~n4699;
  assign n6299 = ~pi150 & ~n3377;
  assign n6300 = n3377 & n6281;
  assign n6301 = ~n6299 & ~n6300;
  assign n6302 = n4699 & n6301;
  assign po195 = n6298 | n6302;
  assign n6304 = pi151 & ~n4699;
  assign n6305 = ~pi151 & ~n3390;
  assign n6306 = n3390 & n6281;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = n4699 & n6307;
  assign po196 = n6304 | n6308;
  assign n6310 = pi152 & ~n4699;
  assign n6311 = ~pi152 & ~n1619;
  assign n6312 = n1619 & n6281;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = n4699 & n6313;
  assign po197 = n6310 | n6314;
  assign n6316 = pi153 & ~n4699;
  assign n6317 = ~pi153 & ~n1600;
  assign n6318 = n1600 & n6281;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = n4699 & n6319;
  assign po198 = n6316 | n6320;
  assign n6322 = pi154 & ~n4699;
  assign n6323 = n1608 & n5690;
  assign n6324 = ~pi154 & ~n1608;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = n4699 & n6325;
  assign po199 = n6322 | n6326;
  assign n6328 = pi155 & ~n4699;
  assign n6329 = n3363 & n5690;
  assign n6330 = ~pi155 & ~n3363;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = n4699 & n6331;
  assign po200 = n6328 | n6332;
  assign n6334 = pi156 & ~n4699;
  assign n6335 = n3370 & n5690;
  assign n6336 = ~pi156 & ~n3370;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = n4699 & n6337;
  assign po201 = n6334 | n6338;
  assign n6340 = pi157 & ~n4699;
  assign n6341 = ~pi157 & ~n3377;
  assign n6342 = n3377 & n5690;
  assign n6343 = ~n6341 & ~n6342;
  assign n6344 = n4699 & n6343;
  assign po202 = n6340 | n6344;
  assign n6346 = pi158 & ~n4699;
  assign n6347 = ~pi158 & ~n3390;
  assign n6348 = n3390 & n5690;
  assign n6349 = ~n6347 & ~n6348;
  assign n6350 = n4699 & n6349;
  assign po203 = n6346 | n6350;
  assign n6352 = pi159 & ~n4699;
  assign n6353 = ~pi159 & ~n1619;
  assign n6354 = n1619 & n5690;
  assign n6355 = ~n6353 & ~n6354;
  assign n6356 = n4699 & n6355;
  assign po204 = n6352 | n6356;
  assign n6358 = pi160 & ~n4699;
  assign n6359 = ~pi160 & ~n1600;
  assign n6360 = n1600 & n5690;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = n4699 & n6361;
  assign po205 = n6358 | n6362;
  assign n6364 = pi264 & ~n5696;
  assign n6365 = pi197 & n5696;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n5695 & ~n6366;
  assign n6368 = pi270 & n5695;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = n3256 & ~n6369;
  assign n6371 = pi161 & ~n3256;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = ~n3262 & ~n6372;
  assign n6374 = ~n5707 & n6372;
  assign n6375 = n4834 & n5707;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = n3262 & n6376;
  assign n6378 = ~n6373 & ~n6377;
  assign n6379 = ~pi247 & ~n6378;
  assign n6380 = pi161 & pi247;
  assign n6381 = ~n6379 & ~n6380;
  assign po206 = pi359 & ~n6381;
  assign n6383 = pi271 & ~n5696;
  assign n6384 = pi225 & n5696;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n5695 & ~n6385;
  assign n6387 = pi273 & n5695;
  assign n6388 = ~n6386 & ~n6387;
  assign n6389 = n3256 & ~n6388;
  assign n6390 = pi162 & ~n3256;
  assign n6391 = ~n6389 & ~n6390;
  assign n6392 = ~n3262 & ~n6391;
  assign n6393 = ~n5707 & n6391;
  assign n6394 = n4667 & n5707;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = n3262 & n6395;
  assign n6397 = ~n6392 & ~n6396;
  assign n6398 = ~pi247 & ~n6397;
  assign n6399 = pi162 & pi247;
  assign n6400 = ~n6398 & ~n6399;
  assign po207 = pi359 & ~n6400;
  assign n6402 = pi274 & ~n5696;
  assign n6403 = pi215 & n5696;
  assign n6404 = ~n6402 & ~n6403;
  assign n6405 = ~n5695 & ~n6404;
  assign n6406 = pi269 & n5695;
  assign n6407 = ~n6405 & ~n6406;
  assign n6408 = n3256 & ~n6407;
  assign n6409 = pi163 & ~n3256;
  assign n6410 = ~n6408 & ~n6409;
  assign n6411 = ~n3262 & ~n6410;
  assign n6412 = ~n5707 & n6410;
  assign n6413 = n3541 & n5707;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = n3262 & n6414;
  assign n6416 = ~n6411 & ~n6415;
  assign n6417 = ~pi247 & ~n6416;
  assign n6418 = pi163 & pi247;
  assign n6419 = ~n6417 & ~n6418;
  assign po208 = pi359 & ~n6419;
  assign n6421 = pi272 & ~n5696;
  assign n6422 = pi202 & n5696;
  assign n6423 = ~n6421 & ~n6422;
  assign n6424 = ~n5695 & ~n6423;
  assign n6425 = pi275 & n5695;
  assign n6426 = ~n6424 & ~n6425;
  assign n6427 = n3256 & ~n6426;
  assign n6428 = pi164 & ~n3256;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n3262 & ~n6429;
  assign n6431 = ~n5707 & n6429;
  assign n6432 = n4591 & n5707;
  assign n6433 = ~n6431 & ~n6432;
  assign n6434 = n3262 & n6433;
  assign n6435 = ~n6430 & ~n6434;
  assign n6436 = ~pi247 & ~n6435;
  assign n6437 = pi164 & pi247;
  assign n6438 = ~n6436 & ~n6437;
  assign po209 = pi359 & ~n6438;
  assign n6440 = pi165 & ~n4699;
  assign n6441 = n1780 & n3310;
  assign n6442 = ~pi235 & n1566;
  assign n6443 = ~n6441 & ~n6442;
  assign n6444 = ~n4835 & n6443;
  assign n6445 = ~n1563 & ~n6444;
  assign n6446 = pi170 & n3280;
  assign n6447 = pi169 & n3283;
  assign n6448 = ~n6446 & ~n6447;
  assign n6449 = pi176 & n3293;
  assign n6450 = pi171 & n3295;
  assign n6451 = ~n6449 & ~n6450;
  assign n6452 = pi165 & n3298;
  assign n6453 = pi166 & n3300;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = pi167 & n3287;
  assign n6456 = pi168 & n3290;
  assign n6457 = ~n6455 & ~n6456;
  assign n6458 = n6454 & n6457;
  assign n6459 = n6451 & n6458;
  assign n6460 = n6448 & n6459;
  assign n6461 = n1563 & ~n6460;
  assign n6462 = ~n6445 & ~n6461;
  assign n6463 = n1608 & n6462;
  assign n6464 = ~pi165 & ~n1608;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = n4699 & n6465;
  assign po210 = n6440 | n6466;
  assign n6468 = pi166 & ~n4699;
  assign n6469 = n3363 & n6462;
  assign n6470 = ~pi166 & ~n3363;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = n4699 & n6471;
  assign po211 = n6468 | n6472;
  assign n6474 = pi167 & ~n4699;
  assign n6475 = n3370 & n6462;
  assign n6476 = ~pi167 & ~n3370;
  assign n6477 = ~n6475 & ~n6476;
  assign n6478 = n4699 & n6477;
  assign po212 = n6474 | n6478;
  assign n6480 = pi168 & ~n4699;
  assign n6481 = ~pi168 & ~n3377;
  assign n6482 = n3377 & n6462;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = n4699 & n6483;
  assign po213 = n6480 | n6484;
  assign n6486 = pi169 & ~n4699;
  assign n6487 = ~pi169 & ~n1603;
  assign n6488 = n1603 & n6462;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = n4699 & n6489;
  assign po214 = n6486 | n6490;
  assign n6492 = pi170 & ~n4699;
  assign n6493 = ~pi170 & ~n3390;
  assign n6494 = n3390 & n6462;
  assign n6495 = ~n6493 & ~n6494;
  assign n6496 = n4699 & n6495;
  assign po215 = n6492 | n6496;
  assign n6498 = pi171 & ~n4699;
  assign n6499 = ~pi171 & ~n1600;
  assign n6500 = n1600 & n6462;
  assign n6501 = ~n6499 & ~n6500;
  assign n6502 = n4699 & n6501;
  assign po216 = n6498 | n6502;
  assign n6504 = pi172 & n2070;
  assign n6505 = pi172 & ~n5400;
  assign n6506 = ~n5447 & ~n5471;
  assign n6507 = ~n5461 & ~n6506;
  assign n6508 = n5461 & n6506;
  assign n6509 = ~n6507 & ~n6508;
  assign n6510 = n5400 & ~n6509;
  assign n6511 = ~n6505 & ~n6510;
  assign n6512 = ~n5529 & ~n6511;
  assign n6513 = pi172 & n5529;
  assign n6514 = ~n6512 & ~n6513;
  assign n6515 = ~n5394 & ~n6514;
  assign n6516 = ~n3066 & n5394;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = ~n2070 & ~n6517;
  assign n6519 = ~n6504 & ~n6518;
  assign n6520 = ~n3262 & ~n6519;
  assign n6521 = ~n3541 & n5541;
  assign n6522 = ~n5774 & ~n6519;
  assign n6523 = ~n6521 & ~n6522;
  assign n6524 = n3262 & ~n6523;
  assign n6525 = ~n6520 & ~n6524;
  assign n6526 = ~pi247 & ~n6525;
  assign n6527 = pi172 & pi247;
  assign n6528 = ~n6526 & ~n6527;
  assign po217 = ~pi359 | ~n6528;
  assign n6530 = pi173 & n2070;
  assign n6531 = pi173 & ~n5400;
  assign n6532 = ~n5467 & ~n5470;
  assign n6533 = n5926 & n6532;
  assign n6534 = ~n5926 & ~n6532;
  assign n6535 = ~n6533 & ~n6534;
  assign n6536 = n5400 & ~n6535;
  assign n6537 = ~n6531 & ~n6536;
  assign n6538 = ~n5529 & ~n6537;
  assign n6539 = pi173 & n5529;
  assign n6540 = ~n6538 & ~n6539;
  assign n6541 = ~n5394 & ~n6540;
  assign n6542 = ~n4079 & n5394;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = ~n2070 & ~n6543;
  assign n6545 = ~n6530 & ~n6544;
  assign n6546 = ~n3262 & ~n6545;
  assign n6547 = ~n5774 & ~n6545;
  assign n6548 = ~n4591 & n5541;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = n3262 & ~n6549;
  assign n6551 = ~n6546 & ~n6550;
  assign n6552 = ~pi247 & ~n6551;
  assign n6553 = pi173 & pi247;
  assign n6554 = ~n6552 & ~n6553;
  assign po218 = ~pi359 | ~n6554;
  assign n6556 = pi174 & n2070;
  assign n6557 = pi174 & ~n5400;
  assign n6558 = ~n5450 & n5451;
  assign n6559 = n5450 & ~n5451;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = n5400 & ~n6560;
  assign n6562 = ~n6557 & ~n6561;
  assign n6563 = ~n5529 & ~n6562;
  assign n6564 = pi174 & n5529;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = ~n5394 & ~n6565;
  assign n6567 = ~n4017 & n5394;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = ~n2070 & ~n6568;
  assign n6570 = ~n6556 & ~n6569;
  assign n6571 = ~n3262 & ~n6570;
  assign n6572 = ~n4834 & n5541;
  assign n6573 = ~n5774 & ~n6570;
  assign n6574 = ~n6572 & ~n6573;
  assign n6575 = n3262 & ~n6574;
  assign n6576 = ~n6571 & ~n6575;
  assign n6577 = ~pi247 & ~n6576;
  assign n6578 = pi174 & pi247;
  assign n6579 = ~n6577 & ~n6578;
  assign po219 = ~pi359 | ~n6579;
  assign n6581 = pi175 & ~n4699;
  assign n6582 = ~pi175 & ~n1603;
  assign n6583 = n1603 & n6281;
  assign n6584 = ~n6582 & ~n6583;
  assign n6585 = n4699 & n6584;
  assign po220 = n6581 | n6585;
  assign n6587 = pi176 & ~n4699;
  assign n6588 = ~pi176 & ~n1619;
  assign n6589 = n1619 & n6462;
  assign n6590 = ~n6588 & ~n6589;
  assign n6591 = n4699 & n6590;
  assign po221 = n6587 | n6591;
  assign n6593 = ~n3447 & n5542;
  assign n6594 = pi177 & ~n5400;
  assign n6595 = ~n5417 & ~n5520;
  assign n6596 = n5487 & n5495;
  assign n6597 = ~n5474 & n5499;
  assign n6598 = n6596 & n6597;
  assign n6599 = n5510 & n6598;
  assign n6600 = ~n5492 & n5495;
  assign n6601 = n5441 & ~n6600;
  assign n6602 = n5499 & ~n6601;
  assign n6603 = n5428 & ~n6602;
  assign n6604 = n5510 & ~n6603;
  assign n6605 = n5518 & ~n6604;
  assign n6606 = ~n6599 & n6605;
  assign n6607 = n6595 & n6606;
  assign n6608 = ~n6595 & ~n6606;
  assign n6609 = ~n6607 & ~n6608;
  assign n6610 = n5400 & ~n6609;
  assign n6611 = ~n6594 & ~n6610;
  assign n6612 = ~n5529 & ~n6611;
  assign n6613 = pi177 & n5529;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = ~n5394 & ~n6614;
  assign n6616 = ~n3684 & n5394;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = ~n2070 & ~n6617;
  assign n6619 = pi177 & n2070;
  assign n6620 = ~n6618 & ~n6619;
  assign n6621 = ~n5544 & ~n6620;
  assign n6622 = ~n6593 & ~n6621;
  assign n6623 = n3262 & ~n6622;
  assign n6624 = ~n3262 & ~n6620;
  assign n6625 = ~n6623 & ~n6624;
  assign n6626 = ~pi247 & ~n6625;
  assign n6627 = pi177 & pi247;
  assign n6628 = ~n6626 & ~n6627;
  assign po222 = ~pi359 | ~n6628;
  assign n6630 = ~n4400 & n5298;
  assign n6631 = pi318 & n5247;
  assign n6632 = pi178 & ~n5247;
  assign n6633 = ~n6631 & ~n6632;
  assign n6634 = ~n2070 & ~n6633;
  assign n6635 = pi178 & n2070;
  assign n6636 = ~n6634 & ~n6635;
  assign n6637 = n5099 & ~n6636;
  assign n6638 = ~pi344 & ~n1254;
  assign n6639 = pi178 & pi344;
  assign n6640 = ~n6638 & ~n6639;
  assign n6641 = ~pi243 & ~n6640;
  assign n6642 = pi178 & n1090;
  assign n6643 = ~n6641 & ~n6642;
  assign n6644 = pi178 & n787;
  assign n6645 = ~n787 & ~n1040;
  assign n6646 = ~n6644 & ~n6645;
  assign n6647 = n977 & ~n6646;
  assign n6648 = ~n4386 & n4393;
  assign n6649 = ~n6647 & n6648;
  assign n6650 = n6643 & n6649;
  assign n6651 = ~n5099 & ~n6650;
  assign n6652 = ~n6637 & ~n6651;
  assign n6653 = ~n5266 & ~n6652;
  assign n6654 = pi350 & n5266;
  assign n6655 = ~n6653 & ~n6654;
  assign n6656 = ~n5298 & ~n6655;
  assign n6657 = ~n6630 & ~n6656;
  assign n6658 = n3262 & ~n6657;
  assign n6659 = ~n3262 & ~n6655;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = ~pi247 & ~n6660;
  assign n6662 = pi178 & pi247;
  assign n6663 = ~n6661 & ~n6662;
  assign po223 = ~pi359 | ~n6663;
  assign n6665 = ~n4400 & n5542;
  assign n6666 = n2648 & n4142;
  assign n6667 = n5393 & n6666;
  assign n6668 = pi179 & n5529;
  assign n6669 = ~n5394 & ~n6668;
  assign n6670 = pi179 & ~n5400;
  assign n6671 = n782 & ~n4142;
  assign n6672 = pi179 & ~n782;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = ~n5406 & ~n6673;
  assign n6675 = n5406 & n6673;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = n5406 & ~n5514;
  assign n6678 = ~n5407 & n5408;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = n5403 & ~n5514;
  assign n6681 = n6679 & ~n6680;
  assign n6682 = ~n5408 & ~n5413;
  assign n6683 = ~n5417 & n5515;
  assign n6684 = ~n5520 & ~n6683;
  assign n6685 = n6682 & ~n6684;
  assign n6686 = ~n6681 & ~n6685;
  assign n6687 = ~n5417 & ~n5505;
  assign n6688 = n6682 & n6687;
  assign n6689 = n5421 & ~n5509;
  assign n6690 = ~n5516 & ~n6689;
  assign n6691 = ~n5433 & ~n5498;
  assign n6692 = ~n5422 & ~n5509;
  assign n6693 = ~n5930 & n6692;
  assign n6694 = n6691 & n6693;
  assign n6695 = n5432 & ~n5498;
  assign n6696 = ~n5426 & ~n6695;
  assign n6697 = n6692 & ~n6696;
  assign n6698 = ~n6694 & ~n6697;
  assign n6699 = n6690 & n6698;
  assign n6700 = n6688 & ~n6699;
  assign n6701 = n6686 & ~n6700;
  assign n6702 = ~n6676 & ~n6701;
  assign n6703 = n6676 & n6701;
  assign n6704 = ~n6702 & ~n6703;
  assign n6705 = n5400 & ~n6704;
  assign n6706 = ~n6670 & ~n6705;
  assign n6707 = ~n5529 & ~n6706;
  assign n6708 = n6669 & ~n6707;
  assign n6709 = ~n6667 & ~n6708;
  assign n6710 = ~n2070 & n6709;
  assign n6711 = pi179 & n2070;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~n5544 & ~n6712;
  assign n6714 = ~n6665 & ~n6713;
  assign n6715 = n3262 & ~n6714;
  assign n6716 = ~n3262 & ~n6712;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = ~pi247 & ~n6717;
  assign n6719 = pi179 & pi247;
  assign n6720 = ~n6718 & ~n6719;
  assign po224 = ~pi359 | ~n6720;
  assign n6722 = pi321 & n5247;
  assign n6723 = pi138 & n5727;
  assign n6724 = pi138 & n5723;
  assign n6725 = ~pi180 & ~n5630;
  assign n6726 = ~n6002 & ~n6725;
  assign n6727 = ~n5723 & ~n6726;
  assign n6728 = ~n6724 & ~n6727;
  assign n6729 = ~n5727 & ~n6728;
  assign n6730 = ~n6723 & ~n6729;
  assign n6731 = n2633 & ~n6730;
  assign n6732 = ~pi180 & ~n2633;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = ~n5247 & ~n6733;
  assign n6735 = ~n6722 & ~n6734;
  assign n6736 = ~n2070 & ~n6735;
  assign n6737 = ~pi180 & n2070;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = n5099 & ~n6738;
  assign n6740 = pi272 & n3259;
  assign n6741 = ~n1325 & ~n3259;
  assign n6742 = ~n6740 & ~n6741;
  assign n6743 = ~pi243 & ~n6742;
  assign n6744 = pi272 & ~n2793;
  assign n6745 = n1084 & n6744;
  assign n6746 = ~pi180 & n1090;
  assign n6747 = ~n6745 & ~n6746;
  assign n6748 = n4580 & ~n4583;
  assign n6749 = n6747 & n6748;
  assign n6750 = ~n6743 & n6749;
  assign n6751 = ~n5099 & ~n6750;
  assign n6752 = ~n6739 & ~n6751;
  assign n6753 = ~n5717 & ~n6752;
  assign n6754 = ~n4587 & n5717;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = ~n5298 & ~n6755;
  assign n6757 = ~n4591 & n5298;
  assign n6758 = ~n6756 & ~n6757;
  assign n6759 = n3262 & ~n6758;
  assign n6760 = ~n3262 & ~n6755;
  assign n6761 = ~n6759 & ~n6760;
  assign n6762 = ~pi247 & ~n6761;
  assign n6763 = ~pi180 & pi247;
  assign n6764 = ~n6762 & ~n6763;
  assign po225 = ~pi359 | ~n6764;
  assign n6766 = pi315 & n5247;
  assign n6767 = pi139 & n5727;
  assign n6768 = pi139 & n5723;
  assign n6769 = ~pi181 & ~n5630;
  assign n6770 = ~n6031 & ~n6769;
  assign n6771 = ~n5723 & ~n6770;
  assign n6772 = ~n6768 & ~n6771;
  assign n6773 = ~n5727 & ~n6772;
  assign n6774 = ~n6767 & ~n6773;
  assign n6775 = n2633 & ~n6774;
  assign n6776 = ~pi181 & ~n2633;
  assign n6777 = ~n6775 & ~n6776;
  assign n6778 = ~n5247 & ~n6777;
  assign n6779 = ~n6766 & ~n6778;
  assign n6780 = ~n2070 & ~n6779;
  assign n6781 = ~pi181 & n2070;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = n5099 & ~n6782;
  assign n6784 = pi273 & n3259;
  assign n6785 = ~n1217 & ~n3259;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = ~pi243 & ~n6786;
  assign n6788 = pi273 & ~n2793;
  assign n6789 = n1084 & n6788;
  assign n6790 = ~pi181 & n1090;
  assign n6791 = ~n6789 & ~n6790;
  assign n6792 = ~n4463 & n4470;
  assign n6793 = n6791 & n6792;
  assign n6794 = ~n6787 & n6793;
  assign n6795 = ~n5099 & ~n6794;
  assign n6796 = ~n6783 & ~n6795;
  assign n6797 = ~n5717 & ~n6796;
  assign n6798 = ~n4663 & n5717;
  assign n6799 = ~n6797 & ~n6798;
  assign n6800 = ~n5298 & ~n6799;
  assign n6801 = ~n4477 & n5298;
  assign n6802 = ~n6800 & ~n6801;
  assign n6803 = n3262 & ~n6802;
  assign n6804 = ~n3262 & ~n6799;
  assign n6805 = ~n6803 & ~n6804;
  assign n6806 = ~pi247 & ~n6805;
  assign n6807 = ~pi181 & pi247;
  assign n6808 = ~n6806 & ~n6807;
  assign po226 = ~pi359 | ~n6808;
  assign n6810 = ~n3541 & n5542;
  assign n6811 = n2648 & n3893;
  assign n6812 = n5393 & n6811;
  assign n6813 = pi182 & n5529;
  assign n6814 = ~n5394 & ~n6813;
  assign n6815 = pi182 & ~n5400;
  assign n6816 = ~n5509 & ~n5516;
  assign n6817 = n5501 & n6816;
  assign n6818 = ~n5501 & ~n6816;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = n5400 & ~n6819;
  assign n6821 = ~n6815 & ~n6820;
  assign n6822 = ~n5529 & ~n6821;
  assign n6823 = n6814 & ~n6822;
  assign n6824 = ~n6812 & ~n6823;
  assign n6825 = ~n2070 & n6824;
  assign n6826 = pi182 & n2070;
  assign n6827 = ~n6825 & ~n6826;
  assign n6828 = ~n5544 & ~n6827;
  assign n6829 = ~n6810 & ~n6828;
  assign n6830 = n3262 & ~n6829;
  assign n6831 = ~n3262 & ~n6827;
  assign n6832 = ~n6830 & ~n6831;
  assign n6833 = ~pi247 & ~n6832;
  assign n6834 = pi182 & pi247;
  assign n6835 = ~n6833 & ~n6834;
  assign po227 = ~pi359 | ~n6835;
  assign n6837 = ~n4477 & n5542;
  assign n6838 = n2648 & n3754;
  assign n6839 = n5393 & n6838;
  assign n6840 = pi183 & n5529;
  assign n6841 = ~n5394 & ~n6840;
  assign n6842 = pi183 & ~n5400;
  assign n6843 = ~n5413 & ~n5514;
  assign n6844 = n5918 & n6691;
  assign n6845 = ~n6189 & n6687;
  assign n6846 = n6844 & n6845;
  assign n6847 = n6692 & n6846;
  assign n6848 = ~n5917 & n6691;
  assign n6849 = n6696 & ~n6848;
  assign n6850 = n6692 & ~n6849;
  assign n6851 = n6690 & ~n6850;
  assign n6852 = n6687 & ~n6851;
  assign n6853 = n6684 & ~n6852;
  assign n6854 = ~n6847 & n6853;
  assign n6855 = n6843 & n6854;
  assign n6856 = ~n6843 & ~n6854;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = n5400 & ~n6857;
  assign n6859 = ~n6842 & ~n6858;
  assign n6860 = ~n5529 & ~n6859;
  assign n6861 = n6841 & ~n6860;
  assign n6862 = ~n6839 & ~n6861;
  assign n6863 = ~n2070 & n6862;
  assign n6864 = pi183 & n2070;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = ~n5544 & ~n6865;
  assign n6867 = ~n6837 & ~n6866;
  assign n6868 = n3262 & ~n6867;
  assign n6869 = ~n3262 & ~n6865;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = ~pi247 & ~n6870;
  assign n6872 = pi183 & pi247;
  assign n6873 = ~n6871 & ~n6872;
  assign po228 = ~pi359 | ~n6873;
  assign n6875 = ~n3447 & n5298;
  assign n6876 = pi324 & n5247;
  assign n6877 = ~pi184 & ~n5630;
  assign n6878 = ~n5723 & ~n6877;
  assign n6879 = ~n5814 & ~n6878;
  assign n6880 = ~n5727 & ~n6879;
  assign n6881 = n2633 & n6880;
  assign n6882 = pi184 & ~n2633;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n5247 & ~n6883;
  assign n6885 = ~n6876 & ~n6884;
  assign n6886 = n5733 & ~n6885;
  assign n6887 = n1093 & n1178;
  assign n6888 = n975 & ~n1178;
  assign n6889 = ~n6887 & ~n6888;
  assign n6890 = ~n1195 & n6889;
  assign n6891 = ~pi243 & ~n6890;
  assign n6892 = pi184 & n1381;
  assign n6893 = n1380 & ~n1381;
  assign n6894 = ~n6892 & ~n6893;
  assign n6895 = ~pi129 & ~n6894;
  assign n6896 = ~n1381 & ~n1388;
  assign n6897 = ~pi202 & n6896;
  assign n6898 = pi184 & n6897;
  assign n6899 = ~n6892 & ~n6898;
  assign n6900 = pi129 & ~n6899;
  assign n6901 = ~n6895 & ~n6900;
  assign n6902 = n1087 & ~n6901;
  assign n6903 = pi184 & n1090;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = ~n1084 & n6904;
  assign n6906 = ~n6891 & n6905;
  assign n6907 = ~n5099 & ~n6906;
  assign n6908 = pi184 & n2070;
  assign n6909 = n5099 & n6908;
  assign n6910 = ~n6907 & ~n6909;
  assign n6911 = ~n6886 & n6910;
  assign n6912 = n5718 & ~n6911;
  assign n6913 = ~n5298 & n6912;
  assign n6914 = ~n6875 & ~n6913;
  assign n6915 = n3262 & ~n6914;
  assign n6916 = ~n3262 & n6912;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = ~pi247 & ~n6917;
  assign n6919 = pi184 & pi247;
  assign n6920 = ~n6918 & ~n6919;
  assign po229 = ~pi359 | ~n6920;
  assign n6922 = ~n4667 & n5542;
  assign n6923 = pi185 & ~n5400;
  assign n6924 = ~n5421 & ~n5422;
  assign n6925 = ~n6189 & n6844;
  assign n6926 = n6849 & ~n6925;
  assign n6927 = ~n6924 & ~n6926;
  assign n6928 = n6924 & n6926;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = n5400 & ~n6929;
  assign n6931 = ~n6923 & ~n6930;
  assign n6932 = ~n5529 & ~n6931;
  assign n6933 = pi185 & n5529;
  assign n6934 = ~n6932 & ~n6933;
  assign n6935 = ~n5394 & ~n6934;
  assign n6936 = ~n4334 & n5394;
  assign n6937 = ~n6935 & ~n6936;
  assign n6938 = ~n2070 & ~n6937;
  assign n6939 = pi185 & n2070;
  assign n6940 = ~n6938 & ~n6939;
  assign n6941 = ~n5544 & ~n6940;
  assign n6942 = ~n6922 & ~n6941;
  assign n6943 = n3262 & ~n6942;
  assign n6944 = ~n3262 & ~n6940;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = ~pi247 & ~n6945;
  assign n6947 = pi185 & pi247;
  assign n6948 = ~n6946 & ~n6947;
  assign po230 = ~pi359 | ~n6948;
  assign n6950 = ~n4591 & n5542;
  assign n6951 = n2648 & n3612;
  assign n6952 = n5393 & n6951;
  assign n6953 = pi186 & n5529;
  assign n6954 = ~n5394 & ~n6953;
  assign n6955 = pi186 & ~n5400;
  assign n6956 = ~n5505 & ~n5515;
  assign n6957 = n6699 & n6956;
  assign n6958 = ~n6699 & ~n6956;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = n5400 & ~n6959;
  assign n6961 = ~n6955 & ~n6960;
  assign n6962 = ~n5529 & ~n6961;
  assign n6963 = n6954 & ~n6962;
  assign n6964 = ~n6952 & ~n6963;
  assign n6965 = ~n2070 & n6964;
  assign n6966 = pi186 & n2070;
  assign n6967 = ~n6965 & ~n6966;
  assign n6968 = ~n5544 & ~n6967;
  assign n6969 = ~n6950 & ~n6968;
  assign n6970 = n3262 & ~n6969;
  assign n6971 = ~n3262 & ~n6967;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = ~pi247 & ~n6972;
  assign n6974 = pi186 & pi247;
  assign n6975 = ~n6973 & ~n6974;
  assign po231 = ~pi359 | ~n6975;
  assign n6977 = ~n4834 & n5542;
  assign n6978 = pi187 & ~n5400;
  assign n6979 = ~n5426 & ~n5498;
  assign n6980 = ~n5474 & n6596;
  assign n6981 = n6601 & ~n6980;
  assign n6982 = ~n6979 & ~n6981;
  assign n6983 = n6979 & n6981;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = n5400 & ~n6984;
  assign n6986 = ~n6978 & ~n6985;
  assign n6987 = ~n5529 & ~n6986;
  assign n6988 = pi187 & n5529;
  assign n6989 = ~n6987 & ~n6988;
  assign n6990 = ~n5394 & ~n6989;
  assign n6991 = ~n4208 & n5394;
  assign n6992 = ~n6990 & ~n6991;
  assign n6993 = ~n2070 & ~n6992;
  assign n6994 = pi187 & n2070;
  assign n6995 = ~n6993 & ~n6994;
  assign n6996 = ~n5544 & ~n6995;
  assign n6997 = ~n6977 & ~n6996;
  assign n6998 = n3262 & ~n6997;
  assign n6999 = ~n3262 & ~n6995;
  assign n7000 = ~n6998 & ~n6999;
  assign n7001 = ~pi247 & ~n7000;
  assign n7002 = pi187 & pi247;
  assign n7003 = ~n7001 & ~n7002;
  assign po232 = ~pi359 | ~n7003;
  assign n7005 = pi188 & n5005;
  assign n7006 = pi359 & n7005;
  assign n7007 = ~pi188 & pi190;
  assign n7008 = pi188 & ~pi190;
  assign n7009 = ~n7007 & ~n7008;
  assign n7010 = n2077 & ~n2109;
  assign n7011 = ~n2785 & ~n7010;
  assign n7012 = pi000 & n1529;
  assign n7013 = pi188 & n7012;
  assign n7014 = n2749 & n7013;
  assign n7015 = pi345 & ~n7014;
  assign n7016 = ~n3026 & n7015;
  assign n7017 = n7011 & n7016;
  assign n7018 = ~pi356 & n7017;
  assign n7019 = ~n7009 & n7018;
  assign n7020 = ~pi356 & n2978;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = ~pi213 & pi214;
  assign n7023 = pi213 & ~pi214;
  assign n7024 = ~n7022 & ~n7023;
  assign n7025 = ~pi356 & ~n7011;
  assign n7026 = ~n7024 & n7025;
  assign n7027 = n7021 & ~n7026;
  assign n7028 = pi188 & pi356;
  assign n7029 = n7027 & ~n7028;
  assign n7030 = n2633 & ~n7029;
  assign n7031 = ~n5003 & n7030;
  assign n7032 = pi188 & ~n5003;
  assign n7033 = ~n2633 & n7032;
  assign n7034 = ~n7031 & ~n7033;
  assign n7035 = pi188 & n5003;
  assign n7036 = n7034 & ~n7035;
  assign n7037 = ~n5005 & ~n7036;
  assign n7038 = pi359 & n7037;
  assign po233 = n7006 | n7038;
  assign n7040 = pi189 & n5005;
  assign n7041 = pi359 & n7040;
  assign n7042 = ~pi356 & n7011;
  assign n7043 = n7016 & n7042;
  assign n7044 = ~n2785 & n7043;
  assign n7045 = ~n2682 & n7044;
  assign n7046 = ~n7020 & ~n7045;
  assign n7047 = ~pi213 & ~pi214;
  assign n7048 = ~pi201 & ~n7047;
  assign n7049 = pi201 & n7047;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = n7025 & ~n7050;
  assign n7052 = n7046 & ~n7051;
  assign n7053 = pi189 & pi356;
  assign n7054 = n7052 & ~n7053;
  assign n7055 = n2633 & ~n7054;
  assign n7056 = ~n5003 & n7055;
  assign n7057 = pi189 & ~n5003;
  assign n7058 = ~n2633 & n7057;
  assign n7059 = ~n7056 & ~n7058;
  assign n7060 = pi189 & n5003;
  assign n7061 = n7059 & ~n7060;
  assign n7062 = ~n5005 & ~n7061;
  assign n7063 = pi359 & n7062;
  assign po234 = n7041 | n7063;
  assign n7065 = pi190 & n5003;
  assign n7066 = pi190 & pi356;
  assign n7067 = ~n2978 & ~n7011;
  assign n7068 = pi213 & ~pi356;
  assign n7069 = n7067 & n7068;
  assign n7070 = pi190 & n7016;
  assign n7071 = ~n2978 & ~n7070;
  assign n7072 = n7042 & n7071;
  assign n7073 = ~n7069 & ~n7072;
  assign n7074 = ~n7066 & n7073;
  assign n7075 = n2633 & ~n7074;
  assign n7076 = ~n5003 & n7075;
  assign n7077 = pi190 & ~n5003;
  assign n7078 = ~n2633 & n7077;
  assign n7079 = ~n7076 & ~n7078;
  assign n7080 = ~n7065 & n7079;
  assign n7081 = ~n5005 & ~n7080;
  assign n7082 = pi190 & n5005;
  assign n7083 = ~n7081 & ~n7082;
  assign po235 = ~pi359 | ~n7083;
  assign n7085 = n804 & n809;
  assign n7086 = ~n838 & ~n2136;
  assign n7087 = n804 & ~n7086;
  assign n7088 = n804 & n2238;
  assign n7089 = ~n7087 & ~n7088;
  assign n7090 = ~n7085 & n7089;
  assign n7091 = n787 & ~n7090;
  assign n7092 = n2634 & ~n2994;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = pi347 & ~n7093;
  assign n7095 = n2071 & n3009;
  assign n7096 = n782 & n2077;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = pi191 & n7097;
  assign n7099 = ~n5527 & n7096;
  assign n7100 = ~n7098 & ~n7099;
  assign n7101 = ~n2070 & ~n7100;
  assign n7102 = pi191 & n2070;
  assign n7103 = ~n7101 & ~n7102;
  assign n7104 = n7093 & ~n7103;
  assign n7105 = ~n7094 & ~n7104;
  assign n7106 = n782 & ~n7105;
  assign n7107 = ~n782 & ~n7103;
  assign n7108 = ~n7106 & ~n7107;
  assign n7109 = ~pi247 & ~n7108;
  assign n7110 = pi191 & pi247;
  assign n7111 = ~n7109 & ~n7110;
  assign po236 = pi359 & ~n7111;
  assign n7113 = ~pi192 & ~n785;
  assign n7114 = pi193 & n2635;
  assign n7115 = n1557 & n5393;
  assign n7116 = ~n2635 & ~n7115;
  assign n7117 = pi192 & n7116;
  assign n7118 = ~n7114 & ~n7117;
  assign n7119 = n785 & n7118;
  assign n7120 = ~n7113 & ~n7119;
  assign n7121 = pi302 & n823;
  assign n7122 = n883 & n7121;
  assign n7123 = n1559 & n7122;
  assign n7124 = n787 & n7123;
  assign n7125 = n782 & n7124;
  assign n7126 = ~n7120 & ~n7125;
  assign n7127 = ~n5007 & n7126;
  assign n7128 = ~pi356 & n2633;
  assign n7129 = n7126 & ~n7128;
  assign n7130 = ~n2978 & n7011;
  assign n7131 = pi300 & n792;
  assign n7132 = ~pi302 & n7131;
  assign n7133 = pi303 & n2787;
  assign n7134 = pi296 & n787;
  assign n7135 = n7133 & n7134;
  assign n7136 = n7132 & n7135;
  assign n7137 = ~pi297 & n1558;
  assign n7138 = n787 & n7137;
  assign n7139 = n2218 & n7138;
  assign n7140 = pi296 & n7139;
  assign n7141 = pi302 & n7140;
  assign n7142 = ~n7136 & ~n7141;
  assign n7143 = ~pi297 & n1559;
  assign n7144 = pi302 & n7137;
  assign n7145 = ~n7143 & ~n7144;
  assign n7146 = n787 & ~n7145;
  assign n7147 = pi296 & n7146;
  assign n7148 = n2218 & n7147;
  assign n7149 = n7142 & ~n7148;
  assign n7150 = ~pi192 & pi358;
  assign n7151 = n7149 & n7150;
  assign n7152 = ~n7115 & n7151;
  assign n7153 = pi355 & n7149;
  assign n7154 = ~n7152 & ~n7153;
  assign n7155 = ~n7016 & ~n7154;
  assign n7156 = n7126 & ~n7155;
  assign n7157 = n7130 & n7156;
  assign n7158 = n7126 & ~n7130;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = ~pi356 & ~n7159;
  assign n7161 = n2633 & n7160;
  assign n7162 = ~n7129 & ~n7161;
  assign n7163 = ~n5003 & ~n7162;
  assign n7164 = ~n5005 & n7163;
  assign n7165 = ~n7127 & ~n7164;
  assign po237 = pi359 & ~n7165;
  assign n7167 = n785 & n7115;
  assign n7168 = pi193 & ~n7167;
  assign n7169 = ~n7125 & ~n7168;
  assign n7170 = ~n7128 & n7169;
  assign n7171 = ~n7130 & n7169;
  assign n7172 = n7152 & ~n7153;
  assign n7173 = ~n7016 & n7172;
  assign n7174 = n7130 & ~n7173;
  assign n7175 = n7169 & n7174;
  assign n7176 = ~n7171 & ~n7175;
  assign n7177 = ~pi356 & ~n7176;
  assign n7178 = n2633 & n7177;
  assign n7179 = ~n7170 & ~n7178;
  assign n7180 = ~n5005 & ~n7179;
  assign n7181 = ~n5003 & n7180;
  assign n7182 = ~n5007 & n7169;
  assign n7183 = ~n7181 & ~n7182;
  assign po238 = pi359 & ~n7183;
  assign n7185 = ~pi099 & n1564;
  assign n7186 = n780 & n2071;
  assign n7187 = ~pi194 & ~n7186;
  assign n7188 = ~n7128 & ~n7187;
  assign n7189 = ~n7016 & n7130;
  assign n7190 = n2633 & ~n7189;
  assign n7191 = ~n7187 & n7190;
  assign n7192 = ~pi356 & n7191;
  assign n7193 = ~n7188 & ~n7192;
  assign n7194 = ~n5003 & ~n7193;
  assign n7195 = ~n5005 & n7194;
  assign n7196 = ~n5007 & ~n7187;
  assign n7197 = ~n7195 & ~n7196;
  assign n7198 = ~n7185 & ~n7197;
  assign po239 = ~pi359 | n7198;
  assign n7200 = pi195 & n7016;
  assign n7201 = ~n7173 & ~n7200;
  assign n7202 = n7011 & ~n7201;
  assign n7203 = ~n2978 & n7202;
  assign n7204 = pi195 & ~n7130;
  assign n7205 = ~n7203 & ~n7204;
  assign n7206 = n2633 & ~n7205;
  assign n7207 = ~pi356 & n7206;
  assign n7208 = pi195 & ~n7128;
  assign n7209 = ~n7207 & ~n7208;
  assign n7210 = ~n5003 & ~n7209;
  assign n7211 = ~n5005 & n7210;
  assign n7212 = pi195 & ~n5007;
  assign n7213 = ~n7211 & ~n7212;
  assign po240 = pi359 & ~n7213;
  assign n7215 = pi196 & n7016;
  assign n7216 = ~n7016 & n7153;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = n7130 & ~n7217;
  assign n7219 = pi196 & ~n7130;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = n7128 & ~n7220;
  assign n7222 = pi196 & ~n7128;
  assign n7223 = ~n7221 & ~n7222;
  assign n7224 = ~n5003 & ~n7223;
  assign n7225 = ~n5005 & n7224;
  assign n7226 = pi196 & ~n5007;
  assign n7227 = ~n7225 & ~n7226;
  assign po241 = pi359 & ~n7227;
  assign n7229 = pi303 & n2147;
  assign n7230 = ~n2223 & ~n2226;
  assign n7231 = n1536 & ~n7230;
  assign n7232 = n811 & n2196;
  assign n7233 = ~n2116 & ~n7232;
  assign n7234 = n811 & n2140;
  assign n7235 = n804 & n849;
  assign n7236 = n811 & ~n849;
  assign n7237 = ~n7235 & ~n7236;
  assign n7238 = n2192 & ~n7237;
  assign n7239 = pi303 & n2173;
  assign n7240 = ~n7238 & ~n7239;
  assign n7241 = ~n2991 & n7240;
  assign n7242 = ~n7234 & n7241;
  assign n7243 = n7233 & n7242;
  assign n7244 = pi303 & n2250;
  assign n7245 = n7243 & ~n7244;
  assign n7246 = n811 & n887;
  assign n7247 = n811 & n2252;
  assign n7248 = ~n7246 & ~n7247;
  assign n7249 = n7245 & n7248;
  assign n7250 = ~n7231 & n7249;
  assign n7251 = ~n811 & ~n7235;
  assign n7252 = n873 & ~n7251;
  assign n7253 = n7250 & ~n7252;
  assign n7254 = ~n2112 & ~n2154;
  assign n7255 = n7253 & n7254;
  assign n7256 = ~n7229 & n7255;
  assign n7257 = n787 & ~n7256;
  assign n7258 = n803 & ~n849;
  assign n7259 = n2343 & n7258;
  assign n7260 = ~n850 & n2360;
  assign n7261 = n1536 & n7260;
  assign n7262 = ~n7259 & ~n7261;
  assign n7263 = n1546 & n2343;
  assign n7264 = n849 & n7263;
  assign n7265 = n804 & n2364;
  assign n7266 = n804 & n2313;
  assign n7267 = ~n7265 & ~n7266;
  assign n7268 = n937 & n7267;
  assign n7269 = ~n2355 & ~n2376;
  assign n7270 = n811 & ~n7269;
  assign n7271 = n7268 & ~n7270;
  assign n7272 = ~n7264 & n7271;
  assign n7273 = n7262 & n7272;
  assign n7274 = pi301 & ~n7273;
  assign n7275 = ~n7257 & ~n7274;
  assign n7276 = pi296 & n2109;
  assign n7277 = n7275 & ~n7276;
  assign n7278 = ~n803 & ~n1546;
  assign n7279 = pi298 & ~n849;
  assign n7280 = ~n7278 & n7279;
  assign n7281 = n2343 & n7280;
  assign n7282 = pi298 & n811;
  assign n7283 = n7260 & n7282;
  assign n7284 = ~n7281 & ~n7283;
  assign n7285 = n788 & n2355;
  assign n7286 = n788 & n2376;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = n7267 & n7287;
  assign n7289 = n937 & n7288;
  assign n7290 = n7284 & n7289;
  assign n7291 = pi301 & ~n7290;
  assign n7292 = n2223 & n7282;
  assign n7293 = n811 & n2236;
  assign n7294 = pi298 & n7293;
  assign n7295 = ~n7292 & ~n7294;
  assign n7296 = n2226 & n7282;
  assign n7297 = pi298 & n2250;
  assign n7298 = ~n7296 & ~n7297;
  assign n7299 = n788 & n2196;
  assign n7300 = ~n2116 & ~n7299;
  assign n7301 = n811 & n2197;
  assign n7302 = pi298 & n7301;
  assign n7303 = n7300 & ~n7302;
  assign n7304 = n7298 & n7303;
  assign n7305 = ~n7234 & n7304;
  assign n7306 = pi298 & n2173;
  assign n7307 = ~n804 & ~n811;
  assign n7308 = n7279 & ~n7307;
  assign n7309 = n2192 & n7308;
  assign n7310 = ~n7306 & ~n7309;
  assign n7311 = n802 & n2136;
  assign n7312 = n7310 & ~n7311;
  assign n7313 = n7305 & n7312;
  assign n7314 = n7295 & n7313;
  assign n7315 = ~n7247 & n7314;
  assign n7316 = n811 & n7279;
  assign n7317 = ~pi298 & ~n849;
  assign n7318 = n804 & ~n7317;
  assign n7319 = ~n7316 & ~n7318;
  assign n7320 = n873 & ~n7319;
  assign n7321 = n7315 & ~n7320;
  assign n7322 = ~pi190 & ~n888;
  assign n7323 = n887 & n7322;
  assign n7324 = pi298 & n2147;
  assign n7325 = n7254 & ~n7324;
  assign n7326 = ~n7323 & n7325;
  assign n7327 = n7321 & n7326;
  assign n7328 = n787 & ~n7327;
  assign n7329 = ~n7291 & ~n7328;
  assign n7330 = pi291 & n2109;
  assign n7331 = n7329 & ~n7330;
  assign n7332 = n849 & ~n7307;
  assign n7333 = n2192 & n7332;
  assign n7334 = n849 & n873;
  assign n7335 = n811 & n7334;
  assign n7336 = ~n7333 & ~n7335;
  assign n7337 = n787 & ~n7336;
  assign n7338 = n803 & n849;
  assign n7339 = n2343 & n7338;
  assign n7340 = ~n2340 & ~n7339;
  assign n7341 = ~n7264 & n7340;
  assign n7342 = pi301 & ~n7341;
  assign n7343 = ~n7337 & ~n7342;
  assign n7344 = pi302 & n2147;
  assign n7345 = ~n7293 & ~n7301;
  assign n7346 = pi302 & ~n7345;
  assign n7347 = ~n7234 & ~n7247;
  assign n7348 = ~n2116 & n7347;
  assign n7349 = ~n7346 & n7348;
  assign n7350 = n2192 & ~n7307;
  assign n7351 = pi302 & ~n849;
  assign n7352 = n7350 & n7351;
  assign n7353 = pi302 & n811;
  assign n7354 = n2226 & n7353;
  assign n7355 = ~n2173 & ~n2250;
  assign n7356 = pi302 & ~n7355;
  assign n7357 = ~n7354 & ~n7356;
  assign n7358 = n2223 & n7353;
  assign n7359 = n7357 & ~n7358;
  assign n7360 = ~n7352 & n7359;
  assign n7361 = n7349 & n7360;
  assign n7362 = pi302 & ~n7307;
  assign n7363 = ~n7332 & ~n7362;
  assign n7364 = n873 & ~n7363;
  assign n7365 = n7361 & ~n7364;
  assign n7366 = ~n7344 & n7365;
  assign n7367 = n7254 & n7366;
  assign n7368 = n787 & ~n7367;
  assign n7369 = ~n935 & ~n7265;
  assign n7370 = ~n7278 & n7351;
  assign n7371 = n2343 & n7370;
  assign n7372 = n7260 & n7353;
  assign n7373 = ~n7371 & ~n7372;
  assign n7374 = ~n936 & n7373;
  assign n7375 = ~n2340 & n7374;
  assign n7376 = ~n7266 & n7375;
  assign n7377 = n7369 & n7376;
  assign n7378 = pi301 & ~n7377;
  assign n7379 = ~n7368 & ~n7378;
  assign n7380 = pi297 & n2109;
  assign n7381 = n7379 & ~n7380;
  assign n7382 = ~n7343 & n7381;
  assign n7383 = n7331 & n7382;
  assign n7384 = ~n7277 & n7383;
  assign n7385 = ~n7331 & ~n7381;
  assign n7386 = n7343 & ~n7385;
  assign n7387 = ~n7384 & ~n7386;
  assign n7388 = n7277 & n7331;
  assign n7389 = n7382 & n7388;
  assign n7390 = n7343 & n7385;
  assign n7391 = ~n7277 & n7390;
  assign n7392 = n7277 & n7390;
  assign n7393 = ~n7343 & ~n7381;
  assign n7394 = n7388 & n7393;
  assign n7395 = ~n7392 & ~n7394;
  assign n7396 = ~n7391 & n7395;
  assign n7397 = ~n7389 & n7396;
  assign n7398 = n7387 & n7397;
  assign n7399 = pi197 & n7398;
  assign n7400 = ~n1660 & n7277;
  assign n7401 = ~n1780 & ~n7277;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = n7386 & ~n7402;
  assign n7404 = ~n7399 & ~n7403;
  assign n7405 = pi187 & n7384;
  assign n7406 = pi354 & n7392;
  assign n7407 = pi174 & n7389;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = pi126 & n7391;
  assign n7410 = n7408 & ~n7409;
  assign n7411 = ~n7405 & n7410;
  assign n7412 = n7404 & n7411;
  assign n7413 = ~pi247 & ~n7412;
  assign n7414 = pi197 & pi247;
  assign po242 = n7413 | n7414;
  assign n7416 = pi198 & n7398;
  assign n7417 = ~n1857 & n7277;
  assign n7418 = ~n1709 & ~n7277;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = n7386 & ~n7419;
  assign n7421 = ~n7416 & ~n7420;
  assign n7422 = pi183 & n7384;
  assign n7423 = pi353 & n7392;
  assign n7424 = pi144 & n7389;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = pi139 & n7391;
  assign n7427 = n7425 & ~n7426;
  assign n7428 = ~n7422 & n7427;
  assign n7429 = n7421 & n7428;
  assign n7430 = ~pi247 & ~n7429;
  assign n7431 = pi198 & pi247;
  assign po243 = n7430 | n7431;
  assign n7433 = ~n1527 & ~n2202;
  assign n7434 = ~n2289 & n7433;
  assign n7435 = n804 & ~n7434;
  assign n7436 = ~n2243 & ~n2288;
  assign n7437 = ~n2274 & n7436;
  assign n7438 = n804 & ~n7437;
  assign n7439 = ~n7435 & ~n7438;
  assign n7440 = n787 & ~n7439;
  assign n7441 = pi350 & n7440;
  assign n7442 = pi228 & ~n7440;
  assign n7443 = ~n7441 & ~n7442;
  assign n7444 = ~pi199 & n7443;
  assign n7445 = pi199 & ~n7443;
  assign n7446 = ~n7444 & ~n7445;
  assign n7447 = pi212 & ~n7443;
  assign n7448 = ~pi212 & n7443;
  assign n7449 = pi200 & ~n7443;
  assign n7450 = ~n7448 & n7449;
  assign n7451 = ~n7447 & ~n7450;
  assign n7452 = ~pi200 & n7443;
  assign n7453 = ~n7448 & ~n7452;
  assign n7454 = pi347 & n7440;
  assign n7455 = ~n7442 & ~n7454;
  assign n7456 = pi211 & ~n7455;
  assign n7457 = ~pi211 & n7455;
  assign n7458 = pi353 & n7440;
  assign n7459 = ~n7442 & ~n7458;
  assign n7460 = pi210 & ~n7459;
  assign n7461 = ~n7457 & n7460;
  assign n7462 = ~n7456 & ~n7461;
  assign n7463 = n7453 & ~n7462;
  assign n7464 = n7451 & ~n7463;
  assign n7465 = pi348 & n7440;
  assign n7466 = ~n7442 & ~n7465;
  assign n7467 = ~pi208 & n7466;
  assign n7468 = pi352 & n7440;
  assign n7469 = ~n7442 & ~n7468;
  assign n7470 = ~pi209 & n7469;
  assign n7471 = ~n7467 & ~n7470;
  assign n7472 = pi351 & n7440;
  assign n7473 = ~n7442 & ~n7472;
  assign n7474 = ~pi207 & n7473;
  assign n7475 = n7471 & ~n7474;
  assign n7476 = ~pi228 & ~n7440;
  assign n7477 = pi354 & n7440;
  assign n7478 = ~n7476 & ~n7477;
  assign n7479 = pi220 & ~n7478;
  assign n7480 = pi349 & n7440;
  assign n7481 = ~n7442 & ~n7480;
  assign n7482 = ~pi206 & n7481;
  assign n7483 = n7479 & ~n7482;
  assign n7484 = n7475 & n7483;
  assign n7485 = pi206 & ~n7481;
  assign n7486 = ~n7474 & n7485;
  assign n7487 = pi207 & ~n7473;
  assign n7488 = ~n7486 & ~n7487;
  assign n7489 = n7471 & ~n7488;
  assign n7490 = ~n7484 & ~n7489;
  assign n7491 = pi209 & ~n7469;
  assign n7492 = pi208 & ~n7466;
  assign n7493 = ~n7470 & n7492;
  assign n7494 = ~n7491 & ~n7493;
  assign n7495 = n7490 & n7494;
  assign n7496 = ~pi210 & n7459;
  assign n7497 = ~n7457 & ~n7496;
  assign n7498 = n7453 & n7497;
  assign n7499 = ~n7495 & n7498;
  assign n7500 = n7464 & ~n7499;
  assign n7501 = ~n7446 & n7500;
  assign n7502 = n7446 & ~n7500;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = ~pi296 & ~pi303;
  assign n7505 = n2792 & n7504;
  assign n7506 = n3322 & n7505;
  assign n7507 = n787 & n7506;
  assign n7508 = n849 & n7507;
  assign n7509 = ~pi196 & pi230;
  assign n7510 = ~pi195 & n7509;
  assign n7511 = n2647 & n7510;
  assign n7512 = ~n7508 & n7511;
  assign n7513 = ~n3011 & n7512;
  assign n7514 = n7503 & n7513;
  assign n7515 = pi199 & ~n7513;
  assign n7516 = ~n7514 & ~n7515;
  assign n7517 = n2071 & ~n7516;
  assign n7518 = pi199 & ~n2071;
  assign n7519 = ~n7517 & ~n7518;
  assign n7520 = n2070 & ~n7519;
  assign n7521 = ~n7476 & n7503;
  assign n7522 = pi199 & ~n2653;
  assign n7523 = ~n4319 & ~n7522;
  assign n7524 = n3646 & ~n7523;
  assign n7525 = ~n4362 & ~n7524;
  assign n7526 = ~n2650 & ~n7525;
  assign n7527 = ~n4365 & ~n7526;
  assign n7528 = n2647 & ~n7527;
  assign n7529 = ~n4368 & ~n7528;
  assign n7530 = n2633 & ~n7529;
  assign n7531 = pi199 & ~n2633;
  assign n7532 = ~n7530 & ~n7531;
  assign n7533 = n788 & ~n2994;
  assign n7534 = pi301 & n7533;
  assign n7535 = n811 & n2215;
  assign n7536 = ~n838 & ~n2133;
  assign n7537 = n788 & ~n7536;
  assign n7538 = n788 & n2192;
  assign n7539 = ~n7537 & ~n7538;
  assign n7540 = n811 & n2119;
  assign n7541 = n788 & n809;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = n811 & n2226;
  assign n7544 = n7542 & ~n7543;
  assign n7545 = ~n2136 & ~n2193;
  assign n7546 = n788 & ~n7545;
  assign n7547 = n7544 & ~n7546;
  assign n7548 = ~n7234 & n7547;
  assign n7549 = n7539 & n7548;
  assign n7550 = ~n2182 & ~n2238;
  assign n7551 = n788 & ~n7550;
  assign n7552 = n7549 & ~n7551;
  assign n7553 = n788 & n2280;
  assign n7554 = n811 & n2241;
  assign n7555 = ~n7553 & ~n7554;
  assign n7556 = n7552 & n7555;
  assign n7557 = ~n2289 & n7436;
  assign n7558 = ~n2274 & n7557;
  assign n7559 = n811 & ~n7558;
  assign n7560 = n7556 & ~n7559;
  assign n7561 = n811 & ~n7433;
  assign n7562 = n803 & n2636;
  assign n7563 = n826 & n7562;
  assign n7564 = ~n7561 & ~n7563;
  assign n7565 = n7560 & n7564;
  assign n7566 = ~n7535 & n7565;
  assign n7567 = n787 & ~n7566;
  assign n7568 = ~n2109 & ~n2796;
  assign n7569 = n2785 & ~n7568;
  assign n7570 = ~n2077 & ~n7569;
  assign n7571 = ~n7567 & n7570;
  assign n7572 = ~n7534 & n7571;
  assign n7573 = n7532 & n7572;
  assign n7574 = ~n7503 & ~n7572;
  assign n7575 = ~n7573 & ~n7574;
  assign n7576 = n7476 & n7575;
  assign n7577 = ~n7521 & ~n7576;
  assign n7578 = n2071 & n7577;
  assign n7579 = ~n2071 & n7532;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = ~n2070 & n7580;
  assign n7582 = ~n7520 & ~n7581;
  assign n7583 = ~pi247 & ~n7582;
  assign n7584 = pi199 & pi247;
  assign n7585 = ~n7583 & ~n7584;
  assign po244 = pi359 & ~n7585;
  assign n7587 = ~n7449 & ~n7452;
  assign n7588 = ~n7494 & n7497;
  assign n7589 = n7462 & ~n7588;
  assign n7590 = ~n7474 & ~n7482;
  assign n7591 = n7479 & n7590;
  assign n7592 = n7488 & ~n7591;
  assign n7593 = n7471 & n7497;
  assign n7594 = ~n7592 & n7593;
  assign n7595 = n7589 & ~n7594;
  assign n7596 = ~n7587 & n7595;
  assign n7597 = n7587 & ~n7595;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = n7513 & n7598;
  assign n7600 = pi200 & ~n7513;
  assign n7601 = ~n7599 & ~n7600;
  assign n7602 = n2071 & ~n7601;
  assign n7603 = pi200 & ~n2071;
  assign n7604 = ~n7602 & ~n7603;
  assign n7605 = n2070 & ~n7604;
  assign n7606 = ~n7476 & n7598;
  assign n7607 = pi200 & ~n2653;
  assign n7608 = ~n4256 & ~n7607;
  assign n7609 = n3646 & ~n7608;
  assign n7610 = ~n4298 & ~n7609;
  assign n7611 = ~n2650 & ~n7610;
  assign n7612 = ~n4301 & ~n7611;
  assign n7613 = n2647 & ~n7612;
  assign n7614 = ~n4304 & ~n7613;
  assign n7615 = n2633 & ~n7614;
  assign n7616 = pi200 & ~n2633;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = n7572 & n7617;
  assign n7619 = ~n7572 & ~n7598;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = n7476 & n7620;
  assign n7622 = ~n7606 & ~n7621;
  assign n7623 = n2071 & n7622;
  assign n7624 = ~n2071 & n7617;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n2070 & n7625;
  assign n7627 = ~n7605 & ~n7626;
  assign n7628 = ~pi247 & ~n7627;
  assign n7629 = pi200 & pi247;
  assign n7630 = ~n7628 & ~n7629;
  assign po245 = pi359 & ~n7630;
  assign n7632 = ~pi201 & ~n7128;
  assign n7633 = pi189 & n2978;
  assign n7634 = ~pi201 & ~n2978;
  assign n7635 = ~n7633 & ~n7634;
  assign n7636 = n7128 & ~n7635;
  assign n7637 = ~n7632 & ~n7636;
  assign n7638 = ~n5003 & ~n7637;
  assign n7639 = ~n5005 & n7638;
  assign n7640 = ~pi201 & ~n5007;
  assign n7641 = ~n7639 & ~n7640;
  assign po246 = pi359 & ~n7641;
  assign n7643 = pi202 & pi247;
  assign n7644 = pi202 & n7398;
  assign n7645 = ~n1822 & n7277;
  assign n7646 = ~n1744 & ~n7277;
  assign n7647 = ~n7645 & ~n7646;
  assign n7648 = n7386 & ~n7647;
  assign n7649 = ~n7644 & ~n7648;
  assign n7650 = pi186 & n7384;
  assign n7651 = pi348 & n7392;
  assign n7652 = pi173 & n7389;
  assign n7653 = ~n7651 & ~n7652;
  assign n7654 = pi138 & n7391;
  assign n7655 = n7653 & ~n7654;
  assign n7656 = ~n7650 & n7655;
  assign n7657 = n7649 & n7656;
  assign n7658 = ~pi247 & ~n7657;
  assign po247 = n7643 | n7658;
  assign n7660 = ~pi203 & n7443;
  assign n7661 = pi203 & ~n7443;
  assign n7662 = ~n7660 & ~n7661;
  assign n7663 = ~pi221 & n7443;
  assign n7664 = ~n7444 & ~n7663;
  assign n7665 = ~n7595 & n7664;
  assign n7666 = n7453 & n7665;
  assign n7667 = pi221 & ~n7443;
  assign n7668 = n7445 & ~n7663;
  assign n7669 = ~n7667 & ~n7668;
  assign n7670 = ~n7451 & n7664;
  assign n7671 = n7669 & ~n7670;
  assign n7672 = ~n7666 & n7671;
  assign n7673 = ~n7662 & n7672;
  assign n7674 = n7662 & ~n7672;
  assign n7675 = ~n7673 & ~n7674;
  assign n7676 = n7513 & n7675;
  assign n7677 = pi203 & ~n7513;
  assign n7678 = ~n7676 & ~n7677;
  assign n7679 = n2071 & ~n7678;
  assign n7680 = pi203 & ~n2071;
  assign n7681 = ~n7679 & ~n7680;
  assign n7682 = n2070 & ~n7681;
  assign n7683 = ~n7476 & n7675;
  assign n7684 = pi203 & ~n2653;
  assign n7685 = ~n3597 & ~n7684;
  assign n7686 = n3646 & ~n7685;
  assign n7687 = ~n3648 & ~n7686;
  assign n7688 = ~n2650 & ~n7687;
  assign n7689 = ~n3651 & ~n7688;
  assign n7690 = n2647 & ~n7689;
  assign n7691 = ~n3654 & ~n7690;
  assign n7692 = n2633 & ~n7691;
  assign n7693 = pi203 & ~n2633;
  assign n7694 = ~n7692 & ~n7693;
  assign n7695 = n7572 & n7694;
  assign n7696 = ~n7572 & ~n7675;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = n7476 & n7697;
  assign n7699 = ~n7683 & ~n7698;
  assign n7700 = n2071 & n7699;
  assign n7701 = ~n2071 & n7694;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = ~n2070 & n7702;
  assign n7704 = ~n7682 & ~n7703;
  assign n7705 = ~pi247 & ~n7704;
  assign n7706 = pi203 & pi247;
  assign n7707 = ~n7705 & ~n7706;
  assign po248 = pi359 & ~n7707;
  assign n7709 = pi204 & ~n7443;
  assign n7710 = ~pi204 & n7443;
  assign n7711 = ~n7709 & ~n7710;
  assign n7712 = ~n7452 & ~n7457;
  assign n7713 = ~n7470 & ~n7496;
  assign n7714 = n7712 & n7713;
  assign n7715 = ~n7660 & ~n7663;
  assign n7716 = ~n7444 & ~n7448;
  assign n7717 = ~n7467 & n7487;
  assign n7718 = ~n7492 & ~n7717;
  assign n7719 = ~n7483 & ~n7485;
  assign n7720 = ~n7467 & ~n7474;
  assign n7721 = ~n7719 & n7720;
  assign n7722 = n7718 & ~n7721;
  assign n7723 = n7716 & ~n7722;
  assign n7724 = n7715 & n7723;
  assign n7725 = n7714 & n7724;
  assign n7726 = ~n7660 & n7667;
  assign n7727 = ~n7661 & ~n7726;
  assign n7728 = ~n7444 & n7447;
  assign n7729 = ~n7445 & ~n7728;
  assign n7730 = ~n7452 & n7456;
  assign n7731 = ~n7449 & ~n7730;
  assign n7732 = n7491 & ~n7496;
  assign n7733 = ~n7460 & ~n7732;
  assign n7734 = n7712 & ~n7733;
  assign n7735 = n7731 & ~n7734;
  assign n7736 = n7716 & ~n7735;
  assign n7737 = n7729 & ~n7736;
  assign n7738 = n7715 & ~n7737;
  assign n7739 = n7727 & ~n7738;
  assign n7740 = ~n7725 & n7739;
  assign n7741 = ~n7711 & n7740;
  assign n7742 = n7711 & ~n7740;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = n7513 & n7743;
  assign n7745 = pi204 & ~n7513;
  assign n7746 = ~n7744 & ~n7745;
  assign n7747 = n2071 & ~n7746;
  assign n7748 = pi204 & ~n2071;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = n2070 & ~n7749;
  assign n7751 = ~n7476 & n7743;
  assign n7752 = pi204 & ~n2653;
  assign n7753 = ~n3669 & ~n7752;
  assign n7754 = n3646 & ~n7753;
  assign n7755 = ~n3718 & ~n7754;
  assign n7756 = ~n2650 & ~n7755;
  assign n7757 = ~n3721 & ~n7756;
  assign n7758 = n2647 & ~n7757;
  assign n7759 = ~n3724 & ~n7758;
  assign n7760 = n2633 & ~n7759;
  assign n7761 = pi204 & ~n2633;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = n7572 & n7762;
  assign n7764 = ~n7572 & ~n7743;
  assign n7765 = ~n7763 & ~n7764;
  assign n7766 = n7476 & n7765;
  assign n7767 = ~n7751 & ~n7766;
  assign n7768 = n2071 & n7767;
  assign n7769 = ~n2071 & n7762;
  assign n7770 = ~n7768 & ~n7769;
  assign n7771 = ~n2070 & n7770;
  assign n7772 = ~n7750 & ~n7771;
  assign n7773 = ~pi247 & ~n7772;
  assign n7774 = pi204 & pi247;
  assign n7775 = ~n7773 & ~n7774;
  assign po249 = pi359 & ~n7775;
  assign n7777 = pi205 & pi247;
  assign n7778 = pi205 & ~n7443;
  assign n7779 = ~pi205 & n7443;
  assign n7780 = ~n7778 & ~n7779;
  assign n7781 = ~n7660 & ~n7710;
  assign n7782 = ~n7495 & n7781;
  assign n7783 = n7498 & n7782;
  assign n7784 = n7664 & n7783;
  assign n7785 = n7661 & ~n7710;
  assign n7786 = ~n7709 & ~n7785;
  assign n7787 = ~n7464 & n7664;
  assign n7788 = n7669 & ~n7787;
  assign n7789 = n7781 & ~n7788;
  assign n7790 = n7786 & ~n7789;
  assign n7791 = ~n7784 & n7790;
  assign n7792 = ~n7780 & n7791;
  assign n7793 = n7780 & ~n7791;
  assign n7794 = ~n7792 & ~n7793;
  assign n7795 = n7513 & n7794;
  assign n7796 = pi205 & ~n7513;
  assign n7797 = ~n7795 & ~n7796;
  assign n7798 = n2071 & ~n7797;
  assign n7799 = pi205 & ~n2071;
  assign n7800 = ~n7798 & ~n7799;
  assign n7801 = n2070 & n7800;
  assign n7802 = ~pi247 & ~n7801;
  assign n7803 = ~n7777 & ~n7802;
  assign n7804 = pi205 & ~n2653;
  assign n7805 = ~n3739 & ~n7804;
  assign n7806 = n3646 & ~n7805;
  assign n7807 = ~n3788 & ~n7806;
  assign n7808 = ~n2650 & ~n7807;
  assign n7809 = ~n3791 & ~n7808;
  assign n7810 = n2647 & ~n7809;
  assign n7811 = ~n3794 & ~n7810;
  assign n7812 = n2633 & ~n7811;
  assign n7813 = pi205 & ~n2633;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = ~n2071 & n7814;
  assign n7816 = ~n7476 & n7794;
  assign n7817 = n7572 & n7814;
  assign n7818 = ~n7572 & ~n7794;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = n7476 & n7819;
  assign n7821 = ~n7816 & ~n7820;
  assign n7822 = n2071 & n7821;
  assign n7823 = ~n7815 & ~n7822;
  assign n7824 = ~pi247 & ~n2070;
  assign n7825 = ~n7823 & n7824;
  assign n7826 = ~n7803 & ~n7825;
  assign po250 = pi359 & n7826;
  assign n7828 = ~n7482 & ~n7485;
  assign n7829 = n7479 & n7828;
  assign n7830 = ~n7479 & ~n7828;
  assign n7831 = ~n7829 & ~n7830;
  assign n7832 = n7513 & n7831;
  assign n7833 = pi206 & ~n7513;
  assign n7834 = ~n7832 & ~n7833;
  assign n7835 = n2071 & ~n7834;
  assign n7836 = pi206 & ~n2071;
  assign n7837 = ~n7835 & ~n7836;
  assign n7838 = n2070 & ~n7837;
  assign n7839 = ~n7476 & n7831;
  assign n7840 = pi206 & ~n2653;
  assign n7841 = ~n3015 & ~n7840;
  assign n7842 = ~n3027 & n7841;
  assign n7843 = n3012 & ~n7842;
  assign n7844 = ~n3030 & ~n7843;
  assign n7845 = ~n2650 & ~n7844;
  assign n7846 = ~n3034 & ~n7845;
  assign n7847 = n2647 & ~n7846;
  assign n7848 = ~n3037 & ~n7847;
  assign n7849 = n2633 & ~n7848;
  assign n7850 = pi206 & ~n2633;
  assign n7851 = ~n7849 & ~n7850;
  assign n7852 = n7572 & n7851;
  assign n7853 = ~n7572 & ~n7831;
  assign n7854 = ~n7852 & ~n7853;
  assign n7855 = n7476 & n7854;
  assign n7856 = ~n7839 & ~n7855;
  assign n7857 = n2071 & n7856;
  assign n7858 = ~n2071 & n7851;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n2070 & n7859;
  assign n7861 = ~n7838 & ~n7860;
  assign n7862 = ~pi247 & ~n7861;
  assign n7863 = pi206 & pi247;
  assign n7864 = ~n7862 & ~n7863;
  assign po251 = pi359 & ~n7864;
  assign n7866 = ~n7474 & ~n7487;
  assign n7867 = n7719 & ~n7866;
  assign n7868 = ~n7719 & n7866;
  assign n7869 = ~n7867 & ~n7868;
  assign n7870 = n7513 & n7869;
  assign n7871 = pi207 & ~n7513;
  assign n7872 = ~n7870 & ~n7871;
  assign n7873 = n2071 & ~n7872;
  assign n7874 = pi207 & ~n2071;
  assign n7875 = ~n7873 & ~n7874;
  assign n7876 = n2070 & ~n7875;
  assign n7877 = ~n7476 & n7869;
  assign n7878 = pi207 & ~n2653;
  assign n7879 = ~n3093 & ~n7878;
  assign n7880 = ~n3027 & n7879;
  assign n7881 = n3012 & ~n7880;
  assign n7882 = ~n3096 & ~n7881;
  assign n7883 = ~n2650 & ~n7882;
  assign n7884 = ~n3100 & ~n7883;
  assign n7885 = n2647 & ~n7884;
  assign n7886 = ~n3103 & ~n7885;
  assign n7887 = n2633 & ~n7886;
  assign n7888 = pi207 & ~n2633;
  assign n7889 = ~n7887 & ~n7888;
  assign n7890 = n7572 & n7889;
  assign n7891 = ~n7572 & ~n7869;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = n7476 & n7892;
  assign n7894 = ~n7877 & ~n7893;
  assign n7895 = n2071 & n7894;
  assign n7896 = ~n2071 & n7889;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = ~n2070 & n7897;
  assign n7899 = ~n7876 & ~n7898;
  assign n7900 = ~pi247 & ~n7899;
  assign n7901 = pi207 & pi247;
  assign n7902 = ~n7900 & ~n7901;
  assign po252 = pi359 & ~n7902;
  assign n7904 = ~n7467 & ~n7492;
  assign n7905 = ~n7592 & n7904;
  assign n7906 = n7592 & ~n7904;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = n7513 & n7907;
  assign n7909 = pi208 & ~n7513;
  assign n7910 = ~n7908 & ~n7909;
  assign n7911 = n2071 & ~n7910;
  assign n7912 = pi208 & ~n2071;
  assign n7913 = ~n7911 & ~n7912;
  assign n7914 = n2070 & ~n7913;
  assign n7915 = ~n7476 & n7907;
  assign n7916 = pi208 & ~n2653;
  assign n7917 = ~n4064 & ~n7916;
  assign n7918 = n3646 & ~n7917;
  assign n7919 = ~n4106 & ~n7918;
  assign n7920 = ~n2650 & ~n7919;
  assign n7921 = ~n4109 & ~n7920;
  assign n7922 = n2647 & ~n7921;
  assign n7923 = ~n4112 & ~n7922;
  assign n7924 = n2633 & ~n7923;
  assign n7925 = pi208 & ~n2633;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = n7572 & n7926;
  assign n7928 = ~n7572 & ~n7907;
  assign n7929 = ~n7927 & ~n7928;
  assign n7930 = n7476 & n7929;
  assign n7931 = ~n7915 & ~n7930;
  assign n7932 = n2071 & n7931;
  assign n7933 = ~n2071 & n7926;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = ~n2070 & n7934;
  assign n7936 = ~n7914 & ~n7935;
  assign n7937 = ~pi247 & ~n7936;
  assign n7938 = pi208 & pi247;
  assign n7939 = ~n7937 & ~n7938;
  assign po253 = pi359 & ~n7939;
  assign n7941 = ~n7470 & ~n7491;
  assign n7942 = ~n7722 & n7941;
  assign n7943 = n7722 & ~n7941;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = n7513 & n7944;
  assign n7946 = pi209 & ~n7513;
  assign n7947 = ~n7945 & ~n7946;
  assign n7948 = n2071 & ~n7947;
  assign n7949 = pi209 & ~n2071;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = n2070 & ~n7950;
  assign n7952 = ~n7476 & n7944;
  assign n7953 = pi209 & ~n2653;
  assign n7954 = ~n3941 & ~n7953;
  assign n7955 = n3646 & ~n7954;
  assign n7956 = ~n3982 & ~n7955;
  assign n7957 = ~n2650 & ~n7956;
  assign n7958 = ~n3985 & ~n7957;
  assign n7959 = n2647 & ~n7958;
  assign n7960 = ~n3988 & ~n7959;
  assign n7961 = n2633 & ~n7960;
  assign n7962 = pi209 & ~n2633;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = n7572 & n7963;
  assign n7965 = ~n7572 & ~n7944;
  assign n7966 = ~n7964 & ~n7965;
  assign n7967 = n7476 & n7966;
  assign n7968 = ~n7952 & ~n7967;
  assign n7969 = n2071 & n7968;
  assign n7970 = ~n2071 & n7963;
  assign n7971 = ~n7969 & ~n7970;
  assign n7972 = ~n2070 & n7971;
  assign n7973 = ~n7951 & ~n7972;
  assign n7974 = ~pi247 & ~n7973;
  assign n7975 = pi209 & pi247;
  assign n7976 = ~n7974 & ~n7975;
  assign po254 = pi359 & ~n7976;
  assign n7978 = ~n7460 & ~n7496;
  assign n7979 = n7495 & ~n7978;
  assign n7980 = ~n7495 & n7978;
  assign n7981 = ~n7979 & ~n7980;
  assign n7982 = n7513 & n7981;
  assign n7983 = pi210 & ~n7513;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = n2071 & ~n7984;
  assign n7986 = pi210 & ~n2071;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = n2070 & ~n7987;
  assign n7989 = ~n7476 & n7981;
  assign n7990 = pi210 & ~n2653;
  assign n7991 = ~n3161 & ~n7990;
  assign n7992 = ~n3027 & n7991;
  assign n7993 = n3012 & ~n7992;
  assign n7994 = ~n3164 & ~n7993;
  assign n7995 = ~n2650 & ~n7994;
  assign n7996 = ~n3168 & ~n7995;
  assign n7997 = n2647 & ~n7996;
  assign n7998 = ~n3171 & ~n7997;
  assign n7999 = n2633 & ~n7998;
  assign n8000 = pi210 & ~n2633;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = n7572 & n8001;
  assign n8003 = ~n7572 & ~n7981;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = n7476 & n8004;
  assign n8006 = ~n7989 & ~n8005;
  assign n8007 = n2071 & n8006;
  assign n8008 = ~n2071 & n8001;
  assign n8009 = ~n8007 & ~n8008;
  assign n8010 = ~n2070 & n8009;
  assign n8011 = ~n7988 & ~n8010;
  assign n8012 = ~pi247 & ~n8011;
  assign n8013 = pi210 & pi247;
  assign n8014 = ~n8012 & ~n8013;
  assign po255 = pi359 & ~n8014;
  assign n8016 = ~n7456 & ~n7457;
  assign n8017 = n7713 & ~n7722;
  assign n8018 = n7733 & ~n8017;
  assign n8019 = ~n8016 & n8018;
  assign n8020 = n8016 & ~n8018;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = n7513 & n8021;
  assign n8023 = pi211 & ~n7513;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = n2071 & ~n8024;
  assign n8026 = pi211 & ~n2071;
  assign n8027 = ~n8025 & ~n8026;
  assign n8028 = n2070 & ~n8027;
  assign n8029 = ~n7476 & n8021;
  assign n8030 = pi211 & ~n2653;
  assign n8031 = ~n3230 & ~n8030;
  assign n8032 = ~n3027 & n8031;
  assign n8033 = n3012 & ~n8032;
  assign n8034 = ~n3233 & ~n8033;
  assign n8035 = ~n2650 & ~n8034;
  assign n8036 = ~n3237 & ~n8035;
  assign n8037 = n2647 & ~n8036;
  assign n8038 = ~n3240 & ~n8037;
  assign n8039 = n2633 & ~n8038;
  assign n8040 = pi211 & ~n2633;
  assign n8041 = ~n8039 & ~n8040;
  assign n8042 = n7572 & n8041;
  assign n8043 = ~n7572 & ~n8021;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = n7476 & n8044;
  assign n8046 = ~n8029 & ~n8045;
  assign n8047 = n2071 & n8046;
  assign n8048 = ~n2071 & n8041;
  assign n8049 = ~n8047 & ~n8048;
  assign n8050 = ~n2070 & n8049;
  assign n8051 = ~n8028 & ~n8050;
  assign n8052 = ~pi247 & ~n8051;
  assign n8053 = pi211 & pi247;
  assign n8054 = ~n8052 & ~n8053;
  assign po256 = pi359 & ~n8054;
  assign n8056 = ~n7447 & ~n7448;
  assign n8057 = n7714 & ~n7722;
  assign n8058 = n7735 & ~n8057;
  assign n8059 = ~n8056 & n8058;
  assign n8060 = n8056 & ~n8058;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = n7513 & n8061;
  assign n8063 = pi212 & ~n7513;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = n2071 & ~n8064;
  assign n8066 = pi212 & ~n2071;
  assign n8067 = ~n8065 & ~n8066;
  assign n8068 = n2070 & ~n8067;
  assign n8069 = ~n7476 & n8061;
  assign n8070 = pi212 & ~n2653;
  assign n8071 = ~n4193 & ~n8070;
  assign n8072 = n3646 & ~n8071;
  assign n8073 = ~n4235 & ~n8072;
  assign n8074 = ~n2650 & ~n8073;
  assign n8075 = ~n4238 & ~n8074;
  assign n8076 = n2647 & ~n8075;
  assign n8077 = ~n4241 & ~n8076;
  assign n8078 = n2633 & ~n8077;
  assign n8079 = pi212 & ~n2633;
  assign n8080 = ~n8078 & ~n8079;
  assign n8081 = n7572 & n8080;
  assign n8082 = ~n7572 & ~n8061;
  assign n8083 = ~n8081 & ~n8082;
  assign n8084 = n7476 & n8083;
  assign n8085 = ~n8069 & ~n8084;
  assign n8086 = n2071 & n8085;
  assign n8087 = ~n2071 & n8080;
  assign n8088 = ~n8086 & ~n8087;
  assign n8089 = ~n2070 & n8088;
  assign n8090 = ~n8068 & ~n8089;
  assign n8091 = ~pi247 & ~n8090;
  assign n8092 = pi212 & pi247;
  assign n8093 = ~n8091 & ~n8092;
  assign po257 = pi359 & ~n8093;
  assign n8095 = ~pi213 & ~n7128;
  assign n8096 = pi190 & n2978;
  assign n8097 = ~pi213 & ~n2978;
  assign n8098 = ~n8096 & ~n8097;
  assign n8099 = n7128 & ~n8098;
  assign n8100 = ~n8095 & ~n8099;
  assign n8101 = ~n5003 & ~n8100;
  assign n8102 = ~n5005 & n8101;
  assign n8103 = ~pi213 & ~n5007;
  assign n8104 = ~n8102 & ~n8103;
  assign po258 = pi359 & ~n8104;
  assign n8106 = ~pi214 & ~n7128;
  assign n8107 = pi188 & n2978;
  assign n8108 = ~pi214 & ~n2978;
  assign n8109 = ~n8107 & ~n8108;
  assign n8110 = n7128 & ~n8109;
  assign n8111 = ~n8106 & ~n8110;
  assign n8112 = ~n5003 & ~n8111;
  assign n8113 = ~n5005 & n8112;
  assign n8114 = ~pi214 & ~n5007;
  assign n8115 = ~n8113 & ~n8114;
  assign po259 = pi359 & ~n8115;
  assign n8117 = pi215 & n7398;
  assign n8118 = ~n1643 & n7277;
  assign n8119 = ~n1764 & ~n7277;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = n7386 & ~n8120;
  assign n8122 = ~n8117 & ~n8121;
  assign n8123 = pi182 & n7384;
  assign n8124 = pi351 & n7392;
  assign n8125 = pi172 & n7389;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = pi141 & n7391;
  assign n8128 = n8126 & ~n8127;
  assign n8129 = ~n8123 & n8128;
  assign n8130 = n8122 & n8129;
  assign n8131 = ~pi247 & ~n8130;
  assign n8132 = pi215 & pi247;
  assign po260 = n8131 | n8132;
  assign n8134 = pi216 & n7398;
  assign n8135 = ~n1838 & n7277;
  assign n8136 = ~n1727 & ~n7277;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = n7386 & ~n8137;
  assign n8139 = ~n8134 & ~n8138;
  assign n8140 = pi177 & n7384;
  assign n8141 = pi352 & n7392;
  assign n8142 = pi146 & n7389;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = pi143 & n7391;
  assign n8145 = n8143 & ~n8144;
  assign n8146 = ~n8140 & n8145;
  assign n8147 = n8139 & n8146;
  assign n8148 = ~pi247 & ~n8147;
  assign n8149 = pi216 & pi247;
  assign po261 = n8148 | n8149;
  assign n8151 = pi217 & n7398;
  assign n8152 = ~n2006 & n7277;
  assign n8153 = ~n1693 & ~n7277;
  assign n8154 = ~n8152 & ~n8153;
  assign n8155 = n7386 & ~n8154;
  assign n8156 = ~n8151 & ~n8155;
  assign n8157 = pi117 & n7384;
  assign n8158 = pi347 & n7392;
  assign n8159 = pi137 & n7389;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = pi140 & n7391;
  assign n8162 = n8160 & ~n8161;
  assign n8163 = ~n8157 & n8162;
  assign n8164 = n8156 & n8163;
  assign n8165 = ~pi247 & ~n8164;
  assign n8166 = pi217 & pi247;
  assign po262 = n8165 | n8166;
  assign n8168 = pi218 & ~n7443;
  assign n8169 = ~pi218 & n7443;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = ~pi219 & n7443;
  assign n8172 = ~n7779 & ~n8171;
  assign n8173 = ~n7672 & n7781;
  assign n8174 = n8172 & n8173;
  assign n8175 = ~n7786 & n8172;
  assign n8176 = n7443 & ~n7778;
  assign n8177 = ~pi219 & n8171;
  assign n8178 = ~n8176 & ~n8177;
  assign n8179 = n7443 & n8171;
  assign n8180 = ~pi219 & ~n7778;
  assign n8181 = ~n8179 & ~n8180;
  assign n8182 = n8178 & n8181;
  assign n8183 = ~n8175 & ~n8182;
  assign n8184 = ~n8174 & n8183;
  assign n8185 = ~n8170 & n8184;
  assign n8186 = n8170 & ~n8184;
  assign n8187 = ~n8185 & ~n8186;
  assign n8188 = ~n7476 & n8187;
  assign n8189 = pi218 & ~n2653;
  assign n8190 = ~n4127 & ~n8189;
  assign n8191 = n3646 & ~n8190;
  assign n8192 = ~n4172 & ~n8191;
  assign n8193 = ~n2650 & ~n8192;
  assign n8194 = ~n4175 & ~n8193;
  assign n8195 = n2647 & ~n8194;
  assign n8196 = ~n4178 & ~n8195;
  assign n8197 = n2633 & ~n8196;
  assign n8198 = pi218 & ~n2633;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = n7572 & n8199;
  assign n8201 = ~n7572 & ~n8187;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = n7476 & n8202;
  assign n8204 = ~n8188 & ~n8203;
  assign n8205 = n2071 & n8204;
  assign n8206 = ~n2071 & n8199;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 = ~n2070 & ~n8207;
  assign n8209 = n7513 & n8187;
  assign n8210 = pi218 & ~n7513;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = n2071 & ~n8211;
  assign n8213 = pi218 & ~n2071;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = n2070 & n8214;
  assign n8216 = ~n8208 & ~n8215;
  assign n8217 = ~pi247 & n8216;
  assign n8218 = pi218 & pi247;
  assign n8219 = ~n8217 & ~n8218;
  assign po263 = pi359 & ~n8219;
  assign n8221 = pi219 & ~n7443;
  assign n8222 = ~n8171 & ~n8221;
  assign n8223 = n7712 & ~n8018;
  assign n8224 = n7731 & ~n8223;
  assign n8225 = n7716 & ~n8224;
  assign n8226 = n7729 & ~n8225;
  assign n8227 = n7715 & ~n8226;
  assign n8228 = ~n7710 & n8227;
  assign n8229 = ~n7779 & n8228;
  assign n8230 = ~n7710 & ~n7727;
  assign n8231 = ~n7709 & ~n8230;
  assign n8232 = ~n7779 & ~n8231;
  assign n8233 = ~n7778 & ~n8232;
  assign n8234 = ~n8229 & n8233;
  assign n8235 = n8222 & n8234;
  assign n8236 = ~n8222 & ~n8234;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = n7513 & ~n8237;
  assign n8239 = pi219 & ~n7513;
  assign n8240 = ~n8238 & ~n8239;
  assign n8241 = n2071 & ~n8240;
  assign n8242 = pi219 & ~n2071;
  assign n8243 = ~n8241 & ~n8242;
  assign n8244 = n2070 & ~n8243;
  assign n8245 = pi219 & ~n2653;
  assign n8246 = ~n3809 & ~n8245;
  assign n8247 = n3646 & ~n8246;
  assign n8248 = ~n3857 & ~n8247;
  assign n8249 = ~n2650 & ~n8248;
  assign n8250 = ~n3860 & ~n8249;
  assign n8251 = n2647 & ~n8250;
  assign n8252 = ~n3863 & ~n8251;
  assign n8253 = n2633 & ~n8252;
  assign n8254 = pi219 & ~n2633;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = n7572 & n8255;
  assign n8257 = ~n7572 & n8237;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = n7476 & n8258;
  assign n8260 = ~n7476 & ~n8237;
  assign n8261 = ~n8259 & ~n8260;
  assign n8262 = n2071 & n8261;
  assign n8263 = ~n2071 & n8255;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = ~n2070 & n8264;
  assign n8266 = ~n8244 & ~n8265;
  assign n8267 = ~pi247 & ~n8266;
  assign n8268 = pi219 & pi247;
  assign n8269 = ~n8267 & ~n8268;
  assign po264 = pi359 & ~n8269;
  assign n8271 = ~pi220 & n7478;
  assign n8272 = ~n7479 & ~n8271;
  assign n8273 = ~n7476 & n8272;
  assign n8274 = pi220 & ~n2653;
  assign n8275 = ~n4041 & ~n8274;
  assign n8276 = n3646 & ~n8275;
  assign n8277 = ~n4040 & ~n8276;
  assign n8278 = ~n2650 & ~n8277;
  assign n8279 = ~n4046 & ~n8278;
  assign n8280 = n2647 & ~n8279;
  assign n8281 = ~n4049 & ~n8280;
  assign n8282 = n2633 & ~n8281;
  assign n8283 = pi220 & ~n2633;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = n7572 & n8284;
  assign n8286 = ~n7572 & ~n8272;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = n7476 & n8287;
  assign n8289 = ~n8273 & ~n8288;
  assign n8290 = n2071 & n8289;
  assign n8291 = ~n2071 & n8284;
  assign n8292 = ~n8290 & ~n8291;
  assign n8293 = ~n2070 & ~n8292;
  assign n8294 = n7513 & n8272;
  assign n8295 = pi220 & ~n7513;
  assign n8296 = ~n8294 & ~n8295;
  assign n8297 = n2071 & ~n8296;
  assign n8298 = pi220 & ~n2071;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = n2070 & n8299;
  assign n8301 = ~n8293 & ~n8300;
  assign n8302 = ~pi247 & n8301;
  assign n8303 = pi220 & pi247;
  assign n8304 = ~n8302 & ~n8303;
  assign po265 = pi359 & ~n8304;
  assign n8306 = pi221 & ~n7513;
  assign n8307 = ~n7663 & ~n7667;
  assign n8308 = ~n8226 & n8307;
  assign n8309 = n8226 & ~n8307;
  assign n8310 = ~n8308 & ~n8309;
  assign n8311 = n7513 & n8310;
  assign n8312 = ~n8306 & ~n8311;
  assign n8313 = n2071 & ~n8312;
  assign n8314 = pi221 & ~n2071;
  assign n8315 = ~n8313 & ~n8314;
  assign n8316 = n2070 & ~n8315;
  assign n8317 = ~n7476 & n8310;
  assign n8318 = pi221 & ~n2653;
  assign n8319 = ~n3878 & ~n8318;
  assign n8320 = n3646 & ~n8319;
  assign n8321 = ~n3920 & ~n8320;
  assign n8322 = ~n2650 & ~n8321;
  assign n8323 = ~n3923 & ~n8322;
  assign n8324 = n2647 & ~n8323;
  assign n8325 = ~n3926 & ~n8324;
  assign n8326 = n2633 & ~n8325;
  assign n8327 = pi221 & ~n2633;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = n7572 & n8328;
  assign n8330 = ~n7572 & ~n8310;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = n7476 & n8331;
  assign n8333 = ~n8317 & ~n8332;
  assign n8334 = n2071 & n8333;
  assign n8335 = ~n2071 & n8328;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n2070 & n8336;
  assign n8338 = ~n8316 & ~n8337;
  assign n8339 = ~pi247 & ~n8338;
  assign n8340 = pi221 & pi247;
  assign n8341 = ~n8339 & ~n8340;
  assign po266 = pi359 & ~n8341;
  assign n8343 = pi351 & ~n7093;
  assign n8344 = pi222 & n7097;
  assign n8345 = ~n6819 & n7096;
  assign n8346 = ~n8344 & ~n8345;
  assign n8347 = ~n2070 & ~n8346;
  assign n8348 = pi222 & n2070;
  assign n8349 = ~n8347 & ~n8348;
  assign n8350 = n7093 & ~n8349;
  assign n8351 = ~n8343 & ~n8350;
  assign n8352 = n782 & ~n8351;
  assign n8353 = ~n782 & ~n8349;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = ~pi247 & ~n8354;
  assign n8356 = pi222 & pi247;
  assign n8357 = ~n8355 & ~n8356;
  assign po267 = pi359 & ~n8357;
  assign n8359 = pi223 & pi247;
  assign n8360 = pi223 & n7398;
  assign n8361 = ~n1988 & n7277;
  assign n8362 = ~n1676 & ~n7277;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = n7386 & ~n8363;
  assign n8365 = ~n8360 & ~n8364;
  assign n8366 = pi179 & n7384;
  assign n8367 = pi350 & n7392;
  assign n8368 = pi135 & n7389;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = pi133 & n7391;
  assign n8371 = n8369 & ~n8370;
  assign n8372 = ~n8366 & n8371;
  assign n8373 = n8365 & n8372;
  assign n8374 = ~pi247 & ~n8373;
  assign po268 = n8359 | n8374;
  assign n8376 = pi350 & ~n7093;
  assign n8377 = ~pi224 & n7097;
  assign n8378 = ~n6704 & n7096;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = ~n2070 & ~n8379;
  assign n8381 = ~pi224 & n2070;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = n7093 & ~n8382;
  assign n8384 = ~n8376 & ~n8383;
  assign n8385 = n782 & ~n8384;
  assign n8386 = ~n782 & ~n8382;
  assign n8387 = ~n8385 & ~n8386;
  assign n8388 = ~pi247 & ~n8387;
  assign n8389 = ~pi224 & pi247;
  assign n8390 = ~n8388 & ~n8389;
  assign po269 = pi359 & ~n8390;
  assign n8392 = pi225 & n7398;
  assign n8393 = ~n1627 & n7277;
  assign n8394 = ~n1796 & ~n7277;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = n7386 & ~n8395;
  assign n8397 = ~n8392 & ~n8396;
  assign n8398 = pi185 & n7384;
  assign n8399 = pi349 & n7392;
  assign n8400 = pi130 & n7389;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = pi142 & n7391;
  assign n8403 = n8401 & ~n8402;
  assign n8404 = ~n8398 & n8403;
  assign n8405 = n8397 & n8404;
  assign n8406 = ~pi247 & ~n8405;
  assign n8407 = pi225 & pi247;
  assign po270 = n8406 | n8407;
  assign n8409 = pi352 & ~n7093;
  assign n8410 = pi226 & n7097;
  assign n8411 = ~n6609 & n7096;
  assign n8412 = ~n8410 & ~n8411;
  assign n8413 = ~n2070 & ~n8412;
  assign n8414 = pi226 & n2070;
  assign n8415 = ~n8413 & ~n8414;
  assign n8416 = n7093 & ~n8415;
  assign n8417 = ~n8409 & ~n8416;
  assign n8418 = n782 & ~n8417;
  assign n8419 = ~n782 & ~n8415;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~pi247 & ~n8420;
  assign n8422 = pi226 & pi247;
  assign n8423 = ~n8421 & ~n8422;
  assign po271 = pi359 & ~n8423;
  assign n8425 = pi353 & ~n7093;
  assign n8426 = pi227 & n7097;
  assign n8427 = ~n6857 & n7096;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = ~n2070 & ~n8428;
  assign n8430 = pi227 & n2070;
  assign n8431 = ~n8429 & ~n8430;
  assign n8432 = n7093 & ~n8431;
  assign n8433 = ~n8425 & ~n8432;
  assign n8434 = n782 & ~n8433;
  assign n8435 = ~n782 & ~n8431;
  assign n8436 = ~n8434 & ~n8435;
  assign n8437 = ~pi247 & ~n8436;
  assign n8438 = pi227 & pi247;
  assign n8439 = ~n8437 & ~n8438;
  assign po272 = pi359 & ~n8439;
  assign n8441 = pi228 & ~n2633;
  assign n8442 = ~n2070 & n8441;
  assign n8443 = pi345 & ~n2070;
  assign n8444 = pi301 & ~n934;
  assign n8445 = n5096 & ~n8444;
  assign n8446 = n2633 & ~n8445;
  assign n8447 = n8443 & n8446;
  assign n8448 = ~n8442 & ~n8447;
  assign n8449 = ~pi247 & ~n8448;
  assign n8450 = ~pi247 & n2070;
  assign n8451 = pi228 & n8450;
  assign n8452 = ~n8449 & ~n8451;
  assign n8453 = pi359 & ~n8452;
  assign n8454 = pi247 & pi359;
  assign n8455 = pi228 & n8454;
  assign po273 = n8453 | n8455;
  assign n8457 = pi348 & ~n7093;
  assign n8458 = pi229 & n7097;
  assign n8459 = ~n6959 & n7096;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = ~n2070 & ~n8460;
  assign n8462 = pi229 & n2070;
  assign n8463 = ~n8461 & ~n8462;
  assign n8464 = n7093 & ~n8463;
  assign n8465 = ~n8457 & ~n8464;
  assign n8466 = n782 & ~n8465;
  assign n8467 = ~n782 & ~n8463;
  assign n8468 = ~n8466 & ~n8467;
  assign n8469 = ~pi247 & ~n8468;
  assign n8470 = pi229 & pi247;
  assign n8471 = ~n8469 & ~n8470;
  assign po274 = pi359 & ~n8471;
  assign n8473 = ~pi230 & n827;
  assign n8474 = n5005 & n8473;
  assign n8475 = pi359 & n8474;
  assign n8476 = ~n2633 & n8473;
  assign n8477 = ~n5003 & n8476;
  assign n8478 = ~n7508 & ~n8473;
  assign n8479 = n2633 & ~n8478;
  assign n8480 = ~n5003 & n8479;
  assign n8481 = ~n8477 & ~n8480;
  assign n8482 = ~n5005 & ~n8481;
  assign n8483 = n5003 & ~n5005;
  assign n8484 = n8473 & n8483;
  assign n8485 = ~n8482 & ~n8484;
  assign n8486 = pi359 & ~n8485;
  assign po275 = n8475 | n8486;
  assign n8488 = ~n2176 & ~n2256;
  assign n8489 = n811 & ~n8488;
  assign n8490 = n803 & n2280;
  assign n8491 = ~n8489 & ~n8490;
  assign n8492 = ~n4984 & n8491;
  assign n8493 = n787 & ~n8492;
  assign n8494 = ~pi297 & n2087;
  assign n8495 = pi301 & n3322;
  assign n8496 = n8494 & n8495;
  assign n8497 = ~n8493 & ~n8496;
  assign n8498 = ~pi247 & ~n8497;
  assign n8499 = n2633 & n8498;
  assign n8500 = ~n2116 & ~n2173;
  assign n8501 = ~n7299 & n8500;
  assign n8502 = ~n7301 & n8501;
  assign n8503 = ~n7543 & n8502;
  assign n8504 = ~n7538 & n8503;
  assign n8505 = ~n7234 & n8504;
  assign n8506 = ~n7311 & n8505;
  assign n8507 = n811 & n2223;
  assign n8508 = n8506 & ~n8507;
  assign n8509 = ~n874 & ~n2112;
  assign n8510 = ~n2147 & n8509;
  assign n8511 = n8508 & n8510;
  assign n8512 = n780 & n1527;
  assign n8513 = ~n7247 & ~n8512;
  assign n8514 = ~n7323 & n8513;
  assign n8515 = ~n7293 & n8514;
  assign n8516 = n8511 & n8515;
  assign n8517 = ~n2250 & n8516;
  assign n8518 = ~n2154 & n8517;
  assign n8519 = n787 & ~n8518;
  assign n8520 = n811 & n7260;
  assign n8521 = n802 & n2343;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = n780 & n932;
  assign n8524 = n780 & n929;
  assign n8525 = ~n8523 & ~n8524;
  assign n8526 = n8522 & n8525;
  assign n8527 = n7288 & n8526;
  assign n8528 = pi301 & ~n8527;
  assign n8529 = ~n8519 & ~n8528;
  assign n8530 = n811 & ~n2810;
  assign n8531 = n811 & n2096;
  assign n8532 = ~n2489 & ~n8531;
  assign n8533 = ~n2496 & n8532;
  assign n8534 = ~n8530 & n8533;
  assign n8535 = n2109 & ~n8534;
  assign n8536 = n8529 & ~n8535;
  assign n8537 = n2633 & ~n8536;
  assign n8538 = ~pi247 & n8537;
  assign n8539 = ~n8499 & ~n8538;
  assign n8540 = pi359 & ~n8539;
  assign n8541 = ~pi231 & n8454;
  assign po276 = n8540 | n8541;
  assign n8543 = pi349 & ~n7093;
  assign n8544 = ~n6929 & n7096;
  assign n8545 = pi232 & ~n7096;
  assign n8546 = ~n7095 & n8545;
  assign n8547 = ~n8544 & ~n8546;
  assign n8548 = ~n2070 & ~n8547;
  assign n8549 = pi232 & n2070;
  assign n8550 = ~n8548 & ~n8549;
  assign n8551 = n7093 & ~n8550;
  assign n8552 = ~n8543 & ~n8551;
  assign n8553 = n782 & ~n8552;
  assign n8554 = ~n782 & ~n8550;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = ~pi247 & ~n8555;
  assign n8557 = pi232 & pi247;
  assign n8558 = ~n8556 & ~n8557;
  assign po277 = pi359 & ~n8558;
  assign n8560 = n780 & n2636;
  assign n8561 = ~n7562 & ~n8560;
  assign n8562 = n826 & ~n8561;
  assign n8563 = n2712 & n7550;
  assign n8564 = ~n799 & n8563;
  assign n8565 = n811 & ~n8564;
  assign n8566 = ~n8562 & ~n8565;
  assign n8567 = ~n809 & ~n2193;
  assign n8568 = ~n2280 & n8567;
  assign n8569 = ~n838 & n8568;
  assign n8570 = ~n795 & n8569;
  assign n8571 = n811 & ~n8570;
  assign n8572 = n8566 & ~n8571;
  assign n8573 = n787 & ~n8572;
  assign n8574 = ~n909 & n2994;
  assign n8575 = n811 & ~n8574;
  assign n8576 = pi301 & n8575;
  assign n8577 = ~n8573 & ~n8576;
  assign n8578 = pi347 & ~n8577;
  assign n8579 = pi233 & n7097;
  assign n8580 = ~n5978 & n7096;
  assign n8581 = ~n8579 & ~n8580;
  assign n8582 = ~n2070 & ~n8581;
  assign n8583 = pi233 & n2070;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n8577 & ~n8584;
  assign n8586 = ~n8578 & ~n8585;
  assign n8587 = n782 & ~n8586;
  assign n8588 = ~n782 & ~n8584;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 = ~pi247 & ~n8589;
  assign n8591 = pi233 & pi247;
  assign n8592 = ~n8590 & ~n8591;
  assign po278 = pi359 & ~n8592;
  assign n8594 = ~pi247 & ~n7331;
  assign n8595 = n2633 & n8594;
  assign n8596 = ~n8499 & ~n8595;
  assign n8597 = pi359 & ~n8596;
  assign n8598 = ~pi234 & n8454;
  assign po279 = n8597 | n8598;
  assign n8600 = ~pi247 & ~n1780;
  assign n8601 = ~pi235 & pi247;
  assign po280 = n8600 | n8601;
  assign n8603 = ~pi247 & ~n1857;
  assign n8604 = ~pi236 & pi247;
  assign po281 = n8603 | n8604;
  assign po282 = pi252 & pi359;
  assign n8607 = pi354 & ~n7093;
  assign n8608 = pi238 & n7097;
  assign n8609 = ~n6984 & n7096;
  assign n8610 = ~n8608 & ~n8609;
  assign n8611 = ~n2070 & ~n8610;
  assign n8612 = pi238 & n2070;
  assign n8613 = ~n8611 & ~n8612;
  assign n8614 = n7093 & ~n8613;
  assign n8615 = ~n8607 & ~n8614;
  assign n8616 = n782 & ~n8615;
  assign n8617 = ~n782 & ~n8613;
  assign n8618 = ~n8616 & ~n8617;
  assign n8619 = ~pi247 & ~n8618;
  assign n8620 = pi238 & pi247;
  assign n8621 = ~n8619 & ~n8620;
  assign po283 = pi359 & ~n8621;
  assign n8623 = ~pi247 & ~n7277;
  assign n8624 = n2633 & n8623;
  assign n8625 = ~n8499 & ~n8624;
  assign n8626 = pi359 & ~n8625;
  assign n8627 = ~pi239 & n8454;
  assign po284 = n8626 | n8627;
  assign n8629 = ~pi247 & ~n7381;
  assign n8630 = n2633 & n8629;
  assign n8631 = ~n8499 & ~n8630;
  assign n8632 = pi359 & ~n8631;
  assign n8633 = ~pi240 & n8454;
  assign po285 = n8632 | n8633;
  assign n8635 = ~n2162 & ~n2266;
  assign n8636 = ~n2156 & n8635;
  assign n8637 = pi302 & ~n8636;
  assign n8638 = ~n2163 & ~n2270;
  assign n8639 = ~n2274 & n8638;
  assign n8640 = pi302 & ~n8639;
  assign n8641 = ~n7344 & ~n8640;
  assign n8642 = ~n811 & n2236;
  assign n8643 = ~n1527 & ~n8642;
  assign n8644 = pi302 & ~n8643;
  assign n8645 = ~n8512 & ~n8644;
  assign n8646 = pi302 & ~n2543;
  assign n8647 = ~n2223 & ~n2241;
  assign n8648 = ~n2226 & n8647;
  assign n8649 = pi302 & ~n8648;
  assign n8650 = ~n8646 & ~n8649;
  assign n8651 = ~n2250 & n8650;
  assign n8652 = ~n879 & ~n2243;
  assign n8653 = ~n2254 & ~n2256;
  assign n8654 = n2741 & n8653;
  assign n8655 = n2730 & n8654;
  assign n8656 = n8652 & n8655;
  assign n8657 = pi302 & ~n8656;
  assign n8658 = n8651 & ~n8657;
  assign n8659 = ~n2170 & ~n2176;
  assign n8660 = ~n2140 & ~n2179;
  assign n8661 = n8567 & n8660;
  assign n8662 = n2839 & n8661;
  assign n8663 = n8659 & n8662;
  assign n8664 = pi302 & ~n8663;
  assign n8665 = ~n2119 & n2139;
  assign n8666 = ~n838 & n8665;
  assign n8667 = pi302 & ~n8666;
  assign n8668 = ~n8664 & ~n8667;
  assign n8669 = pi302 & n2196;
  assign n8670 = n7307 & n8669;
  assign n8671 = ~pi302 & ~n811;
  assign n8672 = n2197 & ~n8671;
  assign n8673 = ~n8670 & ~n8672;
  assign n8674 = n8668 & n8673;
  assign n8675 = n8658 & n8674;
  assign n8676 = n8645 & n8675;
  assign n8677 = n2911 & n2912;
  assign n8678 = n2916 & n8677;
  assign n8679 = n800 & n8678;
  assign n8680 = pi302 & ~n8679;
  assign n8681 = n8676 & ~n8680;
  assign n8682 = ~n2280 & n2920;
  assign n8683 = ~n2286 & n8682;
  assign n8684 = pi302 & ~n8683;
  assign n8685 = n8681 & ~n8684;
  assign n8686 = n8641 & n8685;
  assign n8687 = ~n8637 & n8686;
  assign n8688 = n787 & ~n8687;
  assign n8689 = ~pi302 & ~n780;
  assign n8690 = ~n2806 & ~n8689;
  assign n8691 = pi302 & ~n780;
  assign n8692 = ~n2807 & n8691;
  assign n8693 = ~n8690 & ~n8692;
  assign n8694 = pi302 & ~n811;
  assign n8695 = ~n2089 & ~n2101;
  assign n8696 = n8694 & ~n8695;
  assign n8697 = ~n2099 & ~n8671;
  assign n8698 = ~n8696 & ~n8697;
  assign n8699 = n8693 & n8698;
  assign n8700 = n2109 & ~n8699;
  assign n8701 = pi302 & n2358;
  assign n8702 = pi302 & n905;
  assign n8703 = ~n8701 & ~n8702;
  assign n8704 = ~n804 & n8671;
  assign n8705 = n2355 & ~n8704;
  assign n8706 = pi302 & n2364;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = ~n7265 & n8707;
  assign n8709 = n2376 & n7307;
  assign n8710 = ~n2329 & ~n8709;
  assign n8711 = n2318 & n8710;
  assign n8712 = pi302 & ~n8711;
  assign n8713 = pi302 & n2348;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = pi302 & n909;
  assign n8716 = n929 & ~n8689;
  assign n8717 = ~n8715 & ~n8716;
  assign n8718 = ~n2343 & ~n2380;
  assign n8719 = pi302 & ~n8718;
  assign n8720 = n8717 & ~n8719;
  assign n8721 = n932 & ~n8689;
  assign n8722 = pi302 & n2337;
  assign n8723 = ~n8721 & ~n8722;
  assign n8724 = ~n2340 & n8723;
  assign n8725 = n8720 & n8724;
  assign n8726 = n8714 & n8725;
  assign n8727 = n8708 & n8726;
  assign n8728 = ~n2472 & ~n2701;
  assign n8729 = pi302 & ~n8728;
  assign n8730 = ~n2360 & ~n2474;
  assign n8731 = pi302 & ~n8730;
  assign n8732 = ~n8729 & ~n8731;
  assign n8733 = n8727 & n8732;
  assign n8734 = ~n935 & n8733;
  assign n8735 = n8703 & n8734;
  assign n8736 = pi301 & ~n8735;
  assign n8737 = ~n8700 & ~n8736;
  assign n8738 = ~n8688 & n8737;
  assign n8739 = n2633 & ~n8738;
  assign n8740 = ~pi247 & pi359;
  assign n8741 = ~n2070 & n8740;
  assign n8742 = n8739 & n8741;
  assign n8743 = pi241 & n8454;
  assign po286 = n8742 | n8743;
  assign n8745 = n787 & n2154;
  assign n8746 = n7345 & n7355;
  assign n8747 = ~n7234 & n8513;
  assign n8748 = ~n2112 & n8747;
  assign n8749 = n7300 & n8748;
  assign n8750 = n8746 & n8749;
  assign n8751 = n787 & ~n8750;
  assign n8752 = ~n8745 & ~n8751;
  assign n8753 = ~n8535 & n8752;
  assign n8754 = ~n2340 & n7369;
  assign n8755 = ~n8523 & n8754;
  assign n8756 = n7287 & ~n8524;
  assign n8757 = ~n7266 & n8756;
  assign n8758 = n8755 & n8757;
  assign n8759 = pi301 & ~n8758;
  assign n8760 = n8753 & ~n8759;
  assign n8761 = n2633 & ~n8760;
  assign n8762 = n8741 & n8761;
  assign n8763 = pi242 & n8454;
  assign po287 = n8762 | n8763;
  assign n8765 = n811 & n2089;
  assign n8766 = n8534 & ~n8765;
  assign n8767 = ~n2490 & n8766;
  assign n8768 = n2109 & ~n8767;
  assign n8769 = ~n2313 & ~n2364;
  assign n8770 = n2634 & ~n8769;
  assign n8771 = ~n8768 & ~n8770;
  assign n8772 = ~n8745 & n8771;
  assign n8773 = n787 & n2116;
  assign n8774 = n8772 & ~n8773;
  assign n8775 = n2633 & ~n8774;
  assign n8776 = n8741 & n8775;
  assign n8777 = pi243 & n8454;
  assign po288 = n8776 | n8777;
  assign n8779 = pi350 & ~n8577;
  assign n8780 = pi244 & n7097;
  assign n8781 = ~n5933 & n7096;
  assign n8782 = ~n8780 & ~n8781;
  assign n8783 = ~n2070 & ~n8782;
  assign n8784 = pi244 & n2070;
  assign n8785 = ~n8783 & ~n8784;
  assign n8786 = n8577 & ~n8785;
  assign n8787 = ~n8779 & ~n8786;
  assign n8788 = n782 & ~n8787;
  assign n8789 = ~n782 & ~n8785;
  assign n8790 = ~n8788 & ~n8789;
  assign n8791 = ~pi247 & ~n8790;
  assign n8792 = pi244 & pi247;
  assign n8793 = ~n8791 & ~n8792;
  assign po289 = pi359 & ~n8793;
  assign n8795 = ~pi247 & ~n1822;
  assign n8796 = ~pi245 & pi247;
  assign po290 = n8795 | n8796;
  assign n8798 = pi298 & n3009;
  assign n8799 = pi246 & ~n3009;
  assign n8800 = ~n8798 & ~n8799;
  assign n8801 = n2071 & ~n8800;
  assign n8802 = pi246 & ~n2071;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = ~n7096 & ~n8803;
  assign n8805 = ~n6192 & n7096;
  assign n8806 = ~n8804 & ~n8805;
  assign n8807 = ~n2070 & ~n8806;
  assign n8808 = pi246 & n2070;
  assign n8809 = ~n8807 & ~n8808;
  assign n8810 = n8577 & ~n8809;
  assign n8811 = pi353 & ~n8577;
  assign n8812 = ~n8810 & ~n8811;
  assign n8813 = n782 & ~n8812;
  assign n8814 = ~n782 & ~n8809;
  assign n8815 = ~n8813 & ~n8814;
  assign n8816 = ~pi247 & ~n8815;
  assign n8817 = pi246 & pi247;
  assign n8818 = ~n8816 & ~n8817;
  assign po291 = pi359 & ~n8818;
  assign n8820 = n2633 & ~n5005;
  assign n8821 = pi356 & n8820;
  assign n8822 = pi359 & n8821;
  assign n8823 = ~n5003 & n8822;
  assign n8824 = n5005 & n8454;
  assign po292 = n8823 | n8824;
  assign n8826 = ~pi247 & ~n1643;
  assign n8827 = pi247 & ~pi248;
  assign po293 = n8826 | n8827;
  assign n8829 = ~pi247 & ~n1838;
  assign n8830 = pi247 & ~pi249;
  assign po294 = n8829 | n8830;
  assign n8832 = ~pi247 & ~n2006;
  assign n8833 = pi247 & ~pi250;
  assign po295 = n8832 | n8833;
  assign n8835 = n2633 & n8497;
  assign n8836 = n8740 & n8835;
  assign n8837 = ~n7343 & n8836;
  assign n8838 = ~pi251 & n8454;
  assign po296 = n8837 | n8838;
  assign n8840 = ~n2633 & ~n4996;
  assign po297 = pi359 & n8840;
  assign n8842 = ~pi247 & ~n1988;
  assign n8843 = pi247 & ~pi253;
  assign po298 = n8842 | n8843;
  assign n8845 = ~pi247 & ~n1676;
  assign n8846 = pi247 & ~pi254;
  assign po299 = n8845 | n8846;
  assign n8848 = ~pi247 & ~n1627;
  assign n8849 = pi247 & ~pi255;
  assign po300 = n8848 | n8849;
  assign n8851 = pi256 & n8454;
  assign n8852 = n2543 & n2730;
  assign n8853 = pi298 & ~n8852;
  assign n8854 = pi298 & ~n811;
  assign n8855 = n2236 & n8854;
  assign n8856 = ~n780 & n1527;
  assign n8857 = pi298 & n8856;
  assign n8858 = ~n8855 & ~n8857;
  assign n8859 = pi298 & ~n8647;
  assign n8860 = n8858 & ~n8859;
  assign n8861 = ~n2226 & n8654;
  assign n8862 = n8652 & n8861;
  assign n8863 = pi298 & ~n8862;
  assign n8864 = pi298 & ~n8663;
  assign n8865 = ~n8863 & ~n8864;
  assign n8866 = pi298 & n7307;
  assign n8867 = n2196 & n8866;
  assign n8868 = n2197 & n8854;
  assign n8869 = ~n8867 & ~n8868;
  assign n8870 = pi298 & ~n8666;
  assign n8871 = n8869 & ~n8870;
  assign n8872 = n8865 & n8871;
  assign n8873 = n8860 & n8872;
  assign n8874 = ~n8853 & n8873;
  assign n8875 = pi298 & n2150;
  assign n8876 = ~n2154 & ~n8875;
  assign n8877 = ~n7324 & n8876;
  assign n8878 = ~n2156 & ~n2263;
  assign n8879 = pi298 & ~n8878;
  assign n8880 = n8877 & ~n8879;
  assign n8881 = pi298 & ~n8683;
  assign n8882 = pi298 & ~n8679;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = n2272 & ~n2274;
  assign n8885 = ~n2163 & n8884;
  assign n8886 = pi298 & ~n8885;
  assign n8887 = pi298 & ~n8635;
  assign n8888 = ~n8886 & ~n8887;
  assign n8889 = n8883 & n8888;
  assign n8890 = n8880 & n8889;
  assign n8891 = n8874 & n8890;
  assign n8892 = n787 & ~n8891;
  assign n8893 = ~n2493 & n8854;
  assign n8894 = pi298 & ~n780;
  assign n8895 = ~n2808 & n8894;
  assign n8896 = ~n8893 & ~n8895;
  assign n8897 = n2109 & ~n8896;
  assign n8898 = pi298 & ~n8718;
  assign n8899 = pi298 & n909;
  assign n8900 = n929 & n8894;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = pi298 & n2358;
  assign n8903 = pi298 & n2329;
  assign n8904 = ~n2360 & ~n2701;
  assign n8905 = pi298 & ~n8904;
  assign n8906 = ~n8903 & ~n8905;
  assign n8907 = ~n8902 & n8906;
  assign n8908 = pi298 & n905;
  assign n8909 = n2355 & n8866;
  assign n8910 = ~n8908 & ~n8909;
  assign n8911 = pi298 & n2364;
  assign n8912 = ~n7265 & ~n8911;
  assign n8913 = ~n935 & n8912;
  assign n8914 = n8910 & n8913;
  assign n8915 = n8907 & n8914;
  assign n8916 = n2376 & n8866;
  assign n8917 = pi298 & ~n2318;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = n8915 & n8918;
  assign n8920 = n8901 & n8919;
  assign n8921 = ~n8898 & n8920;
  assign n8922 = pi298 & n2313;
  assign n8923 = n8921 & ~n8922;
  assign n8924 = pi298 & ~n2525;
  assign n8925 = n932 & n8894;
  assign n8926 = pi298 & n2384;
  assign n8927 = ~n8925 & ~n8926;
  assign n8928 = ~n8924 & n8927;
  assign n8929 = ~n7266 & n8928;
  assign n8930 = n8923 & n8929;
  assign n8931 = pi301 & ~n8930;
  assign n8932 = ~n8897 & ~n8931;
  assign n8933 = ~n8892 & n8932;
  assign n8934 = n8741 & ~n8933;
  assign n8935 = n2633 & n8934;
  assign po301 = n8851 | n8935;
  assign n8937 = pi257 & n8454;
  assign n8938 = pi303 & ~n8666;
  assign n8939 = pi303 & n7307;
  assign n8940 = ~n804 & ~n8939;
  assign n8941 = n2196 & ~n8940;
  assign n8942 = pi303 & ~n811;
  assign n8943 = n2197 & n8942;
  assign n8944 = ~n8941 & ~n8943;
  assign n8945 = pi303 & ~n8862;
  assign n8946 = pi303 & ~n8663;
  assign n8947 = ~n8945 & ~n8946;
  assign n8948 = pi303 & n8856;
  assign n8949 = pi303 & ~n8647;
  assign n8950 = n2236 & n8942;
  assign n8951 = ~n8949 & ~n8950;
  assign n8952 = ~n8948 & n8951;
  assign n8953 = pi303 & ~n8852;
  assign n8954 = n8952 & ~n8953;
  assign n8955 = n8947 & n8954;
  assign n8956 = n8944 & n8955;
  assign n8957 = ~n8938 & n8956;
  assign n8958 = ~n2150 & n8878;
  assign n8959 = pi303 & ~n8958;
  assign n8960 = ~n7229 & ~n8959;
  assign n8961 = ~n2266 & ~n2270;
  assign n8962 = ~n2271 & n8961;
  assign n8963 = ~n2163 & n8962;
  assign n8964 = pi303 & ~n8963;
  assign n8965 = pi303 & ~n8683;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = pi303 & ~n8679;
  assign n8968 = n8966 & ~n8967;
  assign n8969 = n8960 & n8968;
  assign n8970 = n8957 & n8969;
  assign n8971 = n787 & ~n8970;
  assign n8972 = ~n2084 & ~n2103;
  assign n8973 = pi303 & ~n8972;
  assign n8974 = ~n2489 & ~n8973;
  assign n8975 = pi303 & ~n780;
  assign n8976 = ~n2495 & n8975;
  assign n8977 = ~n2810 & n8942;
  assign n8978 = ~n8976 & ~n8977;
  assign n8979 = ~n2089 & ~n2096;
  assign n8980 = pi303 & ~n8979;
  assign n8981 = ~n8765 & ~n8980;
  assign n8982 = ~n8531 & n8981;
  assign n8983 = n8978 & n8982;
  assign n8984 = ~n2490 & n8983;
  assign n8985 = n8974 & n8984;
  assign n8986 = n2109 & ~n8985;
  assign n8987 = n7307 & ~n8939;
  assign n8988 = n2376 & ~n8987;
  assign n8989 = n2318 & ~n2329;
  assign n8990 = pi303 & ~n8989;
  assign n8991 = ~n8988 & ~n8990;
  assign n8992 = pi303 & n2451;
  assign n8993 = n929 & n8975;
  assign n8994 = ~n8992 & ~n8993;
  assign n8995 = ~n909 & ~n2343;
  assign n8996 = pi303 & ~n8995;
  assign n8997 = n8994 & ~n8996;
  assign n8998 = ~n2474 & n8904;
  assign n8999 = pi303 & ~n8998;
  assign n9000 = ~n7266 & ~n8999;
  assign n9001 = pi303 & n905;
  assign n9002 = n2355 & ~n8987;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = pi303 & n2358;
  assign n9005 = n9003 & ~n9004;
  assign n9006 = ~n935 & n9005;
  assign n9007 = pi303 & n2313;
  assign n9008 = n9006 & ~n9007;
  assign n9009 = n9000 & n9008;
  assign n9010 = n8997 & n9009;
  assign n9011 = n8991 & n9010;
  assign n9012 = pi303 & n2348;
  assign n9013 = n9011 & ~n9012;
  assign n9014 = n932 & n8975;
  assign n9015 = pi303 & n2384;
  assign n9016 = ~n9014 & ~n9015;
  assign n9017 = n9013 & n9016;
  assign n9018 = pi301 & ~n9017;
  assign n9019 = ~n8986 & ~n9018;
  assign n9020 = ~n8971 & n9019;
  assign n9021 = n8741 & ~n9020;
  assign n9022 = n2633 & n9021;
  assign po302 = n8937 | n9022;
  assign n9024 = pi247 & ~pi258;
  assign n9025 = ~pi247 & ~n1660;
  assign po303 = n9024 | n9025;
  assign n9027 = pi352 & ~n8577;
  assign n9028 = pi302 & n3009;
  assign n9029 = pi259 & ~n3009;
  assign n9030 = ~n9028 & ~n9029;
  assign n9031 = n2071 & ~n9030;
  assign n9032 = pi259 & ~n2071;
  assign n9033 = ~n9031 & ~n9032;
  assign n9034 = ~n7096 & ~n9033;
  assign n9035 = ~n6237 & n7096;
  assign n9036 = ~n9034 & ~n9035;
  assign n9037 = ~n2070 & ~n9036;
  assign n9038 = pi259 & n2070;
  assign n9039 = ~n9037 & ~n9038;
  assign n9040 = n8577 & ~n9039;
  assign n9041 = ~n9027 & ~n9040;
  assign n9042 = n782 & ~n9041;
  assign n9043 = ~n782 & ~n9039;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = ~pi247 & ~n9044;
  assign n9046 = pi247 & pi259;
  assign n9047 = ~n9045 & ~n9046;
  assign po304 = pi359 & ~n9047;
  assign n9049 = ~pi247 & ~n1796;
  assign n9050 = pi247 & ~pi260;
  assign po305 = n9049 | n9050;
  assign n9052 = ~pi247 & ~n1764;
  assign n9053 = pi247 & ~pi261;
  assign po306 = n9052 | n9053;
  assign n9055 = ~pi247 & ~n1709;
  assign n9056 = pi247 & ~pi262;
  assign po307 = n9055 | n9056;
  assign n9058 = pi247 & ~pi263;
  assign n9059 = ~pi247 & ~n1693;
  assign po308 = n9058 | n9059;
  assign n9061 = pi247 & pi264;
  assign n9062 = ~n2077 & ~n2785;
  assign n9063 = n2196 & ~n7237;
  assign n9064 = n804 & n2133;
  assign n9065 = ~n9063 & ~n9064;
  assign n9066 = ~n1549 & ~n2566;
  assign n9067 = ~n7085 & n9066;
  assign n9068 = n9065 & n9067;
  assign n9069 = n780 & n849;
  assign n9070 = ~n811 & ~n9069;
  assign n9071 = n817 & ~n9070;
  assign n9072 = pi296 & n780;
  assign n9073 = n2286 & n9072;
  assign n9074 = ~n9071 & ~n9073;
  assign n9075 = n826 & ~n827;
  assign n9076 = n780 & n9075;
  assign n9077 = n9074 & ~n9076;
  assign n9078 = ~n2112 & ~n2147;
  assign n9079 = pi296 & ~n9078;
  assign n9080 = ~n7246 & ~n9079;
  assign n9081 = n9077 & n9080;
  assign n9082 = n780 & n833;
  assign n9083 = n9081 & ~n9082;
  assign n9084 = ~n2574 & ~n7088;
  assign n9085 = ~n7535 & n9084;
  assign n9086 = n9083 & n9085;
  assign n9087 = n9068 & n9086;
  assign n9088 = n787 & ~n9087;
  assign n9089 = n2355 & ~n7237;
  assign n9090 = n804 & ~n849;
  assign n9091 = ~n7338 & ~n9090;
  assign n9092 = n2337 & ~n9091;
  assign n9093 = n2376 & ~n7237;
  assign n9094 = n780 & n9004;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = ~n2340 & n9095;
  assign n9097 = ~n9092 & n9096;
  assign n9098 = ~n9089 & n9097;
  assign n9099 = pi301 & ~n9098;
  assign n9100 = ~n9088 & ~n9099;
  assign n9101 = ~n7276 & n9100;
  assign n9102 = n9062 & ~n9101;
  assign n9103 = pi296 & ~n9062;
  assign n9104 = ~n9102 & ~n9103;
  assign n9105 = pi297 & n2594;
  assign n9106 = pi297 & n811;
  assign n9107 = n2140 & n9106;
  assign n9108 = ~n7301 & ~n9107;
  assign n9109 = ~n2173 & n9108;
  assign n9110 = ~n7307 & n7351;
  assign n9111 = n2196 & n9110;
  assign n9112 = n9109 & ~n9111;
  assign n9113 = ~n9105 & n9112;
  assign n9114 = ~n2566 & n9113;
  assign n9115 = ~n9064 & n9114;
  assign n9116 = ~pi302 & ~n849;
  assign n9117 = n818 & ~n9116;
  assign n9118 = n9115 & ~n9117;
  assign n9119 = n2252 & n9106;
  assign n9120 = ~n7293 & ~n8512;
  assign n9121 = ~n2250 & n9120;
  assign n9122 = ~n9119 & n9121;
  assign n9123 = n2241 & n9106;
  assign n9124 = n9122 & ~n9123;
  assign n9125 = n9118 & n9124;
  assign n9126 = ~n2574 & n9125;
  assign n9127 = ~n7535 & n9126;
  assign n9128 = pi297 & ~n9078;
  assign n9129 = n9127 & ~n9128;
  assign n9130 = n787 & ~n9129;
  assign n9131 = ~n812 & ~n1541;
  assign n9132 = n2355 & n9110;
  assign n9133 = ~n805 & n2337;
  assign n9134 = n7351 & n9133;
  assign n9135 = ~n9132 & ~n9134;
  assign n9136 = ~n2340 & n7268;
  assign n9137 = n2376 & n9110;
  assign n9138 = n780 & n8701;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = n9136 & n9139;
  assign n9141 = n9135 & n9140;
  assign n9142 = ~n9131 & n9141;
  assign n9143 = pi301 & ~n9142;
  assign n9144 = ~n9130 & ~n9143;
  assign n9145 = ~n7380 & n9144;
  assign n9146 = n9062 & ~n9145;
  assign n9147 = pi297 & ~n9062;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n7269 & n7332;
  assign n9150 = n849 & n9133;
  assign n9151 = ~n9149 & ~n9150;
  assign n9152 = n850 & n2506;
  assign n9153 = n9151 & ~n9152;
  assign n9154 = n8525 & n9153;
  assign n9155 = pi301 & ~n9154;
  assign n9156 = n2196 & n7332;
  assign n9157 = ~n8512 & n8746;
  assign n9158 = n1551 & n9157;
  assign n9159 = ~n9156 & n9158;
  assign n9160 = ~n810 & ~n834;
  assign n9161 = n9159 & n9160;
  assign n9162 = ~n829 & n9161;
  assign n9163 = n787 & ~n9162;
  assign n9164 = n817 & n849;
  assign n9165 = n787 & n811;
  assign n9166 = n9164 & n9165;
  assign n9167 = ~n9163 & ~n9166;
  assign n9168 = ~n9155 & n9167;
  assign n9169 = n9062 & ~n9168;
  assign n9170 = n7279 & n9133;
  assign n9171 = n2355 & n7308;
  assign n9172 = ~n9170 & ~n9171;
  assign n9173 = n811 & n929;
  assign n9174 = n9172 & ~n9173;
  assign n9175 = n2376 & n7308;
  assign n9176 = n780 & n8902;
  assign n9177 = ~n9175 & ~n9176;
  assign n9178 = n9136 & n9177;
  assign n9179 = ~n4979 & n9178;
  assign n9180 = n9174 & n9179;
  assign n9181 = pi301 & ~n9180;
  assign n9182 = ~n7330 & ~n9181;
  assign n9183 = n780 & ~n7317;
  assign n9184 = ~n7316 & ~n9183;
  assign n9185 = n817 & ~n9184;
  assign n9186 = pi291 & n780;
  assign n9187 = n2286 & n9186;
  assign n9188 = ~n9185 & ~n9187;
  assign n9189 = ~n834 & ~n2574;
  assign n9190 = pi291 & n811;
  assign n9191 = n2241 & n9190;
  assign n9192 = n2252 & n9190;
  assign n9193 = ~n805 & n2238;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = ~n9191 & n9194;
  assign n9196 = ~n7535 & n9195;
  assign n9197 = n2140 & n9190;
  assign n9198 = n2196 & n7308;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = n1551 & n9199;
  assign n9201 = n9196 & n9200;
  assign n9202 = n9189 & n9201;
  assign n9203 = ~n810 & ~n9064;
  assign n9204 = ~n2566 & n9203;
  assign n9205 = n9202 & n9204;
  assign n9206 = pi291 & ~n9078;
  assign n9207 = ~n7323 & ~n9206;
  assign n9208 = n9205 & n9207;
  assign n9209 = ~n829 & n9208;
  assign n9210 = n9188 & n9209;
  assign n9211 = n787 & ~n9210;
  assign n9212 = n9182 & ~n9211;
  assign n9213 = ~n2077 & ~n9212;
  assign n9214 = ~n2785 & n9213;
  assign n9215 = pi291 & ~n9062;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = n9169 & n9216;
  assign n9218 = ~n9148 & n9217;
  assign n9219 = n9104 & n9218;
  assign n9220 = n9148 & n9169;
  assign n9221 = ~n9216 & n9220;
  assign n9222 = ~n9104 & n9221;
  assign n9223 = pi212 & n9222;
  assign n9224 = ~n9219 & ~n9223;
  assign n9225 = n9104 & n9221;
  assign n9226 = pi220 & n9225;
  assign n9227 = n9224 & ~n9226;
  assign n9228 = ~n9169 & ~n9216;
  assign n9229 = ~n9148 & n9228;
  assign n9230 = n9104 & n9229;
  assign n9231 = pi354 & n9230;
  assign n9232 = ~n9104 & n9229;
  assign n9233 = pi126 & n9232;
  assign n9234 = ~n9231 & ~n9233;
  assign n9235 = ~n9104 & n9218;
  assign n9236 = pi132 & n9235;
  assign n9237 = n9148 & n9217;
  assign n9238 = ~n9104 & n9237;
  assign n9239 = pi187 & n9238;
  assign n9240 = ~n9236 & ~n9239;
  assign n9241 = ~n9148 & ~n9216;
  assign n9242 = ~n9169 & ~n9241;
  assign n9243 = ~n6460 & ~n9104;
  assign n9244 = ~n4855 & n9104;
  assign n9245 = ~n9243 & ~n9244;
  assign n9246 = n9242 & ~n9245;
  assign n9247 = n9104 & n9237;
  assign n9248 = pi174 & n9247;
  assign n9249 = ~n9246 & ~n9248;
  assign n9250 = n9240 & n9249;
  assign n9251 = n9234 & n9250;
  assign n9252 = n9227 & n9251;
  assign n9253 = ~pi247 & ~n9252;
  assign po309 = n9061 | n9253;
  assign n9255 = pi348 & ~n8577;
  assign n9256 = pi303 & n3009;
  assign n9257 = pi265 & ~n3009;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = n2071 & ~n9258;
  assign n9260 = pi265 & ~n2071;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = ~n7096 & ~n9261;
  assign n9263 = ~n6535 & n7096;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = ~n2070 & ~n9264;
  assign n9266 = pi265 & n2070;
  assign n9267 = ~n9265 & ~n9266;
  assign n9268 = n8577 & ~n9267;
  assign n9269 = ~n9255 & ~n9268;
  assign n9270 = n782 & ~n9269;
  assign n9271 = ~n782 & ~n9267;
  assign n9272 = ~n9270 & ~n9271;
  assign n9273 = ~pi247 & ~n9272;
  assign n9274 = pi247 & pi265;
  assign n9275 = ~n9273 & ~n9274;
  assign po310 = pi359 & ~n9275;
  assign n9277 = ~pi247 & ~n1727;
  assign n9278 = pi247 & ~pi266;
  assign po311 = n9277 | n9278;
  assign n9280 = pi247 & ~pi267;
  assign n9281 = ~pi247 & ~n1744;
  assign po312 = n9280 | n9281;
  assign n9283 = pi351 & ~n8577;
  assign n9284 = pi268 & n7097;
  assign n9285 = ~n6509 & n7096;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = ~n2070 & ~n9286;
  assign n9288 = pi268 & n2070;
  assign n9289 = ~n9287 & ~n9288;
  assign n9290 = n8577 & ~n9289;
  assign n9291 = ~n9283 & ~n9290;
  assign n9292 = n782 & ~n9291;
  assign n9293 = ~n782 & ~n9289;
  assign n9294 = ~n9292 & ~n9293;
  assign n9295 = ~pi247 & ~n9294;
  assign n9296 = pi247 & pi268;
  assign n9297 = ~n9295 & ~n9296;
  assign po313 = pi359 & ~n9297;
  assign n9299 = pi247 & pi269;
  assign n9300 = pi347 & n9230;
  assign n9301 = pi140 & n9232;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = pi219 & n9222;
  assign n9304 = pi211 & n9225;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 = pi131 & n9235;
  assign n9307 = pi117 & n9238;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = ~n4715 & ~n9104;
  assign n9310 = ~n3305 & n9104;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = n9242 & ~n9311;
  assign n9313 = pi137 & n9247;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = n9308 & n9314;
  assign n9316 = n9305 & n9315;
  assign n9317 = n9302 & n9316;
  assign n9318 = ~pi247 & ~n9317;
  assign po314 = n9299 | n9318;
  assign n9320 = pi247 & pi270;
  assign n9321 = pi204 & n9222;
  assign n9322 = pi209 & n9225;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = pi352 & n9230;
  assign n9325 = pi143 & n9232;
  assign n9326 = ~n9324 & ~n9325;
  assign n9327 = pi184 & n9235;
  assign n9328 = pi177 & n9238;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = ~n5053 & ~n9104;
  assign n9331 = ~n3423 & n9104;
  assign n9332 = ~n9330 & ~n9331;
  assign n9333 = n9242 & ~n9332;
  assign n9334 = pi146 & n9247;
  assign n9335 = ~n9333 & ~n9334;
  assign n9336 = n9329 & n9335;
  assign n9337 = n9326 & n9336;
  assign n9338 = n9323 & n9337;
  assign n9339 = ~pi247 & ~n9338;
  assign po315 = n9320 | n9339;
  assign n9341 = pi247 & pi271;
  assign n9342 = pi199 & n9222;
  assign n9343 = pi206 & n9225;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = pi349 & n9230;
  assign n9346 = pi142 & n9232;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = pi129 & n9235;
  assign n9349 = pi185 & n9238;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n5688 & ~n9104;
  assign n9352 = ~n4687 & n9104;
  assign n9353 = ~n9351 & ~n9352;
  assign n9354 = n9242 & ~n9353;
  assign n9355 = pi130 & n9247;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = n9350 & n9356;
  assign n9358 = n9347 & n9357;
  assign n9359 = n9344 & n9358;
  assign n9360 = ~pi247 & ~n9359;
  assign po316 = n9341 | n9360;
  assign n9362 = pi247 & pi272;
  assign n9363 = pi203 & n9222;
  assign n9364 = pi208 & n9225;
  assign n9365 = ~n9363 & ~n9364;
  assign n9366 = pi348 & n9230;
  assign n9367 = pi138 & n9232;
  assign n9368 = ~n9366 & ~n9367;
  assign n9369 = ~pi180 & n9235;
  assign n9370 = pi186 & n9238;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = ~n5569 & ~n9104;
  assign n9373 = ~n4569 & n9104;
  assign n9374 = ~n9372 & ~n9373;
  assign n9375 = n9242 & ~n9374;
  assign n9376 = pi173 & n9247;
  assign n9377 = ~n9375 & ~n9376;
  assign n9378 = n9371 & n9377;
  assign n9379 = n9368 & n9378;
  assign n9380 = n9365 & n9379;
  assign n9381 = ~pi247 & ~n9380;
  assign po317 = n9362 | n9381;
  assign n9383 = pi247 & pi273;
  assign n9384 = pi205 & n9222;
  assign n9385 = pi210 & n9225;
  assign n9386 = ~n9384 & ~n9385;
  assign n9387 = pi353 & n9230;
  assign n9388 = pi139 & n9232;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n5081 & ~n9104;
  assign n9391 = ~n4496 & n9104;
  assign n9392 = ~n9390 & ~n9391;
  assign n9393 = n9242 & ~n9392;
  assign n9394 = pi144 & n9247;
  assign n9395 = ~n9393 & ~n9394;
  assign n9396 = ~pi181 & n9235;
  assign n9397 = pi183 & n9238;
  assign n9398 = ~n9396 & ~n9397;
  assign n9399 = n9395 & n9398;
  assign n9400 = n9389 & n9399;
  assign n9401 = n9386 & n9400;
  assign n9402 = ~pi247 & ~n9401;
  assign po318 = n9383 | n9402;
  assign n9404 = pi247 & pi274;
  assign n9405 = pi351 & n9230;
  assign n9406 = pi141 & n9232;
  assign n9407 = ~n9405 & ~n9406;
  assign n9408 = pi221 & n9222;
  assign n9409 = pi207 & n9225;
  assign n9410 = ~n9408 & ~n9409;
  assign n9411 = pi102 & n9235;
  assign n9412 = pi182 & n9238;
  assign n9413 = ~n9411 & ~n9412;
  assign n9414 = ~n6279 & ~n9104;
  assign n9415 = ~n3518 & n9104;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = n9242 & ~n9416;
  assign n9418 = pi172 & n9247;
  assign n9419 = ~n9417 & ~n9418;
  assign n9420 = n9413 & n9419;
  assign n9421 = n9410 & n9420;
  assign n9422 = n9407 & n9421;
  assign n9423 = ~pi247 & ~n9422;
  assign po319 = n9404 | n9423;
  assign n9425 = pi247 & pi275;
  assign n9426 = pi350 & n9230;
  assign n9427 = pi133 & n9232;
  assign n9428 = ~n9426 & ~n9427;
  assign n9429 = pi218 & n9222;
  assign n9430 = pi200 & n9225;
  assign n9431 = ~n9429 & ~n9430;
  assign n9432 = pi178 & n9235;
  assign n9433 = pi179 & n9238;
  assign n9434 = ~n9432 & ~n9433;
  assign n9435 = ~n4877 & ~n9104;
  assign n9436 = ~n4420 & n9104;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = n9242 & ~n9437;
  assign n9439 = pi135 & n9247;
  assign n9440 = ~n9438 & ~n9439;
  assign n9441 = n9434 & n9440;
  assign n9442 = n9431 & n9441;
  assign n9443 = n9428 & n9442;
  assign n9444 = ~pi247 & ~n9443;
  assign po320 = n9425 | n9444;
  assign n9446 = pi349 & ~n8577;
  assign n9447 = pi276 & n7097;
  assign n9448 = ~n5762 & n7096;
  assign n9449 = ~n9447 & ~n9448;
  assign n9450 = ~n2070 & ~n9449;
  assign n9451 = pi276 & n2070;
  assign n9452 = ~n9450 & ~n9451;
  assign n9453 = n8577 & ~n9452;
  assign n9454 = ~n9446 & ~n9453;
  assign n9455 = n782 & ~n9454;
  assign n9456 = ~n782 & ~n9452;
  assign n9457 = ~n9455 & ~n9456;
  assign n9458 = ~pi247 & ~n9457;
  assign n9459 = pi247 & pi276;
  assign n9460 = ~n9458 & ~n9459;
  assign po321 = pi359 & ~n9460;
  assign n9462 = ~n2650 & ~n5394;
  assign n9463 = n2784 & n9462;
  assign n9464 = ~pi247 & ~n9463;
  assign n9465 = pi247 & pi277;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = ~n1575 & ~n9462;
  assign n9468 = ~n2077 & ~n9467;
  assign n9469 = ~pi247 & ~n9468;
  assign po322 = ~n9466 | n9469;
  assign n9471 = pi247 & pi278;
  assign n9472 = ~pi294 & n804;
  assign n9473 = ~pi247 & pi301;
  assign n9474 = n8933 & ~n9020;
  assign n9475 = n9473 & n9474;
  assign n9476 = n9472 & n9475;
  assign n9477 = ~n9471 & ~n9476;
  assign po323 = pi359 & ~n9477;
  assign n9479 = n2099 & ~n2101;
  assign n9480 = n804 & ~n9479;
  assign n9481 = n2109 & n9480;
  assign n9482 = pi196 & n826;
  assign n9483 = n788 & n9482;
  assign n9484 = pi195 & n826;
  assign n9485 = n788 & n9484;
  assign n9486 = ~pi196 & n9485;
  assign n9487 = n803 & n2133;
  assign n9488 = n802 & n2238;
  assign n9489 = ~n9487 & ~n9488;
  assign n9490 = ~n2197 & ~n2236;
  assign n9491 = n804 & ~n9490;
  assign n9492 = n9489 & ~n9491;
  assign n9493 = n788 & n833;
  assign n9494 = n9492 & ~n9493;
  assign n9495 = n811 & n2286;
  assign n9496 = n804 & n2241;
  assign n9497 = ~n2170 & ~n2254;
  assign n9498 = n811 & ~n9497;
  assign n9499 = ~n9496 & ~n9498;
  assign n9500 = n802 & ~n2827;
  assign n9501 = n9499 & ~n9500;
  assign n9502 = ~n9495 & n9501;
  assign n9503 = ~n4985 & n9502;
  assign n9504 = n9494 & n9503;
  assign n9505 = n788 & n817;
  assign n9506 = n9504 & ~n9505;
  assign n9507 = ~n890 & n9506;
  assign n9508 = ~n9486 & n9507;
  assign n9509 = ~n9483 & n9508;
  assign n9510 = n787 & ~n9509;
  assign n9511 = n803 & ~n8769;
  assign n9512 = n802 & n2337;
  assign n9513 = ~n9511 & ~n9512;
  assign n9514 = ~n933 & ~n4977;
  assign n9515 = ~n930 & n9514;
  assign n9516 = ~n912 & n9515;
  assign n9517 = n9513 & n9516;
  assign n9518 = pi301 & ~n9517;
  assign n9519 = ~n9510 & ~n9518;
  assign n9520 = ~n9481 & n9519;
  assign n9521 = n785 & ~n9520;
  assign n9522 = n4988 & ~n9521;
  assign n9523 = ~n3255 & ~n5003;
  assign n9524 = ~n7299 & n7439;
  assign n9525 = n787 & ~n9524;
  assign n9526 = ~n805 & n905;
  assign n9527 = ~n7285 & ~n9526;
  assign n9528 = n803 & ~n1541;
  assign n9529 = n803 & n901;
  assign n9530 = n811 & n2313;
  assign n9531 = ~n9529 & ~n9530;
  assign n9532 = ~n9528 & n9531;
  assign n9533 = ~n7286 & n9532;
  assign n9534 = n9527 & n9533;
  assign n9535 = pi301 & ~n9534;
  assign n9536 = ~n9525 & ~n9535;
  assign n9537 = n2785 & n7568;
  assign n9538 = n9520 & ~n9537;
  assign n9539 = n9536 & n9538;
  assign n9540 = ~n9523 & n9539;
  assign n9541 = ~n9521 & ~n9540;
  assign n9542 = ~n9522 & ~n9541;
  assign n9543 = ~n780 & ~n9542;
  assign n9544 = ~n780 & n9521;
  assign n9545 = n4988 & n9544;
  assign n9546 = ~n9543 & ~n9545;
  assign n9547 = n780 & n9523;
  assign n9548 = pi359 & ~n9547;
  assign n9549 = ~n2603 & n9548;
  assign po324 = ~n9546 | ~n9549;
  assign n9551 = n9148 & ~n9216;
  assign n9552 = n2977 & n9551;
  assign n9553 = pi314 & n9552;
  assign n9554 = pi304 & ~n9552;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = ~pi247 & ~n9555;
  assign n9557 = pi247 & pi280;
  assign po325 = n9556 | n9557;
  assign n9559 = ~n4988 & ~n9521;
  assign n9560 = ~n9541 & ~n9559;
  assign n9561 = ~n780 & ~n9560;
  assign n9562 = ~n4988 & n9544;
  assign n9563 = ~n9561 & ~n9562;
  assign n9564 = ~pi195 & ~n9523;
  assign n9565 = ~n782 & ~n9564;
  assign n9566 = n780 & n9565;
  assign n9567 = n9563 & ~n9566;
  assign po326 = ~pi359 | ~n9567;
  assign n9569 = pi354 & ~n8577;
  assign n9570 = pi282 & n7097;
  assign n9571 = ~n6560 & n7096;
  assign n9572 = ~n9570 & ~n9571;
  assign n9573 = ~n2070 & ~n9572;
  assign n9574 = pi282 & n2070;
  assign n9575 = ~n9573 & ~n9574;
  assign n9576 = n8577 & ~n9575;
  assign n9577 = ~n9569 & ~n9576;
  assign n9578 = n782 & ~n9577;
  assign n9579 = ~n782 & ~n9575;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = ~pi247 & ~n9580;
  assign n9582 = pi247 & pi282;
  assign n9583 = ~n9581 & ~n9582;
  assign po327 = pi359 & ~n9583;
  assign n9585 = ~pi247 & ~n9148;
  assign n9586 = pi247 & pi283;
  assign n9587 = ~n9585 & ~n9586;
  assign n9588 = ~pi247 & n9552;
  assign po328 = ~n9587 | n9588;
  assign n9590 = ~pi247 & ~n9216;
  assign n9591 = pi247 & pi284;
  assign n9592 = ~n9590 & ~n9591;
  assign po329 = n9588 | ~n9592;
  assign n9594 = ~pi247 & n9462;
  assign n9595 = n2958 & n9594;
  assign n9596 = pi247 & pi285;
  assign n9597 = ~n9595 & ~n9596;
  assign po330 = n9469 | ~n9597;
  assign n9599 = n5242 & n5643;
  assign n9600 = pi140 & n9599;
  assign n9601 = n2070 & n2071;
  assign n9602 = pi292 & pi295;
  assign n9603 = pi289 & n9602;
  assign n9604 = pi290 & n9603;
  assign n9605 = pi288 & n9604;
  assign n9606 = pi287 & n9605;
  assign n9607 = pi286 & n9606;
  assign n9608 = ~pi286 & ~n9606;
  assign n9609 = ~n9607 & ~n9608;
  assign n9610 = n9601 & n9609;
  assign n9611 = pi286 & ~n9601;
  assign n9612 = ~n9610 & ~n9611;
  assign n9613 = n5242 & ~n5643;
  assign n9614 = n5242 & ~n9613;
  assign n9615 = ~n9612 & ~n9614;
  assign n9616 = ~n9600 & ~n9615;
  assign n9617 = n5258 & ~n9616;
  assign n9618 = n782 & n9617;
  assign n9619 = ~n5259 & ~n9612;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = ~pi247 & ~n9620;
  assign n9622 = pi247 & pi286;
  assign n9623 = ~n9621 & ~n9622;
  assign po331 = pi359 & ~n9623;
  assign n9625 = pi139 & n9599;
  assign n9626 = pi288 & pi290;
  assign n9627 = n9603 & n9626;
  assign n9628 = pi287 & ~n9627;
  assign n9629 = ~pi287 & n9627;
  assign n9630 = ~n9628 & ~n9629;
  assign n9631 = n9601 & ~n9630;
  assign n9632 = pi287 & ~n9601;
  assign n9633 = ~n9631 & ~n9632;
  assign n9634 = ~n9614 & ~n9633;
  assign n9635 = ~n9625 & ~n9634;
  assign n9636 = n5258 & ~n9635;
  assign n9637 = n782 & n9636;
  assign n9638 = ~n5259 & ~n9633;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = ~pi247 & ~n9639;
  assign n9641 = pi247 & pi287;
  assign n9642 = ~n9640 & ~n9641;
  assign po332 = pi359 & ~n9642;
  assign n9644 = pi138 & n9599;
  assign n9645 = pi288 & ~n9603;
  assign n9646 = ~pi288 & n9603;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = n9601 & ~n9647;
  assign n9649 = pi288 & ~n9601;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = ~n9614 & ~n9650;
  assign n9652 = ~n9644 & ~n9651;
  assign n9653 = n5258 & ~n9652;
  assign n9654 = n782 & n9653;
  assign n9655 = ~n5259 & ~n9650;
  assign n9656 = ~n9654 & ~n9655;
  assign n9657 = ~pi247 & ~n9656;
  assign n9658 = pi247 & pi288;
  assign n9659 = ~n9657 & ~n9658;
  assign po333 = pi359 & ~n9659;
  assign n9661 = pi141 & n9599;
  assign n9662 = pi289 & ~n9602;
  assign n9663 = ~pi289 & n9602;
  assign n9664 = ~n9662 & ~n9663;
  assign n9665 = n9601 & ~n9664;
  assign n9666 = pi289 & ~n9601;
  assign n9667 = ~n9665 & ~n9666;
  assign n9668 = ~n9614 & ~n9667;
  assign n9669 = ~n9661 & ~n9668;
  assign n9670 = n5258 & ~n9669;
  assign n9671 = n782 & n9670;
  assign n9672 = ~n5259 & ~n9667;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = ~pi247 & ~n9673;
  assign n9675 = pi247 & pi289;
  assign n9676 = ~n9674 & ~n9675;
  assign po334 = pi359 & ~n9676;
  assign n9678 = pi143 & n9599;
  assign n9679 = pi288 & pi289;
  assign n9680 = n9602 & n9679;
  assign n9681 = pi290 & ~n9680;
  assign n9682 = ~pi290 & n9680;
  assign n9683 = ~n9681 & ~n9682;
  assign n9684 = n9601 & ~n9683;
  assign n9685 = pi290 & ~n9601;
  assign n9686 = ~n9684 & ~n9685;
  assign n9687 = ~n9614 & ~n9686;
  assign n9688 = ~n9678 & ~n9687;
  assign n9689 = n5258 & ~n9688;
  assign n9690 = n782 & n9689;
  assign n9691 = ~n5259 & ~n9686;
  assign n9692 = ~n9690 & ~n9691;
  assign n9693 = ~pi247 & ~n9692;
  assign n9694 = pi247 & pi290;
  assign n9695 = ~n9693 & ~n9694;
  assign po335 = pi359 & ~n9695;
  assign n9697 = n2109 & n2785;
  assign n9698 = pi291 & ~n9697;
  assign n9699 = pi367 & n9697;
  assign n9700 = ~n9698 & ~n9699;
  assign n9701 = ~n2070 & n2071;
  assign n9702 = ~n9700 & n9701;
  assign n9703 = ~pi331 & pi333;
  assign n9704 = pi195 & n9703;
  assign n9705 = n2071 & n9704;
  assign n9706 = pi195 & n2651;
  assign n9707 = pi230 & ~n9706;
  assign n9708 = ~pi196 & n9707;
  assign n9709 = pi367 & n2071;
  assign n9710 = n9708 & n9709;
  assign n9711 = ~n9705 & ~n9710;
  assign n9712 = n2070 & ~n9711;
  assign n9713 = pi291 & ~n2071;
  assign n9714 = ~n9712 & ~n9713;
  assign n9715 = ~n9702 & n9714;
  assign n9716 = ~pi247 & ~n9715;
  assign n9717 = pi247 & pi291;
  assign n9718 = ~n9716 & ~n9717;
  assign po336 = pi359 & ~n9718;
  assign n9720 = pi126 & n9599;
  assign n9721 = pi292 & ~n2070;
  assign n9722 = pi292 & ~n2071;
  assign n9723 = ~pi292 & n2071;
  assign n9724 = ~n9722 & ~n9723;
  assign n9725 = n2070 & ~n9724;
  assign n9726 = ~n9721 & ~n9725;
  assign n9727 = ~n9614 & ~n9726;
  assign n9728 = ~n9720 & ~n9727;
  assign n9729 = n5258 & ~n9728;
  assign n9730 = n782 & n9729;
  assign n9731 = ~n5259 & ~n9726;
  assign n9732 = ~n9730 & ~n9731;
  assign n9733 = ~pi247 & ~n9732;
  assign n9734 = pi247 & pi292;
  assign n9735 = ~n9733 & ~n9734;
  assign po337 = pi359 & ~n9735;
  assign n9737 = ~n780 & ~n9540;
  assign n9738 = pi359 & ~n4991;
  assign n9739 = ~n9547 & n9738;
  assign po338 = n9737 | ~n9739;
  assign n9741 = n2070 & ~n2071;
  assign n9742 = pi294 & n9741;
  assign n9743 = ~n7142 & n7148;
  assign n9744 = n9601 & ~n9743;
  assign n9745 = ~n7142 & n9744;
  assign n9746 = ~n7149 & n9745;
  assign n9747 = ~n2070 & ~n2077;
  assign n9748 = pi294 & n9747;
  assign n9749 = ~n7142 & ~n7148;
  assign n9750 = ~pi294 & ~n9749;
  assign n9751 = n2077 & ~n9750;
  assign n9752 = ~n2070 & n9751;
  assign n9753 = ~n9748 & ~n9752;
  assign n9754 = ~n9746 & n9753;
  assign n9755 = ~n9742 & n9754;
  assign n9756 = ~pi247 & ~n9755;
  assign n9757 = pi247 & pi294;
  assign n9758 = ~n9756 & ~n9757;
  assign po339 = pi359 & ~n9758;
  assign n9760 = pi142 & n9599;
  assign n9761 = pi295 & ~n2070;
  assign n9762 = pi292 & ~pi295;
  assign n9763 = ~pi292 & pi295;
  assign n9764 = ~n9762 & ~n9763;
  assign n9765 = n2071 & ~n9764;
  assign n9766 = pi295 & ~n2071;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = n2070 & ~n9767;
  assign n9769 = ~n9761 & ~n9768;
  assign n9770 = ~n9614 & ~n9769;
  assign n9771 = ~n9760 & ~n9770;
  assign n9772 = n5258 & ~n9771;
  assign n9773 = n782 & n9772;
  assign n9774 = ~n5259 & ~n9769;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = ~pi247 & ~n9775;
  assign n9777 = pi247 & pi295;
  assign n9778 = ~n9776 & ~n9777;
  assign po340 = pi359 & ~n9778;
  assign n9780 = pi296 & ~n9697;
  assign n9781 = pi365 & n9697;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = n9701 & ~n9782;
  assign n9784 = pi365 & n2071;
  assign n9785 = n9708 & n9784;
  assign n9786 = ~n9705 & ~n9785;
  assign n9787 = n2070 & ~n9786;
  assign n9788 = pi296 & ~n2071;
  assign n9789 = ~n9787 & ~n9788;
  assign n9790 = ~n9783 & n9789;
  assign n9791 = ~pi247 & ~n9790;
  assign n9792 = pi247 & pi296;
  assign n9793 = ~n9791 & ~n9792;
  assign po341 = pi359 & ~n9793;
  assign n9795 = pi297 & ~n9697;
  assign n9796 = pi366 & n9697;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = n9701 & ~n9797;
  assign n9799 = pi366 & n2071;
  assign n9800 = n9708 & n9799;
  assign n9801 = ~n9705 & ~n9800;
  assign n9802 = n2070 & ~n9801;
  assign n9803 = pi297 & ~n2071;
  assign n9804 = ~n9802 & ~n9803;
  assign n9805 = ~n9798 & n9804;
  assign n9806 = ~pi247 & ~n9805;
  assign n9807 = pi247 & pi297;
  assign n9808 = ~n9806 & ~n9807;
  assign po342 = pi359 & ~n9808;
  assign n9810 = pi298 & ~n9697;
  assign n9811 = pi370 & n9697;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = n9701 & ~n9812;
  assign n9814 = pi370 & n2071;
  assign n9815 = n9708 & n9814;
  assign n9816 = ~n9705 & ~n9815;
  assign n9817 = n2070 & ~n9816;
  assign n9818 = pi298 & ~n2071;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = ~n9813 & n9819;
  assign n9821 = ~pi247 & ~n9820;
  assign n9822 = pi247 & pi298;
  assign n9823 = ~n9821 & ~n9822;
  assign po343 = pi359 & ~n9823;
  assign n9825 = pi299 & ~n9697;
  assign n9826 = pi371 & n9697;
  assign n9827 = ~n9825 & ~n9826;
  assign n9828 = n9701 & ~n9827;
  assign n9829 = pi371 & n2071;
  assign n9830 = n9708 & n9829;
  assign n9831 = ~n9705 & ~n9830;
  assign n9832 = n2070 & ~n9831;
  assign n9833 = pi299 & ~n2071;
  assign n9834 = ~n9832 & ~n9833;
  assign n9835 = ~n9828 & n9834;
  assign n9836 = ~pi247 & ~n9835;
  assign n9837 = pi247 & pi299;
  assign n9838 = ~n9836 & ~n9837;
  assign po344 = pi359 & ~n9838;
  assign n9840 = pi300 & ~n9697;
  assign n9841 = pi372 & n9697;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = n9701 & ~n9842;
  assign n9844 = pi372 & n2071;
  assign n9845 = n9708 & n9844;
  assign n9846 = ~n9705 & ~n9845;
  assign n9847 = n2070 & ~n9846;
  assign n9848 = pi300 & ~n2071;
  assign n9849 = ~n9847 & ~n9848;
  assign n9850 = ~n9843 & n9849;
  assign n9851 = ~pi247 & ~n9850;
  assign n9852 = pi247 & pi300;
  assign n9853 = ~n9851 & ~n9852;
  assign po345 = pi359 & ~n9853;
  assign n9855 = pi301 & n9741;
  assign n9856 = n7148 & n9744;
  assign n9857 = ~n7149 & n9856;
  assign n9858 = pi301 & n9747;
  assign n9859 = ~n2070 & ~n9749;
  assign n9860 = pi301 & n9859;
  assign n9861 = n2077 & n9860;
  assign n9862 = ~n9858 & ~n9861;
  assign n9863 = ~n9857 & n9862;
  assign n9864 = ~n9855 & n9863;
  assign n9865 = ~pi247 & ~n9864;
  assign n9866 = pi247 & pi301;
  assign n9867 = ~n9865 & ~n9866;
  assign po346 = pi359 & ~n9867;
  assign n9869 = pi302 & ~n9697;
  assign n9870 = pi369 & n9697;
  assign n9871 = ~n9869 & ~n9870;
  assign n9872 = n9701 & ~n9871;
  assign n9873 = pi369 & n2071;
  assign n9874 = n9708 & n9873;
  assign n9875 = ~n9705 & ~n9874;
  assign n9876 = n2070 & ~n9875;
  assign n9877 = pi302 & ~n2071;
  assign n9878 = ~n9876 & ~n9877;
  assign n9879 = ~n9872 & n9878;
  assign n9880 = ~pi247 & ~n9879;
  assign n9881 = pi247 & pi302;
  assign n9882 = ~n9880 & ~n9881;
  assign po347 = pi359 & ~n9882;
  assign n9884 = pi303 & ~n9697;
  assign n9885 = pi368 & n9697;
  assign n9886 = ~n9884 & ~n9885;
  assign n9887 = n9701 & ~n9886;
  assign n9888 = pi368 & n2071;
  assign n9889 = n9708 & n9888;
  assign n9890 = ~n9705 & ~n9889;
  assign n9891 = n2070 & ~n9890;
  assign n9892 = pi303 & ~n2071;
  assign n9893 = ~n9891 & ~n9892;
  assign n9894 = ~n9887 & n9893;
  assign n9895 = ~pi247 & ~n9894;
  assign n9896 = pi247 & pi303;
  assign n9897 = ~n9895 & ~n9896;
  assign po348 = pi359 & ~n9897;
  assign n9899 = pi304 & n2070;
  assign n9900 = pi302 & n7131;
  assign n9901 = n870 & n9900;
  assign n9902 = n787 & n9901;
  assign n9903 = pi296 & n9902;
  assign n9904 = pi303 & n9903;
  assign n9905 = pi304 & n9904;
  assign n9906 = ~pi304 & ~n9904;
  assign n9907 = ~n9905 & ~n9906;
  assign n9908 = ~n2070 & n9907;
  assign n9909 = ~n9899 & ~n9908;
  assign n9910 = ~pi247 & ~n9909;
  assign n9911 = pi247 & pi304;
  assign n9912 = ~n9910 & ~n9911;
  assign po349 = pi359 & ~n9912;
  assign n9914 = ~n7149 & n9743;
  assign n9915 = n7142 & n7148;
  assign n9916 = ~n7149 & ~n9915;
  assign n9917 = ~n9743 & n9916;
  assign n9918 = ~n9914 & ~n9917;
  assign n9919 = pi305 & ~n9918;
  assign n9920 = n2071 & ~n9919;
  assign n9921 = ~pi305 & ~n2071;
  assign n9922 = ~n9920 & ~n9921;
  assign n9923 = n2070 & n9922;
  assign n9924 = ~pi305 & ~n2077;
  assign n9925 = ~n2070 & ~n9924;
  assign n9926 = ~n9923 & ~n9925;
  assign n9927 = ~pi247 & ~n9926;
  assign n9928 = pi247 & pi305;
  assign n9929 = ~n9927 & ~n9928;
  assign po350 = pi359 & ~n9929;
  assign po351 = ~pi359 | ~n9544;
  assign n9932 = n870 & n5721;
  assign n9933 = ~n7137 & ~n9932;
  assign n9934 = ~pi296 & ~n9933;
  assign n9935 = ~pi302 & n5626;
  assign n9936 = ~pi291 & n9935;
  assign n9937 = ~n1558 & ~n9936;
  assign n9938 = n821 & ~n9937;
  assign n9939 = ~pi296 & n1558;
  assign n9940 = n870 & n9939;
  assign n9941 = ~pi303 & n5626;
  assign n9942 = n852 & n2091;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = n870 & ~n9943;
  assign n9945 = ~pi296 & n9944;
  assign n9946 = ~n9940 & ~n9945;
  assign n9947 = ~n9938 & ~n9946;
  assign n9948 = ~n9934 & n9947;
  assign n9949 = n9938 & n9946;
  assign n9950 = n9934 & n9949;
  assign n9951 = ~n9948 & ~n9950;
  assign n9952 = n9938 & ~n9946;
  assign n9953 = n9934 & n9952;
  assign n9954 = ~pi300 & n849;
  assign n9955 = n7505 & n9954;
  assign n9956 = n981 & n3322;
  assign n9957 = pi296 & ~n9956;
  assign n9958 = ~n9955 & ~n9957;
  assign n9959 = n2151 & n5721;
  assign n9960 = ~n1358 & ~n2309;
  assign n9961 = ~pi300 & n9960;
  assign n9962 = ~n792 & n9961;
  assign n9963 = ~pi291 & ~n9962;
  assign n9964 = ~n9959 & ~n9963;
  assign n9965 = ~pi300 & n850;
  assign n9966 = ~pi297 & ~n9965;
  assign n9967 = n9964 & ~n9966;
  assign n9968 = n9958 & n9967;
  assign n9969 = ~n9938 & n9946;
  assign n9970 = ~n9934 & n9969;
  assign n9971 = ~n9968 & n9970;
  assign n9972 = ~n9953 & ~n9971;
  assign n9973 = ~pi131 & n811;
  assign n9974 = ~n9934 & n9949;
  assign n9975 = ~n9973 & n9974;
  assign n9976 = ~pi132 & n811;
  assign n9977 = n9934 & n9969;
  assign n9978 = ~n9976 & n9977;
  assign n9979 = ~n9975 & ~n9978;
  assign n9980 = n9934 & n9947;
  assign n9981 = pi132 & n811;
  assign n9982 = n9980 & ~n9981;
  assign n9983 = pi131 & n811;
  assign n9984 = ~n9934 & n9952;
  assign n9985 = ~n9983 & n9984;
  assign n9986 = ~n9982 & ~n9985;
  assign n9987 = n9979 & n9986;
  assign n9988 = n9972 & n9987;
  assign n9989 = n9951 & n9988;
  assign n9990 = n787 & ~n9989;
  assign n9991 = ~pi300 & n2787;
  assign n9992 = pi291 & ~pi297;
  assign n9993 = ~n9991 & ~n9992;
  assign n9994 = pi291 & pi302;
  assign n9995 = ~pi298 & pi300;
  assign n9996 = ~n9994 & ~n9995;
  assign n9997 = n9993 & n9996;
  assign n9998 = ~n832 & n9997;
  assign n9999 = ~n2114 & n9998;
  assign n10000 = ~n1558 & n9999;
  assign n10001 = ~n2087 & n10000;
  assign n10002 = ~n2091 & n10001;
  assign n10003 = pi301 & ~n10002;
  assign n10004 = ~n9990 & ~n10003;
  assign n10005 = n813 & n2339;
  assign n10006 = pi297 & n10005;
  assign n10007 = n2109 & ~n10006;
  assign n10008 = n10004 & ~n10007;
  assign n10009 = ~pi247 & ~n10008;
  assign n10010 = pi247 & pi307;
  assign n10011 = ~n10009 & ~n10010;
  assign po352 = pi359 & ~n10011;
  assign n10013 = pi308 & n8454;
  assign n10014 = pi291 & ~n1358;
  assign n10015 = n3322 & ~n10014;
  assign n10016 = n883 & n10015;
  assign n10017 = ~pi291 & pi300;
  assign n10018 = n2130 & n10017;
  assign n10019 = ~n10016 & ~n10018;
  assign n10020 = n9473 & ~n10019;
  assign n10021 = n2218 & n7131;
  assign n10022 = ~pi297 & ~pi302;
  assign n10023 = n10021 & n10022;
  assign n10024 = ~pi291 & ~pi296;
  assign n10025 = n5626 & n10024;
  assign n10026 = ~n10023 & ~n10025;
  assign n10027 = n9970 & ~n10026;
  assign n10028 = n2788 & n9970;
  assign n10029 = n852 & n10028;
  assign n10030 = n1559 & n10029;
  assign n10031 = ~n10027 & ~n10030;
  assign n10032 = n787 & ~n10031;
  assign n10033 = ~n2714 & n9950;
  assign n10034 = n787 & n10033;
  assign n10035 = n2636 & n9948;
  assign n10036 = n787 & n10035;
  assign n10037 = ~n10034 & ~n10036;
  assign n10038 = ~n10032 & n10037;
  assign n10039 = ~pi247 & ~n10038;
  assign n10040 = ~n10020 & ~n10039;
  assign n10041 = pi359 & ~n10040;
  assign po353 = n10013 | n10041;
  assign n10043 = ~n7331 & n7381;
  assign n10044 = n2977 & n10043;
  assign n10045 = ~pi247 & n10044;
  assign n10046 = pi247 & pi309;
  assign n10047 = ~n10045 & ~n10046;
  assign po354 = n8594 | ~n10047;
  assign n10049 = ~pi296 & n2109;
  assign n10050 = n2792 & n10049;
  assign n10051 = pi196 & n9948;
  assign n10052 = n2714 & n9950;
  assign n10053 = ~n10051 & ~n10052;
  assign n10054 = ~n9974 & ~n9977;
  assign n10055 = ~n9984 & n10054;
  assign n10056 = pi291 & ~n9965;
  assign n10057 = ~pi298 & n2091;
  assign n10058 = ~n10056 & ~n10057;
  assign n10059 = pi297 & ~n10058;
  assign n10060 = ~n9959 & ~n10059;
  assign n10061 = ~n1558 & n10060;
  assign n10062 = ~pi296 & ~n10061;
  assign n10063 = n1558 & n2792;
  assign n10064 = pi297 & n9900;
  assign n10065 = ~n10063 & ~n10064;
  assign n10066 = n850 & n3322;
  assign n10067 = ~pi291 & n10066;
  assign n10068 = ~pi303 & n7131;
  assign n10069 = ~n10067 & ~n10068;
  assign n10070 = n870 & n2091;
  assign n10071 = ~n10066 & ~n10070;
  assign n10072 = pi296 & ~n10071;
  assign n10073 = n10069 & ~n10072;
  assign n10074 = pi302 & n2091;
  assign n10075 = ~n7132 & ~n10074;
  assign n10076 = n870 & ~n10075;
  assign n10077 = ~pi303 & n7137;
  assign n10078 = ~n10076 & ~n10077;
  assign n10079 = ~pi297 & ~pi300;
  assign n10080 = n850 & n10079;
  assign n10081 = n10078 & ~n10080;
  assign n10082 = n10073 & n10081;
  assign n10083 = n10065 & n10082;
  assign n10084 = ~n10062 & n10083;
  assign n10085 = n9970 & ~n10084;
  assign n10086 = ~n2767 & n9953;
  assign n10087 = ~n10085 & ~n10086;
  assign n10088 = n10055 & n10087;
  assign n10089 = ~n9980 & n10088;
  assign n10090 = n10053 & n10089;
  assign n10091 = n787 & ~n10090;
  assign n10092 = ~n10050 & ~n10091;
  assign n10093 = pi301 & n789;
  assign n10094 = n3322 & n10093;
  assign n10095 = n8495 & n10024;
  assign n10096 = ~n10094 & ~n10095;
  assign n10097 = n10092 & n10096;
  assign n10098 = ~pi247 & ~n10097;
  assign n10099 = pi247 & pi310;
  assign n10100 = ~n10098 & ~n10099;
  assign po355 = pi359 & ~n10100;
  assign n10102 = pi247 & pi311;
  assign n10103 = pi314 & n10044;
  assign n10104 = pi304 & ~n10044;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = ~pi247 & ~n10105;
  assign po356 = n10102 | n10106;
  assign n10108 = pi247 & pi312;
  assign n10109 = ~n8629 & ~n10108;
  assign po357 = n10045 | ~n10109;
  assign n10111 = pi313 & ~n9601;
  assign n10112 = ~pi298 & n9743;
  assign n10113 = ~n7149 & n10112;
  assign n10114 = pi313 & ~n9743;
  assign n10115 = n9916 & n10114;
  assign n10116 = ~n10113 & ~n10115;
  assign n10117 = n9601 & ~n10116;
  assign n10118 = ~n10111 & ~n10117;
  assign n10119 = ~pi247 & ~n10118;
  assign n10120 = pi247 & pi313;
  assign n10121 = ~n10119 & ~n10120;
  assign po358 = pi359 & ~n10121;
  assign n10123 = pi314 & ~n9601;
  assign n10124 = pi298 & n9914;
  assign n10125 = pi314 & ~n9743;
  assign n10126 = n9916 & n10125;
  assign n10127 = ~n10124 & ~n10126;
  assign n10128 = n9601 & ~n10127;
  assign n10129 = ~n10123 & ~n10128;
  assign n10130 = ~pi247 & ~n10129;
  assign n10131 = pi247 & pi314;
  assign n10132 = ~n10130 & ~n10131;
  assign po359 = pi359 & ~n10132;
  assign n10134 = ~pi181 & n5247;
  assign n10135 = pi315 & ~n5247;
  assign n10136 = ~n10134 & ~n10135;
  assign n10137 = n7824 & ~n10136;
  assign n10138 = pi315 & ~n7824;
  assign n10139 = ~n10137 & ~n10138;
  assign po360 = ~pi359 | ~n10139;
  assign n10141 = pi138 & n5247;
  assign n10142 = pi316 & ~n5247;
  assign n10143 = ~n10141 & ~n10142;
  assign n10144 = n7824 & ~n10143;
  assign n10145 = pi316 & ~n7824;
  assign n10146 = ~n10144 & ~n10145;
  assign po361 = ~pi359 | ~n10146;
  assign n10148 = pi139 & n5247;
  assign n10149 = pi317 & ~n5247;
  assign n10150 = ~n10148 & ~n10149;
  assign n10151 = n7824 & ~n10150;
  assign n10152 = pi317 & ~n7824;
  assign n10153 = ~n10151 & ~n10152;
  assign po362 = ~pi359 | ~n10153;
  assign n10155 = pi178 & n5247;
  assign n10156 = pi318 & ~n5247;
  assign n10157 = ~n10155 & ~n10156;
  assign n10158 = n7824 & ~n10157;
  assign n10159 = pi318 & ~n7824;
  assign n10160 = ~n10158 & ~n10159;
  assign po363 = ~pi359 | ~n10160;
  assign n10162 = pi142 & n5247;
  assign n10163 = pi319 & ~n5247;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = n7824 & ~n10164;
  assign n10166 = pi319 & ~n7824;
  assign n10167 = ~n10165 & ~n10166;
  assign po364 = ~pi359 | ~n10167;
  assign n10169 = pi129 & n5247;
  assign n10170 = pi320 & ~n5247;
  assign n10171 = ~n10169 & ~n10170;
  assign n10172 = n7824 & ~n10171;
  assign n10173 = pi320 & ~n7824;
  assign n10174 = ~n10172 & ~n10173;
  assign po365 = ~pi359 | ~n10174;
  assign n10176 = ~pi180 & n5247;
  assign n10177 = pi321 & ~n5247;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = n7824 & ~n10178;
  assign n10180 = pi321 & ~n7824;
  assign n10181 = ~n10179 & ~n10180;
  assign po366 = ~pi359 | ~n10181;
  assign n10183 = pi132 & n5247;
  assign n10184 = pi322 & ~n5247;
  assign n10185 = ~n10183 & ~n10184;
  assign n10186 = n7824 & ~n10185;
  assign n10187 = pi322 & ~n7824;
  assign n10188 = ~n10186 & ~n10187;
  assign po367 = ~pi359 | ~n10188;
  assign n10190 = pi102 & n5247;
  assign n10191 = pi323 & ~n5247;
  assign n10192 = ~n10190 & ~n10191;
  assign n10193 = n7824 & ~n10192;
  assign n10194 = pi323 & ~n7824;
  assign n10195 = ~n10193 & ~n10194;
  assign po368 = ~pi359 | ~n10195;
  assign n10197 = pi184 & n5247;
  assign n10198 = pi324 & ~n5247;
  assign n10199 = ~n10197 & ~n10198;
  assign n10200 = n7824 & ~n10199;
  assign n10201 = pi324 & ~n7824;
  assign n10202 = ~n10200 & ~n10201;
  assign po369 = ~pi359 | ~n10202;
  assign n10204 = pi131 & n5247;
  assign n10205 = pi325 & ~n5247;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = n7824 & ~n10206;
  assign n10208 = pi325 & ~n7824;
  assign n10209 = ~n10207 & ~n10208;
  assign po370 = ~pi359 | ~n10209;
  assign n10211 = pi126 & n5247;
  assign n10212 = pi326 & ~n5247;
  assign n10213 = ~n10211 & ~n10212;
  assign n10214 = n7824 & ~n10213;
  assign n10215 = pi326 & ~n7824;
  assign n10216 = ~n10214 & ~n10215;
  assign po371 = ~pi359 | ~n10216;
  assign n10218 = pi141 & n5247;
  assign n10219 = pi327 & ~n5247;
  assign n10220 = ~n10218 & ~n10219;
  assign n10221 = n7824 & ~n10220;
  assign n10222 = pi327 & ~n7824;
  assign n10223 = ~n10221 & ~n10222;
  assign po372 = ~pi359 | ~n10223;
  assign n10225 = pi143 & n5247;
  assign n10226 = pi328 & ~n5247;
  assign n10227 = ~n10225 & ~n10226;
  assign n10228 = n7824 & ~n10227;
  assign n10229 = pi328 & ~n7824;
  assign n10230 = ~n10228 & ~n10229;
  assign po373 = ~pi359 | ~n10230;
  assign n10232 = pi140 & n5247;
  assign n10233 = pi329 & ~n5247;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = n7824 & ~n10234;
  assign n10236 = pi329 & ~n7824;
  assign n10237 = ~n10235 & ~n10236;
  assign po374 = ~pi359 | ~n10237;
  assign n10239 = pi133 & n5247;
  assign n10240 = pi330 & ~n5247;
  assign n10241 = ~n10239 & ~n10240;
  assign n10242 = n7824 & ~n10241;
  assign n10243 = pi330 & ~n7824;
  assign n10244 = ~n10242 & ~n10243;
  assign po375 = ~pi359 | ~n10244;
  assign n10246 = ~n844 & n3322;
  assign n10247 = n2793 & n10246;
  assign n10248 = pi301 & ~n10247;
  assign n10249 = ~n787 & ~n10248;
  assign n10250 = ~n2109 & n10249;
  assign n10251 = n2792 & n3322;
  assign n10252 = ~pi296 & n849;
  assign n10253 = pi296 & ~n849;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = n10251 & n10254;
  assign n10256 = ~n859 & n10255;
  assign n10257 = ~n1372 & n10256;
  assign n10258 = pi301 & ~n10257;
  assign n10259 = ~n787 & ~n10258;
  assign n10260 = ~n2109 & n10259;
  assign n10261 = ~n10250 & ~n10260;
  assign n10262 = pi331 & n10261;
  assign n10263 = ~n10250 & ~n10261;
  assign n10264 = ~n10262 & ~n10263;
  assign n10265 = ~pi247 & ~n10264;
  assign n10266 = pi247 & pi331;
  assign n10267 = ~n10265 & ~n10266;
  assign po376 = pi359 & ~n10267;
  assign n10269 = pi133 & n9599;
  assign n10270 = pi332 & ~n9614;
  assign n10271 = ~n10269 & ~n10270;
  assign n10272 = n5258 & ~n10271;
  assign n10273 = n782 & n10272;
  assign n10274 = pi332 & ~n5259;
  assign n10275 = ~n10273 & ~n10274;
  assign n10276 = ~pi247 & ~n10275;
  assign n10277 = pi247 & pi332;
  assign n10278 = ~n10276 & ~n10277;
  assign po377 = pi359 & ~n10278;
  assign n10280 = pi333 & n10261;
  assign n10281 = ~n10260 & ~n10261;
  assign n10282 = ~n10280 & ~n10281;
  assign n10283 = ~pi247 & ~n10282;
  assign n10284 = pi247 & pi333;
  assign n10285 = ~n10283 & ~n10284;
  assign po378 = pi359 & ~n10285;
  assign n10287 = ~n783 & ~n7186;
  assign po379 = ~pi359 | n10287;
  assign n10289 = n787 & ~n8746;
  assign n10290 = pi301 & n935;
  assign n10291 = ~n10289 & ~n10290;
  assign n10292 = ~pi247 & ~n10291;
  assign n10293 = pi247 & pi335;
  assign n10294 = ~n10292 & ~n10293;
  assign po380 = pi359 & ~n10294;
  assign n10296 = pi336 & ~n5259;
  assign n10297 = pi139 & n9613;
  assign n10298 = pi336 & ~n9613;
  assign n10299 = ~n10297 & ~n10298;
  assign n10300 = n5259 & ~n10299;
  assign n10301 = ~n10296 & ~n10300;
  assign n10302 = ~pi247 & ~n10301;
  assign n10303 = pi247 & pi336;
  assign n10304 = ~n10302 & ~n10303;
  assign po381 = pi359 & ~n10304;
  assign n10306 = pi337 & ~n5259;
  assign n10307 = pi141 & n9613;
  assign n10308 = pi337 & ~n9613;
  assign n10309 = ~n10307 & ~n10308;
  assign n10310 = n5259 & ~n10309;
  assign n10311 = ~n10306 & ~n10310;
  assign n10312 = ~pi247 & ~n10311;
  assign n10313 = pi247 & pi337;
  assign n10314 = ~n10312 & ~n10313;
  assign po382 = pi359 & ~n10314;
  assign n10316 = pi338 & ~n5259;
  assign n10317 = pi143 & n9613;
  assign n10318 = pi338 & ~n9613;
  assign n10319 = ~n10317 & ~n10318;
  assign n10320 = n5259 & ~n10319;
  assign n10321 = ~n10316 & ~n10320;
  assign n10322 = ~pi247 & ~n10321;
  assign n10323 = pi247 & pi338;
  assign n10324 = ~n10322 & ~n10323;
  assign po383 = pi359 & ~n10324;
  assign n10326 = pi339 & ~n5259;
  assign n10327 = pi133 & n9613;
  assign n10328 = pi339 & ~n9613;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = n5259 & ~n10329;
  assign n10331 = ~n10326 & ~n10330;
  assign n10332 = ~pi247 & ~n10331;
  assign n10333 = pi247 & pi339;
  assign n10334 = ~n10332 & ~n10333;
  assign po384 = pi359 & ~n10334;
  assign n10336 = pi340 & ~n5259;
  assign n10337 = pi140 & n9613;
  assign n10338 = pi340 & ~n9613;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = n5259 & ~n10339;
  assign n10341 = ~n10336 & ~n10340;
  assign n10342 = ~pi247 & ~n10341;
  assign n10343 = pi247 & pi340;
  assign n10344 = ~n10342 & ~n10343;
  assign po385 = pi359 & ~n10344;
  assign n10346 = pi341 & ~n5259;
  assign n10347 = pi126 & n9613;
  assign n10348 = pi341 & ~n9613;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = n5259 & ~n10349;
  assign n10351 = ~n10346 & ~n10350;
  assign n10352 = ~pi247 & ~n10351;
  assign n10353 = pi247 & pi341;
  assign n10354 = ~n10352 & ~n10353;
  assign po386 = pi359 & ~n10354;
  assign n10356 = pi342 & ~n5259;
  assign n10357 = pi142 & n9613;
  assign n10358 = pi342 & ~n9613;
  assign n10359 = ~n10357 & ~n10358;
  assign n10360 = n5259 & ~n10359;
  assign n10361 = ~n10356 & ~n10360;
  assign n10362 = ~pi247 & ~n10361;
  assign n10363 = pi247 & pi342;
  assign n10364 = ~n10362 & ~n10363;
  assign po387 = pi359 & ~n10364;
  assign n10366 = pi343 & ~n5259;
  assign n10367 = pi138 & n9613;
  assign n10368 = pi343 & ~n9613;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = n5259 & ~n10369;
  assign n10371 = ~n10366 & ~n10370;
  assign n10372 = ~pi247 & ~n10371;
  assign n10373 = pi247 & pi343;
  assign n10374 = ~n10372 & ~n10373;
  assign po388 = pi359 & ~n10374;
  assign n10376 = n7299 & n8740;
  assign n10377 = n787 & n10376;
  assign n10378 = pi344 & n8454;
  assign po389 = n10377 | n10378;
  assign n10380 = ~pi131 & pi302;
  assign n10381 = n8444 & ~n10380;
  assign n10382 = pi102 & pi302;
  assign n10383 = ~pi131 & n10382;
  assign n10384 = n5095 & ~n10383;
  assign n10385 = n5094 & ~n10382;
  assign n10386 = ~n10384 & ~n10385;
  assign n10387 = ~n10381 & n10386;
  assign po390 = pi359 & ~n10387;
  assign n10389 = pi247 & pi346;
  assign n10390 = pi304 & n9468;
  assign n10391 = pi314 & ~n9468;
  assign n10392 = ~n10390 & ~n10391;
  assign n10393 = ~pi247 & ~n10392;
  assign po391 = n10389 | n10393;
  assign n10395 = pi347 & ~n2071;
  assign n10396 = ~n9829 & ~n10395;
  assign po392 = pi359 & ~n10396;
  assign n10398 = pi348 & ~n2071;
  assign n10399 = ~n9888 & ~n10398;
  assign po393 = pi359 & ~n10399;
  assign n10401 = pi349 & ~n2071;
  assign n10402 = ~n9799 & ~n10401;
  assign po394 = pi359 & ~n10402;
  assign n10404 = pi350 & ~n2071;
  assign n10405 = ~n9844 & ~n10404;
  assign po395 = pi359 & ~n10405;
  assign n10407 = pi351 & ~n2071;
  assign n10408 = ~n9709 & ~n10407;
  assign po396 = pi359 & ~n10408;
  assign n10410 = pi352 & ~n2071;
  assign n10411 = ~n9873 & ~n10410;
  assign po397 = pi359 & ~n10411;
  assign n10413 = pi353 & ~n2071;
  assign n10414 = ~n9814 & ~n10413;
  assign po398 = pi359 & ~n10414;
  assign n10416 = pi354 & ~n2071;
  assign n10417 = ~n9784 & ~n10416;
  assign po399 = pi359 & ~n10417;
  assign n10419 = pi357 & ~pi363;
  assign n10420 = ~pi355 & ~n10419;
  assign n10421 = ~pi196 & ~n10420;
  assign po400 = pi359 & n10421;
  assign po401 = pi359 & ~pi364;
  assign po402 = pi359 & pi363;
  assign po403 = pi359 & ~pi362;
  assign po032 = 1'b1;
  assign po007 = ~pi247;
  assign po000 = pi194;
  assign po001 = pi281;
  assign po002 = pi279;
  assign po003 = pi293;
  assign po004 = pi306;
  assign po005 = pi334;
  assign po006 = pi230;
  assign po008 = pi035;
  assign po009 = pi001;
  assign po010 = pi002;
  assign po011 = pi036;
  assign po012 = pi034;
  assign po013 = pi003;
  assign po014 = pi004;
  assign po015 = pi039;
  assign po016 = pi038;
  assign po017 = pi040;
  assign po018 = pi033;
  assign po019 = pi029;
  assign po020 = pi030;
  assign po021 = pi031;
  assign po022 = pi032;
  assign po023 = pi037;
  assign po024 = pi161;
  assign po025 = pi162;
  assign po026 = pi163;
  assign po027 = pi164;
  assign po028 = pi145;
  assign po029 = pi128;
  assign po030 = pi136;
  assign po031 = pi134;
  assign po033 = pi360;
  assign po035 = pi247;
  assign po036 = pi000;
  assign po077 = pi041;
  assign po080 = pi042;
  assign po082 = pi043;
  assign po084 = pi044;
  assign po086 = pi045;
  assign po088 = pi046;
  assign po090 = pi047;
  assign po092 = pi048;
endmodule


