module ac97_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205,
    pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214,
    pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223,
    pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232,
    pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241,
    pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250,
    pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259,
    pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268,
    pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277,
    pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286,
    pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295,
    pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304,
    pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313,
    pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322,
    pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331,
    pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340,
    pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349,
    pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358,
    pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367,
    pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376,
    pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385,
    pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394,
    pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403,
    pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412,
    pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421,
    pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430,
    pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439,
    pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448,
    pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457,
    pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466,
    pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475,
    pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484,
    pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493,
    pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502,
    pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511,
    pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520,
    pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529,
    pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538,
    pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547,
    pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556,
    pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565,
    pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574,
    pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583,
    pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592,
    pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601,
    pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610,
    pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619,
    pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628,
    pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637,
    pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646,
    pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655,
    pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664,
    pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673,
    pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682,
    pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691,
    pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700,
    pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709,
    pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718,
    pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727,
    pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736,
    pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745,
    pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754,
    pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763,
    pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772,
    pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781,
    pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790,
    pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799,
    pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808,
    pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817,
    pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826,
    pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835,
    pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844,
    pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853,
    pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862,
    pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871,
    pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880,
    pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889,
    pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898,
    pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907,
    pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916,
    pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925,
    pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934,
    pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943,
    pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952,
    pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961,
    pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970,
    pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979,
    pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988,
    pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997,
    pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006,
    pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015,
    pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024,
    pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033,
    pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042,
    pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051,
    pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060,
    pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069,
    pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078,
    pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087,
    pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096,
    pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105,
    pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114,
    pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123,
    pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132,
    pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141,
    pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150,
    pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159,
    pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168,
    pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177,
    pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186,
    pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195,
    pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204,
    pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213,
    pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222,
    pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231,
    pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240,
    pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249,
    pi2250, pi2251, pi2252, pi2253, pi2254,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511,
    po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520,
    po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529,
    po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538,
    po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547,
    po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556,
    po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565,
    po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574,
    po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583,
    po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592,
    po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601,
    po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610,
    po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619,
    po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628,
    po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637,
    po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646,
    po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655,
    po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664,
    po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673,
    po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682,
    po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691,
    po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700,
    po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709,
    po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718,
    po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727,
    po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736,
    po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745,
    po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754,
    po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763,
    po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772,
    po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781,
    po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790,
    po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799,
    po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808,
    po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817,
    po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826,
    po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835,
    po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844,
    po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853,
    po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862,
    po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871,
    po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880,
    po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889,
    po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898,
    po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907,
    po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916,
    po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925,
    po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934,
    po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943,
    po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952,
    po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961,
    po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970,
    po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979,
    po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988,
    po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997,
    po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006,
    po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015,
    po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024,
    po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033,
    po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042,
    po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051,
    po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060,
    po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069,
    po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078,
    po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087,
    po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096,
    po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105,
    po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114,
    po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123,
    po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132,
    po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141,
    po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150,
    po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159,
    po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168,
    po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177,
    po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186,
    po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195,
    po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204,
    po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213,
    po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222,
    po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231,
    po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240,
    po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204,
    pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213,
    pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222,
    pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231,
    pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240,
    pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249,
    pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258,
    pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267,
    pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276,
    pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285,
    pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294,
    pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303,
    pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312,
    pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321,
    pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330,
    pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339,
    pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348,
    pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357,
    pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366,
    pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375,
    pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384,
    pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393,
    pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402,
    pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411,
    pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420,
    pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429,
    pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438,
    pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447,
    pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456,
    pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465,
    pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474,
    pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483,
    pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492,
    pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501,
    pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510,
    pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519,
    pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528,
    pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537,
    pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546,
    pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555,
    pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564,
    pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573,
    pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582,
    pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591,
    pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600,
    pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609,
    pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618,
    pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627,
    pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636,
    pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645,
    pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654,
    pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663,
    pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672,
    pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681,
    pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690,
    pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699,
    pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708,
    pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717,
    pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726,
    pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735,
    pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744,
    pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753,
    pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762,
    pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771,
    pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780,
    pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789,
    pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798,
    pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807,
    pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816,
    pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825,
    pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834,
    pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843,
    pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852,
    pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861,
    pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870,
    pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879,
    pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888,
    pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897,
    pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906,
    pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915,
    pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924,
    pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933,
    pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942,
    pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951,
    pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960,
    pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969,
    pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978,
    pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987,
    pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996,
    pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005,
    pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014,
    pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023,
    pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032,
    pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041,
    pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050,
    pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059,
    pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068,
    pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077,
    pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086,
    pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095,
    pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104,
    pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113,
    pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122,
    pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131,
    pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140,
    pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149,
    pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158,
    pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167,
    pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176,
    pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185,
    pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194,
    pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203,
    pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212,
    pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221,
    pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230,
    pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239,
    pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248,
    pi2249, pi2250, pi2251, pi2252, pi2253, pi2254;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510,
    po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519,
    po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528,
    po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537,
    po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546,
    po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555,
    po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564,
    po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573,
    po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582,
    po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591,
    po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600,
    po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609,
    po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618,
    po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627,
    po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636,
    po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645,
    po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654,
    po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663,
    po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672,
    po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681,
    po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690,
    po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699,
    po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708,
    po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717,
    po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726,
    po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735,
    po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744,
    po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753,
    po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762,
    po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771,
    po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780,
    po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789,
    po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798,
    po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807,
    po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816,
    po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825,
    po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834,
    po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843,
    po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852,
    po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861,
    po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870,
    po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879,
    po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888,
    po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897,
    po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906,
    po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915,
    po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924,
    po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933,
    po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942,
    po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951,
    po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960,
    po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969,
    po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978,
    po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987,
    po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996,
    po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005,
    po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014,
    po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023,
    po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032,
    po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041,
    po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050,
    po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059,
    po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068,
    po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077,
    po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086,
    po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095,
    po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104,
    po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113,
    po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122,
    po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131,
    po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140,
    po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149,
    po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158,
    po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167,
    po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176,
    po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185,
    po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194,
    po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203,
    po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212,
    po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221,
    po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230,
    po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239,
    po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248,
    po2249;
  wire n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4520, n4521, n4523, n4524, n4526, n4527, n4529, n4530, n4533,
    n4534, n4536, n4537, n4539, n4540, n4542, n4550, n4551, n4553, n4554,
    n4556, n4557, n4559, n4560, n4562, n4563, n4565, n4566, n4568, n4569,
    n4571, n4572, n4586, n4587, n4589, n4590, n4592, n4593, n4595, n4596,
    n4598, n4599, n4601, n4602, n4604, n4605, n4607, n4608, n4610, n4611,
    n4613, n4614, n4616, n4617, n4619, n4620, n4622, n4623, n4625, n4626,
    n4628, n4629, n4631, n4632, n4638, n4639, n4641, n4642, n4644, n4645,
    n4647, n4648, n4650, n4651, n4653, n4654, n4656, n4657, n4659, n4660,
    n4662, n4663, n4665, n4666, n4668, n4669, n4671, n4672, n4674, n4675,
    n4677, n4678, n4680, n4681, n4683, n4684, n4686, n4687, n4689, n4690,
    n4692, n4693, n4695, n4696, n4698, n4699, n4701, n4702, n4704, n4705,
    n4707, n4708, n4710, n4711, n4713, n4714, n4716, n4717, n4719, n4720,
    n4722, n4723, n4725, n4726, n4728, n4729, n4731, n4732, n4734, n4735,
    n4737, n4738, n4740, n4741, n4743, n4744, n4746, n4747, n4749, n4750,
    n4752, n4753, n4755, n4756, n4778, n4779, n4781, n4782, n4784, n4785,
    n4787, n4788, n4790, n4791, n4793, n4794, n4796, n4797, n4799, n4800,
    n4802, n4803, n4805, n4806, n4808, n4809, n4811, n4812, n4814, n4815,
    n4817, n4818, n4820, n4821, n4823, n4824, n4826, n4827, n4829, n4830,
    n4832, n4833, n4835, n4836, n4838, n4839, n4841, n4842, n4844, n4845,
    n4847, n4848, n4850, n4851, n4853, n4854, n4856, n4857, n4859, n4860,
    n4862, n4863, n4865, n4866, n4868, n4869, n4871, n4872, n4874, n4875,
    n4877, n4878, n4880, n4881, n4883, n4884, n4886, n4887, n4889, n4890,
    n4892, n4893, n4895, n4896, n4898, n4899, n4901, n4902, n4904, n4905,
    n4907, n4908, n4910, n4911, n4913, n4914, n4916, n4917, n4919, n4920,
    n4922, n4923, n4925, n4926, n4928, n4929, n4931, n4932, n4934, n4935,
    n4937, n4938, n4940, n4941, n4943, n4944, n4946, n4947, n4949, n4950,
    n4952, n4953, n4955, n4956, n4958, n4959, n4961, n4962, n4964, n4965,
    n4967, n4968, n4970, n4971, n4973, n4974, n4976, n4977, n4979, n4980,
    n4982, n4983, n4985, n4986, n4988, n4989, n4991, n4992, n4994, n4995,
    n4997, n4998, n5000, n5001, n5003, n5004, n5006, n5007, n5009, n5010,
    n5012, n5013, n5015, n5016, n5018, n5019, n5021, n5022, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5045, n5046,
    n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
    n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
    n5069, n5070, n5072, n5073, n5075, n5076, n5077, n5078, n5079, n5080,
    n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5096, n5097, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
    n5113, n5114, n5115, n5116, n5117, n5118, n5120, n5121, n5123, n5124,
    n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
    n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5144, n5145,
    n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
    n5168, n5169, n5171, n5172, n5174, n5175, n5177, n5178, n5180, n5181,
    n5183, n5184, n5186, n5187, n5189, n5190, n5192, n5193, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
    n5208, n5209, n5210, n5211, n5212, n5215, n5216, n5217, n5218, n5219,
    n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
    n5318, n5319, n5320, n5321, n5322, n5323, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
    n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5393,
    n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5427, n5429, n5430, n5432, n5433, n5435, n5436, n5438, n5439, n5441,
    n5442, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
    n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5480, n5481, n5482, n5483, n5484, n5485,
    n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
    n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5567, n5568, n5569,
    n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5588, n5589, n5590,
    n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
    n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5679, n5681, n5683, n5685, n5687, n5688,
    n5689, n5690, n5691, n5693, n5694, n5696, n5697, n5698, n5699, n5700,
    n5702, n5703, n5705, n5706, n5707, n5708, n5709, n5711, n5712, n5713,
    n5714, n5715, n5717, n5718, n5720, n5721, n5723, n5724, n5725, n5727,
    n5728, n5729, n5731, n5732, n5733, n5735, n5736, n5737, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
    n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
    n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
    n5843, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
    n5864, n5865, n5866, n5867, n5868, n5869, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
    n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5956, n5957,
    n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
    n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
    n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
    n6020, n6021, n6022, n6023, n6024, n6025, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
    n6041, n6042, n6043, n6044, n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
    n6062, n6063, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
    n6084, n6085, n6086, n6087, n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
    n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
    n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
    n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6286, n6287, n6288, n6289, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
    n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6315, n6316, n6317, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6338, n6339, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6364,
    n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6390, n6391, n6392, n6393, n6394, n6395,
    n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6435, n6436, n6437,
    n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
    n6448, n6449, n6450, n6451, n6452, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
    n6491, n6492, n6493, n6494, n6495, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
    n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
    n6677, n6678, n6679, n6680, n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
    n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6708,
    n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
    n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
    n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
    n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6759, n6760,
    n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
    n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
    n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
    n6822, n6823, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
    n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7008, n7009,
    n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
    n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7072,
    n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
    n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
    n7146, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
    n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
    n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
    n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7293, n7294,
    n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
    n7316, n7317, n7318, n7320, n7321, n7323, n7324, n7326, n7327, n7329,
    n7330, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7356, n7357, n7358, n7359, n7360, n7361,
    n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7402, n7403,
    n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
    n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
    n7488, n7489, n7490, n7491, n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7517, n7518, n7519,
    n7520, n7521, n7523, n7524, n7526, n7527, n7528, n7529, n7530, n7532,
    n7533, n7535, n7536, n7537, n7539, n7540, n7541, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7565, n7566, n7567,
    n7568, n7569, n7570, n7572, n7573, n7574, n7575, n7576, n7578, n7579,
    n7580, n7581, n7582, n7583, n7585, n7586, n7587, n7588, n7589, n7590,
    n7592, n7593, n7594, n7595, n7596, n7597, n7599, n7600, n7601, n7602,
    n7603, n7604, n7606, n7607, n7608, n7609, n7610, n7611, n7613, n7614,
    n7615, n7616, n7617, n7618, n7620, n7621, n7622, n7623, n7624, n7625,
    n7627, n7628, n7629, n7630, n7631, n7632, n7634, n7635, n7636, n7637,
    n7638, n7639, n7641, n7642, n7643, n7644, n7645, n7646, n7648, n7649,
    n7650, n7651, n7652, n7653, n7655, n7656, n7657, n7658, n7659, n7660,
    n7662, n7663, n7664, n7665, n7666, n7667, n7669, n7670, n7671, n7672,
    n7673, n7675, n7676, n7677, n7678, n7679, n7681, n7682, n7683, n7684,
    n7685, n7687, n7688, n7689, n7690, n7691, n7693, n7694, n7695, n7696,
    n7697, n7699, n7700, n7701, n7702, n7703, n7705, n7706, n7707, n7708,
    n7709, n7711, n7712, n7713, n7714, n7715, n7717, n7718, n7719, n7720,
    n7721, n7723, n7724, n7725, n7726, n7727, n7729, n7730, n7731, n7732,
    n7733, n7735, n7736, n7737, n7738, n7739, n7741, n7742, n7743, n7744,
    n7745, n7747, n7748, n7749, n7750, n7751, n7753, n7754, n7755, n7756,
    n7757, n7759, n7760, n7761, n7762, n7763, n7765, n7766, n7767, n7768,
    n7769, n7771, n7772, n7773, n7774, n7775, n7777, n7778, n7779, n7780,
    n7781, n7783, n7784, n7785, n7786, n7787, n7789, n7790, n7791, n7792,
    n7793, n7795, n7796, n7797, n7798, n7799, n7801, n7802, n7803, n7804,
    n7805, n7807, n7808, n7809, n7810, n7811, n7813, n7814, n7815, n7816,
    n7817, n7819, n7820, n7821, n7822, n7823, n7825, n7826, n7827, n7828,
    n7829, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
    n7862, n7863, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
    n7884, n7885, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7898, n7899, n7900, n7901, n7902, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7915, n7916, n7917,
    n7918, n7919, n7921, n7922, n7923, n7924, n7925, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7949, n7950, n7951,
    n7952, n7953, n7954, n7955, n7956, n7957, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968, n7970, n7971, n7972, n7973,
    n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
    n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
    n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
    n8004, n8005, n8006, n8007, n8008, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
    n8076, n8077, n8078, n8079, n8080, n8081, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8154, n8155, n8156, n8157, n8158, n8159,
    n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
    n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8199, n8200, n8201,
    n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
    n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8232,
    n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8282, n8283, n8284, n8285,
    n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
    n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
    n8410, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
    n8462, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
    n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
    n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
    n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
    n8576, n8577, n8578, n8579, n8580, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
    n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
    n8618, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8692, n8693,
    n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8703, n8704,
    n8705, n8706, n8707, n8709, n8710, n8711, n8712, n8713, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8737, n8738,
    n8739, n8740, n8741, n8743, n8744, n8745, n8746, n8748, n8750, n8752,
    n8754, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
    n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
    n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8806, n8807,
    n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8830,
    n8831, n8832, n8833, n8834, n8835, n8837, n8838, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848, n8850, n8851, n8852, n8853,
    n8854, n8855, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870, n8872, n8873, n8874, n8875,
    n8876, n8877, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8887,
    n8888, n8889, n8890, n8891, n8892, n8894, n8895, n8896, n8897, n8898,
    n8899, n8901, n8902, n8903, n8904, n8905, n8906, n8908, n8909, n8910,
    n8911, n8912, n8913, n8915, n8916, n8917, n8918, n8919, n8921, n8922,
    n8923, n8924, n8925, n8926, n8928, n8929, n8930, n8931, n8932, n8934,
    n8935, n8936, n8937, n8938, n8940, n8941, n8942, n8943, n8944, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
    n8957, n8959, n8960, n8961, n8962, n8963, n8965, n8966, n8967, n8968,
    n8969, n8971, n8972, n8974, n8975, n8977, n8978, n8980, n8981, n8983,
    n8984, n8985, n8986, n8987, n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8998, n8999, n9000, n9001, n9002, n9003, n9005, n9006,
    n9007, n9008, n9009, n9010, n9012, n9013, n9014, n9015, n9016, n9017,
    n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
    n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9039, n9040,
    n9041, n9042, n9043, n9044, n9046, n9047, n9048, n9049, n9050, n9051,
    n9053, n9054, n9055, n9056, n9057, n9058, n9060, n9061, n9062, n9063,
    n9064, n9065, n9067, n9068, n9069, n9070, n9071, n9073, n9074, n9075,
    n9076, n9077, n9079, n9080, n9081, n9082, n9083, n9085, n9086, n9087,
    n9088, n9089, n9090, n9092, n9093, n9094, n9095, n9096, n9098, n9099,
    n9100, n9101, n9102, n9103, n9105, n9106, n9107, n9108, n9109, n9111,
    n9112, n9113, n9114, n9115, n9117, n9118, n9119, n9120, n9121, n9122,
    n9124, n9125, n9126, n9127, n9128, n9129, n9131, n9132, n9133, n9134,
    n9135, n9136, n9138, n9139, n9140, n9141, n9142, n9144, n9145, n9146,
    n9147, n9148, n9149, n9151, n9152, n9153, n9154, n9155, n9156, n9158,
    n9159, n9160, n9161, n9162, n9164, n9165, n9166, n9167, n9168, n9170,
    n9171, n9172, n9173, n9174, n9175, n9177, n9178, n9179, n9180, n9181,
    n9183, n9184, n9185, n9186, n9187, n9189, n9190, n9191, n9192, n9193,
    n9195, n9196, n9197, n9198, n9199, n9201, n9202, n9203, n9204, n9205,
    n9207, n9208, n9209, n9210, n9211, n9213, n9214, n9215, n9216, n9217,
    n9219, n9220, n9221, n9222, n9223, n9225, n9226, n9227, n9228, n9229,
    n9231, n9232, n9233, n9234, n9235, n9237, n9238, n9239, n9240, n9241,
    n9243, n9244, n9245, n9246, n9247, n9249, n9250, n9251, n9252, n9253,
    n9255, n9256, n9257, n9258, n9259, n9261, n9262, n9263, n9264, n9265,
    n9267, n9268, n9269, n9270, n9271, n9273, n9274, n9275, n9276, n9277,
    n9279, n9280, n9281, n9282, n9283, n9285, n9286, n9287, n9288, n9289,
    n9291, n9292, n9293, n9294, n9295, n9297, n9298, n9299, n9300, n9301,
    n9303, n9304, n9305, n9306, n9307, n9309, n9310, n9311, n9312, n9313,
    n9315, n9316, n9317, n9318, n9319, n9321, n9322, n9323, n9324, n9325,
    n9327, n9328, n9329, n9330, n9331, n9333, n9334, n9335, n9336, n9337,
    n9339, n9340, n9341, n9342, n9343, n9345, n9346, n9347, n9348, n9349,
    n9351, n9352, n9353, n9354, n9355, n9357, n9358, n9359, n9360, n9361,
    n9363, n9364, n9365, n9366, n9367, n9369, n9370, n9371, n9372, n9373,
    n9375, n9376, n9377, n9378, n9379, n9381, n9382, n9383, n9384, n9385,
    n9387, n9388, n9389, n9390, n9391, n9393, n9394, n9395, n9396, n9397,
    n9399, n9400, n9401, n9402, n9403, n9405, n9406, n9407, n9408, n9409,
    n9411, n9412, n9413, n9414, n9415, n9417, n9418, n9419, n9420, n9421,
    n9423, n9424, n9425, n9426, n9427, n9429, n9430, n9431, n9432, n9433,
    n9435, n9436, n9437, n9438, n9439, n9441, n9442, n9443, n9444, n9445,
    n9447, n9448, n9449, n9450, n9451, n9453, n9454, n9455, n9456, n9457,
    n9459, n9460, n9461, n9462, n9463, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9498, n9499, n9500, n9501, n9502,
    n9503, n9504, n9505, n9506, n9507, n9509, n9510, n9511, n9512, n9513,
    n9514, n9515, n9516, n9517, n9518, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9531, n9532, n9533, n9534, n9535,
    n9537, n9538, n9539, n9540, n9541, n9543, n9544, n9545, n9546, n9547,
    n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
    n9560, n9561, n9562, n9563, n9564, n9566, n9567, n9568, n9569, n9570,
    n9572, n9573, n9574, n9575, n9576, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9600, n9601, n9602, n9603, n9604,
    n9605, n9606, n9607, n9608, n9609, n9611, n9612, n9613, n9614, n9615,
    n9617, n9618, n9619, n9620, n9621, n9623, n9624, n9625, n9626, n9627,
    n9629, n9630, n9631, n9632, n9633, n9635, n9636, n9637, n9638, n9639,
    n9641, n9642, n9643, n9644, n9645, n9647, n9648, n9649, n9650, n9651,
    n9653, n9654, n9655, n9656, n9657, n9659, n9660, n9661, n9662, n9663,
    n9665, n9666, n9667, n9668, n9669, n9671, n9672, n9673, n9674, n9675,
    n9677, n9678, n9679, n9680, n9681, n9683, n9684, n9685, n9686, n9687,
    n9689, n9690, n9691, n9692, n9693, n9695, n9696, n9697, n9698, n9699,
    n9701, n9702, n9703, n9704, n9705, n9707, n9708, n9709, n9710, n9711,
    n9713, n9714, n9715, n9716, n9717, n9719, n9720, n9721, n9722, n9723,
    n9725, n9726, n9727, n9728, n9729, n9731, n9732, n9733, n9734, n9735,
    n9737, n9738, n9739, n9740, n9741, n9743, n9744, n9745, n9746, n9747,
    n9749, n9750, n9751, n9752, n9753, n9755, n9756, n9757, n9758, n9759,
    n9761, n9762, n9763, n9764, n9765, n9767, n9768, n9769, n9770, n9771,
    n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9783,
    n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9794,
    n9795, n9796, n9797, n9798, n9800, n9801, n9802, n9803, n9804, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9828,
    n9829, n9830, n9831, n9832, n9834, n9835, n9836, n9837, n9838, n9840,
    n9841, n9842, n9843, n9844, n9846, n9847, n9848, n9849, n9850, n9852,
    n9853, n9854, n9855, n9856, n9858, n9859, n9860, n9861, n9862, n9864,
    n9865, n9866, n9867, n9868, n9870, n9871, n9872, n9873, n9874, n9876,
    n9877, n9878, n9879, n9880, n9882, n9883, n9884, n9885, n9886, n9888,
    n9889, n9890, n9891, n9892, n9894, n9895, n9896, n9897, n9898, n9900,
    n9901, n9902, n9903, n9904, n9906, n9907, n9908, n9909, n9910, n9912,
    n9913, n9914, n9915, n9916, n9918, n9919, n9920, n9921, n9922, n9924,
    n9925, n9926, n9927, n9928, n9930, n9931, n9932, n9933, n9934, n9936,
    n9937, n9938, n9939, n9940, n9942, n9943, n9944, n9945, n9946, n9948,
    n9949, n9950, n9951, n9952, n9954, n9955, n9956, n9957, n9958, n9960,
    n9961, n9962, n9963, n9964, n9966, n9967, n9968, n9969, n9970, n9972,
    n9973, n9974, n9975, n9976, n9978, n9979, n9980, n9981, n9982, n9984,
    n9985, n9986, n9987, n9988, n9990, n9991, n9992, n9993, n9994, n9996,
    n9997, n9998, n9999, n10000, n10001, n10003, n10005, n10006, n10007,
    n10008, n10009, n10011, n10012, n10013, n10014, n10015, n10017, n10018,
    n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
    n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
    n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
    n10097, n10099, n10100, n10101, n10102, n10103, n10105, n10106, n10107,
    n10108, n10109, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10120, n10122, n10123, n10124, n10125, n10126, n10127,
    n10128, n10129, n10130, n10131, n10133, n10134, n10135, n10136, n10137,
    n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
    n10148, n10150, n10151, n10152, n10153, n10154, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10167, n10168,
    n10169, n10170, n10171, n10173, n10174, n10175, n10176, n10177, n10179,
    n10180, n10181, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10194, n10195, n10196, n10197, n10198, n10200,
    n10201, n10202, n10203, n10204, n10206, n10207, n10208, n10209, n10210,
    n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10245, n10246, n10247, n10248, n10249, n10251,
    n10252, n10253, n10254, n10255, n10257, n10258, n10259, n10260, n10261,
    n10263, n10264, n10265, n10266, n10267, n10269, n10270, n10271, n10272,
    n10273, n10275, n10276, n10277, n10278, n10279, n10281, n10282, n10283,
    n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10292, n10293,
    n10294, n10295, n10296, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10309, n10310, n10311, n10312, n10313,
    n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
    n10324, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10337, n10338, n10339, n10340, n10341, n10343, n10344,
    n10345, n10346, n10347, n10349, n10350, n10351, n10352, n10353, n10354,
    n10355, n10356, n10357, n10358, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10371, n10372, n10373, n10374,
    n10375, n10377, n10378, n10379, n10380, n10381, n10383, n10384, n10385,
    n10386, n10387, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
    n10396, n10397, n10398, n10400, n10401, n10402, n10403, n10404, n10406,
    n10407, n10408, n10409, n10410, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432, n10434, n10435, n10436,
    n10437, n10438, n10440, n10441, n10442, n10443, n10444, n10446, n10447,
    n10448, n10449, n10450, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10463, n10464, n10465, n10466, n10467,
    n10469, n10470, n10471, n10472, n10473, n10475, n10476, n10477, n10478,
    n10479, n10481, n10482, n10483, n10484, n10485, n10487, n10488, n10489,
    n10490, n10491, n10493, n10494, n10495, n10496, n10497, n10499, n10500,
    n10501, n10502, n10503, n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10516, n10517, n10518, n10519, n10520,
    n10522, n10523, n10524, n10525, n10526, n10528, n10529, n10530, n10531,
    n10532, n10534, n10535, n10536, n10537, n10538, n10540, n10541, n10542,
    n10543, n10544, n10546, n10547, n10548, n10549, n10550, n10552, n10553,
    n10554, n10555, n10556, n10558, n10559, n10560, n10561, n10562, n10564,
    n10565, n10566, n10567, n10568, n10570, n10571, n10572, n10573, n10574,
    n10576, n10577, n10578, n10579, n10580, n10582, n10583, n10584, n10585,
    n10586, n10588, n10589, n10590, n10591, n10592, n10594, n10595, n10596,
    n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10605, n10606,
    n10607, n10608, n10609, n10611, n10612, n10613, n10614, n10615, n10617,
    n10618, n10619, n10620, n10621, n10623, n10624, n10625, n10626, n10627,
    n10629, n10630, n10631, n10632, n10633, n10635, n10636, n10637, n10638,
    n10639, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10652, n10653, n10654, n10655, n10656, n10658, n10659,
    n10660, n10661, n10662, n10664, n10665, n10666, n10667, n10668, n10670,
    n10671, n10672, n10673, n10674, n10676, n10677, n10678, n10679, n10680,
    n10682, n10683, n10684, n10685, n10686, n10688, n10689, n10690, n10691,
    n10692, n10694, n10695, n10696, n10697, n10698, n10700, n10701, n10702,
    n10703, n10704, n10706, n10707, n10708, n10709, n10710, n10712, n10713,
    n10714, n10715, n10716, n10718, n10719, n10720, n10721, n10722, n10724,
    n10725, n10726, n10727, n10728, n10730, n10731, n10732, n10733, n10734,
    n10736, n10737, n10738, n10739, n10740, n10742, n10743, n10744, n10745,
    n10746, n10748, n10749, n10750, n10751, n10752, n10754, n10755, n10756,
    n10757, n10758, n10760, n10761, n10762, n10763, n10764, n10766, n10767,
    n10768, n10769, n10770, n10772, n10773, n10774, n10775, n10776, n10778,
    n10779, n10780, n10781, n10782, n10784, n10785, n10786, n10787, n10788,
    n10790, n10791, n10792, n10793, n10794, n10796, n10797, n10798, n10799,
    n10800, n10801, n10802, n10803, n10804, n10805, n10807, n10808, n10809,
    n10810, n10811, n10813, n10814, n10815, n10816, n10817, n10819, n10820,
    n10821, n10822, n10823, n10825, n10826, n10827, n10828, n10829, n10831,
    n10832, n10834, n10835, n10836, n10837, n10838, n10840, n10841, n10842,
    n10843, n10844, n10846, n10847, n10848, n10849, n10850, n10852, n10853,
    n10854, n10855, n10856, n10858, n10859, n10860, n10861, n10862, n10864,
    n10865, n10866, n10867, n10868, n10870, n10871, n10872, n10873, n10874,
    n10876, n10877, n10878, n10879, n10880, n10882, n10883, n10884, n10885,
    n10886, n10888, n10889, n10890, n10891, n10892, n10894, n10895, n10896,
    n10897, n10898, n10900, n10901, n10902, n10903, n10904, n10906, n10907,
    n10908, n10909, n10910, n10912, n10913, n10914, n10915, n10916, n10918,
    n10919, n10920, n10921, n10922, n10924, n10925, n10926, n10927, n10928,
    n10930, n10931, n10932, n10933, n10934, n10936, n10937, n10938, n10939,
    n10940, n10942, n10943, n10944, n10945, n10946, n10948, n10949, n10950,
    n10951, n10952, n10954, n10955, n10956, n10957, n10958, n10960, n10961,
    n10962, n10963, n10964, n10966, n10967, n10968, n10969, n10970, n10972,
    n10973, n10974, n10975, n10976, n10978, n10979, n10980, n10981, n10982,
    n10984, n10985, n10986, n10987, n10988, n10990, n10991, n10992, n10993,
    n10994, n10996, n10997, n10998, n10999, n11000, n11002, n11003, n11004,
    n11005, n11006, n11008, n11009, n11010, n11011, n11012, n11014, n11015,
    n11016, n11017, n11018, n11020, n11021, n11022, n11023, n11024, n11026,
    n11027, n11028, n11029, n11030, n11032, n11033, n11034, n11035, n11036,
    n11038, n11039, n11040, n11041, n11042, n11044, n11045, n11046, n11047,
    n11048, n11050, n11051, n11052, n11053, n11054, n11056, n11057, n11058,
    n11059, n11060, n11062, n11063, n11064, n11065, n11066, n11067, n11069,
    n11070, n11072, n11073, n11075, n11076, n11078, n11079, n11081, n11082,
    n11084, n11085, n11087, n11088, n11090, n11091, n11093, n11094, n11096,
    n11097, n11099, n11100, n11102, n11103, n11105, n11106, n11108, n11109,
    n11111, n11112, n11113, n11114, n11115, n11117, n11119, n11121, n11123,
    n11124, n11125, n11127, n11128, n11130, n11131, n11132, n11133, n11134,
    n11136, n11137, n11139, n11140, n11141, n11143, n11144, n11146, n11148,
    n11149, n11151, n11152, n11154, n11155, n11157, n11158, n11160, n11161,
    n11163, n11164, n11165, n11166, n11167, n11168, n11170, n11171, n11173,
    n11174, n11176, n11177, n11179, n11180, n11182, n11183, n11185, n11186,
    n11188, n11189, n11191, n11192, n11194, n11195, n11197, n11198, n11200,
    n11201, n11203, n11204, n11206, n11207, n11209, n11210, n11212, n11213,
    n11215, n11216, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
    n11225, n11226, n11227, n11228, n11229, n11230, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11246, n11248, n11250, n11251, n11252, n11253, n11254, n11255,
    n11256, n11257, n11258, n11260, n11261, n11262, n11264, n11265, n11267,
    n11268, n11270, n11271, n11273, n11274, n11276, n11277, n11279, n11280,
    n11282, n11283, n11285, n11286, n11288, n11289, n11291, n11292, n11294,
    n11295, n11297, n11298, n11300, n11301, n11303, n11304, n11306, n11307,
    n11309, n11310, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324, n11326, n11327, n11328,
    n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
    n11338, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
    n11348, n11349, n11350, n11351, n11352, n11354, n11355, n11356, n11357,
    n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
    n11369, n11370, n11372, n11373, n11375, n11376, n11378, n11379, n11381,
    n11382, n11384, n11385, n11387, n11392, n11393, n11395, n11396, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404, n11406, n11407, n11408,
    n11409, n11410, n11412, n11413, n11415, n11416, n11418, n11419, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11462, n11463,
    n11464, n11465, n11467, n11468, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11484,
    n11485, n11486, n11487, n11490, n11491, n11493, n11494, n11495, n11496,
    n11497, n11499, n11500, n11501, n11502, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
    n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11543, n11544,
    n11545, n11546, n11547, n11549, n11550, n11551, n11552, n11553, n11554,
    n11556, n11557, n11558, n11559, n11560, n11562, n11563, n11564, n11565,
    n11566, n11567, n11569, n11570, n11571, n11572, n11573, n11575, n11576,
    n11577, n11578, n11579, n11580, n11582, n11583, n11584, n11585, n11586,
    n11588, n11589, n11590, n11591, n11592, n11593, n11595, n11597, n11598,
    n11599, n11600, n11601, n11603, n11604, n11605, n11606, n11607, n11608,
    n11610, n11611, n11612, n11613, n11614, n11616, n11617, n11618, n11619,
    n11620, n11621, n11623, n11624, n11626, n11627, n11629, n11630, n11631,
    n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
    n11641, n11643, n11644, n11646, n11647, n11649, n11650, n11652, n11653,
    n11655, n11656, n11658, n11659, n11661, n11662, n11664, n11665, n11667,
    n11668, n11669, n11671, n11672, n11673, n11675, n11676, n11677, n11679,
    n11680, n11681, n11683, n11684, n11685, n11687, n11688, n11689, n11691,
    n11692, n11694, n11695, n11696, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11721, n11722,
    n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
    n11732, n11733, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
    n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11751, n11752,
    n11753, n11754, n11755, n11756, n11757, n11759, n11760, n11761, n11763,
    n11764, n11765, n11766, n11767, n11768, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11778, n11779, n11780, n11781, n11782, n11783,
    n11784, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11794,
    n11795, n11796, n11797, n11798, n11799, n11800, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11810, n11811, n11812, n11813, n11814,
    n11815, n11816, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
    n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11834, n11835,
    n11836, n11837, n11838, n11839, n11840, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11850, n11851, n11852, n11853, n11854, n11855,
    n11856, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11866,
    n11867, n11869, n11870, n11872, n11873, n11875, n11876, n11878, n11879,
    n11881, n11882, n11883, n11884, n11885, n11886, n11888, n11889, n11890,
    n11891, n11892, n11894, n11895, n11896, n11897, n11898, n11900, n11901,
    n11902, n11903, n11904, n11906, n11907, n11908, n11909, n11910, n11912,
    n11913, n11914, n11915, n11916, n11918, n11919, n11920, n11921, n11922,
    n11924, n11925, n11926, n11927, n11928, n11930, n11931, n11932, n11933,
    n11934, n11936, n11937, n11938, n11939, n11940, n11942, n11943, n11944,
    n11945, n11946, n11947, n11949, n11950, n11951, n11952, n11953, n11955,
    n11956, n11957, n11958, n11959, n11961, n11962, n11963, n11964, n11965,
    n11967, n11968, n11969, n11970, n11971, n11973, n11974, n11975, n11976,
    n11977, n11979, n11980, n11981, n11982, n11983, n11985, n11986, n11987,
    n11988, n11989, n11991, n11992, n11993, n11994, n11995, n11997, n11998,
    n11999, n12000, n12001, n12003, n12004, n12005, n12006, n12007, n12008,
    n12010, n12011, n12012, n12013, n12014, n12016, n12017, n12018, n12019,
    n12020, n12022, n12023, n12024, n12025, n12026, n12028, n12029, n12030,
    n12031, n12032, n12034, n12035, n12036, n12037, n12038, n12040, n12041,
    n12042, n12043, n12044, n12046, n12047, n12048, n12049, n12050, n12052,
    n12053, n12054, n12055, n12056, n12058, n12059, n12060, n12061, n12062,
    n12064, n12065, n12066, n12067, n12068, n12069, n12071, n12072, n12073,
    n12074, n12075, n12077, n12078, n12079, n12080, n12081, n12083, n12084,
    n12085, n12086, n12087, n12089, n12090, n12091, n12092, n12093, n12095,
    n12096, n12097, n12098, n12099, n12101, n12102, n12103, n12104, n12105,
    n12107, n12108, n12109, n12110, n12111, n12113, n12114, n12115, n12116,
    n12117, n12119, n12120, n12121, n12122, n12123, n12125, n12126, n12127,
    n12128, n12129, n12130, n12132, n12133, n12134, n12135, n12136, n12138,
    n12139, n12140, n12141, n12142, n12144, n12145, n12146, n12147, n12148,
    n12149, n12151, n12152, n12153, n12154, n12155, n12157, n12158, n12159,
    n12160, n12161, n12163, n12164, n12165, n12166, n12167, n12169, n12170,
    n12171, n12172, n12173, n12175, n12176, n12177, n12178, n12179, n12181,
    n12182, n12183, n12184, n12185, n12187, n12188, n12189, n12190, n12191,
    n12193, n12194, n12195, n12196, n12197, n12199, n12200, n12201, n12202,
    n12203, n12205, n12206, n12207, n12208, n12209, n12211, n12212, n12213,
    n12214, n12215, n12217, n12218, n12219, n12220, n12221, n12223, n12224,
    n12225, n12226, n12227, n12229, n12230, n12231, n12232, n12233, n12235,
    n12236, n12237, n12238, n12239, n12241, n12242, n12243, n12244, n12245,
    n12247, n12249, n12250, n12252, n12253, n12254, n12255, n12256, n12258,
    n12259, n12260, n12261, n12262, n12264, n12265, n12266, n12267, n12268,
    n12270, n12271, n12272, n12273, n12274, n12276, n12277, n12278, n12279,
    n12280, n12282, n12283, n12284, n12285, n12286, n12288, n12289, n12290,
    n12291, n12292, n12294, n12295, n12296, n12297, n12299, n12300, n12301,
    n12302, n12303, n12305, n12306, n12307, n12308, n12309, n12311, n12312,
    n12313, n12314, n12315, n12317, n12318, n12319, n12320, n12321, n12323,
    n12324, n12325, n12326, n12327, n12329, n12330, n12331, n12332, n12333,
    n12335, n12336, n12337, n12338, n12339, n12341, n12342, n12343, n12344,
    n12345, n12347, n12348, n12349, n12350, n12351, n12353, n12354, n12355,
    n12356, n12357, n12359, n12360, n12361, n12362, n12363, n12365, n12366,
    n12367, n12368, n12369, n12371, n12372, n12373, n12374, n12375, n12377,
    n12378, n12379, n12380, n12381, n12383, n12384, n12386, n12387, n12388,
    n12389, n12391, n12392, n12393, n12394, n12395, n12397, n12398, n12399,
    n12400, n12401, n12403, n12404, n12405, n12406, n12407, n12409, n12410,
    n12411, n12412, n12413, n12415, n12416, n12417, n12418, n12419, n12421,
    n12422, n12423, n12424, n12425, n12427, n12428, n12429, n12430, n12431,
    n12433, n12434, n12435, n12436, n12437, n12439, n12440, n12441, n12442,
    n12443, n12445, n12446, n12447, n12448, n12449, n12451, n12452, n12453,
    n12454, n12455, n12457, n12458, n12459, n12460, n12461, n12463, n12464,
    n12465, n12466, n12467, n12469, n12470, n12471, n12472, n12473, n12475,
    n12476, n12477, n12478, n12479, n12481, n12482, n12483, n12484, n12485,
    n12487, n12488, n12489, n12490, n12491, n12493, n12494, n12495, n12496,
    n12497, n12499, n12500, n12501, n12502, n12503, n12505, n12506, n12507,
    n12508, n12509, n12511, n12512, n12513, n12514, n12515, n12517, n12518,
    n12519, n12520, n12521, n12523, n12524, n12525, n12526, n12527, n12529,
    n12530, n12531, n12532, n12533, n12535, n12536, n12537, n12538, n12539,
    n12541, n12542, n12543, n12544, n12545, n12547, n12548, n12549, n12550,
    n12551, n12553, n12554, n12555, n12556, n12557, n12559, n12560, n12561,
    n12562, n12563, n12565, n12566, n12567, n12568, n12569, n12571, n12572,
    n12573, n12574, n12575, n12577, n12578, n12579, n12580, n12581, n12583,
    n12584, n12585, n12586, n12587, n12589, n12590, n12591, n12592, n12593,
    n12595, n12596, n12597, n12598, n12599, n12601, n12602, n12603, n12604,
    n12605, n12607, n12608, n12609, n12610, n12611, n12613, n12614, n12615,
    n12616, n12617, n12619, n12620, n12621, n12622, n12623, n12625, n12626,
    n12627, n12628, n12629, n12631, n12632, n12633, n12634, n12635, n12637,
    n12638, n12639, n12640, n12641, n12643, n12644, n12645, n12646, n12647,
    n12649, n12650, n12651, n12652, n12653, n12655, n12656, n12657, n12658,
    n12659, n12661, n12662, n12663, n12664, n12665, n12667, n12668, n12669,
    n12670, n12671, n12673, n12674, n12675, n12676, n12677, n12679, n12680,
    n12681, n12682, n12683, n12685, n12686, n12687, n12688, n12689, n12691,
    n12692, n12693, n12694, n12695, n12697, n12698, n12699, n12700, n12701,
    n12703, n12704, n12705, n12706, n12707, n12709, n12710, n12711, n12712,
    n12713, n12715, n12716, n12717, n12718, n12719, n12721, n12722, n12723,
    n12724, n12725, n12727, n12728, n12729, n12730, n12731, n12733, n12734,
    n12735, n12736, n12737, n12739, n12740, n12741, n12742, n12743, n12745,
    n12746, n12747, n12748, n12749, n12751, n12752, n12753, n12754, n12755,
    n12757, n12758, n12759, n12760, n12761, n12763, n12764, n12765, n12766,
    n12767, n12769, n12770, n12771, n12772, n12773, n12775, n12776, n12777,
    n12778, n12779, n12781, n12782, n12783, n12784, n12785, n12787, n12788,
    n12789, n12790, n12791, n12793, n12794, n12795, n12796, n12797, n12799,
    n12800, n12801, n12802, n12803, n12805, n12806, n12807, n12808, n12809,
    n12811, n12812, n12813, n12814, n12815, n12817, n12818, n12819, n12820,
    n12821, n12823, n12824, n12825, n12826, n12827, n12829, n12830, n12831,
    n12832, n12833, n12835, n12836, n12837, n12838, n12839, n12841, n12842,
    n12843, n12844, n12845, n12847, n12848, n12849, n12850, n12851, n12853,
    n12854, n12855, n12856, n12857, n12859, n12860, n12861, n12862, n12863,
    n12865, n12866, n12867, n12868, n12869, n12871, n12872, n12873, n12874,
    n12875, n12877, n12878, n12879, n12880, n12881, n12883, n12884, n12886,
    n12887, n12889, n12890, n12891, n12892, n12893, n12895, n12896, n12898,
    n12899, n12901, n12902, n12904, n12905, n12907, n12908, n12909, n12911,
    n12912, n12914, n12915, n12917, n12918, n12919, n12920, n12921, n12923,
    n12924, n12925, n12926, n12927, n12929, n12930, n12932, n12933, n12935,
    n12936, n12938, n12939, n12941, n12942, n12944, n12945, n12947, n12948,
    n12950, n12951, n12953, n12954, n12956, n12957, n12959, n12960, n12962,
    n12963, n12965, n12966, n12968, n12969, n12971, n12972, n12974, n12975,
    n12977, n12978, n12980, n12981, n12983, n12984, n12986, n12987, n12989,
    n12990, n12992, n12993, n12995, n12996, n12998, n12999, n13001, n13002,
    n13004, n13005, n13007, n13008, n13010, n13011, n13013, n13014, n13016,
    n13017, n13019, n13020, n13022, n13023, n13025, n13026, n13028, n13029,
    n13031, n13032, n13034, n13035, n13037, n13038, n13040, n13041, n13043,
    n13044, n13046, n13047, n13049, n13050, n13052, n13053, n13055, n13056,
    n13058, n13059, n13061, n13062, n13064, n13065, n13067, n13068, n13070,
    n13071, n13073, n13074, n13076, n13077, n13079, n13080, n13082, n13083,
    n13085, n13086, n13088, n13089, n13091, n13092, n13094, n13095, n13097,
    n13098, n13100, n13101, n13103, n13104, n13106, n13107, n13109, n13110,
    n13112, n13113, n13115, n13116, n13118, n13119, n13121, n13122, n13124,
    n13125, n13127, n13128, n13130, n13131, n13133, n13134, n13136, n13137,
    n13139, n13140, n13142, n13143, n13145, n13146, n13148, n13149, n13151,
    n13152, n13154, n13155, n13157, n13158, n13160, n13161, n13163, n13164,
    n13166, n13167, n13169, n13170, n13172, n13173, n13175, n13176, n13178,
    n13179, n13181, n13182, n13184, n13185, n13187, n13188, n13190, n13191,
    n13192, n13193, n13194, n13196, n13197, n13198, n13199, n13200, n13202,
    n13203, n13204, n13205, n13206, n13208, n13209, n13210, n13211, n13212,
    n13214, n13215, n13216, n13217, n13218, n13220, n13221, n13222, n13223,
    n13224, n13226, n13227, n13228, n13229, n13230, n13232, n13233, n13234,
    n13235, n13236, n13238, n13239, n13240, n13241, n13242, n13244, n13245,
    n13246, n13247, n13248, n13250, n13251, n13252, n13253, n13254, n13256,
    n13257, n13258, n13259, n13260, n13262, n13263, n13264, n13265, n13266,
    n13268, n13269, n13270, n13271, n13272, n13274, n13275, n13276, n13277,
    n13278, n13280, n13281, n13282, n13283, n13284, n13286, n13287, n13288,
    n13289, n13290, n13292, n13293, n13294, n13295, n13296, n13298, n13299,
    n13300, n13301, n13302, n13304, n13305, n13306, n13307, n13308, n13310,
    n13311, n13312, n13313, n13314, n13316, n13317, n13318, n13319, n13320,
    n13322, n13323, n13324, n13325, n13326, n13328, n13329, n13330, n13331,
    n13332, n13334, n13335, n13336, n13337, n13338, n13340, n13341, n13342,
    n13343, n13344, n13346, n13347, n13348, n13349, n13350, n13352, n13353,
    n13354, n13355, n13356, n13358, n13359, n13360, n13361, n13362, n13364,
    n13365, n13366, n13367, n13368, n13370, n13371, n13372, n13373, n13374,
    n13376, n13377, n13378, n13379, n13380, n13382, n13383, n13384, n13385,
    n13386, n13388, n13389, n13390, n13391, n13392, n13394, n13395, n13396,
    n13397, n13398, n13400, n13401, n13402, n13403, n13404, n13406, n13407,
    n13408, n13409, n13410, n13412, n13413, n13414, n13415, n13416, n13418,
    n13419, n13420, n13421, n13422, n13424, n13425, n13426, n13427, n13428,
    n13430, n13431, n13432, n13433, n13434, n13436, n13437, n13438, n13439,
    n13440, n13442, n13443, n13444, n13445, n13446, n13448, n13449, n13450,
    n13451, n13452, n13454, n13455, n13456, n13457, n13458, n13460, n13461,
    n13462, n13463, n13464, n13466, n13467, n13468, n13469, n13470, n13472,
    n13473, n13474, n13475, n13476, n13478, n13479, n13480, n13481, n13482,
    n13484, n13485, n13486, n13487, n13488, n13490, n13491, n13492, n13493,
    n13494, n13496, n13497, n13498, n13499, n13500, n13502, n13503, n13504,
    n13505, n13506, n13508, n13509, n13510, n13511, n13512, n13514, n13515,
    n13516, n13517, n13518, n13520, n13521, n13522, n13523, n13524, n13526,
    n13527, n13528, n13529, n13530, n13532, n13533, n13534, n13535, n13536,
    n13538, n13539, n13540, n13541, n13542, n13544, n13545, n13546, n13547,
    n13548, n13550, n13551, n13552, n13553, n13554, n13556, n13557, n13558,
    n13559, n13560, n13562, n13563, n13564, n13565, n13566, n13568, n13569,
    n13570, n13571, n13572, n13574, n13575, n13576, n13577, n13578, n13580,
    n13581, n13582, n13583, n13584, n13586, n13587, n13588, n13589, n13590,
    n13592, n13593, n13594, n13595, n13596, n13598, n13599, n13600, n13601,
    n13602, n13604, n13605, n13606, n13607, n13608, n13610, n13611, n13612,
    n13613, n13614, n13616, n13617, n13618, n13619, n13620, n13622, n13623,
    n13624, n13625, n13626, n13628, n13629, n13630, n13631, n13632, n13634,
    n13635, n13636, n13637, n13638, n13640, n13641, n13642, n13643, n13644,
    n13646, n13647, n13648, n13649, n13650, n13652, n13653, n13654, n13655,
    n13656, n13658, n13659, n13660, n13661, n13662, n13664, n13665, n13666,
    n13667, n13668, n13670, n13671, n13672, n13673, n13674, n13676, n13677,
    n13678, n13679, n13680, n13682, n13683, n13684, n13685, n13686, n13688,
    n13689, n13690, n13691, n13692, n13694, n13695, n13696, n13697, n13698,
    n13700, n13701, n13702, n13703, n13704, n13706, n13707, n13708, n13709,
    n13710, n13712, n13713, n13714, n13715, n13716, n13718, n13719, n13720,
    n13721, n13722, n13724, n13725, n13726, n13727, n13728, n13730, n13731,
    n13732, n13733, n13734, n13736, n13737, n13738, n13739, n13740, n13742,
    n13743, n13744, n13745, n13746, n13748, n13749, n13750, n13751, n13752,
    n13754, n13755, n13756, n13757, n13758, n13760, n13761, n13762, n13763,
    n13764, n13766, n13767, n13768, n13769, n13770, n13772, n13773, n13774,
    n13775, n13776, n13778, n13779, n13780, n13781, n13782, n13784, n13785,
    n13786, n13787, n13788, n13790, n13791, n13792, n13793, n13794, n13796,
    n13797, n13798, n13799, n13800, n13802, n13803, n13804, n13805, n13806,
    n13808, n13809, n13810, n13811, n13812, n13814, n13815, n13816, n13817,
    n13818, n13820, n13821, n13822, n13823, n13824, n13826, n13827, n13828,
    n13829, n13830, n13832, n13833, n13834, n13835, n13836, n13838, n13839,
    n13840, n13841, n13842, n13844, n13845, n13846, n13847, n13848, n13850,
    n13851, n13852, n13853, n13854, n13856, n13857, n13858, n13859, n13860,
    n13862, n13863, n13864, n13865, n13866, n13868, n13869, n13870, n13871,
    n13872, n13874, n13875, n13876, n13877, n13878, n13880, n13881, n13882,
    n13883, n13884, n13886, n13887, n13888, n13889, n13890, n13892, n13893,
    n13894, n13895, n13896, n13898, n13899, n13900, n13901, n13902, n13904,
    n13905, n13906, n13907, n13908, n13910, n13911, n13912, n13913, n13914,
    n13916, n13917, n13918, n13919, n13920, n13922, n13923, n13924, n13925,
    n13926, n13928, n13929, n13930, n13931, n13932, n13934, n13935, n13936,
    n13937, n13938, n13940, n13941, n13942, n13943, n13944, n13946, n13947,
    n13948, n13949, n13950, n13952, n13953, n13954, n13955, n13956, n13958,
    n13959, n13960, n13961, n13962, n13964, n13965, n13966, n13967, n13968,
    n13970, n13971, n13972, n13973, n13974, n13976, n13977, n13978, n13979,
    n13980, n13982, n13983, n13984, n13985, n13986, n13988, n13989, n13990,
    n13991, n13992, n13994, n13995, n13996, n13997, n13998, n14000, n14001,
    n14002, n14003, n14004, n14006, n14007, n14008, n14009, n14010, n14012,
    n14013, n14014, n14015, n14016, n14018, n14019, n14020, n14021, n14022,
    n14024, n14025, n14026, n14027, n14028, n14030, n14031, n14032, n14033,
    n14034, n14036, n14037, n14038, n14039, n14040, n14042, n14043, n14044,
    n14045, n14046, n14048, n14049, n14050, n14051, n14052, n14054, n14055,
    n14056, n14057, n14058, n14060, n14061, n14062, n14063, n14064, n14066,
    n14067, n14068, n14069, n14070, n14072, n14073, n14074, n14075, n14076,
    n14078, n14079, n14080, n14081, n14082, n14084, n14085, n14086, n14087,
    n14088, n14090, n14091, n14092, n14093, n14094, n14096, n14097, n14098,
    n14099, n14100, n14102, n14103, n14104, n14105, n14106, n14108, n14109,
    n14110, n14111, n14112, n14114, n14115, n14116, n14117, n14118, n14120,
    n14121, n14122, n14123, n14124, n14126, n14127, n14128, n14129, n14130,
    n14132, n14133, n14134, n14135, n14136, n14138, n14139, n14140, n14141,
    n14142, n14144, n14145, n14146, n14147, n14148, n14150, n14151, n14152,
    n14153, n14154, n14156, n14157, n14158, n14159, n14160, n14162, n14163,
    n14164, n14165, n14166, n14168, n14169, n14170, n14171, n14172, n14174,
    n14175, n14176, n14177, n14178, n14180, n14181, n14182, n14183, n14184,
    n14186, n14187, n14188, n14189, n14190, n14192, n14193, n14194, n14195,
    n14196, n14198, n14199, n14200, n14201, n14202, n14204, n14205, n14206,
    n14207, n14208, n14210, n14211, n14212, n14213, n14214, n14216, n14217,
    n14218, n14219, n14220, n14222, n14223, n14224, n14225, n14226, n14228,
    n14229, n14230, n14231, n14232, n14234, n14235, n14236, n14237, n14238,
    n14240, n14241, n14242, n14243, n14244, n14246, n14247, n14248, n14249,
    n14250, n14252, n14253, n14254, n14255, n14256, n14258, n14259, n14260,
    n14261, n14262, n14264, n14265, n14266, n14267, n14268, n14270, n14271,
    n14272, n14273, n14274, n14276, n14277, n14278, n14279, n14280, n14282,
    n14283, n14284, n14285, n14286, n14288, n14289, n14290, n14291, n14292,
    n14294, n14295, n14296, n14297, n14298, n14300, n14301, n14302, n14303,
    n14304, n14306, n14307, n14308, n14309, n14310, n14312, n14313, n14314,
    n14315, n14316, n14318, n14319, n14320, n14321, n14322, n14324, n14325,
    n14326, n14327, n14328, n14330, n14331, n14332, n14333, n14334, n14336,
    n14337, n14338, n14339, n14340, n14342, n14343, n14344, n14345, n14346,
    n14348, n14349, n14350, n14351, n14352, n14354, n14355, n14356, n14357,
    n14358, n14360, n14361, n14362, n14363, n14364, n14366, n14367, n14368,
    n14369, n14370, n14372, n14373, n14374, n14375, n14376, n14378, n14379,
    n14380, n14381, n14382, n14384, n14385, n14386, n14387, n14388, n14390,
    n14391, n14392, n14393, n14394, n14396, n14397, n14398, n14399, n14400,
    n14402, n14403, n14404, n14405, n14406, n14408, n14409, n14410, n14411,
    n14412, n14414, n14415, n14416, n14417, n14418, n14420, n14421, n14422,
    n14423, n14424, n14426, n14427, n14428, n14429, n14430, n14432, n14433,
    n14434, n14435, n14436, n14438, n14439, n14440, n14441, n14442, n14444,
    n14445, n14446, n14447, n14448, n14450, n14451, n14452, n14453, n14454,
    n14456, n14457, n14458, n14459, n14460, n14462, n14463, n14464, n14465,
    n14466, n14468, n14469, n14470, n14471, n14472, n14474, n14475, n14476,
    n14477, n14478, n14480, n14481, n14482, n14483, n14484, n14486, n14487,
    n14488, n14489, n14490, n14492, n14493, n14494, n14495, n14496, n14498,
    n14499, n14500, n14501, n14502, n14504, n14505, n14506, n14507, n14508,
    n14510, n14511, n14512, n14513, n14514, n14516, n14517, n14518, n14519,
    n14520, n14522, n14523, n14524, n14525, n14526, n14528, n14529, n14530,
    n14531, n14532, n14534, n14535, n14536, n14537, n14538, n14540, n14541,
    n14542, n14543, n14544, n14546, n14547, n14548, n14549, n14550, n14552,
    n14553, n14554, n14555, n14556, n14558, n14559, n14560, n14561, n14562,
    n14564, n14565, n14566, n14567, n14568, n14570, n14571, n14572, n14573,
    n14574, n14576, n14577, n14578, n14579, n14580, n14582, n14583, n14584,
    n14585, n14586, n14588, n14589, n14590, n14591, n14592, n14594, n14595,
    n14596, n14597, n14598, n14600, n14601, n14602, n14603, n14604, n14606,
    n14607, n14608, n14609, n14610, n14612, n14613, n14614, n14615, n14616,
    n14618, n14619, n14620, n14621, n14622, n14624, n14625, n14626, n14627,
    n14628, n14630, n14631, n14632, n14633, n14634, n14636, n14637, n14638,
    n14639, n14640, n14642, n14643, n14644, n14645, n14646, n14648, n14649,
    n14650, n14651, n14652, n14654, n14655, n14656, n14657, n14658, n14660,
    n14661, n14662, n14663, n14664, n14666, n14667, n14668, n14669, n14670,
    n14672, n14673, n14674, n14675, n14676, n14678, n14679, n14680, n14681,
    n14682, n14684, n14685, n14686, n14687, n14688, n14690, n14691, n14692,
    n14693, n14694, n14696, n14697, n14698, n14699, n14700, n14702, n14703,
    n14704, n14705, n14706, n14708, n14709, n14710, n14711, n14712, n14714,
    n14715, n14716, n14717, n14718, n14720, n14721, n14722, n14723, n14724,
    n14726, n14727, n14728, n14729, n14730, n14732, n14733, n14734, n14735,
    n14736, n14738, n14739, n14740, n14741, n14742, n14744, n14745, n14746,
    n14747, n14748, n14750, n14751, n14752, n14753, n14754, n14756, n14757,
    n14758, n14759, n14760, n14762, n14763, n14764, n14765, n14766, n14768,
    n14769, n14770, n14771, n14772, n14774, n14775, n14776, n14777, n14778,
    n14780, n14781, n14782, n14783, n14784, n14786, n14787, n14788, n14789,
    n14790, n14792, n14793, n14794, n14795, n14796, n14798, n14799, n14800,
    n14801, n14802, n14804, n14805, n14806, n14807, n14808, n14810, n14811,
    n14812, n14813, n14814, n14816, n14817, n14818, n14819, n14820, n14822,
    n14823, n14824, n14825, n14826, n14828, n14829, n14830, n14831, n14832,
    n14834, n14835, n14836, n14837, n14838, n14840, n14841, n14842, n14843,
    n14844, n14846, n14847, n14848, n14849, n14850, n14852, n14853, n14854,
    n14855, n14856, n14858, n14859, n14860, n14861, n14862, n14864, n14865,
    n14866, n14867, n14868, n14870, n14871, n14872, n14873, n14874, n14876,
    n14877, n14878, n14879, n14880, n14882, n14883, n14884, n14885, n14886,
    n14888, n14889, n14890, n14891, n14892, n14894, n14895, n14896, n14897,
    n14898, n14900, n14901, n14902, n14903, n14904, n14906, n14907, n14908,
    n14909, n14910, n14912, n14913, n14914, n14915, n14916, n14918, n14919,
    n14920, n14921, n14922, n14924, n14925, n14926, n14927, n14928, n14930,
    n14931, n14932, n14933, n14934, n14936, n14937, n14938, n14939, n14940,
    n14942, n14943, n14944, n14945, n14946, n14948, n14949, n14950, n14951,
    n14952, n14954, n14955, n14956, n14957, n14958, n14960, n14961, n14962,
    n14963, n14964, n14966, n14967, n14968, n14969, n14970, n14972, n14973,
    n14974, n14975, n14976, n14978, n14979, n14980, n14981, n14982, n14984,
    n14985, n14986, n14987, n14988, n14990, n14991, n14992, n14993, n14994,
    n14996, n14997, n14998, n14999, n15000, n15002, n15003, n15004, n15005,
    n15006, n15008, n15009, n15010, n15011, n15012, n15014, n15015, n15016,
    n15017, n15018, n15020, n15021, n15022, n15023, n15024, n15026, n15027,
    n15028, n15029, n15030, n15032, n15033, n15034, n15035, n15036, n15038,
    n15039, n15040, n15041, n15042, n15044, n15045, n15046, n15047, n15048,
    n15050, n15051, n15052, n15053, n15054, n15056, n15057, n15058, n15059,
    n15060, n15062, n15063, n15064, n15065, n15066, n15068, n15069, n15070,
    n15071, n15072, n15074, n15075, n15076, n15077, n15078, n15080, n15081,
    n15082, n15083, n15084, n15086, n15087, n15088, n15089, n15090, n15092,
    n15093, n15094, n15095, n15096, n15098, n15099, n15100, n15101, n15102,
    n15104, n15105, n15106, n15107, n15108, n15110, n15111, n15112, n15113,
    n15114, n15116, n15117, n15118, n15119, n15120, n15122, n15123, n15124,
    n15125, n15126, n15128, n15129, n15130, n15131, n15132, n15134, n15135,
    n15136, n15137, n15138, n15140, n15141, n15142, n15143, n15144, n15146,
    n15147, n15148, n15149, n15150, n15152, n15153, n15154, n15155, n15156,
    n15158, n15159, n15160, n15161, n15162, n15164, n15165, n15166, n15167,
    n15168, n15170, n15171, n15172, n15173, n15174, n15176, n15177, n15178,
    n15179, n15180, n15182, n15183, n15184, n15185, n15186, n15188, n15189,
    n15190, n15191, n15192, n15194, n15195, n15196, n15197, n15198, n15200,
    n15201, n15202, n15203, n15204, n15206, n15207, n15208, n15209, n15210,
    n15212, n15213, n15214, n15215, n15216, n15218, n15219, n15220, n15221,
    n15222, n15224, n15225, n15226, n15227, n15228, n15230, n15231, n15232,
    n15233, n15234, n15236, n15237, n15238, n15239, n15240, n15242, n15243,
    n15244, n15245, n15246, n15248, n15249, n15250, n15251, n15252, n15254,
    n15255, n15256, n15257, n15258, n15260, n15261, n15262, n15263, n15264,
    n15266, n15267, n15268, n15269, n15270, n15272, n15273, n15274, n15275,
    n15276, n15278, n15279, n15280, n15281, n15282, n15284, n15285, n15286,
    n15287, n15288, n15290, n15291, n15292, n15293, n15294, n15296, n15297,
    n15298, n15299, n15300, n15302, n15303, n15304, n15305, n15306, n15308,
    n15309, n15310, n15311, n15312, n15314, n15315, n15316, n15317, n15318,
    n15320, n15321, n15322, n15323, n15324, n15326, n15327, n15328, n15329,
    n15330, n15332, n15333, n15334, n15335, n15336, n15338, n15339, n15340,
    n15341, n15342, n15344, n15345, n15346, n15347, n15348, n15350, n15351,
    n15352, n15353, n15354, n15356, n15357, n15358, n15359, n15360, n15362,
    n15363, n15364, n15365, n15366, n15368, n15369, n15370, n15371, n15372,
    n15374, n15375, n15376, n15377, n15378, n15380, n15381, n15382, n15383,
    n15384, n15386, n15387, n15388, n15389, n15390, n15392, n15393, n15394,
    n15395, n15396, n15398, n15399, n15400, n15401, n15402, n15404, n15405,
    n15406, n15407, n15408, n15410, n15411, n15412, n15413, n15414, n15416,
    n15417, n15418, n15419, n15420, n15422, n15423, n15424, n15425, n15426,
    n15428, n15429, n15430, n15431, n15432, n15434, n15435, n15436, n15437,
    n15438, n15440, n15441, n15442, n15443, n15444, n15446, n15447, n15448,
    n15449, n15450, n15452, n15453, n15454, n15455, n15456, n15458, n15459,
    n15460, n15461, n15462, n15464, n15465, n15466, n15467, n15468, n15470,
    n15471, n15472, n15473, n15474, n15476, n15477, n15478, n15479, n15480,
    n15482, n15483, n15484, n15485, n15486, n15488, n15489, n15490, n15491,
    n15492, n15494, n15495, n15496, n15497, n15498, n15500, n15501, n15502,
    n15503, n15504, n15506, n15507, n15508, n15509, n15510, n15512, n15513,
    n15514, n15515, n15516, n15518, n15519, n15520, n15521, n15522, n15524,
    n15525, n15526, n15527, n15528, n15530, n15531, n15532, n15533, n15534,
    n15536, n15537, n15538, n15539, n15540, n15542, n15543, n15544, n15545,
    n15546, n15548, n15549, n15550, n15551, n15552, n15554, n15555, n15556,
    n15557, n15558, n15560, n15561, n15562, n15563, n15564, n15566, n15567,
    n15568, n15569, n15570, n15572, n15573, n15574, n15575, n15576, n15578,
    n15579, n15580, n15581, n15582, n15584, n15585, n15586, n15587, n15588,
    n15590, n15591, n15592, n15593, n15594, n15596, n15597, n15598, n15599,
    n15600, n15602, n15603, n15604, n15605, n15606, n15608, n15609, n15610,
    n15611, n15612, n15614, n15615, n15616, n15617, n15618, n15620, n15621,
    n15622, n15623, n15624, n15626, n15627, n15628, n15629, n15630, n15632,
    n15633, n15634, n15635, n15636, n15638, n15639, n15640, n15641, n15642,
    n15644, n15645, n15646, n15647, n15648, n15650, n15651, n15652, n15653,
    n15654, n15656, n15657, n15658, n15659, n15660, n15662, n15663, n15664,
    n15665, n15666, n15668, n15669, n15670, n15671, n15672, n15674, n15675,
    n15676, n15677, n15678, n15680, n15681, n15682, n15683, n15684, n15686,
    n15687, n15688, n15689, n15690, n15692, n15693, n15694, n15695, n15696,
    n15698, n15699, n15700, n15701, n15702, n15704, n15705, n15706, n15707,
    n15708, n15710, n15711, n15712, n15713, n15714, n15716, n15717, n15718,
    n15719, n15720, n15722, n15723, n15724, n15725, n15726, n15728, n15729,
    n15730, n15731, n15732, n15734, n15735, n15736, n15737, n15738, n15740,
    n15741, n15742, n15743, n15744, n15746, n15747, n15748, n15749, n15750,
    n15752, n15753, n15754, n15755, n15756, n15758, n15759, n15760, n15761,
    n15762, n15764, n15765, n15766, n15767, n15768, n15770, n15771, n15772,
    n15773, n15774, n15776, n15777, n15778, n15779, n15780, n15782, n15783,
    n15784, n15785, n15786, n15788, n15789, n15790, n15791, n15792, n15794,
    n15795, n15796, n15797, n15798, n15800, n15801, n15802, n15803, n15804,
    n15806, n15807, n15808, n15809, n15810, n15812, n15813, n15814, n15815,
    n15816, n15818, n15819, n15820, n15821, n15822, n15824, n15825, n15826,
    n15827, n15828, n15830, n15831, n15832, n15833, n15834, n15836, n15837,
    n15838, n15839, n15840, n15842, n15843, n15844, n15845, n15846, n15848,
    n15849, n15850, n15851, n15852, n15854, n15855, n15856, n15857, n15858,
    n15860, n15861, n15862, n15863, n15864, n15866, n15867, n15868, n15869,
    n15870, n15872, n15873, n15874, n15875, n15876, n15878, n15879, n15880,
    n15881, n15882, n15884, n15885, n15886, n15887, n15888, n15890, n15891,
    n15892, n15893, n15894, n15896, n15897, n15898, n15899, n15900, n15902,
    n15903, n15904, n15905, n15906, n15908, n15909, n15910, n15911, n15912,
    n15914, n15915, n15916, n15917, n15918, n15920, n15921, n15922, n15923,
    n15924, n15926, n15927, n15928, n15929, n15930, n15932, n15933, n15934,
    n15935, n15936, n15938, n15939, n15940, n15941, n15942, n15944, n15945,
    n15946, n15947, n15948, n15950, n15951, n15952, n15953, n15954, n15956,
    n15957, n15958, n15959, n15960, n15962, n15963, n15964, n15965, n15966,
    n15968, n15969, n15970, n15971, n15972, n15974, n15975, n15976, n15977,
    n15978, n15980, n15981, n15982, n15983, n15984, n15986, n15987, n15989,
    n15990, n15991, n15992, n15993, n15995, n15996, n15997, n15998, n15999,
    n16001, n16002, n16003, n16004, n16005, n16007, n16008, n16009, n16010,
    n16011, n16013, n16014, n16015, n16016, n16017, n16019, n16020, n16021,
    n16022, n16023, n16025, n16026, n16027, n16028, n16029, n16031, n16032,
    n16033, n16034, n16035, n16037, n16038, n16039, n16040, n16041, n16043,
    n16044, n16045, n16046, n16047, n16049, n16050, n16051, n16052, n16053,
    n16055, n16056, n16057, n16058, n16059, n16061, n16062, n16063, n16064,
    n16065, n16067, n16068, n16069, n16070, n16071, n16073, n16074, n16075,
    n16076, n16077, n16079, n16080, n16081, n16082, n16083, n16085, n16086,
    n16087, n16088, n16089, n16091, n16092, n16093, n16094, n16095, n16097,
    n16098, n16099, n16100, n16101, n16103, n16104, n16105, n16106, n16107,
    n16109, n16110, n16111, n16112, n16113, n16115, n16116, n16117, n16118,
    n16119, n16121, n16122, n16123, n16124, n16125, n16127, n16128, n16129,
    n16130, n16131, n16133, n16134, n16135, n16136, n16137, n16139, n16140,
    n16141, n16142, n16143, n16145, n16146, n16147, n16148, n16149, n16151,
    n16152, n16153, n16154, n16155, n16157, n16158, n16159, n16160, n16161,
    n16163, n16164, n16165, n16166, n16167, n16169, n16170, n16171, n16172,
    n16173, n16175, n16176, n16177, n16178, n16179, n16181, n16182, n16183,
    n16184, n16185, n16187, n16188, n16189, n16190, n16191, n16193, n16194,
    n16195, n16196, n16197, n16199, n16200, n16201, n16202, n16203, n16205,
    n16206, n16207, n16208, n16209, n16211, n16212, n16213, n16214, n16215,
    n16217, n16218, n16219, n16220, n16221, n16223, n16224, n16225, n16226,
    n16227, n16229, n16230, n16231, n16232, n16233, n16235, n16236, n16237,
    n16238, n16239, n16241, n16242, n16243, n16244, n16245, n16247, n16248,
    n16249, n16250, n16251, n16253, n16254, n16255, n16256, n16257, n16259,
    n16260, n16261, n16262, n16263, n16265, n16266, n16267, n16268, n16269,
    n16271, n16272, n16273, n16274, n16275, n16277, n16278, n16279, n16280,
    n16281, n16283, n16284, n16285, n16286, n16287, n16289, n16290, n16291,
    n16292, n16293, n16295, n16296, n16297, n16298, n16299, n16301, n16302,
    n16303, n16304, n16305, n16307, n16308, n16309, n16310, n16311, n16313,
    n16314, n16315, n16316, n16317, n16319, n16320, n16321, n16322, n16323,
    n16325, n16326, n16327, n16328, n16329, n16331, n16332, n16333, n16334,
    n16335, n16337, n16338, n16339, n16340, n16341, n16343, n16344, n16345,
    n16346, n16347, n16349, n16350, n16351, n16352, n16353, n16355, n16356,
    n16357, n16358, n16359, n16361, n16362, n16363, n16364, n16365, n16367,
    n16368, n16369, n16370, n16371, n16373, n16374, n16375, n16376, n16377,
    n16379, n16380, n16382, n16383, n16384, n16385, n16386, n16388, n16389,
    n16390, n16391, n16392, n16394, n16395, n16396, n16397, n16398, n16400,
    n16401, n16403, n16404, n16405, n16406, n16407, n16409, n16410, n16412,
    n16413, n16414, n16415, n16416, n16418, n16419, n16420, n16421, n16422,
    n16424, n16425, n16426, n16427, n16428, n16430, n16431, n16432, n16433,
    n16434, n16436, n16437, n16438, n16439, n16440, n16442, n16443, n16444,
    n16445, n16446, n16448, n16449, n16450, n16451, n16452, n16454, n16455,
    n16457, n16458, n16459, n16460, n16461, n16463, n16464, n16465, n16466,
    n16467, n16469, n16470, n16471, n16472, n16473, n16475, n16476, n16477,
    n16478, n16479, n16481, n16482, n16483, n16484, n16485, n16487, n16488,
    n16490, n16491, n16492, n16493, n16494, n16496, n16497, n16499, n16500,
    n16501, n16502, n16503, n16505, n16506, n16507, n16508, n16509, n16511,
    n16512, n16513, n16514, n16515, n16517, n16518, n16519, n16520, n16521,
    n16523, n16524, n16525, n16526, n16527, n16529, n16530, n16531, n16532,
    n16533, n16535, n16536, n16537, n16538, n16539, n16541, n16542, n16543,
    n16544, n16545, n16547, n16548, n16549, n16550, n16551, n16553, n16554,
    n16556, n16557, n16558, n16559, n16560, n16562, n16563, n16564, n16565,
    n16566, n16568, n16569, n16570, n16571, n16572, n16574, n16575, n16576,
    n16577, n16578, n16580, n16581, n16582, n16583, n16584, n16586, n16587,
    n16588, n16589, n16590, n16592, n16593, n16594, n16595, n16596, n16598,
    n16599, n16600, n16601, n16602, n16604, n16605, n16606, n16607, n16608,
    n16610, n16611, n16612, n16613, n16614, n16616, n16617, n16618, n16619,
    n16620, n16622, n16623, n16624, n16625, n16626, n16628, n16629, n16630,
    n16631, n16632, n16634, n16635, n16636, n16637, n16638, n16640, n16641,
    n16642, n16643, n16644, n16646, n16647, n16648, n16649, n16650, n16652,
    n16653, n16654, n16655, n16656, n16658, n16659, n16660, n16661, n16662,
    n16664, n16665, n16666, n16667, n16668, n16670, n16671, n16672, n16673,
    n16674, n16676, n16677, n16678, n16679, n16680, n16682, n16683, n16684,
    n16685, n16686, n16688, n16689, n16690, n16691, n16692, n16694, n16695,
    n16696, n16697, n16698, n16700, n16701, n16702, n16703, n16704, n16706,
    n16707, n16708, n16709, n16710, n16712, n16713, n16714, n16715, n16716,
    n16718, n16719, n16720, n16721, n16722, n16724, n16725, n16726, n16727,
    n16728, n16730, n16731, n16732, n16733, n16734, n16736, n16737, n16738,
    n16739, n16740, n16742, n16743, n16745, n16746, n16747, n16748, n16749,
    n16751, n16752, n16753, n16754, n16755, n16757, n16758, n16759, n16760,
    n16761, n16763, n16764, n16765, n16766, n16767, n16769, n16770, n16771,
    n16772, n16773, n16775, n16776, n16777, n16778, n16779, n16781, n16782,
    n16783, n16784, n16785, n16787, n16788, n16789, n16790, n16791, n16793,
    n16794, n16795, n16796, n16797, n16799, n16800, n16801, n16802, n16803,
    n16805, n16806, n16807, n16809, n16810, n16811, n16812, n16813, n16815,
    n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
    n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16833, n16834,
    n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
    n16844, n16845, n16846, n16847, n16848, n16849, n16851, n16852, n16853,
    n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16869, n16870, n16872, n16873,
    n16875, n16876, n16878, n16879, n16881, n16882, n16884, n16885, n16887,
    n16888, n16890, n16891, n16893, n16894, n16896, n16897, n16899, n16900,
    n16902, n16903, n16905, n16906, n16908, n16909, n16911, n16912, n16914,
    n16915, n16917, n16918, n16919, n16920, n16921, n16923, n16924, n16925,
    n16926, n16927, n16929, n16930, n16932, n16933, n16935, n16936, n16937,
    n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16953, n16954, n16955, n16956,
    n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
    n16966, n16967, n16968, n16969, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
    n17004, n17005, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
    n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
    n17023, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
    n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
    n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
    n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17061,
    n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
    n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17079, n17080,
    n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
    n17090, n17091, n17092, n17093, n17094, n17095, n17097, n17098, n17099,
    n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17115, n17116, n17117, n17118,
    n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17133, n17134, n17135, n17136, n17137,
    n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
    n17147, n17148, n17149, n17151, n17152, n17154, n17155, n17157, n17158,
    n17159, n17160, n17161, n17163, n17164, n17166, n17167, n17169, n17170,
    n17172, n17173, n17175, n17176, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17189, n17190, n17192, n17193, n17195,
    n17196, n17198, n17199, n17201, n17202, n17203, n17204, n17205, n17206,
    n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17231, n17232, n17233, n17234, n17235,
    n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
    n17245, n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
    n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
    n17293, n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
    n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
    n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17331, n17332,
    n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
    n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17367, n17368, n17369, n17370, n17371,
    n17372, n17373, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
    n17382, n17383, n17384, n17385, n17387, n17388, n17390, n17391, n17392,
    n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
    n17402, n17403, n17404, n17406, n17407, n17408, n17409, n17410, n17411,
    n17412, n17413, n17414, n17415, n17416, n17417, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
    n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
    n17441, n17442, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17457, n17458, n17459, n17460,
    n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17469, n17470,
    n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
    n17480, n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17490,
    n17491, n17492, n17493, n17494, n17495, n17496, n17498, n17500, n17502,
    n17503, n17504, n17505, n17506, n17507, n17509, n17510, n17511, n17512,
    n17513, n17514, n17516, n17517, n17518, n17519, n17520, n17521, n17523,
    n17524, n17525, n17527, n17528, n17529, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17539, n17540, n17541, n17543, n17544, n17546,
    n17547, n17549, n17550, n17552, n17553, n17555, n17556, n17558, n17561,
    n17562, n17564, n17565, n17567, n17568, n17570, n17571, n17573, n17574,
    n17575, n17576, n17577, n17578, n17579, n17581, n17583, n17587, n17589,
    n17590, n17591, n17592, n17594, n17595, n17596, n17597, n17598, n17599,
    n17600, n17601, n17602, n17603, n17605, n17606, n17607, n17608, n17609,
    n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
    n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
    n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660, n17662, n17664, n17665,
    n17667, n17669, n17671, n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17683, n17684, n17685, n17686, n17687, n17688,
    n17689, n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
    n17700, n17701, n17702, n17703, n17704, n17705, n17707, n17708, n17710,
    n17711, n17713, n17714, n17716, n17717, n17719, n17720, n17722, n17723,
    n17724, n17726, n17728, n17730, n17732, n17734, n17736, n17738, n17740,
    n17742, n17744, n17746, n17748, n17750, n17752, n17754, n17755, n17757,
    n17758, n17760, n17761, n17763, n17764, n17766, n17768, n17769, n17771,
    n17772, n17774, n17775, n17776, n17778, n17779, n17780, n17781, n17782,
    n17783, n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
    n17803, n17805, n17807, n17808, n17809, n17811, n17812, n17813, n17815,
    n17816, n17818, n17819, n17820, n17822, n17823, n17824, n17825, n17826,
    n17827, n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17837,
    n17838, n17839, n17840, n17841, n17842, n17845, n17846, n17848, n17849,
    n17850, n17851, n17852, n17853, n17855, n17856, n17857, n17858, n17859,
    n17860, n17862, n17863, n17864, n17865, n17866, n17867, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17879, n17880,
    n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17889, n17890,
    n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17909, n17910,
    n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
    n17922, n17923, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17934, n17935, n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17946, n17947, n17948, n17950, n17951, n17952, n17954,
    n17955, n17956, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
    n17965, n17966, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
    n17997, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18007,
    n18008, n18009, n18010, n18011, n18012, n18014, n18015, n18016, n18017,
    n18018, n18019, n18021, n18022, n18023, n18024, n18025, n18026, n18028,
    n18029, n18030, n18031, n18032, n18033, n18035, n18036, n18037, n18038,
    n18039, n18040, n18042, n18043, n18044, n18045, n18046, n18047, n18049,
    n18050, n18051, n18052, n18053, n18054, n18056, n18057, n18058, n18059,
    n18060, n18061, n18063, n18064, n18065, n18066, n18067, n18068, n18070,
    n18071, n18073, n18075, n18076, n18077, n18079, n18080, n18081, n18082,
    n18084, n18086, n18087, n18088, n18090, n18091, n18092, n18093, n18094,
    n18095, n18097, n18098, n18099, n18100, n18101, n18102, n18104, n18105,
    n18106, n18107, n18108, n18109, n18111, n18112, n18113, n18114, n18115,
    n18116, n18118, n18119, n18120, n18121, n18122, n18123, n18125, n18126,
    n18127, n18128, n18129, n18130, n18132, n18133, n18134, n18135, n18136,
    n18137, n18139, n18140, n18141, n18142, n18143, n18144, n18146, n18147,
    n18148, n18149, n18150, n18151, n18153, n18154, n18155, n18156, n18157,
    n18158, n18160, n18161, n18162, n18163, n18164, n18165, n18167, n18168,
    n18169, n18170, n18171, n18172, n18174, n18175, n18176, n18177, n18178,
    n18179, n18181, n18182, n18183, n18184, n18185, n18186, n18188, n18189,
    n18190, n18191, n18192, n18193, n18195, n18196, n18197, n18198, n18199,
    n18200, n18202, n18203, n18204, n18205, n18206, n18207, n18209, n18211,
    n18212, n18213, n18214, n18216, n18217, n18218, n18219, n18220, n18222,
    n18223, n18224, n18226, n18227, n18228, n18230, n18231, n18233, n18234,
    n18235, n18236, n18237, n18238, n18239, n18241, n18242, n18243, n18244,
    n18245, n18246, n18248, n18249, n18250, n18251, n18252, n18253, n18255,
    n18256, n18257, n18258, n18259, n18260, n18262, n18263, n18264, n18265,
    n18266, n18267, n18269, n18270, n18271, n18272, n18273, n18274, n18276,
    n18277, n18278, n18279, n18280, n18281, n18283, n18284, n18285, n18286,
    n18287, n18288, n18290, n18291, n18292, n18293, n18294, n18295, n18297,
    n18298, n18299, n18300, n18301, n18302, n18304, n18305, n18306, n18307,
    n18308, n18309, n18311, n18312, n18313, n18314, n18315, n18316, n18318,
    n18319, n18320, n18321, n18322, n18323, n18325, n18326, n18327, n18328,
    n18329, n18330, n18332, n18333, n18334, n18335, n18336, n18337, n18339,
    n18340, n18341, n18342, n18343, n18344, n18346, n18347, n18348, n18349,
    n18350, n18351, n18353, n18354, n18355, n18356, n18357, n18358, n18360,
    n18361, n18362, n18363, n18364, n18365, n18367, n18368, n18369, n18370,
    n18371, n18372, n18374, n18375, n18376, n18377, n18378, n18379, n18381,
    n18382, n18383, n18384, n18385, n18386, n18388, n18389, n18390, n18391,
    n18392, n18393, n18395, n18396, n18397, n18398, n18399, n18400, n18402,
    n18403, n18404, n18405, n18406, n18407, n18409, n18410, n18411, n18412,
    n18413, n18414, n18416, n18417, n18418, n18419, n18420, n18421, n18423,
    n18424, n18425, n18426, n18427, n18428, n18430, n18431, n18432, n18433,
    n18434, n18435, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
    n18445, n18446, n18447, n18448, n18449, n18450, n18452, n18453, n18454,
    n18455, n18456, n18457, n18459, n18460, n18461, n18462, n18463, n18464,
    n18466, n18467, n18468, n18469, n18470, n18471, n18473, n18474, n18475,
    n18476, n18477, n18478, n18480, n18481, n18482, n18483, n18484, n18485,
    n18487, n18488, n18489, n18490, n18491, n18492, n18494, n18495, n18496,
    n18497, n18498, n18499, n18501, n18502, n18503, n18504, n18505, n18506,
    n18508, n18509, n18510, n18511, n18512, n18513, n18515, n18516, n18517,
    n18518, n18519, n18520, n18522, n18523, n18524, n18525, n18526, n18527,
    n18529, n18530, n18531, n18532, n18533, n18534, n18536, n18537, n18538,
    n18539, n18540, n18541, n18543, n18544, n18545, n18546, n18547, n18548,
    n18550, n18551, n18552, n18553, n18554, n18555, n18557, n18558, n18559,
    n18560, n18561, n18562, n18564, n18565, n18566, n18567, n18568, n18569,
    n18571, n18572, n18573, n18574, n18575, n18576, n18578, n18579, n18580,
    n18581, n18582, n18583, n18585, n18586, n18587, n18588, n18589, n18590,
    n18592, n18593, n18594, n18595, n18596, n18597, n18599, n18600, n18601,
    n18602, n18603, n18604, n18606, n18607, n18608, n18609, n18610, n18611,
    n18613, n18614, n18615, n18616, n18617, n18618, n18620, n18621, n18622,
    n18623, n18624, n18625, n18627, n18628, n18629, n18630, n18631, n18632,
    n18634, n18635, n18636, n18637, n18638, n18639, n18641, n18642, n18643,
    n18644, n18645, n18646, n18648, n18649, n18650, n18651, n18652, n18653,
    n18655, n18656, n18657, n18658, n18659, n18660, n18662, n18663, n18664,
    n18665, n18666, n18667, n18669, n18670, n18671, n18672, n18673, n18674,
    n18676, n18677, n18678, n18679, n18680, n18681, n18683, n18684, n18685,
    n18686, n18687, n18688, n18690, n18691, n18692, n18693, n18694, n18695,
    n18697, n18698, n18699, n18700, n18701, n18702, n18704, n18705, n18706,
    n18707, n18708, n18709, n18711, n18712, n18713, n18714, n18715, n18716,
    n18718, n18720, n18722, n18723, n18725, n18726, n18728, n18729, n18731,
    n18732, n18734, n18735, n18737, n18738, n18740, n18741, n18743, n18744,
    n18746, n18747, n18749, n18750, n18752, n18753, n18755, n18756, n18758,
    n18759, n18761, n18762, n18764, n18765, n18767, n18768, n18770, n18771,
    n18773;
  assign po0035 = pi0880 | pi2019;
  assign n4508 = pi0888 & ~pi2032;
  assign n4509 = ~pi0889 & ~pi0903;
  assign n4510 = ~pi0884 & ~pi0885;
  assign n4511 = n4509 & n4510;
  assign n4512 = ~pi2032 & ~n4511;
  assign n4513 = pi0001 & pi2032;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~pi0879 & ~pi0887;
  assign n4516 = ~pi0886 & n4515;
  assign n4517 = ~pi2032 & ~n4516;
  assign n4518 = n4514 & ~n4517;
  assign po0048 = n4508 | ~n4518;
  assign n4520 = pi0889 & ~pi2032;
  assign n4521 = pi0002 & pi2032;
  assign po0049 = n4520 | n4521;
  assign n4523 = pi0903 & ~pi2032;
  assign n4524 = pi0003 & pi2032;
  assign po0050 = n4523 | n4524;
  assign n4526 = pi0884 & ~pi2032;
  assign n4527 = pi0004 & pi2032;
  assign po0051 = n4526 | n4527;
  assign n4529 = pi0885 & ~pi2032;
  assign n4530 = pi0005 & pi2032;
  assign po0052 = n4529 | n4530;
  assign po0053 = pi0006 & pi2032;
  assign n4533 = pi0886 & ~pi2032;
  assign n4534 = pi0007 & pi2032;
  assign po0054 = n4533 | n4534;
  assign n4536 = pi0887 & ~pi2032;
  assign n4537 = pi0008 & pi2032;
  assign po0055 = n4536 | n4537;
  assign n4539 = pi0879 & ~pi2032;
  assign n4540 = pi0009 & pi2032;
  assign po0056 = n4539 | n4540;
  assign n4542 = pi0010 & pi2032;
  assign po0057 = n4508 | n4542;
  assign po0058 = pi0011 & pi2032;
  assign po0059 = pi0012 & pi2032;
  assign po0060 = pi0013 & pi2032;
  assign po0061 = pi0014 & pi2032;
  assign po0062 = pi0015 & pi2032;
  assign po0063 = pi0016 & pi2032;
  assign n4550 = pi1144 & ~pi2032;
  assign n4551 = pi0017 & pi2032;
  assign po0064 = n4550 | n4551;
  assign n4553 = pi1012 & ~pi2032;
  assign n4554 = pi0018 & pi2032;
  assign po0065 = n4553 | n4554;
  assign n4556 = pi1143 & ~pi2032;
  assign n4557 = pi0019 & pi2032;
  assign po0066 = n4556 | n4557;
  assign n4559 = pi1142 & ~pi2032;
  assign n4560 = pi0020 & pi2032;
  assign po0067 = n4559 | n4560;
  assign n4562 = pi1141 & ~pi2032;
  assign n4563 = pi0021 & pi2032;
  assign po0068 = n4562 | n4563;
  assign n4565 = pi1771 & ~pi2032;
  assign n4566 = pi0022 & pi2032;
  assign po0069 = n4565 | n4566;
  assign n4568 = pi1140 & ~pi2032;
  assign n4569 = pi0023 & pi2032;
  assign po0070 = n4568 | n4569;
  assign n4571 = pi1139 & ~pi2032;
  assign n4572 = pi0024 & pi2032;
  assign po0071 = n4571 | n4572;
  assign po0072 = pi0025 & pi2032;
  assign po0073 = pi0026 & pi2032;
  assign po0074 = pi0027 & pi2032;
  assign po0075 = pi0028 & pi2032;
  assign po0076 = pi0029 & pi2032;
  assign po0077 = pi0030 & pi2032;
  assign po0078 = pi0031 & pi2032;
  assign po0079 = pi0032 & pi2032;
  assign po0080 = pi0033 & pi2032;
  assign po0081 = pi0034 & pi2032;
  assign po0082 = pi0035 & pi2032;
  assign po0083 = pi0036 & pi2032;
  assign n4586 = ~pi1217 & ~pi2032;
  assign n4587 = pi0037 & pi2032;
  assign po0084 = n4586 | n4587;
  assign n4589 = ~pi1129 & ~pi2032;
  assign n4590 = pi0038 & pi2032;
  assign po0085 = n4589 | n4590;
  assign n4592 = ~pi1216 & ~pi2032;
  assign n4593 = pi0039 & pi2032;
  assign po0086 = n4592 | n4593;
  assign n4595 = ~pi1215 & ~pi2032;
  assign n4596 = pi0040 & pi2032;
  assign po0087 = n4595 | n4596;
  assign n4598 = ~pi1214 & ~pi2032;
  assign n4599 = pi0041 & pi2032;
  assign po0088 = n4598 | n4599;
  assign n4601 = ~pi1213 & ~pi2032;
  assign n4602 = pi0042 & pi2032;
  assign po0089 = n4601 | n4602;
  assign n4604 = ~pi1126 & ~pi2032;
  assign n4605 = pi0043 & pi2032;
  assign po0090 = n4604 | n4605;
  assign n4607 = ~pi1223 & ~pi2032;
  assign n4608 = pi0044 & pi2032;
  assign po0091 = n4607 | n4608;
  assign n4610 = ~pi1756 & ~pi2032;
  assign n4611 = pi0045 & pi2032;
  assign po0092 = n4610 | n4611;
  assign n4613 = ~pi1222 & ~pi2032;
  assign n4614 = pi0046 & pi2032;
  assign po0093 = n4613 | n4614;
  assign n4616 = ~pi1221 & ~pi2032;
  assign n4617 = pi0047 & pi2032;
  assign po0094 = n4616 | n4617;
  assign n4619 = ~pi1220 & ~pi2032;
  assign n4620 = pi0048 & pi2032;
  assign po0095 = n4619 | n4620;
  assign n4622 = ~pi1125 & ~pi2032;
  assign n4623 = pi0049 & pi2032;
  assign po0096 = n4622 | n4623;
  assign n4625 = ~pi1219 & ~pi2032;
  assign n4626 = pi0050 & pi2032;
  assign po0097 = n4625 | n4626;
  assign n4628 = ~pi1218 & ~pi2032;
  assign n4629 = pi0051 & pi2032;
  assign po0098 = n4628 | n4629;
  assign n4631 = ~pi1212 & ~pi2032;
  assign n4632 = pi0052 & pi2032;
  assign po0099 = n4631 | n4632;
  assign po0100 = pi0053 & pi2032;
  assign po0101 = pi0054 & pi2032;
  assign po0102 = pi0055 & pi2032;
  assign po0103 = pi0056 & pi2032;
  assign n4638 = ~pi0305 & ~pi2032;
  assign n4639 = pi0057 & pi2032;
  assign po0104 = n4638 | n4639;
  assign n4641 = ~pi0303 & ~pi2032;
  assign n4642 = pi0058 & pi2032;
  assign po0105 = n4641 | n4642;
  assign n4644 = ~pi0302 & ~pi2032;
  assign n4645 = pi0059 & pi2032;
  assign po0106 = n4644 | n4645;
  assign n4647 = ~pi0301 & ~pi2032;
  assign n4648 = pi0060 & pi2032;
  assign po0107 = n4647 | n4648;
  assign n4650 = ~pi0300 & ~pi2032;
  assign n4651 = pi0061 & pi2032;
  assign po0108 = n4650 | n4651;
  assign n4653 = ~pi0299 & ~pi2032;
  assign n4654 = pi0062 & pi2032;
  assign po0109 = n4653 | n4654;
  assign n4656 = ~pi0298 & ~pi2032;
  assign n4657 = pi0063 & pi2032;
  assign po0110 = n4656 | n4657;
  assign n4659 = ~pi0308 & ~pi2032;
  assign n4660 = pi0064 & pi2032;
  assign po0111 = n4659 | n4660;
  assign n4662 = ~pi0297 & ~pi2032;
  assign n4663 = pi0065 & pi2032;
  assign po0112 = n4662 | n4663;
  assign n4665 = ~pi0296 & ~pi2032;
  assign n4666 = pi0066 & pi2032;
  assign po0113 = n4665 | n4666;
  assign n4668 = ~pi0321 & ~pi2032;
  assign n4669 = pi0067 & pi2032;
  assign po0114 = n4668 | n4669;
  assign n4671 = ~pi0317 & ~pi2032;
  assign n4672 = pi0068 & pi2032;
  assign po0115 = n4671 | n4672;
  assign n4674 = ~pi0315 & ~pi2032;
  assign n4675 = pi0069 & pi2032;
  assign po0116 = n4674 | n4675;
  assign n4677 = ~pi0313 & ~pi2032;
  assign n4678 = pi0070 & pi2032;
  assign po0117 = n4677 | n4678;
  assign n4680 = ~pi0319 & ~pi2032;
  assign n4681 = pi0071 & pi2032;
  assign po0118 = n4680 | n4681;
  assign n4683 = ~pi0311 & ~pi2032;
  assign n4684 = pi0072 & pi2032;
  assign po0119 = n4683 | n4684;
  assign n4686 = ~pi0245 & ~pi2032;
  assign n4687 = pi0073 & pi2032;
  assign po0120 = n4686 | n4687;
  assign n4689 = ~pi0244 & ~pi2032;
  assign n4690 = pi0074 & pi2032;
  assign po0121 = n4689 | n4690;
  assign n4692 = ~pi0258 & ~pi2032;
  assign n4693 = pi0075 & pi2032;
  assign po0122 = n4692 | n4693;
  assign n4695 = ~pi0256 & ~pi2032;
  assign n4696 = pi0076 & pi2032;
  assign po0123 = n4695 | n4696;
  assign n4698 = ~pi0421 & ~pi2032;
  assign n4699 = pi0077 & pi2032;
  assign po0124 = n4698 | n4699;
  assign n4701 = ~pi0419 & ~pi2032;
  assign n4702 = pi0078 & pi2032;
  assign po0125 = n4701 | n4702;
  assign n4704 = ~pi0422 & ~pi2032;
  assign n4705 = pi0079 & pi2032;
  assign po0126 = n4704 | n4705;
  assign n4707 = ~pi0417 & ~pi2032;
  assign n4708 = pi0080 & pi2032;
  assign po0127 = n4707 | n4708;
  assign n4710 = ~pi0416 & ~pi2032;
  assign n4711 = pi0081 & pi2032;
  assign po0128 = n4710 | n4711;
  assign n4713 = ~pi0415 & ~pi2032;
  assign n4714 = pi0082 & pi2032;
  assign po0129 = n4713 | n4714;
  assign n4716 = ~pi0414 & ~pi2032;
  assign n4717 = pi0083 & pi2032;
  assign po0130 = n4716 | n4717;
  assign n4719 = ~pi0420 & ~pi2032;
  assign n4720 = pi0084 & pi2032;
  assign po0131 = n4719 | n4720;
  assign n4722 = ~pi0418 & ~pi2032;
  assign n4723 = pi0085 & pi2032;
  assign po0132 = n4722 | n4723;
  assign n4725 = ~pi0413 & ~pi2032;
  assign n4726 = pi0086 & pi2032;
  assign po0133 = n4725 | n4726;
  assign n4728 = ~pi0427 & ~pi2032;
  assign n4729 = pi0087 & pi2032;
  assign po0134 = n4728 | n4729;
  assign n4731 = ~pi0426 & ~pi2032;
  assign n4732 = pi0088 & pi2032;
  assign po0135 = n4731 | n4732;
  assign n4734 = ~pi0425 & ~pi2032;
  assign n4735 = pi0089 & pi2032;
  assign po0136 = n4734 | n4735;
  assign n4737 = ~pi0424 & ~pi2032;
  assign n4738 = pi0090 & pi2032;
  assign po0137 = n4737 | n4738;
  assign n4740 = ~pi0423 & ~pi2032;
  assign n4741 = pi0091 & pi2032;
  assign po0138 = n4740 | n4741;
  assign n4743 = ~pi0345 & ~pi2032;
  assign n4744 = pi0092 & pi2032;
  assign po0139 = n4743 | n4744;
  assign n4746 = ~pi0337 & ~pi2032;
  assign n4747 = pi0093 & pi2032;
  assign po0140 = n4746 | n4747;
  assign n4749 = ~pi0340 & ~pi2032;
  assign n4750 = pi0094 & pi2032;
  assign po0141 = n4749 | n4750;
  assign n4752 = ~pi0351 & ~pi2032;
  assign n4753 = pi0095 & pi2032;
  assign po0142 = n4752 | n4753;
  assign n4755 = ~pi0352 & ~pi2032;
  assign n4756 = pi0096 & pi2032;
  assign po0143 = n4755 | n4756;
  assign po0144 = pi0097 & pi2032;
  assign po0145 = pi0098 & pi2032;
  assign po0146 = pi0099 & pi2032;
  assign po0147 = pi0100 & pi2032;
  assign po0148 = pi0101 & pi2032;
  assign po0149 = pi0102 & pi2032;
  assign po0150 = pi0103 & pi2032;
  assign po0151 = pi0104 & pi2032;
  assign po0152 = pi0105 & pi2032;
  assign po0153 = pi0106 & pi2032;
  assign po0154 = pi0107 & pi2032;
  assign po0155 = pi0108 & pi2032;
  assign po0156 = pi0109 & pi2032;
  assign po0157 = pi0110 & pi2032;
  assign po0158 = pi0111 & pi2032;
  assign po0159 = pi0112 & pi2032;
  assign po0160 = pi0113 & pi2032;
  assign po0161 = pi0114 & pi2032;
  assign po0162 = pi0115 & pi2032;
  assign po0163 = pi0116 & pi2032;
  assign n4778 = ~pi0435 & ~pi2032;
  assign n4779 = pi0117 & pi2032;
  assign po0164 = n4778 | n4779;
  assign n4781 = ~pi0434 & ~pi2032;
  assign n4782 = pi0118 & pi2032;
  assign po0165 = n4781 | n4782;
  assign n4784 = ~pi0455 & ~pi2032;
  assign n4785 = pi0119 & pi2032;
  assign po0166 = n4784 | n4785;
  assign n4787 = ~pi0433 & ~pi2032;
  assign n4788 = pi0120 & pi2032;
  assign po0167 = n4787 | n4788;
  assign n4790 = ~pi0432 & ~pi2032;
  assign n4791 = pi0121 & pi2032;
  assign po0168 = n4790 | n4791;
  assign n4793 = ~pi0431 & ~pi2032;
  assign n4794 = pi0122 & pi2032;
  assign po0169 = n4793 | n4794;
  assign n4796 = ~pi0457 & ~pi2032;
  assign n4797 = pi0123 & pi2032;
  assign po0170 = n4796 | n4797;
  assign n4799 = ~pi0430 & ~pi2032;
  assign n4800 = pi0124 & pi2032;
  assign po0171 = n4799 | n4800;
  assign n4802 = ~pi0429 & ~pi2032;
  assign n4803 = pi0125 & pi2032;
  assign po0172 = n4802 | n4803;
  assign n4805 = ~pi0428 & ~pi2032;
  assign n4806 = pi0126 & pi2032;
  assign po0173 = n4805 | n4806;
  assign n4808 = ~pi0440 & ~pi2032;
  assign n4809 = pi0127 & pi2032;
  assign po0174 = n4808 | n4809;
  assign n4811 = ~pi0439 & ~pi2032;
  assign n4812 = pi0128 & pi2032;
  assign po0175 = n4811 | n4812;
  assign n4814 = ~pi0454 & ~pi2032;
  assign n4815 = pi0129 & pi2032;
  assign po0176 = n4814 | n4815;
  assign n4817 = ~pi0438 & ~pi2032;
  assign n4818 = pi0130 & pi2032;
  assign po0177 = n4817 | n4818;
  assign n4820 = ~pi0437 & ~pi2032;
  assign n4821 = pi0131 & pi2032;
  assign po0178 = n4820 | n4821;
  assign n4823 = ~pi0436 & ~pi2032;
  assign n4824 = pi0132 & pi2032;
  assign po0179 = n4823 | n4824;
  assign n4826 = ~pi0338 & ~pi2032;
  assign n4827 = pi0133 & pi2032;
  assign po0180 = n4826 | n4827;
  assign n4829 = ~pi0339 & ~pi2032;
  assign n4830 = pi0134 & pi2032;
  assign po0181 = n4829 | n4830;
  assign n4832 = ~pi0350 & ~pi2032;
  assign n4833 = pi0135 & pi2032;
  assign po0182 = n4832 | n4833;
  assign n4835 = ~pi0349 & ~pi2032;
  assign n4836 = pi0136 & pi2032;
  assign po0183 = n4835 | n4836;
  assign n4838 = ~pi0271 & ~pi2032;
  assign n4839 = pi0137 & pi2032;
  assign po0184 = n4838 | n4839;
  assign n4841 = ~pi0270 & ~pi2032;
  assign n4842 = pi0138 & pi2032;
  assign po0185 = n4841 | n4842;
  assign n4844 = ~pi0273 & ~pi2032;
  assign n4845 = pi0139 & pi2032;
  assign po0186 = n4844 | n4845;
  assign n4847 = ~pi0272 & ~pi2032;
  assign n4848 = pi0140 & pi2032;
  assign po0187 = n4847 | n4848;
  assign n4850 = ~pi0267 & ~pi2032;
  assign n4851 = pi0141 & pi2032;
  assign po0188 = n4850 | n4851;
  assign n4853 = ~pi0266 & ~pi2032;
  assign n4854 = pi0142 & pi2032;
  assign po0189 = n4853 | n4854;
  assign n4856 = ~pi0265 & ~pi2032;
  assign n4857 = pi0143 & pi2032;
  assign po0190 = n4856 | n4857;
  assign n4859 = ~pi0264 & ~pi2032;
  assign n4860 = pi0144 & pi2032;
  assign po0191 = n4859 | n4860;
  assign n4862 = ~pi0269 & ~pi2032;
  assign n4863 = pi0145 & pi2032;
  assign po0192 = n4862 | n4863;
  assign n4865 = ~pi0268 & ~pi2032;
  assign n4866 = pi0146 & pi2032;
  assign po0193 = n4865 | n4866;
  assign n4868 = ~pi0279 & ~pi2032;
  assign n4869 = pi0147 & pi2032;
  assign po0194 = n4868 | n4869;
  assign n4871 = ~pi0278 & ~pi2032;
  assign n4872 = pi0148 & pi2032;
  assign po0195 = n4871 | n4872;
  assign n4874 = ~pi0277 & ~pi2032;
  assign n4875 = pi0149 & pi2032;
  assign po0196 = n4874 | n4875;
  assign n4877 = ~pi0276 & ~pi2032;
  assign n4878 = pi0150 & pi2032;
  assign po0197 = n4877 | n4878;
  assign n4880 = ~pi0275 & ~pi2032;
  assign n4881 = pi0151 & pi2032;
  assign po0198 = n4880 | n4881;
  assign n4883 = ~pi0274 & ~pi2032;
  assign n4884 = pi0152 & pi2032;
  assign po0199 = n4883 | n4884;
  assign n4886 = ~pi0241 & ~pi2032;
  assign n4887 = pi0153 & pi2032;
  assign po0200 = n4886 | n4887;
  assign n4889 = ~pi0240 & ~pi2032;
  assign n4890 = pi0154 & pi2032;
  assign po0201 = n4889 | n4890;
  assign n4892 = ~pi0253 & ~pi2032;
  assign n4893 = pi0155 & pi2032;
  assign po0202 = n4892 | n4893;
  assign n4895 = ~pi0252 & ~pi2032;
  assign n4896 = pi0156 & pi2032;
  assign po0203 = n4895 | n4896;
  assign n4898 = ~pi0287 & ~pi2032;
  assign n4899 = pi0157 & pi2032;
  assign po0204 = n4898 | n4899;
  assign n4901 = ~pi0289 & ~pi2032;
  assign n4902 = pi0158 & pi2032;
  assign po0205 = n4901 | n4902;
  assign n4904 = ~pi0285 & ~pi2032;
  assign n4905 = pi0159 & pi2032;
  assign po0206 = n4904 | n4905;
  assign n4907 = ~pi0288 & ~pi2032;
  assign n4908 = pi0160 & pi2032;
  assign po0207 = n4907 | n4908;
  assign n4910 = ~pi0286 & ~pi2032;
  assign n4911 = pi0161 & pi2032;
  assign po0208 = n4910 | n4911;
  assign n4913 = ~pi0284 & ~pi2032;
  assign n4914 = pi0162 & pi2032;
  assign po0209 = n4913 | n4914;
  assign n4916 = ~pi0283 & ~pi2032;
  assign n4917 = pi0163 & pi2032;
  assign po0210 = n4916 | n4917;
  assign n4919 = ~pi0282 & ~pi2032;
  assign n4920 = pi0164 & pi2032;
  assign po0211 = n4919 | n4920;
  assign n4922 = ~pi0281 & ~pi2032;
  assign n4923 = pi0165 & pi2032;
  assign po0212 = n4922 | n4923;
  assign n4925 = ~pi0280 & ~pi2032;
  assign n4926 = pi0166 & pi2032;
  assign po0213 = n4925 | n4926;
  assign n4928 = ~pi0295 & ~pi2032;
  assign n4929 = pi0167 & pi2032;
  assign po0214 = n4928 | n4929;
  assign n4931 = ~pi0294 & ~pi2032;
  assign n4932 = pi0168 & pi2032;
  assign po0215 = n4931 | n4932;
  assign n4934 = ~pi0293 & ~pi2032;
  assign n4935 = pi0169 & pi2032;
  assign po0216 = n4934 | n4935;
  assign n4937 = ~pi0292 & ~pi2032;
  assign n4938 = pi0170 & pi2032;
  assign po0217 = n4937 | n4938;
  assign n4940 = ~pi0291 & ~pi2032;
  assign n4941 = pi0171 & pi2032;
  assign po0218 = n4940 | n4941;
  assign n4943 = ~pi0290 & ~pi2032;
  assign n4944 = pi0172 & pi2032;
  assign po0219 = n4943 | n4944;
  assign n4946 = ~pi0243 & ~pi2032;
  assign n4947 = pi0173 & pi2032;
  assign po0220 = n4946 | n4947;
  assign n4949 = ~pi0242 & ~pi2032;
  assign n4950 = pi0174 & pi2032;
  assign po0221 = n4949 | n4950;
  assign n4952 = ~pi0255 & ~pi2032;
  assign n4953 = pi0175 & pi2032;
  assign po0222 = n4952 | n4953;
  assign n4955 = ~pi0254 & ~pi2032;
  assign n4956 = pi0176 & pi2032;
  assign po0223 = n4955 | n4956;
  assign n4958 = ~pi0320 & ~pi2032;
  assign n4959 = pi0177 & pi2032;
  assign po0224 = n4958 | n4959;
  assign n4961 = ~pi0316 & ~pi2032;
  assign n4962 = pi0178 & pi2032;
  assign po0225 = n4961 | n4962;
  assign n4964 = ~pi0314 & ~pi2032;
  assign n4965 = pi0179 & pi2032;
  assign po0226 = n4964 | n4965;
  assign n4967 = ~pi0312 & ~pi2032;
  assign n4968 = pi0180 & pi2032;
  assign po0227 = n4967 | n4968;
  assign n4970 = ~pi0318 & ~pi2032;
  assign n4971 = pi0181 & pi2032;
  assign po0228 = n4970 | n4971;
  assign n4973 = ~pi0310 & ~pi2032;
  assign n4974 = pi0182 & pi2032;
  assign po0229 = n4973 | n4974;
  assign n4976 = ~pi0309 & ~pi2032;
  assign n4977 = pi0183 & pi2032;
  assign po0230 = n4976 | n4977;
  assign n4979 = ~pi0307 & ~pi2032;
  assign n4980 = pi0184 & pi2032;
  assign po0231 = n4979 | n4980;
  assign n4982 = ~pi0306 & ~pi2032;
  assign n4983 = pi0185 & pi2032;
  assign po0232 = n4982 | n4983;
  assign n4985 = ~pi0304 & ~pi2032;
  assign n4986 = pi0186 & pi2032;
  assign po0233 = n4985 | n4986;
  assign n4988 = ~pi0327 & ~pi2032;
  assign n4989 = pi0187 & pi2032;
  assign po0234 = n4988 | n4989;
  assign n4991 = ~pi0326 & ~pi2032;
  assign n4992 = pi0188 & pi2032;
  assign po0235 = n4991 | n4992;
  assign n4994 = ~pi0325 & ~pi2032;
  assign n4995 = pi0189 & pi2032;
  assign po0236 = n4994 | n4995;
  assign n4997 = ~pi0324 & ~pi2032;
  assign n4998 = pi0200 & pi2032;
  assign po0237 = n4997 | n4998;
  assign n5000 = pi0209 & ~pi2056;
  assign n5001 = pi0190 & pi2056;
  assign po0238 = n5000 | n5001;
  assign n5003 = pi0209 & ~pi2059;
  assign n5004 = pi0191 & pi2059;
  assign po0239 = n5003 | n5004;
  assign n5006 = pi0209 & ~pi2057;
  assign n5007 = pi0192 & pi2057;
  assign po0240 = n5006 | n5007;
  assign n5009 = pi0209 & ~pi2058;
  assign n5010 = pi0193 & pi2058;
  assign po0241 = n5009 | n5010;
  assign n5012 = pi0228 & ~pi2056;
  assign n5013 = pi0194 & pi2056;
  assign po0242 = n5012 | n5013;
  assign n5015 = pi0228 & ~pi2059;
  assign n5016 = pi0195 & pi2059;
  assign po0243 = n5015 | n5016;
  assign n5018 = pi0228 & ~pi2057;
  assign n5019 = pi0196 & pi2057;
  assign po0244 = n5018 | n5019;
  assign n5021 = pi0228 & ~pi2058;
  assign n5022 = pi0197 & pi2058;
  assign po0245 = n5021 | n5022;
  assign n5024 = pi1035 & pi1168;
  assign n5025 = ~pi1903 & n5024;
  assign n5026 = ~pi1987 & n5024;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = ~pi2140 & n5024;
  assign n5029 = n5027 & ~n5028;
  assign n5030 = ~pi1166 & ~pi1167;
  assign n5031 = ~n5029 & n5030;
  assign n5032 = pi1166 & pi1167;
  assign n5033 = n5025 & n5032;
  assign n5034 = ~n5031 & ~n5033;
  assign n5035 = ~pi1987 & ~pi2140;
  assign n5036 = n5024 & n5035;
  assign n5037 = ~n5025 & ~n5036;
  assign n5038 = ~pi1166 & pi1167;
  assign n5039 = ~n5037 & n5038;
  assign n5040 = n5034 & ~n5039;
  assign n5041 = pi1166 & ~pi1167;
  assign n5042 = ~n5027 & n5041;
  assign n5043 = n5040 & ~n5042;
  assign po0380 = ~pi2247 & ~n5043;
  assign n5045 = pi0329 & po0380;
  assign n5046 = pi0198 & ~pi2247;
  assign po0249 = n5045 | n5046;
  assign n5048 = pi1176 & pi1181;
  assign n5049 = ~pi1904 & n5048;
  assign n5050 = ~pi2005 & n5048;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = ~pi2138 & n5048;
  assign n5053 = n5051 & ~n5052;
  assign n5054 = ~pi1179 & ~pi1180;
  assign n5055 = ~n5053 & n5054;
  assign n5056 = pi1179 & pi1180;
  assign n5057 = n5049 & n5056;
  assign n5058 = ~n5055 & ~n5057;
  assign n5059 = ~pi2005 & ~pi2138;
  assign n5060 = n5048 & n5059;
  assign n5061 = ~n5049 & ~n5060;
  assign n5062 = ~pi1179 & pi1180;
  assign n5063 = ~n5061 & n5062;
  assign n5064 = n5058 & ~n5063;
  assign n5065 = pi1179 & ~pi1180;
  assign n5066 = ~n5051 & n5065;
  assign n5067 = n5064 & ~n5066;
  assign po0381 = ~pi2249 & ~n5067;
  assign n5069 = pi0330 & po0381;
  assign n5070 = pi0199 & ~pi2249;
  assign po0250 = n5069 | n5070;
  assign n5072 = ~pi0323 & ~pi2032;
  assign n5073 = pi0328 & pi2032;
  assign po0251 = n5072 | n5073;
  assign n5075 = pi1164 & pi1185;
  assign n5076 = ~pi1907 & n5075;
  assign n5077 = ~pi2004 & n5075;
  assign n5078 = ~n5076 & ~n5077;
  assign n5079 = ~pi2139 & n5075;
  assign n5080 = n5078 & ~n5079;
  assign n5081 = ~pi1131 & ~pi1184;
  assign n5082 = ~n5080 & n5081;
  assign n5083 = pi1131 & pi1184;
  assign n5084 = n5076 & n5083;
  assign n5085 = ~n5082 & ~n5084;
  assign n5086 = ~pi2004 & ~pi2139;
  assign n5087 = n5075 & n5086;
  assign n5088 = ~n5076 & ~n5087;
  assign n5089 = ~pi1131 & pi1184;
  assign n5090 = ~n5088 & n5089;
  assign n5091 = n5085 & ~n5090;
  assign n5092 = pi1131 & ~pi1184;
  assign n5093 = ~n5078 & n5092;
  assign n5094 = n5091 & ~n5093;
  assign po0392 = ~pi2246 & ~n5094;
  assign n5096 = pi0341 & po0392;
  assign n5097 = pi0201 & ~pi2246;
  assign po0252 = n5096 | n5097;
  assign n5099 = pi1169 & pi1762;
  assign n5100 = ~pi1908 & n5099;
  assign n5101 = ~pi1988 & n5099;
  assign n5102 = ~n5100 & ~n5101;
  assign n5103 = ~pi2158 & n5099;
  assign n5104 = n5102 & ~n5103;
  assign n5105 = ~pi1173 & ~pi1174;
  assign n5106 = ~n5104 & n5105;
  assign n5107 = pi1173 & pi1174;
  assign n5108 = n5100 & n5107;
  assign n5109 = ~n5106 & ~n5108;
  assign n5110 = ~pi1988 & ~pi2158;
  assign n5111 = n5099 & n5110;
  assign n5112 = ~n5100 & ~n5111;
  assign n5113 = ~pi1173 & pi1174;
  assign n5114 = ~n5112 & n5113;
  assign n5115 = n5109 & ~n5114;
  assign n5116 = pi1173 & ~pi1174;
  assign n5117 = ~n5102 & n5116;
  assign n5118 = n5115 & ~n5117;
  assign po0393 = ~pi2248 & ~n5118;
  assign n5120 = pi0342 & po0393;
  assign n5121 = pi0202 & ~pi2248;
  assign po0253 = n5120 | n5121;
  assign n5123 = pi1839 & pi1848;
  assign n5124 = ~pi1909 & n5123;
  assign n5125 = ~pi2006 & n5123;
  assign n5126 = ~n5124 & ~n5125;
  assign n5127 = ~pi2141 & n5123;
  assign n5128 = n5126 & ~n5127;
  assign n5129 = ~pi1847 & ~pi1873;
  assign n5130 = ~n5128 & n5129;
  assign n5131 = pi1847 & pi1873;
  assign n5132 = n5124 & n5131;
  assign n5133 = ~n5130 & ~n5132;
  assign n5134 = ~pi2006 & ~pi2141;
  assign n5135 = n5123 & n5134;
  assign n5136 = ~n5124 & ~n5135;
  assign n5137 = pi1847 & ~pi1873;
  assign n5138 = ~n5136 & n5137;
  assign n5139 = n5133 & ~n5138;
  assign n5140 = ~pi1847 & pi1873;
  assign n5141 = ~n5126 & n5140;
  assign n5142 = n5139 & ~n5141;
  assign po0394 = ~pi2250 & ~n5142;
  assign n5144 = pi0343 & po0394;
  assign n5145 = pi0203 & ~pi2250;
  assign po0254 = n5144 | n5145;
  assign n5147 = pi1838 & pi1843;
  assign n5148 = ~pi1910 & n5147;
  assign n5149 = ~pi2007 & n5147;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~pi2159 & n5147;
  assign n5152 = n5150 & ~n5151;
  assign n5153 = ~pi1841 & ~pi1842;
  assign n5154 = ~n5152 & n5153;
  assign n5155 = pi1841 & pi1842;
  assign n5156 = n5148 & n5155;
  assign n5157 = ~n5154 & ~n5156;
  assign n5158 = ~pi2007 & ~pi2159;
  assign n5159 = n5147 & n5158;
  assign n5160 = ~n5148 & ~n5159;
  assign n5161 = ~pi1841 & pi1842;
  assign n5162 = ~n5160 & n5161;
  assign n5163 = n5157 & ~n5162;
  assign n5164 = pi1841 & ~pi1842;
  assign n5165 = ~n5150 & n5164;
  assign n5166 = n5163 & ~n5165;
  assign po0395 = ~pi2251 & ~n5166;
  assign n5168 = pi0344 & po0395;
  assign n5169 = pi0204 & ~pi2251;
  assign po0255 = n5168 | n5169;
  assign n5171 = pi0331 & ~pi2056;
  assign n5172 = pi0205 & pi2056;
  assign po0256 = n5171 | n5172;
  assign n5174 = pi0331 & ~pi2059;
  assign n5175 = pi0206 & pi2059;
  assign po0257 = n5174 | n5175;
  assign n5177 = pi0331 & ~pi2057;
  assign n5178 = pi0207 & pi2057;
  assign po0258 = n5177 | n5178;
  assign n5180 = pi0331 & ~pi2058;
  assign n5181 = pi0208 & pi2058;
  assign po0259 = n5180 | n5181;
  assign n5183 = pi0456 & ~pi2056;
  assign n5184 = pi0210 & pi2056;
  assign po0261 = n5183 | n5184;
  assign n5186 = pi0456 & ~pi2059;
  assign n5187 = pi0211 & pi2059;
  assign po0262 = n5186 | n5187;
  assign n5189 = pi0456 & ~pi2057;
  assign n5190 = pi0212 & pi2057;
  assign po0263 = n5189 | n5190;
  assign n5192 = pi0456 & ~pi2058;
  assign n5193 = pi0213 & pi2058;
  assign po0264 = n5192 | n5193;
  assign po1127 = pi0885 & pi1930;
  assign n5196 = ~pi1076 & po1127;
  assign n5197 = ~pi1020 & ~pi1165;
  assign n5198 = n5196 & ~n5197;
  assign n5199 = ~pi0214 & pi0236;
  assign n5200 = pi0214 & ~pi0236;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = n5198 & n5201;
  assign n5203 = n5196 & n5197;
  assign n5204 = ~pi0214 & ~n5198;
  assign n5205 = ~n5203 & ~n5204;
  assign n5206 = ~n5202 & n5205;
  assign n5207 = pi0214 & ~pi0353;
  assign n5208 = pi0353 & n5199;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = ~n5200 & n5209;
  assign n5211 = n5203 & ~n5210;
  assign n5212 = ~n5206 & ~n5211;
  assign po0265 = pi1035 & ~n5212;
  assign po1128 = pi0886 & pi1930;
  assign n5215 = ~pi1077 & po1128;
  assign n5216 = ~pi1171 & ~pi1789;
  assign n5217 = n5215 & ~n5216;
  assign n5218 = ~pi0215 & pi0238;
  assign n5219 = pi0215 & ~pi0238;
  assign n5220 = ~n5218 & ~n5219;
  assign n5221 = n5217 & n5220;
  assign n5222 = n5215 & n5216;
  assign n5223 = ~pi0215 & ~n5217;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5221 & n5224;
  assign n5226 = pi0215 & ~pi0354;
  assign n5227 = pi0354 & n5218;
  assign n5228 = ~n5226 & ~n5227;
  assign n5229 = ~n5219 & n5228;
  assign n5230 = n5222 & ~n5229;
  assign n5231 = ~n5225 & ~n5230;
  assign po0266 = pi1169 & ~n5231;
  assign po1131 = pi0888 & pi1930;
  assign n5234 = ~pi1080 & po1131;
  assign n5235 = ~pi1832 & ~pi1840;
  assign n5236 = n5234 & n5235;
  assign n5237 = n5234 & ~n5235;
  assign n5238 = ~pi0216 & pi0224;
  assign n5239 = pi0216 & ~pi0224;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241 = n5237 & ~n5240;
  assign n5242 = pi0216 & ~n5237;
  assign n5243 = ~n5241 & ~n5242;
  assign n5244 = ~n5236 & ~n5243;
  assign n5245 = pi0260 & n5238;
  assign n5246 = pi0216 & ~pi0260;
  assign n5247 = ~n5245 & ~n5246;
  assign n5248 = ~n5239 & n5247;
  assign n5249 = n5236 & ~n5248;
  assign n5250 = ~n5244 & ~n5249;
  assign po0267 = pi1838 & ~n5250;
  assign n5252 = pi0884 & ~pi1075;
  assign n5253 = pi1930 & n5252;
  assign n5254 = ~pi1130 & ~pi1183;
  assign n5255 = n5253 & n5254;
  assign n5256 = n5253 & ~n5254;
  assign n5257 = ~pi0217 & pi0225;
  assign n5258 = pi0217 & ~pi0225;
  assign n5259 = ~n5257 & ~n5258;
  assign n5260 = n5256 & ~n5259;
  assign n5261 = pi0217 & ~n5256;
  assign n5262 = ~n5260 & ~n5261;
  assign n5263 = ~n5255 & ~n5262;
  assign n5264 = pi0261 & n5257;
  assign n5265 = pi0217 & ~pi0261;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = ~n5258 & n5266;
  assign n5268 = n5255 & ~n5267;
  assign n5269 = ~n5263 & ~n5268;
  assign po0268 = pi1164 & ~n5269;
  assign po1129 = pi0887 & pi1930;
  assign n5272 = ~pi1078 & po1129;
  assign n5273 = ~pi1178 & ~pi1777;
  assign n5274 = n5272 & n5273;
  assign n5275 = n5272 & ~n5273;
  assign n5276 = ~pi0218 & pi0227;
  assign n5277 = pi0218 & ~pi0227;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = n5275 & ~n5278;
  assign n5280 = pi0218 & ~n5275;
  assign n5281 = ~n5279 & ~n5280;
  assign n5282 = ~n5274 & ~n5281;
  assign n5283 = pi0262 & n5276;
  assign n5284 = pi0218 & ~pi0262;
  assign n5285 = ~n5283 & ~n5284;
  assign n5286 = ~n5277 & n5285;
  assign n5287 = n5274 & ~n5286;
  assign n5288 = ~n5282 & ~n5287;
  assign po0269 = pi1176 & ~n5288;
  assign po1130 = pi0879 & pi1930;
  assign n5291 = ~pi1079 & po1130;
  assign n5292 = ~pi1845 & ~pi1846;
  assign n5293 = n5291 & n5292;
  assign n5294 = n5291 & ~n5292;
  assign n5295 = ~pi0219 & pi0226;
  assign n5296 = pi0219 & ~pi0226;
  assign n5297 = ~n5295 & ~n5296;
  assign n5298 = n5294 & ~n5297;
  assign n5299 = pi0219 & ~n5294;
  assign n5300 = ~n5298 & ~n5299;
  assign n5301 = ~n5293 & ~n5300;
  assign n5302 = pi0263 & n5295;
  assign n5303 = pi0219 & ~pi0263;
  assign n5304 = ~n5302 & ~n5303;
  assign n5305 = ~n5296 & n5304;
  assign n5306 = n5293 & ~n5305;
  assign n5307 = ~n5301 & ~n5306;
  assign po0270 = pi1839 & ~n5307;
  assign n5309 = pi0216 & pi0224;
  assign n5310 = pi0220 & ~n5309;
  assign n5311 = ~pi0220 & n5309;
  assign n5312 = ~n5310 & ~n5311;
  assign n5313 = n5237 & ~n5312;
  assign n5314 = pi0220 & ~n5237;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = ~n5236 & ~n5315;
  assign n5317 = ~pi0220 & pi0260;
  assign n5318 = n5309 & n5317;
  assign n5319 = pi0220 & ~pi0260;
  assign n5320 = ~n5318 & ~n5319;
  assign n5321 = ~n5310 & n5320;
  assign n5322 = n5236 & ~n5321;
  assign n5323 = ~n5316 & ~n5322;
  assign po0271 = pi1838 & ~n5323;
  assign n5325 = pi0217 & pi0225;
  assign n5326 = pi0221 & ~n5325;
  assign n5327 = ~pi0221 & n5325;
  assign n5328 = ~n5326 & ~n5327;
  assign n5329 = n5256 & ~n5328;
  assign n5330 = pi0221 & ~n5256;
  assign n5331 = ~n5329 & ~n5330;
  assign n5332 = ~n5255 & ~n5331;
  assign n5333 = ~pi0221 & pi0261;
  assign n5334 = n5325 & n5333;
  assign n5335 = pi0221 & ~pi0261;
  assign n5336 = ~n5334 & ~n5335;
  assign n5337 = ~n5326 & n5336;
  assign n5338 = n5255 & ~n5337;
  assign n5339 = ~n5332 & ~n5338;
  assign po0272 = pi1164 & ~n5339;
  assign n5341 = pi0218 & pi0227;
  assign n5342 = pi0222 & ~n5341;
  assign n5343 = ~pi0222 & n5341;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = n5275 & ~n5344;
  assign n5346 = pi0222 & ~n5275;
  assign n5347 = ~n5345 & ~n5346;
  assign n5348 = ~n5274 & ~n5347;
  assign n5349 = ~pi0222 & pi0262;
  assign n5350 = n5341 & n5349;
  assign n5351 = pi0222 & ~pi0262;
  assign n5352 = ~n5350 & ~n5351;
  assign n5353 = ~n5342 & n5352;
  assign n5354 = n5274 & ~n5353;
  assign n5355 = ~n5348 & ~n5354;
  assign po0273 = pi1176 & ~n5355;
  assign n5357 = pi0219 & pi0226;
  assign n5358 = pi0223 & ~n5357;
  assign n5359 = ~pi0223 & n5357;
  assign n5360 = ~n5358 & ~n5359;
  assign n5361 = n5294 & ~n5360;
  assign n5362 = pi0223 & ~n5294;
  assign n5363 = ~n5361 & ~n5362;
  assign n5364 = ~n5293 & ~n5363;
  assign n5365 = ~pi0223 & pi0263;
  assign n5366 = n5357 & n5365;
  assign n5367 = pi0223 & ~pi0263;
  assign n5368 = ~n5366 & ~n5367;
  assign n5369 = ~n5358 & n5368;
  assign n5370 = n5293 & ~n5369;
  assign n5371 = ~n5364 & ~n5370;
  assign po0274 = pi1839 & ~n5371;
  assign n5373 = ~pi0224 & n5237;
  assign n5374 = pi0224 & ~n5237;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = ~n5236 & ~n5375;
  assign n5377 = ~pi0224 & pi0260;
  assign n5378 = pi0224 & ~pi0260;
  assign n5379 = ~n5377 & ~n5378;
  assign n5380 = n5236 & ~n5379;
  assign n5381 = ~n5376 & ~n5380;
  assign po0275 = pi1838 & ~n5381;
  assign n5383 = pi0225 & ~pi0261;
  assign n5384 = ~pi0225 & pi0261;
  assign n5385 = ~n5383 & ~n5384;
  assign n5386 = n5255 & ~n5385;
  assign n5387 = ~pi0225 & n5256;
  assign n5388 = pi0225 & ~n5256;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = ~n5255 & ~n5389;
  assign n5391 = ~n5386 & ~n5390;
  assign po0276 = pi1164 & ~n5391;
  assign n5393 = ~pi0226 & n5294;
  assign n5394 = pi0226 & ~n5294;
  assign n5395 = ~n5393 & ~n5394;
  assign n5396 = ~n5293 & ~n5395;
  assign n5397 = pi0226 & ~pi0263;
  assign n5398 = ~pi0226 & pi0263;
  assign n5399 = ~n5397 & ~n5398;
  assign n5400 = n5293 & ~n5399;
  assign n5401 = ~n5396 & ~n5400;
  assign po0277 = pi1839 & ~n5401;
  assign n5403 = ~pi0227 & n5275;
  assign n5404 = pi0227 & ~n5275;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~n5274 & ~n5405;
  assign n5407 = pi0227 & ~pi0262;
  assign n5408 = ~pi0227 & pi0262;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = n5274 & ~n5409;
  assign n5411 = ~n5406 & ~n5410;
  assign po0278 = pi1176 & ~n5411;
  assign n5413 = ~pi0229 & ~pi0838;
  assign n5414 = pi2202 & pi2203;
  assign n5415 = ~pi2131 & ~pi2201;
  assign n5416 = n5414 & n5415;
  assign n5417 = pi2132 & n5416;
  assign n5418 = ~pi2239 & ~pi2240;
  assign n5419 = pi2241 & ~n5418;
  assign n5420 = ~pi2242 & ~n5419;
  assign n5421 = n5417 & n5420;
  assign n5422 = ~pi2238 & pi2239;
  assign n5423 = pi2240 & n5422;
  assign n5424 = ~pi2241 & n5423;
  assign n5425 = n5421 & n5424;
  assign po0280 = ~n5413 & ~n5425;
  assign n5427 = ~pi0230 & ~pi0839;
  assign po0281 = ~n5425 & ~n5427;
  assign n5429 = pi0640 & ~pi2059;
  assign n5430 = pi0231 & pi2059;
  assign po0282 = n5429 | n5430;
  assign n5432 = pi0232 & ~pi2060;
  assign n5433 = pi0640 & pi2060;
  assign po0283 = n5432 | n5433;
  assign n5435 = pi0640 & ~pi2058;
  assign n5436 = pi0233 & pi2058;
  assign po0284 = n5435 | n5436;
  assign n5438 = pi0640 & ~pi2056;
  assign n5439 = pi0234 & pi2056;
  assign po0285 = n5438 | n5439;
  assign n5441 = pi0640 & ~pi2057;
  assign n5442 = pi0235 & pi2057;
  assign po0286 = n5441 | n5442;
  assign n5444 = ~pi0236 & pi0353;
  assign n5445 = pi0236 & ~pi0353;
  assign n5446 = ~n5444 & ~n5445;
  assign n5447 = n5203 & ~n5446;
  assign n5448 = pi0236 & ~n5198;
  assign n5449 = ~pi0236 & n5198;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = ~n5203 & ~n5450;
  assign n5452 = ~n5447 & ~n5451;
  assign po0287 = pi1035 & ~n5452;
  assign n5454 = ~pi0237 & pi0353;
  assign n5455 = pi0214 & pi0236;
  assign n5456 = n5454 & n5455;
  assign n5457 = pi0237 & ~pi0353;
  assign n5458 = ~n5456 & ~n5457;
  assign n5459 = pi0237 & ~n5455;
  assign n5460 = n5458 & ~n5459;
  assign n5461 = n5203 & ~n5460;
  assign n5462 = pi0237 & ~n5198;
  assign n5463 = ~pi0237 & n5455;
  assign n5464 = ~n5459 & ~n5463;
  assign n5465 = n5198 & ~n5464;
  assign n5466 = ~n5462 & ~n5465;
  assign n5467 = ~n5203 & ~n5466;
  assign n5468 = ~n5461 & ~n5467;
  assign po0288 = pi1035 & ~n5468;
  assign n5470 = ~pi0238 & pi0354;
  assign n5471 = pi0238 & ~pi0354;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = n5222 & ~n5472;
  assign n5474 = pi0238 & ~n5217;
  assign n5475 = ~pi0238 & n5217;
  assign n5476 = ~n5474 & ~n5475;
  assign n5477 = ~n5222 & ~n5476;
  assign n5478 = ~n5473 & ~n5477;
  assign po0289 = pi1169 & ~n5478;
  assign n5480 = ~pi0239 & pi0354;
  assign n5481 = pi0215 & pi0238;
  assign n5482 = n5480 & n5481;
  assign n5483 = pi0239 & ~pi0354;
  assign n5484 = ~n5482 & ~n5483;
  assign n5485 = pi0239 & ~n5481;
  assign n5486 = n5484 & ~n5485;
  assign n5487 = n5222 & ~n5486;
  assign n5488 = pi0239 & ~n5217;
  assign n5489 = ~pi0239 & n5481;
  assign n5490 = ~n5485 & ~n5489;
  assign n5491 = n5217 & ~n5490;
  assign n5492 = ~n5488 & ~n5491;
  assign n5493 = ~n5222 & ~n5492;
  assign n5494 = ~n5487 & ~n5493;
  assign po0290 = pi1169 & ~n5494;
  assign n5496 = pi1761 & n5341;
  assign n5497 = pi1775 & n5277;
  assign n5498 = pi1795 & n5276;
  assign n5499 = ~pi0218 & ~pi0227;
  assign n5500 = pi1709 & n5499;
  assign n5501 = ~n5498 & ~n5500;
  assign n5502 = ~n5497 & n5501;
  assign n5503 = ~n5496 & n5502;
  assign n5504 = pi1178 & ~pi1777;
  assign n5505 = ~n5503 & n5504;
  assign n5506 = pi1510 & n5341;
  assign n5507 = pi1486 & n5277;
  assign n5508 = pi1758 & n5499;
  assign n5509 = pi1461 & n5276;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = ~n5507 & n5510;
  assign n5512 = ~n5506 & n5511;
  assign n5513 = ~pi1178 & pi1777;
  assign n5514 = ~n5512 & n5513;
  assign n5515 = ~n5505 & ~n5514;
  assign n5516 = n5272 & ~n5515;
  assign n5517 = ~pi0240 & ~n5272;
  assign n5518 = ~n5516 & ~n5517;
  assign po0291 = pi1176 & ~n5518;
  assign n5520 = pi1529 & n5341;
  assign n5521 = pi1481 & n5276;
  assign n5522 = pi1505 & n5277;
  assign n5523 = pi1711 & n5499;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~n5521 & n5524;
  assign n5526 = ~n5520 & n5525;
  assign n5527 = n5504 & ~n5526;
  assign n5528 = pi1518 & n5341;
  assign n5529 = pi1470 & n5276;
  assign n5530 = pi1494 & n5277;
  assign n5531 = ~pi0218 & pi1704;
  assign n5532 = ~pi0227 & n5531;
  assign n5533 = ~n5530 & ~n5532;
  assign n5534 = ~n5529 & n5533;
  assign n5535 = ~n5528 & n5534;
  assign n5536 = n5513 & ~n5535;
  assign n5537 = ~n5527 & ~n5536;
  assign n5538 = n5272 & ~n5537;
  assign n5539 = ~pi0241 & ~n5272;
  assign n5540 = ~n5538 & ~n5539;
  assign po0292 = pi1176 & ~n5540;
  assign n5542 = pi1601 & n5357;
  assign n5543 = pi1576 & n5296;
  assign n5544 = pi1552 & n5295;
  assign n5545 = ~pi0219 & pi1724;
  assign n5546 = ~pi0226 & n5545;
  assign n5547 = ~n5544 & ~n5546;
  assign n5548 = ~n5543 & n5547;
  assign n5549 = ~n5542 & n5548;
  assign n5550 = ~pi1845 & pi1846;
  assign n5551 = ~n5549 & n5550;
  assign n5552 = pi1584 & n5357;
  assign n5553 = pi1560 & n5296;
  assign n5554 = pi1535 & n5295;
  assign n5555 = ~pi0219 & ~pi0226;
  assign n5556 = pi1102 & n5555;
  assign n5557 = ~n5554 & ~n5556;
  assign n5558 = ~n5553 & n5557;
  assign n5559 = ~n5552 & n5558;
  assign n5560 = pi1845 & ~pi1846;
  assign n5561 = ~n5559 & n5560;
  assign n5562 = ~n5551 & ~n5561;
  assign n5563 = n5291 & ~n5562;
  assign n5564 = ~pi0242 & ~n5291;
  assign n5565 = ~n5563 & ~n5564;
  assign po0293 = pi1839 & ~n5565;
  assign n5567 = pi1592 & n5357;
  assign n5568 = pi1568 & n5296;
  assign n5569 = pi1544 & n5295;
  assign n5570 = pi1718 & n5555;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = ~n5568 & n5571;
  assign n5573 = ~n5567 & n5572;
  assign n5574 = n5560 & ~n5573;
  assign n5575 = pi1066 & n5357;
  assign n5576 = pi1112 & n5296;
  assign n5577 = pi1127 & n5295;
  assign n5578 = pi1726 & n5555;
  assign n5579 = ~n5577 & ~n5578;
  assign n5580 = ~n5576 & n5579;
  assign n5581 = ~n5575 & n5580;
  assign n5582 = n5550 & ~n5581;
  assign n5583 = ~n5574 & ~n5582;
  assign n5584 = n5291 & ~n5583;
  assign n5585 = ~pi0243 & ~n5291;
  assign n5586 = ~n5584 & ~n5585;
  assign po0294 = pi1839 & ~n5586;
  assign n5588 = pi1303 & n5325;
  assign n5589 = pi1048 & n5258;
  assign n5590 = pi1114 & n5257;
  assign n5591 = ~pi0217 & ~pi0225;
  assign n5592 = pi1008 & n5591;
  assign n5593 = ~n5590 & ~n5592;
  assign n5594 = ~n5589 & n5593;
  assign n5595 = ~n5588 & n5594;
  assign n5596 = ~pi1130 & pi1183;
  assign n5597 = ~n5595 & n5596;
  assign n5598 = pi1287 & n5325;
  assign n5599 = pi1253 & n5258;
  assign n5600 = pi1623 & n5257;
  assign n5601 = pi1833 & n5591;
  assign n5602 = ~n5600 & ~n5601;
  assign n5603 = ~n5599 & n5602;
  assign n5604 = ~n5598 & n5603;
  assign n5605 = pi1130 & ~pi1183;
  assign n5606 = ~n5604 & n5605;
  assign n5607 = ~n5597 & ~n5606;
  assign n5608 = n5253 & ~n5607;
  assign n5609 = ~pi0244 & ~n5253;
  assign n5610 = ~n5608 & ~n5609;
  assign po0295 = pi1164 & ~n5610;
  assign n5612 = pi1064 & n5325;
  assign n5613 = pi1281 & n5258;
  assign n5614 = pi1109 & n5257;
  assign n5615 = pi1753 & n5591;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = ~n5613 & n5616;
  assign n5618 = ~n5612 & n5617;
  assign n5619 = n5596 & ~n5618;
  assign n5620 = pi1295 & n5325;
  assign n5621 = pi1271 & n5258;
  assign n5622 = pi1649 & n5257;
  assign n5623 = ~pi0217 & pi0999;
  assign n5624 = ~pi0225 & n5623;
  assign n5625 = ~n5622 & ~n5624;
  assign n5626 = ~n5621 & n5625;
  assign n5627 = ~n5620 & n5626;
  assign n5628 = n5605 & ~n5627;
  assign n5629 = ~n5619 & ~n5628;
  assign n5630 = n5253 & ~n5629;
  assign n5631 = ~pi0245 & ~n5253;
  assign n5632 = ~n5630 & ~n5631;
  assign po0296 = pi1164 & ~n5632;
  assign n5634 = pi1257 & n5309;
  assign n5635 = ~pi0216 & ~pi0224;
  assign n5636 = pi1804 & n5635;
  assign n5637 = pi1627 & n5238;
  assign n5638 = pi1664 & n5239;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = ~n5636 & n5639;
  assign n5641 = ~n5634 & n5640;
  assign n5642 = pi1832 & ~pi1840;
  assign n5643 = ~n5641 & n5642;
  assign n5644 = pi1231 & n5309;
  assign n5645 = pi1638 & n5239;
  assign n5646 = pi0995 & n5635;
  assign n5647 = pi1609 & n5238;
  assign n5648 = ~n5646 & ~n5647;
  assign n5649 = ~n5645 & n5648;
  assign n5650 = ~n5644 & n5649;
  assign n5651 = ~pi1832 & pi1840;
  assign n5652 = ~n5650 & n5651;
  assign n5653 = ~n5643 & ~n5652;
  assign n5654 = n5234 & ~n5653;
  assign n5655 = ~pi0246 & ~n5234;
  assign n5656 = ~n5654 & ~n5655;
  assign po0297 = pi1838 & ~n5656;
  assign n5658 = pi1098 & n5309;
  assign n5659 = pi1798 & n5635;
  assign n5660 = pi1828 & n5239;
  assign n5661 = pi1051 & n5238;
  assign n5662 = ~n5660 & ~n5661;
  assign n5663 = ~n5659 & n5662;
  assign n5664 = ~n5658 & n5663;
  assign n5665 = n5642 & ~n5664;
  assign n5666 = pi1244 & n5309;
  assign n5667 = pi1831 & n5635;
  assign n5668 = pi1652 & n5239;
  assign n5669 = pi1617 & n5238;
  assign n5670 = ~n5668 & ~n5669;
  assign n5671 = ~n5667 & n5670;
  assign n5672 = ~n5666 & n5671;
  assign n5673 = n5651 & ~n5672;
  assign n5674 = ~n5665 & ~n5673;
  assign n5675 = n5234 & ~n5674;
  assign n5676 = ~pi0247 & ~n5234;
  assign n5677 = ~n5675 & ~n5676;
  assign po0298 = pi1838 & ~n5677;
  assign n5679 = ~pi0248 & ~pi0861;
  assign po0299 = ~n5425 & ~n5679;
  assign n5681 = ~pi0249 & ~pi0862;
  assign po0300 = ~n5425 & ~n5681;
  assign n5683 = ~pi0250 & ~pi0863;
  assign po0301 = ~n5425 & ~n5683;
  assign n5685 = ~pi0251 & ~pi0864;
  assign po0302 = ~n5425 & ~n5685;
  assign n5687 = n5272 & n5504;
  assign n5688 = pi1176 & n5687;
  assign n5689 = ~n5512 & n5688;
  assign n5690 = pi1176 & ~n5272;
  assign n5691 = ~pi0252 & n5690;
  assign po0303 = n5689 | n5691;
  assign n5693 = ~n5535 & n5688;
  assign n5694 = ~pi0253 & n5690;
  assign po0304 = n5693 | n5694;
  assign n5696 = n5291 & n5550;
  assign n5697 = pi1839 & n5696;
  assign n5698 = ~n5559 & n5697;
  assign n5699 = pi1839 & ~n5291;
  assign n5700 = ~pi0254 & n5699;
  assign po0305 = n5698 | n5700;
  assign n5702 = ~n5573 & n5697;
  assign n5703 = ~pi0255 & n5699;
  assign po0306 = n5702 | n5703;
  assign n5705 = n5253 & n5596;
  assign n5706 = pi1164 & n5705;
  assign n5707 = ~n5604 & n5706;
  assign n5708 = pi1164 & ~n5253;
  assign n5709 = ~pi0256 & n5708;
  assign po0307 = n5707 | n5709;
  assign n5711 = n5234 & n5642;
  assign n5712 = pi1838 & n5711;
  assign n5713 = ~n5650 & n5712;
  assign n5714 = pi1838 & ~n5234;
  assign n5715 = ~pi0257 & n5714;
  assign po0308 = n5713 | n5715;
  assign n5717 = ~n5627 & n5706;
  assign n5718 = ~pi0258 & n5708;
  assign po0309 = n5717 | n5718;
  assign n5720 = ~n5672 & n5712;
  assign n5721 = ~pi0259 & n5714;
  assign po0310 = n5720 | n5721;
  assign n5723 = pi0260 & n5236;
  assign n5724 = ~pi0260 & ~n5236;
  assign n5725 = ~n5723 & ~n5724;
  assign po0311 = pi1838 & n5725;
  assign n5727 = pi0261 & n5255;
  assign n5728 = ~pi0261 & ~n5255;
  assign n5729 = ~n5727 & ~n5728;
  assign po0312 = pi1164 & n5729;
  assign n5731 = pi0262 & n5274;
  assign n5732 = ~pi0262 & ~n5274;
  assign n5733 = ~n5731 & ~n5732;
  assign po0313 = pi1176 & n5733;
  assign n5735 = pi0263 & n5293;
  assign n5736 = ~pi0263 & ~n5293;
  assign n5737 = ~n5735 & ~n5736;
  assign po0314 = pi1839 & n5737;
  assign n5739 = pi1124 & n5341;
  assign n5740 = pi1774 & n5277;
  assign n5741 = pi1713 & n5499;
  assign n5742 = pi1794 & n5276;
  assign n5743 = ~n5741 & ~n5742;
  assign n5744 = ~n5740 & n5743;
  assign n5745 = ~n5739 & n5744;
  assign n5746 = ~pi0262 & ~n5745;
  assign n5747 = pi1474 & n5276;
  assign n5748 = pi0977 & n5499;
  assign n5749 = ~n5747 & ~n5748;
  assign n5750 = pi1522 & n5341;
  assign n5751 = pi1498 & n5277;
  assign n5752 = ~n5750 & ~n5751;
  assign n5753 = n5749 & n5752;
  assign n5754 = pi0262 & ~n5753;
  assign n5755 = ~n5746 & ~n5754;
  assign n5756 = n5273 & ~n5755;
  assign n5757 = pi1512 & n5341;
  assign n5758 = pi1463 & n5276;
  assign n5759 = pi1081 & n5499;
  assign n5760 = pi1488 & n5277;
  assign n5761 = ~n5759 & ~n5760;
  assign n5762 = ~n5758 & n5761;
  assign n5763 = ~n5757 & n5762;
  assign n5764 = n5504 & ~n5763;
  assign n5765 = pi1462 & n5276;
  assign n5766 = pi1511 & n5341;
  assign n5767 = pi1699 & n5499;
  assign n5768 = pi1487 & n5277;
  assign n5769 = ~n5767 & ~n5768;
  assign n5770 = ~n5766 & n5769;
  assign n5771 = ~n5765 & n5770;
  assign n5772 = n5513 & ~n5771;
  assign n5773 = ~n5764 & ~n5772;
  assign n5774 = ~n5756 & n5773;
  assign n5775 = n5272 & ~n5774;
  assign n5776 = ~pi0264 & ~n5272;
  assign n5777 = ~n5775 & ~n5776;
  assign po0315 = pi1176 & ~n5777;
  assign n5779 = pi1533 & n5341;
  assign n5780 = pi1485 & n5276;
  assign n5781 = pi1509 & n5277;
  assign n5782 = pi0981 & n5499;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = ~n5780 & n5783;
  assign n5785 = ~n5779 & n5784;
  assign n5786 = ~pi0262 & ~n5785;
  assign n5787 = pi1475 & n5276;
  assign n5788 = pi1708 & n5499;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = pi1523 & n5341;
  assign n5791 = pi1499 & n5277;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = n5789 & n5792;
  assign n5794 = pi0262 & ~n5793;
  assign n5795 = ~n5786 & ~n5794;
  assign n5796 = n5273 & ~n5795;
  assign n5797 = pi1513 & n5341;
  assign n5798 = pi1489 & n5277;
  assign n5799 = pi0972 & n5499;
  assign n5800 = pi1464 & n5276;
  assign n5801 = ~n5799 & ~n5800;
  assign n5802 = ~n5798 & n5801;
  assign n5803 = ~n5797 & n5802;
  assign n5804 = n5504 & ~n5803;
  assign n5805 = pi1773 & n5341;
  assign n5806 = pi1787 & n5277;
  assign n5807 = pi1700 & n5499;
  assign n5808 = pi1802 & n5276;
  assign n5809 = ~n5807 & ~n5808;
  assign n5810 = ~n5806 & n5809;
  assign n5811 = ~n5805 & n5810;
  assign n5812 = n5513 & ~n5811;
  assign n5813 = ~n5804 & ~n5812;
  assign n5814 = ~n5796 & n5813;
  assign n5815 = n5272 & ~n5814;
  assign n5816 = ~pi0265 & ~n5272;
  assign n5817 = ~n5815 & ~n5816;
  assign po0316 = pi1176 & ~n5817;
  assign n5819 = ~pi0262 & ~n5771;
  assign n5820 = pi1791 & n5276;
  assign n5821 = pi1706 & n5499;
  assign n5822 = ~n5820 & ~n5821;
  assign n5823 = pi1763 & n5341;
  assign n5824 = pi1780 & n5277;
  assign n5825 = ~n5823 & ~n5824;
  assign n5826 = n5822 & n5825;
  assign n5827 = pi0262 & ~n5826;
  assign n5828 = ~n5819 & ~n5827;
  assign n5829 = n5273 & ~n5828;
  assign n5830 = pi1465 & n5276;
  assign n5831 = pi1490 & n5277;
  assign n5832 = pi1514 & n5341;
  assign n5833 = ~n5831 & ~n5832;
  assign n5834 = pi0973 & n5499;
  assign n5835 = n5833 & ~n5834;
  assign n5836 = ~n5830 & n5835;
  assign n5837 = n5504 & ~n5836;
  assign n5838 = n5513 & ~n5763;
  assign n5839 = ~n5837 & ~n5838;
  assign n5840 = ~n5829 & n5839;
  assign n5841 = n5272 & ~n5840;
  assign n5842 = ~pi0266 & ~n5272;
  assign n5843 = ~n5841 & ~n5842;
  assign po0317 = pi1176 & ~n5843;
  assign n5845 = ~pi0262 & ~n5811;
  assign n5846 = pi1524 & n5341;
  assign n5847 = pi1500 & n5277;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = pi1476 & n5276;
  assign n5850 = pi1707 & n5499;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = n5848 & n5851;
  assign n5853 = pi0262 & ~n5852;
  assign n5854 = ~n5845 & ~n5853;
  assign n5855 = n5273 & ~n5854;
  assign n5856 = pi1765 & n5341;
  assign n5857 = pi1784 & n5277;
  assign n5858 = pi1701 & n5499;
  assign n5859 = pi1785 & n5276;
  assign n5860 = ~n5858 & ~n5859;
  assign n5861 = ~n5857 & n5860;
  assign n5862 = ~n5856 & n5861;
  assign n5863 = n5504 & ~n5862;
  assign n5864 = n5513 & ~n5803;
  assign n5865 = ~n5863 & ~n5864;
  assign n5866 = ~n5855 & n5865;
  assign n5867 = n5272 & ~n5866;
  assign n5868 = ~pi0267 & ~n5272;
  assign n5869 = ~n5867 & ~n5868;
  assign po0318 = pi1176 & ~n5869;
  assign n5871 = pi1531 & n5341;
  assign n5872 = pi1507 & n5277;
  assign n5873 = pi1118 & n5499;
  assign n5874 = pi1483 & n5276;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n5872 & n5875;
  assign n5877 = ~n5871 & n5876;
  assign n5878 = ~pi0262 & ~n5877;
  assign n5879 = pi1797 & n5276;
  assign n5880 = pi0976 & n5499;
  assign n5881 = ~n5879 & ~n5880;
  assign n5882 = pi1764 & n5341;
  assign n5883 = pi1757 & n5277;
  assign n5884 = ~n5882 & ~n5883;
  assign n5885 = n5881 & n5884;
  assign n5886 = pi0262 & ~n5885;
  assign n5887 = ~n5878 & ~n5886;
  assign n5888 = n5273 & ~n5887;
  assign n5889 = n5504 & ~n5771;
  assign n5890 = n5513 & ~n5745;
  assign n5891 = ~n5889 & ~n5890;
  assign n5892 = ~n5888 & n5891;
  assign n5893 = n5272 & ~n5892;
  assign n5894 = ~pi0268 & ~n5272;
  assign n5895 = ~n5893 & ~n5894;
  assign po0319 = pi1176 & ~n5895;
  assign n5897 = pi1532 & n5341;
  assign n5898 = pi1508 & n5277;
  assign n5899 = pi0980 & n5499;
  assign n5900 = pi1484 & n5276;
  assign n5901 = ~n5899 & ~n5900;
  assign n5902 = ~n5898 & n5901;
  assign n5903 = ~n5897 & n5902;
  assign n5904 = ~pi0262 & ~n5903;
  assign n5905 = pi1473 & n5276;
  assign n5906 = pi1136 & n5499;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = pi1521 & n5341;
  assign n5909 = pi1497 & n5277;
  assign n5910 = ~n5908 & ~n5909;
  assign n5911 = n5907 & n5910;
  assign n5912 = pi0262 & ~n5911;
  assign n5913 = ~n5904 & ~n5912;
  assign n5914 = n5273 & ~n5913;
  assign n5915 = n5504 & ~n5811;
  assign n5916 = n5513 & ~n5785;
  assign n5917 = ~n5915 & ~n5916;
  assign n5918 = ~n5914 & n5917;
  assign n5919 = n5272 & ~n5918;
  assign n5920 = ~pi0269 & ~n5272;
  assign n5921 = ~n5919 & ~n5920;
  assign po0320 = pi1176 & ~n5921;
  assign n5923 = ~pi0270 & ~n5272;
  assign n5924 = ~pi0262 & ~n5836;
  assign n5925 = pi1527 & n5341;
  assign n5926 = pi1503 & n5277;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = pi1479 & n5276;
  assign n5929 = pi1117 & n5499;
  assign n5930 = ~n5928 & ~n5929;
  assign n5931 = n5927 & n5930;
  assign n5932 = pi0262 & ~n5931;
  assign n5933 = ~n5924 & ~n5932;
  assign n5934 = n5273 & ~n5933;
  assign n5935 = pi1517 & n5341;
  assign n5936 = pi1493 & n5277;
  assign n5937 = pi1468 & n5276;
  assign n5938 = pi1703 & n5499;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = ~n5936 & n5939;
  assign n5941 = ~n5935 & n5940;
  assign n5942 = n5504 & ~n5941;
  assign n5943 = pi0974 & n5499;
  assign n5944 = pi1466 & n5276;
  assign n5945 = pi1491 & n5277;
  assign n5946 = pi1515 & n5341;
  assign n5947 = ~n5945 & ~n5946;
  assign n5948 = ~n5944 & n5947;
  assign n5949 = ~n5943 & n5948;
  assign n5950 = n5513 & ~n5949;
  assign n5951 = ~n5942 & ~n5950;
  assign n5952 = ~n5934 & n5951;
  assign n5953 = n5272 & ~n5952;
  assign n5954 = ~n5923 & ~n5953;
  assign po0321 = pi1176 & ~n5954;
  assign n5956 = ~pi0262 & ~n5862;
  assign n5957 = pi1528 & n5341;
  assign n5958 = pi1504 & n5277;
  assign n5959 = ~n5957 & ~n5958;
  assign n5960 = pi1480 & n5276;
  assign n5961 = pi0978 & n5499;
  assign n5962 = ~n5960 & ~n5961;
  assign n5963 = n5959 & n5962;
  assign n5964 = pi0262 & ~n5963;
  assign n5965 = ~n5956 & ~n5964;
  assign n5966 = n5273 & ~n5965;
  assign n5967 = pi1767 & n5341;
  assign n5968 = pi1469 & n5276;
  assign n5969 = pi0975 & n5499;
  assign n5970 = pi1786 & n5277;
  assign n5971 = ~n5969 & ~n5970;
  assign n5972 = ~n5968 & n5971;
  assign n5973 = ~n5967 & n5972;
  assign n5974 = n5504 & ~n5973;
  assign n5975 = pi1516 & n5341;
  assign n5976 = pi1467 & n5276;
  assign n5977 = pi1492 & n5277;
  assign n5978 = pi1447 & n5499;
  assign n5979 = ~n5977 & ~n5978;
  assign n5980 = ~n5976 & n5979;
  assign n5981 = ~n5975 & n5980;
  assign n5982 = n5513 & ~n5981;
  assign n5983 = ~n5974 & ~n5982;
  assign n5984 = ~n5966 & n5983;
  assign n5985 = n5272 & ~n5984;
  assign n5986 = ~pi0271 & ~n5272;
  assign n5987 = ~n5985 & ~n5986;
  assign po0322 = pi1176 & ~n5987;
  assign n5989 = ~pi0262 & ~n5763;
  assign n5990 = pi1477 & n5276;
  assign n5991 = pi1122 & n5499;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = pi1525 & n5341;
  assign n5994 = pi1501 & n5277;
  assign n5995 = ~n5993 & ~n5994;
  assign n5996 = n5992 & n5995;
  assign n5997 = pi0262 & ~n5996;
  assign n5998 = ~n5989 & ~n5997;
  assign n5999 = n5273 & ~n5998;
  assign n6000 = n5504 & ~n5949;
  assign n6001 = n5513 & ~n5836;
  assign n6002 = ~n6000 & ~n6001;
  assign n6003 = ~n5999 & n6002;
  assign n6004 = n5272 & ~n6003;
  assign n6005 = ~pi0272 & ~n5272;
  assign n6006 = ~n6004 & ~n6005;
  assign po0323 = pi1176 & ~n6006;
  assign n6008 = ~pi0262 & ~n5803;
  assign n6009 = pi1526 & n5341;
  assign n6010 = pi1502 & n5277;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = pi1478 & n5276;
  assign n6013 = pi1710 & n5499;
  assign n6014 = ~n6012 & ~n6013;
  assign n6015 = n6011 & n6014;
  assign n6016 = pi0262 & ~n6015;
  assign n6017 = ~n6008 & ~n6016;
  assign n6018 = n5273 & ~n6017;
  assign n6019 = n5504 & ~n5981;
  assign n6020 = n5513 & ~n5862;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = ~n6018 & n6021;
  assign n6023 = n5272 & ~n6022;
  assign n6024 = ~pi0273 & ~n5272;
  assign n6025 = ~n6023 & ~n6024;
  assign po0324 = pi1176 & ~n6025;
  assign n6027 = ~pi0262 & ~n5512;
  assign n6028 = pi0262 & ~n5949;
  assign n6029 = ~n6027 & ~n6028;
  assign n6030 = n5273 & ~n6029;
  assign n6031 = pi1759 & n5341;
  assign n6032 = pi1772 & n5277;
  assign n6033 = pi0979 & n5499;
  assign n6034 = pi1793 & n5276;
  assign n6035 = ~n6033 & ~n6034;
  assign n6036 = ~n6032 & n6035;
  assign n6037 = ~n6031 & n6036;
  assign n6038 = n5504 & ~n6037;
  assign n6039 = ~n5503 & n5513;
  assign n6040 = ~n6038 & ~n6039;
  assign n6041 = ~n6030 & n6040;
  assign n6042 = n5272 & ~n6041;
  assign n6043 = ~pi0274 & ~n5272;
  assign n6044 = ~n6042 & ~n6043;
  assign po0325 = pi1176 & ~n6044;
  assign n6046 = pi0262 & ~n5981;
  assign n6047 = ~pi0262 & ~n5535;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = n5273 & ~n6048;
  assign n6050 = pi1530 & n5341;
  assign n6051 = pi1506 & n5277;
  assign n6052 = pi1712 & n5499;
  assign n6053 = pi1482 & n5276;
  assign n6054 = ~n6052 & ~n6053;
  assign n6055 = ~n6051 & n6054;
  assign n6056 = ~n6050 & n6055;
  assign n6057 = n5504 & ~n6056;
  assign n6058 = n5513 & ~n5526;
  assign n6059 = ~n6057 & ~n6058;
  assign n6060 = ~n6049 & n6059;
  assign n6061 = n5272 & ~n6060;
  assign n6062 = ~pi0275 & ~n5272;
  assign n6063 = ~n6061 & ~n6062;
  assign po0326 = pi1176 & ~n6063;
  assign n6065 = pi0262 & ~n5941;
  assign n6066 = ~pi0262 & ~n5503;
  assign n6067 = ~n6065 & ~n6066;
  assign n6068 = n5273 & ~n6067;
  assign n6069 = n5504 & ~n5877;
  assign n6070 = n5513 & ~n6037;
  assign n6071 = ~n6069 & ~n6070;
  assign n6072 = ~n6068 & n6071;
  assign n6073 = n5272 & ~n6072;
  assign n6074 = ~pi0276 & ~n5272;
  assign n6075 = ~n6073 & ~n6074;
  assign po0327 = pi1176 & ~n6075;
  assign n6077 = pi0262 & ~n5973;
  assign n6078 = ~pi0262 & ~n5526;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = n5273 & ~n6079;
  assign n6081 = n5504 & ~n5903;
  assign n6082 = n5513 & ~n6056;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = ~n6080 & n6083;
  assign n6085 = n5272 & ~n6084;
  assign n6086 = ~pi0277 & ~n5272;
  assign n6087 = ~n6085 & ~n6086;
  assign po0328 = pi1176 & ~n6087;
  assign n6089 = ~pi0262 & ~n6037;
  assign n6090 = pi1519 & n5341;
  assign n6091 = pi1495 & n5277;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = pi1471 & n5276;
  assign n6094 = pi1594 & n5499;
  assign n6095 = ~n6093 & ~n6094;
  assign n6096 = n6092 & n6095;
  assign n6097 = pi0262 & ~n6096;
  assign n6098 = ~n6089 & ~n6097;
  assign n6099 = n5273 & ~n6098;
  assign n6100 = n5504 & ~n5745;
  assign n6101 = n5513 & ~n5877;
  assign n6102 = ~n6100 & ~n6101;
  assign n6103 = ~n6099 & n6102;
  assign n6104 = n5272 & ~n6103;
  assign n6105 = ~pi0278 & ~n5272;
  assign n6106 = ~n6104 & ~n6105;
  assign po0329 = pi1176 & ~n6106;
  assign n6108 = ~pi0262 & ~n6056;
  assign n6109 = pi1472 & n5276;
  assign n6110 = pi1705 & n5499;
  assign n6111 = ~n6109 & ~n6110;
  assign n6112 = pi1520 & n5341;
  assign n6113 = pi1496 & n5277;
  assign n6114 = ~n6112 & ~n6113;
  assign n6115 = n6111 & n6114;
  assign n6116 = pi0262 & ~n6115;
  assign n6117 = ~n6108 & ~n6116;
  assign n6118 = n5273 & ~n6117;
  assign n6119 = n5504 & ~n5785;
  assign n6120 = n5513 & ~n5903;
  assign n6121 = ~n6119 & ~n6120;
  assign n6122 = ~n6118 & n6121;
  assign n6123 = n5272 & ~n6122;
  assign n6124 = ~pi0279 & ~n5272;
  assign n6125 = ~n6123 & ~n6124;
  assign po0330 = pi1176 & ~n6125;
  assign n6127 = ~pi0280 & ~n5291;
  assign n6128 = pi1595 & n5357;
  assign n6129 = pi0986 & n5555;
  assign n6130 = pi1570 & n5296;
  assign n6131 = pi1546 & n5295;
  assign n6132 = ~n6130 & ~n6131;
  assign n6133 = ~n6129 & n6132;
  assign n6134 = ~n6128 & n6133;
  assign n6135 = n5292 & ~n6134;
  assign n6136 = pi0263 & n6135;
  assign n6137 = pi1606 & n5357;
  assign n6138 = pi1557 & n5295;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = pi1581 & n5296;
  assign n6141 = pi1062 & n5555;
  assign n6142 = ~n6140 & ~n6141;
  assign n6143 = n6139 & n6142;
  assign n6144 = ~pi0263 & n5292;
  assign n6145 = ~n6143 & n6144;
  assign n6146 = ~n6136 & ~n6145;
  assign n6147 = pi1107 & n5357;
  assign n6148 = pi1120 & n5296;
  assign n6149 = pi1755 & n5295;
  assign n6150 = pi1714 & n5555;
  assign n6151 = ~n6149 & ~n6150;
  assign n6152 = ~n6148 & n6151;
  assign n6153 = ~n6147 & n6152;
  assign n6154 = n5550 & ~n6153;
  assign n6155 = pi1607 & n5357;
  assign n6156 = pi1582 & n5296;
  assign n6157 = pi1558 & n5295;
  assign n6158 = pi1728 & n5555;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = ~n6156 & n6159;
  assign n6161 = ~n6155 & n6160;
  assign n6162 = n5560 & ~n6161;
  assign n6163 = ~n6154 & ~n6162;
  assign n6164 = n6146 & n6163;
  assign n6165 = n5291 & ~n6164;
  assign n6166 = ~n6127 & ~n6165;
  assign po0331 = pi1839 & ~n6166;
  assign n6168 = ~pi0281 & ~n5291;
  assign n6169 = pi1596 & n5357;
  assign n6170 = pi1073 & n5555;
  assign n6171 = pi1571 & n5296;
  assign n6172 = pi1547 & n5295;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = ~n6170 & n6173;
  assign n6175 = ~n6169 & n6174;
  assign n6176 = n5292 & ~n6175;
  assign n6177 = pi0263 & n6176;
  assign n6178 = pi1083 & n5357;
  assign n6179 = pi0990 & n5555;
  assign n6180 = pi1106 & n5296;
  assign n6181 = pi1123 & n5295;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = ~n6179 & n6182;
  assign n6184 = ~n6178 & n6183;
  assign n6185 = n6144 & ~n6184;
  assign n6186 = ~n6177 & ~n6185;
  assign n6187 = pi1585 & n5357;
  assign n6188 = pi1715 & n5555;
  assign n6189 = pi1536 & n5295;
  assign n6190 = pi1561 & n5296;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = ~n6188 & n6191;
  assign n6193 = ~n6187 & n6192;
  assign n6194 = n5550 & ~n6193;
  assign n6195 = pi1608 & n5357;
  assign n6196 = pi0991 & n5555;
  assign n6197 = pi1583 & n5296;
  assign n6198 = pi1559 & n5295;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = ~n6196 & n6199;
  assign n6201 = ~n6195 & n6200;
  assign n6202 = n5560 & ~n6201;
  assign n6203 = ~n6194 & ~n6202;
  assign n6204 = n6186 & n6203;
  assign n6205 = n5291 & ~n6204;
  assign n6206 = ~n6168 & ~n6205;
  assign po0332 = pi1839 & ~n6206;
  assign n6208 = ~pi0282 & ~n5291;
  assign n6209 = ~pi0263 & ~n6161;
  assign n6210 = pi1597 & n5357;
  assign n6211 = pi1572 & n5296;
  assign n6212 = ~n6210 & ~n6211;
  assign n6213 = pi1548 & n5295;
  assign n6214 = pi0987 & n5555;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = n6212 & n6215;
  assign n6217 = pi0263 & ~n6216;
  assign n6218 = ~n6209 & ~n6217;
  assign n6219 = n5292 & ~n6218;
  assign n6220 = pi1586 & n5357;
  assign n6221 = pi1562 & n5296;
  assign n6222 = pi1537 & n5295;
  assign n6223 = pi1087 & n5555;
  assign n6224 = ~n6222 & ~n6223;
  assign n6225 = ~n6221 & n6224;
  assign n6226 = ~n6220 & n6225;
  assign n6227 = n5550 & ~n6226;
  assign n6228 = n5560 & ~n6153;
  assign n6229 = ~n6227 & ~n6228;
  assign n6230 = ~n6219 & n6229;
  assign n6231 = n5291 & ~n6230;
  assign n6232 = ~n6208 & ~n6231;
  assign po0333 = pi1839 & ~n6232;
  assign n6234 = ~pi0283 & ~n5291;
  assign n6235 = ~pi0263 & ~n6201;
  assign n6236 = pi1089 & n5357;
  assign n6237 = pi1105 & n5296;
  assign n6238 = ~n6236 & ~n6237;
  assign n6239 = pi1063 & n5295;
  assign n6240 = pi1720 & n5555;
  assign n6241 = ~n6239 & ~n6240;
  assign n6242 = n6238 & n6241;
  assign n6243 = pi0263 & ~n6242;
  assign n6244 = ~n6235 & ~n6243;
  assign n6245 = n5292 & ~n6244;
  assign n6246 = pi1587 & n5357;
  assign n6247 = pi1563 & n5296;
  assign n6248 = pi1538 & n5295;
  assign n6249 = pi0982 & n5555;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n6247 & n6250;
  assign n6252 = ~n6246 & n6251;
  assign n6253 = n5550 & ~n6252;
  assign n6254 = n5560 & ~n6193;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6245 & n6255;
  assign n6257 = n5291 & ~n6256;
  assign n6258 = ~n6234 & ~n6257;
  assign po0334 = pi1839 & ~n6258;
  assign n6260 = ~pi0284 & ~n5291;
  assign n6261 = ~pi0263 & ~n6153;
  assign n6262 = pi1598 & n5357;
  assign n6263 = pi1573 & n5296;
  assign n6264 = ~n6262 & ~n6263;
  assign n6265 = pi1549 & n5295;
  assign n6266 = pi1723 & n5555;
  assign n6267 = ~n6265 & ~n6266;
  assign n6268 = n6264 & n6267;
  assign n6269 = pi0263 & ~n6268;
  assign n6270 = ~n6261 & ~n6269;
  assign n6271 = n5292 & ~n6270;
  assign n6272 = pi1088 & n5357;
  assign n6273 = pi1119 & n5296;
  assign n6274 = pi1391 & n5295;
  assign n6275 = pi0983 & n5555;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = ~n6273 & n6276;
  assign n6278 = ~n6272 & n6277;
  assign n6279 = n5550 & ~n6278;
  assign n6280 = n5560 & ~n6226;
  assign n6281 = ~n6279 & ~n6280;
  assign n6282 = ~n6271 & n6281;
  assign n6283 = n5291 & ~n6282;
  assign n6284 = ~n6260 & ~n6283;
  assign po0335 = pi1839 & ~n6284;
  assign n6286 = ~pi0285 & ~n5291;
  assign n6287 = ~pi0263 & ~n6252;
  assign n6288 = pi1090 & n5357;
  assign n6289 = pi1113 & n5296;
  assign n6290 = ~n6288 & ~n6289;
  assign n6291 = pi1135 & n5295;
  assign n6292 = pi1725 & n5555;
  assign n6293 = ~n6291 & ~n6292;
  assign n6294 = n6290 & n6293;
  assign n6295 = pi0263 & ~n6294;
  assign n6296 = ~n6287 & ~n6295;
  assign n6297 = n5292 & ~n6296;
  assign n6298 = pi1590 & n5357;
  assign n6299 = pi1566 & n5296;
  assign n6300 = pi1541 & n5295;
  assign n6301 = pi1101 & n5555;
  assign n6302 = ~n6300 & ~n6301;
  assign n6303 = ~n6299 & n6302;
  assign n6304 = ~n6298 & n6303;
  assign n6305 = n5550 & ~n6304;
  assign n6306 = pi1588 & n5357;
  assign n6307 = pi1564 & n5296;
  assign n6308 = pi1539 & n5295;
  assign n6309 = pi1716 & n5555;
  assign n6310 = ~n6308 & ~n6309;
  assign n6311 = ~n6307 & n6310;
  assign n6312 = ~n6306 & n6311;
  assign n6313 = n5560 & ~n6312;
  assign n6314 = ~n6305 & ~n6313;
  assign n6315 = ~n6297 & n6314;
  assign n6316 = n5291 & ~n6315;
  assign n6317 = ~n6286 & ~n6316;
  assign po0336 = pi1839 & ~n6317;
  assign n6319 = ~pi0286 & ~n5291;
  assign n6320 = pi0263 & n5292;
  assign n6321 = pi1599 & n5357;
  assign n6322 = pi1574 & n5296;
  assign n6323 = ~n6321 & ~n6322;
  assign n6324 = pi1550 & n5295;
  assign n6325 = pi1721 & n5555;
  assign n6326 = ~n6324 & ~n6325;
  assign n6327 = n6323 & n6326;
  assign n6328 = n6320 & ~n6327;
  assign n6329 = n6144 & ~n6193;
  assign n6330 = ~n6328 & ~n6329;
  assign n6331 = n5550 & ~n6312;
  assign n6332 = n5560 & ~n6252;
  assign n6333 = ~n6331 & ~n6332;
  assign n6334 = n6330 & n6333;
  assign n6335 = n5291 & ~n6334;
  assign n6336 = ~n6319 & ~n6335;
  assign po0337 = pi1839 & ~n6336;
  assign n6338 = ~pi0287 & ~n5291;
  assign n6339 = ~pi0263 & ~n6312;
  assign n6340 = pi1603 & n5357;
  assign n6341 = pi1578 & n5296;
  assign n6342 = ~n6340 & ~n6341;
  assign n6343 = pi1554 & n5295;
  assign n6344 = pi0988 & n5555;
  assign n6345 = ~n6343 & ~n6344;
  assign n6346 = n6342 & n6345;
  assign n6347 = pi0263 & ~n6346;
  assign n6348 = ~n6339 & ~n6347;
  assign n6349 = n5292 & ~n6348;
  assign n6350 = pi1567 & n5296;
  assign n6351 = pi1591 & n5357;
  assign n6352 = pi1543 & n5295;
  assign n6353 = pi0985 & n5555;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = ~n6351 & n6354;
  assign n6356 = ~n6350 & n6355;
  assign n6357 = n5550 & ~n6356;
  assign n6358 = n5560 & ~n6304;
  assign n6359 = ~n6357 & ~n6358;
  assign n6360 = ~n6349 & n6359;
  assign n6361 = n5291 & ~n6360;
  assign n6362 = ~n6338 & ~n6361;
  assign po0338 = pi1839 & ~n6362;
  assign n6364 = ~pi0288 & ~n5291;
  assign n6365 = ~pi0263 & ~n6226;
  assign n6366 = pi1600 & n5357;
  assign n6367 = pi1575 & n5296;
  assign n6368 = ~n6366 & ~n6367;
  assign n6369 = pi1551 & n5295;
  assign n6370 = pi1722 & n5555;
  assign n6371 = ~n6369 & ~n6370;
  assign n6372 = n6368 & n6371;
  assign n6373 = pi0263 & ~n6372;
  assign n6374 = ~n6365 & ~n6373;
  assign n6375 = n5292 & ~n6374;
  assign n6376 = pi1589 & n5357;
  assign n6377 = pi1565 & n5296;
  assign n6378 = pi1540 & n5295;
  assign n6379 = pi0984 & n5555;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~n6377 & n6380;
  assign n6382 = ~n6376 & n6381;
  assign n6383 = n5550 & ~n6382;
  assign n6384 = n5560 & ~n6278;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n6375 & n6385;
  assign n6387 = n5291 & ~n6386;
  assign n6388 = ~n6364 & ~n6387;
  assign po0339 = pi1839 & ~n6388;
  assign n6390 = ~pi0289 & ~n5291;
  assign n6391 = ~pi0263 & ~n6278;
  assign n6392 = pi1602 & n5357;
  assign n6393 = pi1577 & n5296;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = pi1553 & n5295;
  assign n6396 = pi1047 & n5555;
  assign n6397 = ~n6395 & ~n6396;
  assign n6398 = n6394 & n6397;
  assign n6399 = pi0263 & ~n6398;
  assign n6400 = ~n6391 & ~n6399;
  assign n6401 = n5292 & ~n6400;
  assign n6402 = pi1097 & n5357;
  assign n6403 = pi1116 & n5296;
  assign n6404 = pi1542 & n5295;
  assign n6405 = pi1717 & n5555;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 = ~n6403 & n6406;
  assign n6408 = ~n6402 & n6407;
  assign n6409 = n5550 & ~n6408;
  assign n6410 = n5560 & ~n6382;
  assign n6411 = ~n6409 & ~n6410;
  assign n6412 = ~n6401 & n6411;
  assign n6413 = n5291 & ~n6412;
  assign n6414 = ~n6390 & ~n6413;
  assign po0340 = pi1839 & ~n6414;
  assign n6416 = pi0263 & ~n6382;
  assign n6417 = ~pi0263 & ~n5559;
  assign n6418 = ~n6416 & ~n6417;
  assign n6419 = n5292 & ~n6418;
  assign n6420 = pi1579 & n5296;
  assign n6421 = pi1604 & n5357;
  assign n6422 = pi1555 & n5295;
  assign n6423 = pi0989 & n5555;
  assign n6424 = ~n6422 & ~n6423;
  assign n6425 = ~n6421 & n6424;
  assign n6426 = ~n6420 & n6425;
  assign n6427 = n5550 & ~n6426;
  assign n6428 = ~n5549 & n5560;
  assign n6429 = ~n6427 & ~n6428;
  assign n6430 = ~n6419 & n6429;
  assign n6431 = n5291 & ~n6430;
  assign n6432 = ~pi0290 & ~n5291;
  assign n6433 = ~n6431 & ~n6432;
  assign po0341 = pi1839 & ~n6433;
  assign n6435 = pi0263 & ~n6304;
  assign n6436 = ~pi0263 & ~n5573;
  assign n6437 = ~n6435 & ~n6436;
  assign n6438 = n5292 & ~n6437;
  assign n6439 = n5560 & ~n5581;
  assign n6440 = pi1605 & n5357;
  assign n6441 = pi1727 & n5555;
  assign n6442 = pi1580 & n5296;
  assign n6443 = pi1556 & n5295;
  assign n6444 = ~n6442 & ~n6443;
  assign n6445 = ~n6441 & n6444;
  assign n6446 = ~n6440 & n6445;
  assign n6447 = n5550 & ~n6446;
  assign n6448 = ~n6439 & ~n6447;
  assign n6449 = ~n6438 & n6448;
  assign n6450 = n5291 & ~n6449;
  assign n6451 = ~pi0291 & ~n5291;
  assign n6452 = ~n6450 & ~n6451;
  assign po0342 = pi1839 & ~n6452;
  assign n6454 = ~pi0263 & ~n5549;
  assign n6455 = pi0263 & ~n6408;
  assign n6456 = ~n6454 & ~n6455;
  assign n6457 = n5292 & ~n6456;
  assign n6458 = n5560 & ~n6426;
  assign n6459 = n5550 & ~n6143;
  assign n6460 = ~n6458 & ~n6459;
  assign n6461 = ~n6457 & n6460;
  assign n6462 = n5291 & ~n6461;
  assign n6463 = ~pi0292 & ~n5291;
  assign n6464 = ~n6462 & ~n6463;
  assign po0343 = pi1839 & ~n6464;
  assign n6466 = ~pi0293 & ~n5291;
  assign n6467 = ~pi0263 & ~n5581;
  assign n6468 = pi0263 & ~n6356;
  assign n6469 = ~n6467 & ~n6468;
  assign n6470 = n5292 & ~n6469;
  assign n6471 = n5550 & ~n6184;
  assign n6472 = n5560 & ~n6446;
  assign n6473 = ~n6471 & ~n6472;
  assign n6474 = ~n6470 & n6473;
  assign n6475 = n5291 & ~n6474;
  assign n6476 = ~n6466 & ~n6475;
  assign po0344 = pi1839 & ~n6476;
  assign n6478 = ~pi0263 & ~n6426;
  assign n6479 = pi1569 & n5296;
  assign n6480 = pi1015 & n5555;
  assign n6481 = pi1593 & n5357;
  assign n6482 = pi1545 & n5295;
  assign n6483 = ~n6481 & ~n6482;
  assign n6484 = ~n6480 & n6483;
  assign n6485 = ~n6479 & n6484;
  assign n6486 = pi0263 & ~n6485;
  assign n6487 = ~n6478 & ~n6486;
  assign n6488 = n5292 & ~n6487;
  assign n6489 = n5560 & ~n6143;
  assign n6490 = n5550 & ~n6161;
  assign n6491 = ~n6489 & ~n6490;
  assign n6492 = ~n6488 & n6491;
  assign n6493 = n5291 & ~n6492;
  assign n6494 = ~pi0294 & ~n5291;
  assign n6495 = ~n6493 & ~n6494;
  assign po0345 = pi1839 & ~n6495;
  assign n6497 = ~pi0295 & ~n5291;
  assign n6498 = ~pi0263 & ~n6446;
  assign n6499 = pi1115 & n5296;
  assign n6500 = pi1702 & n5295;
  assign n6501 = pi1096 & n5357;
  assign n6502 = pi1719 & n5555;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = ~n6500 & n6503;
  assign n6505 = ~n6499 & n6504;
  assign n6506 = pi0263 & ~n6505;
  assign n6507 = ~n6498 & ~n6506;
  assign n6508 = n5292 & ~n6507;
  assign n6509 = n5560 & ~n6184;
  assign n6510 = n5550 & ~n6201;
  assign n6511 = ~n6509 & ~n6510;
  assign n6512 = ~n6508 & n6511;
  assign n6513 = n5291 & ~n6512;
  assign n6514 = ~n6497 & ~n6513;
  assign po0346 = pi1839 & ~n6514;
  assign n6516 = pi1069 & n5325;
  assign n6517 = pi1284 & n5258;
  assign n6518 = pi1243 & n5257;
  assign n6519 = pi1010 & n5591;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = ~n6517 & n6520;
  assign n6522 = ~n6516 & n6521;
  assign n6523 = ~pi0261 & ~n6522;
  assign n6524 = pi1070 & n5325;
  assign n6525 = pi1092 & n5258;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = pi1025 & n5257;
  assign n6528 = pi1740 & n5591;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = n6526 & n6529;
  assign n6531 = pi0261 & ~n6530;
  assign n6532 = ~n6523 & ~n6531;
  assign n6533 = n5254 & ~n6532;
  assign n6534 = pi1288 & n5325;
  assign n6535 = pi1255 & n5258;
  assign n6536 = pi1729 & n5591;
  assign n6537 = pi1625 & n5257;
  assign n6538 = ~n6536 & ~n6537;
  assign n6539 = ~n6535 & n6538;
  assign n6540 = ~n6534 & n6539;
  assign n6541 = n5596 & ~n6540;
  assign n6542 = pi1534 & n5325;
  assign n6543 = pi1086 & n5258;
  assign n6544 = pi1248 & n5257;
  assign n6545 = pi1754 & n5591;
  assign n6546 = ~n6544 & ~n6545;
  assign n6547 = ~n6543 & n6546;
  assign n6548 = ~n6542 & n6547;
  assign n6549 = n5605 & ~n6548;
  assign n6550 = ~n6541 & ~n6549;
  assign n6551 = ~n6533 & n6550;
  assign n6552 = n5253 & ~n6551;
  assign n6553 = ~pi0296 & ~n5253;
  assign n6554 = ~n6552 & ~n6553;
  assign po0347 = pi1164 & ~n6554;
  assign n6556 = pi1085 & n5325;
  assign n6557 = pi1099 & n5258;
  assign n6558 = pi0992 & n5591;
  assign n6559 = pi1050 & n5257;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = ~n6557 & n6560;
  assign n6562 = ~n6556 & n6561;
  assign n6563 = n5596 & ~n6562;
  assign n6564 = pi1308 & n5325;
  assign n6565 = pi1286 & n5258;
  assign n6566 = pi1251 & n5257;
  assign n6567 = pi1776 & n5591;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = ~n6565 & n6568;
  assign n6570 = ~n6564 & n6569;
  assign n6571 = n5605 & ~n6570;
  assign n6572 = ~n6563 & ~n6571;
  assign n6573 = pi0261 & n5254;
  assign n6574 = pi1658 & n5257;
  assign n6575 = pi1807 & n5591;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = pi1298 & n5325;
  assign n6578 = pi1273 & n5258;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = n6576 & n6579;
  assign n6581 = n6573 & ~n6580;
  assign n6582 = pi1307 & n5325;
  assign n6583 = pi1285 & n5258;
  assign n6584 = pi1245 & n5257;
  assign n6585 = pi1855 & n5591;
  assign n6586 = ~n6584 & ~n6585;
  assign n6587 = ~n6583 & n6586;
  assign n6588 = ~n6582 & n6587;
  assign n6589 = ~pi0261 & n5254;
  assign n6590 = ~n6588 & n6589;
  assign n6591 = ~n6581 & ~n6590;
  assign n6592 = n6572 & n6591;
  assign n6593 = n5253 & ~n6592;
  assign n6594 = ~pi0297 & ~n5253;
  assign n6595 = ~n6593 & ~n6594;
  assign po0348 = pi1164 & ~n6595;
  assign n6597 = pi1290 & n5325;
  assign n6598 = pi1262 & n5258;
  assign n6599 = pi1632 & n5257;
  assign n6600 = pi1058 & n5591;
  assign n6601 = ~n6599 & ~n6600;
  assign n6602 = ~n6598 & n6601;
  assign n6603 = ~n6597 & n6602;
  assign n6604 = n5596 & ~n6603;
  assign n6605 = n5605 & ~n6562;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = ~pi0261 & ~n6570;
  assign n6608 = n5254 & n6607;
  assign n6609 = pi1662 & n5257;
  assign n6610 = pi1745 & n5591;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = pi1309 & n5325;
  assign n6613 = pi1275 & n5258;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = n6611 & n6614;
  assign n6616 = n6573 & ~n6615;
  assign n6617 = ~n6608 & ~n6616;
  assign n6618 = n6606 & n6617;
  assign n6619 = n5253 & ~n6618;
  assign n6620 = ~pi0298 & ~n5253;
  assign n6621 = ~n6619 & ~n6620;
  assign po0349 = pi1164 & ~n6621;
  assign n6623 = ~pi0299 & ~n5253;
  assign n6624 = ~pi0261 & ~n6540;
  assign n6625 = pi1300 & n5325;
  assign n6626 = pi1091 & n5258;
  assign n6627 = ~n6625 & ~n6626;
  assign n6628 = pi1824 & n5257;
  assign n6629 = pi1746 & n5591;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = n6627 & n6630;
  assign n6632 = pi0261 & ~n6631;
  assign n6633 = ~n6624 & ~n6632;
  assign n6634 = n5254 & ~n6633;
  assign n6635 = pi1634 & n5257;
  assign n6636 = pi1291 & n5325;
  assign n6637 = pi1854 & n5591;
  assign n6638 = pi1264 & n5258;
  assign n6639 = ~n6637 & ~n6638;
  assign n6640 = ~n6636 & n6639;
  assign n6641 = ~n6635 & n6640;
  assign n6642 = n5596 & ~n6641;
  assign n6643 = pi1260 & n5258;
  assign n6644 = pi1289 & n5325;
  assign n6645 = pi1630 & n5257;
  assign n6646 = pi0993 & n5591;
  assign n6647 = ~n6645 & ~n6646;
  assign n6648 = ~n6644 & n6647;
  assign n6649 = ~n6643 & n6648;
  assign n6650 = n5605 & ~n6649;
  assign n6651 = ~n6642 & ~n6650;
  assign n6652 = ~n6634 & n6651;
  assign n6653 = n5253 & ~n6652;
  assign n6654 = ~n6623 & ~n6653;
  assign po0350 = pi1164 & ~n6654;
  assign n6656 = ~pi0300 & ~n5253;
  assign n6657 = ~pi0261 & ~n6562;
  assign n6658 = pi1072 & n5325;
  assign n6659 = pi1276 & n5258;
  assign n6660 = ~n6658 & ~n6659;
  assign n6661 = pi1667 & n5257;
  assign n6662 = pi1005 & n5591;
  assign n6663 = ~n6661 & ~n6662;
  assign n6664 = n6660 & n6663;
  assign n6665 = pi0261 & ~n6664;
  assign n6666 = ~n6657 & ~n6665;
  assign n6667 = n5254 & ~n6666;
  assign n6668 = n5605 & ~n6603;
  assign n6669 = pi1084 & n5325;
  assign n6670 = pi1266 & n5258;
  assign n6671 = pi1043 & n5257;
  assign n6672 = pi0994 & n5591;
  assign n6673 = ~n6671 & ~n6672;
  assign n6674 = ~n6670 & n6673;
  assign n6675 = ~n6669 & n6674;
  assign n6676 = n5596 & ~n6675;
  assign n6677 = ~n6668 & ~n6676;
  assign n6678 = ~n6667 & n6677;
  assign n6679 = n5253 & ~n6678;
  assign n6680 = ~n6656 & ~n6679;
  assign po0351 = pi1164 & ~n6680;
  assign n6682 = ~pi0301 & ~n5253;
  assign n6683 = ~pi0261 & ~n6649;
  assign n6684 = pi1301 & n5325;
  assign n6685 = pi1277 & n5258;
  assign n6686 = ~n6684 & ~n6685;
  assign n6687 = pi1225 & n5257;
  assign n6688 = pi1747 & n5591;
  assign n6689 = ~n6687 & ~n6688;
  assign n6690 = n6686 & n6689;
  assign n6691 = pi0261 & ~n6690;
  assign n6692 = ~n6683 & ~n6691;
  assign n6693 = n5254 & ~n6692;
  assign n6694 = n5605 & ~n6641;
  assign n6695 = pi1292 & n5325;
  assign n6696 = pi1268 & n5258;
  assign n6697 = pi1639 & n5257;
  assign n6698 = pi1031 & n5591;
  assign n6699 = ~n6697 & ~n6698;
  assign n6700 = ~n6696 & n6699;
  assign n6701 = ~n6695 & n6700;
  assign n6702 = n5596 & ~n6701;
  assign n6703 = ~n6694 & ~n6702;
  assign n6704 = ~n6693 & n6703;
  assign n6705 = n5253 & ~n6704;
  assign n6706 = ~n6682 & ~n6705;
  assign po0352 = pi1164 & ~n6706;
  assign n6708 = pi1293 & n5325;
  assign n6709 = pi1269 & n5258;
  assign n6710 = pi1642 & n5257;
  assign n6711 = pi1013 & n5591;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~n6709 & n6712;
  assign n6714 = ~n6708 & n6713;
  assign n6715 = n5596 & ~n6714;
  assign n6716 = n5605 & ~n6675;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = pi1227 & n5257;
  assign n6719 = pi1009 & n5591;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = pi1302 & n5325;
  assign n6722 = pi1278 & n5258;
  assign n6723 = ~n6721 & ~n6722;
  assign n6724 = n6720 & n6723;
  assign n6725 = n6573 & ~n6724;
  assign n6726 = n6589 & ~n6603;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = n6717 & n6727;
  assign n6729 = n5253 & ~n6728;
  assign n6730 = ~pi0302 & ~n5253;
  assign n6731 = ~n6729 & ~n6730;
  assign po0353 = pi1164 & ~n6731;
  assign n6733 = ~pi0303 & ~n5253;
  assign n6734 = ~pi0261 & ~n6641;
  assign n6735 = pi1071 & n5325;
  assign n6736 = pi1279 & n5258;
  assign n6737 = ~n6735 & ~n6736;
  assign n6738 = pi1232 & n5257;
  assign n6739 = pi1752 & n5591;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = n6737 & n6740;
  assign n6742 = pi0261 & ~n6741;
  assign n6743 = ~n6734 & ~n6742;
  assign n6744 = n5254 & ~n6743;
  assign n6745 = pi1294 & n5325;
  assign n6746 = pi1093 & n5258;
  assign n6747 = pi1644 & n5257;
  assign n6748 = pi1732 & n5591;
  assign n6749 = ~n6747 & ~n6748;
  assign n6750 = ~n6746 & n6749;
  assign n6751 = ~n6745 & n6750;
  assign n6752 = n5596 & ~n6751;
  assign n6753 = n5605 & ~n6701;
  assign n6754 = ~n6752 & ~n6753;
  assign n6755 = ~n6744 & n6754;
  assign n6756 = n5253 & ~n6755;
  assign n6757 = ~n6733 & ~n6756;
  assign po0354 = pi1164 & ~n6757;
  assign n6759 = pi1095 & n5309;
  assign n6760 = pi1121 & n5239;
  assign n6761 = pi1750 & n5635;
  assign n6762 = pi1034 & n5238;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = ~n6760 & n6763;
  assign n6765 = ~n6759 & n6764;
  assign n6766 = ~pi0260 & ~n6765;
  assign n6767 = pi1655 & n5239;
  assign n6768 = pi1619 & n5238;
  assign n6769 = pi1103 & n5309;
  assign n6770 = pi1820 & n5635;
  assign n6771 = ~n6769 & ~n6770;
  assign n6772 = ~n6768 & n6771;
  assign n6773 = ~n6767 & n6772;
  assign n6774 = pi0260 & ~n6773;
  assign n6775 = ~n6766 & ~n6774;
  assign n6776 = n5235 & ~n6775;
  assign n6777 = pi1111 & n5309;
  assign n6778 = pi1640 & n5239;
  assign n6779 = pi1730 & n5635;
  assign n6780 = pi1082 & n5238;
  assign n6781 = ~n6779 & ~n6780;
  assign n6782 = ~n6778 & n6781;
  assign n6783 = ~n6777 & n6782;
  assign n6784 = n5642 & ~n6783;
  assign n6785 = pi1094 & n5309;
  assign n6786 = pi1229 & n5239;
  assign n6787 = pi1749 & n5635;
  assign n6788 = pi1636 & n5238;
  assign n6789 = ~n6787 & ~n6788;
  assign n6790 = ~n6786 & n6789;
  assign n6791 = ~n6785 & n6790;
  assign n6792 = n5651 & ~n6791;
  assign n6793 = ~n6784 & ~n6792;
  assign n6794 = ~n6776 & n6793;
  assign n6795 = n5234 & ~n6794;
  assign n6796 = ~pi0304 & ~n5234;
  assign n6797 = ~n6795 & ~n6796;
  assign po0355 = pi1838 & ~n6797;
  assign n6799 = ~pi0305 & ~n5253;
  assign n6800 = ~pi0261 & ~n6675;
  assign n6801 = pi1304 & n5325;
  assign n6802 = pi1280 & n5258;
  assign n6803 = ~n6801 & ~n6802;
  assign n6804 = pi1234 & n5257;
  assign n6805 = pi1872 & n5591;
  assign n6806 = ~n6804 & ~n6805;
  assign n6807 = n6803 & n6806;
  assign n6808 = pi0261 & ~n6807;
  assign n6809 = ~n6800 & ~n6808;
  assign n6810 = n5254 & ~n6809;
  assign n6811 = pi1074 & n5325;
  assign n6812 = pi1270 & n5258;
  assign n6813 = pi1038 & n5257;
  assign n6814 = pi1734 & n5591;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = ~n6812 & n6815;
  assign n6817 = ~n6811 & n6816;
  assign n6818 = n5596 & ~n6817;
  assign n6819 = n5605 & ~n6714;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = ~n6810 & n6820;
  assign n6822 = n5253 & ~n6821;
  assign n6823 = ~n6799 & ~n6822;
  assign po0356 = pi1164 & ~n6823;
  assign n6825 = pi1265 & n5309;
  assign n6826 = pi1228 & n5239;
  assign n6827 = pi1748 & n5635;
  assign n6828 = pi1635 & n5238;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = ~n6826 & n6829;
  assign n6831 = ~n6825 & n6830;
  assign n6832 = ~pi0260 & ~n6831;
  assign n6833 = pi1249 & n5309;
  assign n6834 = pi1656 & n5239;
  assign n6835 = ~n6833 & ~n6834;
  assign n6836 = pi1620 & n5238;
  assign n6837 = pi1741 & n5635;
  assign n6838 = ~n6836 & ~n6837;
  assign n6839 = n6835 & n6838;
  assign n6840 = pi0260 & ~n6839;
  assign n6841 = ~n6832 & ~n6840;
  assign n6842 = n5235 & ~n6841;
  assign n6843 = pi1233 & n5309;
  assign n6844 = pi1641 & n5239;
  assign n6845 = pi0996 & n5635;
  assign n6846 = pi1610 & n5238;
  assign n6847 = ~n6845 & ~n6846;
  assign n6848 = ~n6844 & n6847;
  assign n6849 = ~n6843 & n6848;
  assign n6850 = n5642 & ~n6849;
  assign n6851 = pi1267 & n5309;
  assign n6852 = pi1637 & n5238;
  assign n6853 = pi1751 & n5635;
  assign n6854 = pi1230 & n5239;
  assign n6855 = ~n6853 & ~n6854;
  assign n6856 = ~n6852 & n6855;
  assign n6857 = ~n6851 & n6856;
  assign n6858 = n5651 & ~n6857;
  assign n6859 = ~n6850 & ~n6858;
  assign n6860 = ~n6842 & n6859;
  assign n6861 = n5234 & ~n6860;
  assign n6862 = ~pi0306 & ~n5234;
  assign n6863 = ~n6861 & ~n6862;
  assign po0357 = pi1838 & ~n6863;
  assign n6865 = ~pi0260 & ~n6791;
  assign n6866 = pi1250 & n5309;
  assign n6867 = pi1657 & n5239;
  assign n6868 = ~n6866 & ~n6867;
  assign n6869 = pi1621 & n5238;
  assign n6870 = pi1742 & n5635;
  assign n6871 = ~n6869 & ~n6870;
  assign n6872 = n6868 & n6871;
  assign n6873 = pi0260 & ~n6872;
  assign n6874 = ~n6865 & ~n6873;
  assign n6875 = n5235 & ~n6874;
  assign n6876 = pi1235 & n5309;
  assign n6877 = pi1611 & n5238;
  assign n6878 = pi0997 & n5635;
  assign n6879 = pi1643 & n5239;
  assign n6880 = ~n6878 & ~n6879;
  assign n6881 = ~n6877 & n6880;
  assign n6882 = ~n6876 & n6881;
  assign n6883 = n5642 & ~n6882;
  assign n6884 = n5651 & ~n6783;
  assign n6885 = ~n6883 & ~n6884;
  assign n6886 = ~n6875 & n6885;
  assign n6887 = n5234 & ~n6886;
  assign n6888 = ~pi0307 & ~n5234;
  assign n6889 = ~n6887 & ~n6888;
  assign po0358 = pi1838 & ~n6889;
  assign n6891 = ~pi0261 & ~n6548;
  assign n6892 = pi1299 & n5325;
  assign n6893 = pi1274 & n5258;
  assign n6894 = ~n6892 & ~n6893;
  assign n6895 = pi1660 & n5257;
  assign n6896 = pi1744 & n5591;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = n6894 & n6897;
  assign n6899 = pi0261 & ~n6898;
  assign n6900 = ~n6891 & ~n6899;
  assign n6901 = n5254 & ~n6900;
  assign n6902 = n5596 & ~n6649;
  assign n6903 = n5605 & ~n6540;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = ~n6901 & n6904;
  assign n6906 = n5253 & ~n6905;
  assign n6907 = ~pi0308 & ~n5253;
  assign n6908 = ~n6906 & ~n6907;
  assign po0359 = pi1164 & ~n6908;
  assign n6910 = ~pi0260 & ~n6857;
  assign n6911 = pi1104 & n5309;
  assign n6912 = pi1016 & n5239;
  assign n6913 = ~n6911 & ~n6912;
  assign n6914 = pi1059 & n5238;
  assign n6915 = pi1743 & n5635;
  assign n6916 = ~n6914 & ~n6915;
  assign n6917 = n6913 & n6916;
  assign n6918 = pi0260 & ~n6917;
  assign n6919 = ~n6910 & ~n6918;
  assign n6920 = n5235 & ~n6919;
  assign n6921 = pi1236 & n5309;
  assign n6922 = pi1037 & n5239;
  assign n6923 = pi1731 & n5635;
  assign n6924 = pi1612 & n5238;
  assign n6925 = ~n6923 & ~n6924;
  assign n6926 = ~n6922 & n6925;
  assign n6927 = ~n6921 & n6926;
  assign n6928 = n5642 & ~n6927;
  assign n6929 = n5651 & ~n6849;
  assign n6930 = ~n6928 & ~n6929;
  assign n6931 = ~n6920 & n6930;
  assign n6932 = n5234 & ~n6931;
  assign n6933 = ~pi0309 & ~n5234;
  assign n6934 = ~n6932 & ~n6933;
  assign po0360 = pi1838 & ~n6934;
  assign n6936 = ~pi0260 & ~n6783;
  assign n6937 = pi1252 & n5309;
  assign n6938 = pi1659 & n5239;
  assign n6939 = ~n6937 & ~n6938;
  assign n6940 = pi1622 & n5238;
  assign n6941 = pi1001 & n5635;
  assign n6942 = ~n6940 & ~n6941;
  assign n6943 = n6939 & n6942;
  assign n6944 = pi0260 & ~n6943;
  assign n6945 = ~n6936 & ~n6944;
  assign n6946 = n5235 & ~n6945;
  assign n6947 = pi1238 & n5309;
  assign n6948 = pi1645 & n5239;
  assign n6949 = pi1733 & n5635;
  assign n6950 = pi1067 & n5238;
  assign n6951 = ~n6949 & ~n6950;
  assign n6952 = ~n6948 & n6951;
  assign n6953 = ~n6947 & n6952;
  assign n6954 = n5642 & ~n6953;
  assign n6955 = n5651 & ~n6882;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~n6946 & n6956;
  assign n6958 = n5234 & ~n6957;
  assign n6959 = ~pi0310 & ~n5234;
  assign n6960 = ~n6958 & ~n6959;
  assign po0361 = pi1838 & ~n6960;
  assign n6962 = pi0261 & ~n6701;
  assign n6963 = ~pi0261 & ~n5604;
  assign n6964 = ~n6962 & ~n6963;
  assign n6965 = n5254 & ~n6964;
  assign n6966 = pi1305 & n5325;
  assign n6967 = pi1282 & n5258;
  assign n6968 = pi1781 & n5591;
  assign n6969 = pi1237 & n5257;
  assign n6970 = ~n6968 & ~n6969;
  assign n6971 = ~n6967 & n6970;
  assign n6972 = ~n6966 & n6971;
  assign n6973 = n5596 & ~n6972;
  assign n6974 = ~n5595 & n5605;
  assign n6975 = ~n6973 & ~n6974;
  assign n6976 = ~n6965 & n6975;
  assign n6977 = n5253 & ~n6976;
  assign n6978 = ~pi0311 & ~n5253;
  assign n6979 = ~n6977 & ~n6978;
  assign po0362 = pi1164 & ~n6979;
  assign n6981 = ~pi0260 & ~n6882;
  assign n6982 = pi1100 & n5309;
  assign n6983 = pi1017 & n5239;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = pi1057 & n5238;
  assign n6986 = pi1002 & n5635;
  assign n6987 = ~n6985 & ~n6986;
  assign n6988 = n6984 & n6987;
  assign n6989 = pi0260 & ~n6988;
  assign n6990 = ~n6981 & ~n6989;
  assign n6991 = n5235 & ~n6990;
  assign n6992 = pi1239 & n5309;
  assign n6993 = pi1614 & n5238;
  assign n6994 = pi1647 & n5239;
  assign n6995 = ~pi0216 & pi1800;
  assign n6996 = ~pi0224 & n6995;
  assign n6997 = ~n6994 & ~n6996;
  assign n6998 = ~n6993 & n6997;
  assign n6999 = ~n6992 & n6998;
  assign n7000 = n5642 & ~n6999;
  assign n7001 = n5651 & ~n6953;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = ~n6991 & n7002;
  assign n7004 = n5234 & ~n7003;
  assign n7005 = ~pi0312 & ~n5234;
  assign n7006 = ~n7004 & ~n7005;
  assign po0363 = pi1838 & ~n7006;
  assign n7008 = pi0261 & ~n6751;
  assign n7009 = ~pi0261 & ~n5595;
  assign n7010 = ~n7008 & ~n7009;
  assign n7011 = n5254 & ~n7010;
  assign n7012 = n5596 & ~n6522;
  assign n7013 = n5605 & ~n6972;
  assign n7014 = ~n7012 & ~n7013;
  assign n7015 = ~n7011 & n7014;
  assign n7016 = n5253 & ~n7015;
  assign n7017 = ~pi0313 & ~n5253;
  assign n7018 = ~n7016 & ~n7017;
  assign po0364 = pi1164 & ~n7018;
  assign n7020 = ~pi0260 & ~n6927;
  assign n7021 = pi1256 & n5309;
  assign n7022 = pi1663 & n5239;
  assign n7023 = ~n7021 & ~n7022;
  assign n7024 = pi1626 & n5238;
  assign n7025 = pi1003 & n5635;
  assign n7026 = ~n7024 & ~n7025;
  assign n7027 = n7023 & n7026;
  assign n7028 = pi0260 & ~n7027;
  assign n7029 = ~n7020 & ~n7028;
  assign n7030 = n5235 & ~n7029;
  assign n7031 = pi1240 & n5309;
  assign n7032 = pi1648 & n5239;
  assign n7033 = pi0998 & n5635;
  assign n7034 = pi1615 & n5238;
  assign n7035 = ~n7033 & ~n7034;
  assign n7036 = ~n7032 & n7035;
  assign n7037 = ~n7031 & n7036;
  assign n7038 = n5642 & ~n7037;
  assign n7039 = pi1110 & n5309;
  assign n7040 = pi1646 & n5239;
  assign n7041 = pi1030 & n5635;
  assign n7042 = pi1613 & n5238;
  assign n7043 = ~n7041 & ~n7042;
  assign n7044 = ~n7040 & n7043;
  assign n7045 = ~n7039 & n7044;
  assign n7046 = n5651 & ~n7045;
  assign n7047 = ~n7038 & ~n7046;
  assign n7048 = ~n7030 & n7047;
  assign n7049 = n5234 & ~n7048;
  assign n7050 = ~pi0314 & ~n5234;
  assign n7051 = ~n7049 & ~n7050;
  assign po0365 = pi1838 & ~n7051;
  assign n7053 = pi0261 & ~n6817;
  assign n7054 = ~pi0261 & ~n5618;
  assign n7055 = ~n7053 & ~n7054;
  assign n7056 = n5254 & ~n7055;
  assign n7057 = n5596 & ~n6588;
  assign n7058 = pi1306 & n5325;
  assign n7059 = pi1283 & n5258;
  assign n7060 = pi1241 & n5257;
  assign n7061 = pi1011 & n5591;
  assign n7062 = ~n7060 & ~n7061;
  assign n7063 = ~n7059 & n7062;
  assign n7064 = ~n7058 & n7063;
  assign n7065 = n5605 & ~n7064;
  assign n7066 = ~n7057 & ~n7065;
  assign n7067 = ~n7056 & n7066;
  assign n7068 = n5253 & ~n7067;
  assign n7069 = ~pi0315 & ~n5253;
  assign n7070 = ~n7068 & ~n7069;
  assign po0366 = pi1164 & ~n7070;
  assign n7072 = ~pi0260 & ~n6953;
  assign n7073 = pi1258 & n5309;
  assign n7074 = pi1665 & n5239;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = pi1628 & n5238;
  assign n7077 = pi1004 & n5635;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = n7075 & n7078;
  assign n7080 = pi0260 & ~n7079;
  assign n7081 = ~n7072 & ~n7080;
  assign n7082 = n5235 & ~n7081;
  assign n7083 = pi1108 & n5309;
  assign n7084 = pi1068 & n5238;
  assign n7085 = pi1014 & n5239;
  assign n7086 = pi1735 & n5635;
  assign n7087 = ~n7085 & ~n7086;
  assign n7088 = ~n7084 & n7087;
  assign n7089 = ~n7083 & n7088;
  assign n7090 = n5642 & ~n7089;
  assign n7091 = n5651 & ~n6999;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = ~n7082 & n7092;
  assign n7094 = n5234 & ~n7093;
  assign n7095 = ~pi0316 & ~n5234;
  assign n7096 = ~n7094 & ~n7095;
  assign po0367 = pi1838 & ~n7096;
  assign n7098 = ~pi0261 & ~n6972;
  assign n7099 = pi1296 & n5325;
  assign n7100 = pi1385 & n5258;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = pi1651 & n5257;
  assign n7103 = pi1737 & n5591;
  assign n7104 = ~n7102 & ~n7103;
  assign n7105 = n7101 & n7104;
  assign n7106 = pi0261 & ~n7105;
  assign n7107 = ~n7098 & ~n7106;
  assign n7108 = n5254 & ~n7107;
  assign n7109 = n5596 & ~n6548;
  assign n7110 = n5605 & ~n6522;
  assign n7111 = ~n7109 & ~n7110;
  assign n7112 = ~n7108 & n7111;
  assign n7113 = n5253 & ~n7112;
  assign n7114 = ~pi0317 & ~n5253;
  assign n7115 = ~n7113 & ~n7114;
  assign po0368 = pi1164 & ~n7115;
  assign n7117 = ~pi0260 & ~n6849;
  assign n7118 = pi1254 & n5309;
  assign n7119 = pi1661 & n5239;
  assign n7120 = ~n7118 & ~n7119;
  assign n7121 = pi1624 & n5238;
  assign n7122 = pi1814 & n5635;
  assign n7123 = ~n7121 & ~n7122;
  assign n7124 = n7120 & n7123;
  assign n7125 = pi0260 & ~n7124;
  assign n7126 = ~n7117 & ~n7125;
  assign n7127 = n5235 & ~n7126;
  assign n7128 = n5642 & ~n7045;
  assign n7129 = n5651 & ~n6927;
  assign n7130 = ~n7128 & ~n7129;
  assign n7131 = ~n7127 & n7130;
  assign n7132 = n5234 & ~n7131;
  assign n7133 = ~pi0318 & ~n5234;
  assign n7134 = ~n7132 & ~n7133;
  assign po0369 = pi1838 & ~n7134;
  assign n7136 = pi0261 & ~n6714;
  assign n7137 = ~pi0261 & ~n5627;
  assign n7138 = ~n7136 & ~n7137;
  assign n7139 = n5254 & ~n7138;
  assign n7140 = n5596 & ~n7064;
  assign n7141 = n5605 & ~n5618;
  assign n7142 = ~n7140 & ~n7141;
  assign n7143 = ~n7139 & n7142;
  assign n7144 = n5253 & ~n7143;
  assign n7145 = ~pi0319 & ~n5253;
  assign n7146 = ~n7144 & ~n7145;
  assign po0370 = pi1164 & ~n7146;
  assign n7148 = ~pi0260 & ~n7045;
  assign n7149 = pi1259 & n5309;
  assign n7150 = pi1666 & n5239;
  assign n7151 = ~n7149 & ~n7150;
  assign n7152 = pi1629 & n5238;
  assign n7153 = pi1783 & n5635;
  assign n7154 = ~n7152 & ~n7153;
  assign n7155 = n7151 & n7154;
  assign n7156 = pi0260 & ~n7155;
  assign n7157 = ~n7148 & ~n7156;
  assign n7158 = n5235 & ~n7157;
  assign n7159 = pi1242 & n5309;
  assign n7160 = pi1650 & n5239;
  assign n7161 = pi1616 & n5238;
  assign n7162 = pi1736 & n5635;
  assign n7163 = ~n7161 & ~n7162;
  assign n7164 = ~n7160 & n7163;
  assign n7165 = ~n7159 & n7164;
  assign n7166 = n5642 & ~n7165;
  assign n7167 = n5651 & ~n7037;
  assign n7168 = ~n7166 & ~n7167;
  assign n7169 = ~n7158 & n7168;
  assign n7170 = n5234 & ~n7169;
  assign n7171 = ~pi0320 & ~n5234;
  assign n7172 = ~n7170 & ~n7171;
  assign po0371 = pi1838 & ~n7172;
  assign n7174 = ~pi0261 & ~n7064;
  assign n7175 = pi1297 & n5325;
  assign n7176 = pi1272 & n5258;
  assign n7177 = ~n7175 & ~n7176;
  assign n7178 = pi1653 & n5257;
  assign n7179 = pi1000 & n5591;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = n7177 & n7180;
  assign n7182 = pi0261 & ~n7181;
  assign n7183 = ~n7174 & ~n7182;
  assign n7184 = n5254 & ~n7183;
  assign n7185 = n5596 & ~n6570;
  assign n7186 = n5605 & ~n6588;
  assign n7187 = ~n7185 & ~n7186;
  assign n7188 = ~n7184 & n7187;
  assign n7189 = n5253 & ~n7188;
  assign n7190 = ~pi0321 & ~n5253;
  assign n7191 = ~n7189 & ~n7190;
  assign po0372 = pi1164 & ~n7191;
  assign n7193 = ~pi0260 & ~n5650;
  assign n7194 = pi0260 & ~n6999;
  assign n7195 = ~n7193 & ~n7194;
  assign n7196 = n5235 & ~n7195;
  assign n7197 = pi1261 & n5309;
  assign n7198 = pi1224 & n5239;
  assign n7199 = pi1006 & n5635;
  assign n7200 = pi1631 & n5238;
  assign n7201 = ~n7199 & ~n7200;
  assign n7202 = ~n7198 & n7201;
  assign n7203 = ~n7197 & n7202;
  assign n7204 = n5642 & ~n7203;
  assign n7205 = ~n5641 & n5651;
  assign n7206 = ~n7204 & ~n7205;
  assign n7207 = ~n7196 & n7206;
  assign n7208 = n5234 & ~n7207;
  assign n7209 = ~pi0322 & ~n5234;
  assign n7210 = ~n7208 & ~n7209;
  assign po0373 = pi1838 & ~n7210;
  assign n7212 = pi0260 & ~n7037;
  assign n7213 = ~pi0260 & ~n5672;
  assign n7214 = ~n7212 & ~n7213;
  assign n7215 = n5235 & ~n7214;
  assign n7216 = pi1263 & n5309;
  assign n7217 = pi1226 & n5239;
  assign n7218 = pi1633 & n5238;
  assign n7219 = pi1007 & n5635;
  assign n7220 = ~n7218 & ~n7219;
  assign n7221 = ~n7217 & n7220;
  assign n7222 = ~n7216 & n7221;
  assign n7223 = n5642 & ~n7222;
  assign n7224 = n5651 & ~n5664;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n7215 & n7225;
  assign n7227 = n5234 & ~n7226;
  assign n7228 = ~pi0323 & ~n5234;
  assign n7229 = ~n7227 & ~n7228;
  assign po0374 = pi1838 & ~n7229;
  assign n7231 = pi0260 & ~n7089;
  assign n7232 = ~pi0260 & ~n5641;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = n5235 & ~n7233;
  assign n7235 = n5642 & ~n6765;
  assign n7236 = n5651 & ~n7203;
  assign n7237 = ~n7235 & ~n7236;
  assign n7238 = ~n7234 & n7237;
  assign n7239 = n5234 & ~n7238;
  assign n7240 = ~pi0324 & ~n5234;
  assign n7241 = ~n7239 & ~n7240;
  assign po0375 = pi1838 & ~n7241;
  assign n7243 = pi0260 & ~n7165;
  assign n7244 = ~pi0260 & ~n5664;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = n5235 & ~n7245;
  assign n7247 = n5642 & ~n6831;
  assign n7248 = n5651 & ~n7222;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = ~n7246 & n7249;
  assign n7251 = n5234 & ~n7250;
  assign n7252 = ~pi0325 & ~n5234;
  assign n7253 = ~n7251 & ~n7252;
  assign po0376 = pi1838 & ~n7253;
  assign n7255 = ~pi0260 & ~n7203;
  assign n7256 = pi1246 & n5309;
  assign n7257 = pi1026 & n5239;
  assign n7258 = ~n7256 & ~n7257;
  assign n7259 = pi1618 & n5238;
  assign n7260 = pi1738 & n5635;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = n7258 & n7261;
  assign n7263 = pi0260 & ~n7262;
  assign n7264 = ~n7255 & ~n7263;
  assign n7265 = n5235 & ~n7264;
  assign n7266 = n5642 & ~n6791;
  assign n7267 = n5651 & ~n6765;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = ~n7265 & n7268;
  assign n7270 = n5234 & ~n7269;
  assign n7271 = ~pi0326 & ~n5234;
  assign n7272 = ~n7270 & ~n7271;
  assign po0377 = pi1838 & ~n7272;
  assign n7274 = ~pi0260 & ~n7222;
  assign n7275 = pi1247 & n5309;
  assign n7276 = pi1654 & n5239;
  assign n7277 = ~n7275 & ~n7276;
  assign n7278 = pi1049 & n5238;
  assign n7279 = pi1739 & n5635;
  assign n7280 = ~n7278 & ~n7279;
  assign n7281 = n7277 & n7280;
  assign n7282 = pi0260 & ~n7281;
  assign n7283 = ~n7274 & ~n7282;
  assign n7284 = n5235 & ~n7283;
  assign n7285 = n5642 & ~n6857;
  assign n7286 = n5651 & ~n6831;
  assign n7287 = ~n7285 & ~n7286;
  assign n7288 = ~n7284 & n7287;
  assign n7289 = n5234 & ~n7288;
  assign n7290 = ~pi0327 & ~n5234;
  assign n7291 = ~n7289 & ~n7290;
  assign po0378 = pi1838 & ~n7291;
  assign n7293 = ~pi0322 & ~pi2032;
  assign n7294 = pi0812 & pi2032;
  assign po0379 = n7293 | n7294;
  assign n7296 = pi0332 & ~pi2254;
  assign n7297 = pi0865 & ~pi2254;
  assign n7298 = pi1128 & pi1150;
  assign n7299 = pi2020 & n7298;
  assign n7300 = ~pi2008 & n7298;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = ~pi2137 & n7298;
  assign n7303 = n7301 & ~n7302;
  assign n7304 = ~pi1154 & ~pi1155;
  assign n7305 = ~n7303 & n7304;
  assign n7306 = pi1154 & pi1155;
  assign n7307 = n7299 & n7306;
  assign n7308 = ~n7305 & ~n7307;
  assign n7309 = ~pi2008 & ~pi2137;
  assign n7310 = n7298 & n7309;
  assign n7311 = ~n7299 & ~n7310;
  assign n7312 = ~pi1154 & pi1155;
  assign n7313 = ~n7311 & n7312;
  assign n7314 = n7308 & ~n7313;
  assign n7315 = pi1154 & ~pi1155;
  assign n7316 = ~n7301 & n7315;
  assign n7317 = n7314 & ~n7316;
  assign n7318 = n7297 & ~n7317;
  assign po0383 = n7296 | n7318;
  assign n7320 = pi0840 & ~pi2059;
  assign n7321 = pi0333 & pi2059;
  assign po0384 = n7320 | n7321;
  assign n7323 = pi0840 & ~pi2057;
  assign n7324 = pi0334 & pi2057;
  assign po0385 = n7323 | n7324;
  assign n7326 = pi0840 & ~pi2058;
  assign n7327 = pi0335 & pi2058;
  assign po0386 = n7326 | n7327;
  assign n7329 = pi0840 & ~pi2056;
  assign n7330 = pi0336 & pi2056;
  assign po0387 = n7329 | n7330;
  assign n7332 = pi1369 & n5455;
  assign n7333 = pi1344 & n5200;
  assign n7334 = pi1319 & n5199;
  assign n7335 = ~pi0214 & ~pi0236;
  assign n7336 = pi1673 & n7335;
  assign n7337 = ~n7334 & ~n7336;
  assign n7338 = ~n7333 & n7337;
  assign n7339 = ~n7332 & n7338;
  assign n7340 = ~pi1020 & pi1165;
  assign n7341 = ~n7339 & n7340;
  assign n7342 = pi1380 & n5455;
  assign n7343 = pi1355 & n5200;
  assign n7344 = pi1330 & n5199;
  assign n7345 = pi1681 & n7335;
  assign n7346 = ~n7344 & ~n7345;
  assign n7347 = ~n7343 & n7346;
  assign n7348 = ~n7342 & n7347;
  assign n7349 = pi1020 & ~pi1165;
  assign n7350 = ~n7348 & n7349;
  assign n7351 = ~n7341 & ~n7350;
  assign n7352 = n5196 & ~n7351;
  assign n7353 = ~pi0337 & ~n5196;
  assign n7354 = ~n7352 & ~n7353;
  assign po0388 = pi1035 & ~n7354;
  assign n7356 = pi1456 & n5481;
  assign n7357 = pi1406 & n5218;
  assign n7358 = pi1430 & n5219;
  assign n7359 = ~pi0215 & ~pi0238;
  assign n7360 = pi1696 & n7359;
  assign n7361 = ~n7358 & ~n7360;
  assign n7362 = ~n7357 & n7361;
  assign n7363 = ~n7356 & n7362;
  assign n7364 = ~pi1171 & pi1789;
  assign n7365 = ~n7363 & n7364;
  assign n7366 = pi1444 & n5481;
  assign n7367 = pi1395 & n5218;
  assign n7368 = pi1419 & n5219;
  assign n7369 = pi1688 & n7359;
  assign n7370 = ~n7368 & ~n7369;
  assign n7371 = ~n7367 & n7370;
  assign n7372 = ~n7366 & n7371;
  assign n7373 = pi1171 & ~pi1789;
  assign n7374 = ~n7372 & n7373;
  assign n7375 = ~n7365 & ~n7374;
  assign n7376 = n5215 & ~n7375;
  assign n7377 = ~pi0338 & ~n5215;
  assign n7378 = ~n7376 & ~n7377;
  assign po0389 = pi1169 & ~n7378;
  assign n7380 = pi1811 & n5481;
  assign n7381 = pi1822 & n5218;
  assign n7382 = pi1817 & n5219;
  assign n7383 = ~pi0215 & pi1694;
  assign n7384 = ~pi0238 & n7383;
  assign n7385 = ~n7382 & ~n7384;
  assign n7386 = ~n7381 & n7385;
  assign n7387 = ~n7380 & n7386;
  assign n7388 = n7364 & ~n7387;
  assign n7389 = pi1436 & n5481;
  assign n7390 = pi1386 & n5218;
  assign n7391 = pi1411 & n5219;
  assign n7392 = pi1796 & n7359;
  assign n7393 = ~n7391 & ~n7392;
  assign n7394 = ~n7390 & n7393;
  assign n7395 = ~n7389 & n7394;
  assign n7396 = n7373 & ~n7395;
  assign n7397 = ~n7388 & ~n7396;
  assign n7398 = n5215 & ~n7397;
  assign n7399 = ~pi0339 & ~n5215;
  assign n7400 = ~n7398 & ~n7399;
  assign po0390 = pi1169 & ~n7400;
  assign n7402 = pi1378 & n5455;
  assign n7403 = pi1353 & n5200;
  assign n7404 = pi1328 & n5199;
  assign n7405 = ~pi0214 & pi1679;
  assign n7406 = ~pi0236 & n7405;
  assign n7407 = ~n7404 & ~n7406;
  assign n7408 = ~n7403 & n7407;
  assign n7409 = ~n7402 & n7408;
  assign n7410 = n7349 & ~n7409;
  assign n7411 = pi1360 & n5455;
  assign n7412 = pi1335 & n5200;
  assign n7413 = pi1668 & n7335;
  assign n7414 = pi1310 & n5199;
  assign n7415 = ~n7413 & ~n7414;
  assign n7416 = ~n7412 & n7415;
  assign n7417 = ~n7411 & n7416;
  assign n7418 = n7340 & ~n7417;
  assign n7419 = ~n7410 & ~n7418;
  assign n7420 = n5196 & ~n7419;
  assign n7421 = ~pi0340 & ~n5196;
  assign n7422 = ~n7420 & ~n7421;
  assign po0391 = pi1035 & ~n7422;
  assign n7424 = ~pi0353 & ~n7417;
  assign n7425 = pi1040 & n5455;
  assign n7426 = pi1018 & n5200;
  assign n7427 = pi0954 & n7335;
  assign n7428 = pi1061 & n5199;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 = ~n7426 & n7429;
  assign n7431 = ~n7425 & n7430;
  assign n7432 = pi0353 & ~n7431;
  assign n7433 = ~n7424 & ~n7432;
  assign n7434 = n5197 & ~n7433;
  assign n7435 = pi1381 & n5455;
  assign n7436 = pi1356 & n5200;
  assign n7437 = pi0959 & n7335;
  assign n7438 = pi1331 & n5199;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = ~n7436 & n7439;
  assign n7441 = ~n7435 & n7440;
  assign n7442 = n7349 & ~n7441;
  assign n7443 = n7340 & ~n7409;
  assign n7444 = ~n7442 & ~n7443;
  assign n7445 = ~n7434 & n7444;
  assign n7446 = n5196 & ~n7445;
  assign n7447 = ~pi0345 & ~n5196;
  assign n7448 = ~n7446 & ~n7447;
  assign po0396 = pi1035 & ~n7448;
  assign po1885 = pi0929 & pi1943;
  assign n7451 = ~pi1834 & po1885;
  assign n7452 = pi0346 & ~n7451;
  assign n7453 = ~pi1138 & ~pi1152;
  assign n7454 = pi0411 & pi0412;
  assign n7455 = pi0346 & n7454;
  assign n7456 = ~pi0346 & ~n7454;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n7453 & n7457;
  assign n7459 = pi0411 & pi0635;
  assign n7460 = pi0412 & n7459;
  assign n7461 = pi0346 & ~n7460;
  assign n7462 = ~pi0346 & n7460;
  assign n7463 = ~n7461 & ~n7462;
  assign n7464 = n7453 & ~n7463;
  assign n7465 = ~n7458 & ~n7464;
  assign n7466 = n7451 & ~n7465;
  assign n7467 = ~n7452 & ~n7466;
  assign po0397 = pi1150 & ~n7467;
  assign n7469 = pi0347 & ~pi2252;
  assign n7470 = pi0874 & ~pi2252;
  assign n7471 = pi1145 & pi1161;
  assign n7472 = pi2033 & n7471;
  assign n7473 = ~pi2017 & n7471;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = ~pi2136 & n7471;
  assign n7476 = n7474 & ~n7475;
  assign n7477 = ~pi1159 & ~pi1160;
  assign n7478 = ~n7476 & n7477;
  assign n7479 = pi1159 & pi1160;
  assign n7480 = n7472 & n7479;
  assign n7481 = ~n7478 & ~n7480;
  assign n7482 = ~pi2017 & ~pi2136;
  assign n7483 = n7471 & n7482;
  assign n7484 = ~n7472 & ~n7483;
  assign n7485 = ~pi1159 & pi1160;
  assign n7486 = ~n7484 & n7485;
  assign n7487 = n7481 & ~n7486;
  assign n7488 = pi1159 & ~pi1160;
  assign n7489 = ~n7474 & n7488;
  assign n7490 = n7487 & ~n7489;
  assign n7491 = n7470 & ~n7490;
  assign po0398 = n7469 | n7491;
  assign n7493 = pi0348 & ~pi2253;
  assign n7494 = pi0875 & ~pi2253;
  assign n7495 = pi1036 & pi1149;
  assign n7496 = pi2055 & n7495;
  assign n7497 = ~pi2016 & n7495;
  assign n7498 = ~n7496 & ~n7497;
  assign n7499 = ~pi2135 & n7495;
  assign n7500 = n7498 & ~n7499;
  assign n7501 = ~pi1147 & ~pi1148;
  assign n7502 = ~n7500 & n7501;
  assign n7503 = pi1147 & pi1148;
  assign n7504 = n7496 & n7503;
  assign n7505 = ~n7502 & ~n7504;
  assign n7506 = ~pi2016 & ~pi2135;
  assign n7507 = n7495 & n7506;
  assign n7508 = ~n7496 & ~n7507;
  assign n7509 = ~pi1147 & pi1148;
  assign n7510 = ~n7508 & n7509;
  assign n7511 = n7505 & ~n7510;
  assign n7512 = pi1147 & ~pi1148;
  assign n7513 = ~n7498 & n7512;
  assign n7514 = n7511 & ~n7513;
  assign n7515 = n7494 & ~n7514;
  assign po0399 = n7493 | n7515;
  assign n7517 = n5215 & n7364;
  assign n7518 = pi1169 & n7517;
  assign n7519 = ~n7395 & n7518;
  assign n7520 = pi1169 & ~n5215;
  assign n7521 = ~pi0349 & n7520;
  assign po0400 = n7519 | n7521;
  assign n7523 = ~n7372 & n7518;
  assign n7524 = ~pi0350 & n7520;
  assign po0401 = n7523 | n7524;
  assign n7526 = n5196 & n7349;
  assign n7527 = pi1035 & n7526;
  assign n7528 = ~n7339 & n7527;
  assign n7529 = pi1035 & ~n5196;
  assign n7530 = ~pi0351 & n7529;
  assign po0402 = n7528 | n7530;
  assign n7532 = ~n7417 & n7527;
  assign n7533 = ~pi0352 & n7529;
  assign po0403 = n7532 | n7533;
  assign n7535 = pi0353 & ~n5203;
  assign n7536 = ~pi0353 & n5203;
  assign n7537 = ~n7535 & ~n7536;
  assign po0404 = pi1035 & ~n7537;
  assign n7539 = pi0354 & ~n5222;
  assign n7540 = ~pi0354 & n5222;
  assign n7541 = ~n7539 & ~n7540;
  assign po0405 = pi1169 & ~n7541;
  assign n7543 = ~pi0635 & n7453;
  assign n7544 = n7451 & ~n7543;
  assign n7545 = ~pi0355 & ~n7544;
  assign n7546 = ~pi0411 & ~pi0412;
  assign n7547 = pi0355 & ~n7546;
  assign n7548 = pi1138 & ~pi1152;
  assign n7549 = pi0197 & n7548;
  assign n7550 = pi1901 & n7453;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = n7546 & n7551;
  assign n7553 = ~n7547 & ~n7552;
  assign n7554 = n7544 & n7553;
  assign po0406 = n7545 | n7554;
  assign n7556 = ~pi0356 & ~n7544;
  assign n7557 = pi0356 & ~n7546;
  assign n7558 = pi0193 & n7548;
  assign n7559 = pi1875 & n7453;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = n7546 & n7560;
  assign n7562 = ~n7557 & ~n7561;
  assign n7563 = n7544 & n7562;
  assign po0407 = n7556 | n7563;
  assign n7565 = ~pi0357 & ~n7544;
  assign n7566 = pi0411 & ~pi0412;
  assign n7567 = pi0357 & ~n7566;
  assign n7568 = n7551 & n7566;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = n7544 & n7569;
  assign po0408 = n7565 | n7570;
  assign n7572 = ~pi0358 & ~n7544;
  assign n7573 = pi0358 & ~n7566;
  assign n7574 = n7560 & n7566;
  assign n7575 = ~n7573 & ~n7574;
  assign n7576 = n7544 & n7575;
  assign po0409 = n7572 | n7576;
  assign n7578 = ~pi0359 & ~n7544;
  assign n7579 = pi0359 & ~n7566;
  assign n7580 = pi0947 & n7453;
  assign n7581 = n7566 & ~n7580;
  assign n7582 = ~n7579 & ~n7581;
  assign n7583 = n7544 & n7582;
  assign po0410 = n7578 | n7583;
  assign n7585 = ~pi0360 & ~n7544;
  assign n7586 = pi0360 & ~n7566;
  assign n7587 = pi0923 & n7453;
  assign n7588 = n7566 & ~n7587;
  assign n7589 = ~n7586 & ~n7588;
  assign n7590 = n7544 & n7589;
  assign po0411 = n7585 | n7590;
  assign n7592 = ~pi0361 & ~n7544;
  assign n7593 = pi0361 & ~n7566;
  assign n7594 = pi0877 & n7453;
  assign n7595 = n7566 & ~n7594;
  assign n7596 = ~n7593 & ~n7595;
  assign n7597 = n7544 & n7596;
  assign po0412 = n7592 | n7597;
  assign n7599 = ~pi0362 & ~n7544;
  assign n7600 = pi0362 & ~n7566;
  assign n7601 = pi0871 & n7453;
  assign n7602 = n7566 & ~n7601;
  assign n7603 = ~n7600 & ~n7602;
  assign n7604 = n7544 & n7603;
  assign po0413 = n7599 | n7604;
  assign n7606 = ~pi0363 & ~n7544;
  assign n7607 = pi0363 & ~n7566;
  assign n7608 = pi0814 & n7453;
  assign n7609 = n7566 & ~n7608;
  assign n7610 = ~n7607 & ~n7609;
  assign n7611 = n7544 & n7610;
  assign po0414 = n7606 | n7611;
  assign n7613 = ~pi0364 & ~n7544;
  assign n7614 = pi0364 & ~n7566;
  assign n7615 = pi0480 & n7453;
  assign n7616 = n7566 & ~n7615;
  assign n7617 = ~n7614 & ~n7616;
  assign n7618 = n7544 & n7617;
  assign po0415 = n7613 | n7618;
  assign n7620 = ~pi0365 & ~n7544;
  assign n7621 = pi0365 & ~n7566;
  assign n7622 = pi0335 & n7453;
  assign n7623 = n7566 & ~n7622;
  assign n7624 = ~n7621 & ~n7623;
  assign n7625 = n7544 & n7624;
  assign po0416 = n7620 | n7625;
  assign n7627 = ~pi0366 & ~n7544;
  assign n7628 = pi0366 & ~n7566;
  assign n7629 = pi0233 & n7453;
  assign n7630 = n7566 & ~n7629;
  assign n7631 = ~n7628 & ~n7630;
  assign n7632 = n7544 & n7631;
  assign po0417 = n7627 | n7632;
  assign n7634 = ~pi0367 & ~n7544;
  assign n7635 = pi0367 & ~n7566;
  assign n7636 = pi0213 & n7453;
  assign n7637 = n7566 & ~n7636;
  assign n7638 = ~n7635 & ~n7637;
  assign n7639 = n7544 & n7638;
  assign po0418 = n7634 | n7639;
  assign n7641 = ~pi0368 & ~n7544;
  assign n7642 = pi0368 & ~n7566;
  assign n7643 = pi0208 & n7453;
  assign n7644 = n7566 & ~n7643;
  assign n7645 = ~n7642 & ~n7644;
  assign n7646 = n7544 & n7645;
  assign po0419 = n7641 | n7646;
  assign n7648 = ~pi0369 & ~n7544;
  assign n7649 = pi0369 & ~n7566;
  assign n7650 = pi0197 & n7453;
  assign n7651 = n7566 & ~n7650;
  assign n7652 = ~n7649 & ~n7651;
  assign n7653 = n7544 & n7652;
  assign po0420 = n7648 | n7653;
  assign n7655 = ~pi0370 & ~n7544;
  assign n7656 = pi0370 & ~n7566;
  assign n7657 = pi0193 & n7453;
  assign n7658 = n7566 & ~n7657;
  assign n7659 = ~n7656 & ~n7658;
  assign n7660 = n7544 & n7659;
  assign po0421 = n7655 | n7660;
  assign n7662 = ~pi0371 & ~n7544;
  assign n7663 = ~pi0411 & pi0412;
  assign n7664 = pi0371 & ~n7663;
  assign n7665 = n7551 & n7663;
  assign n7666 = ~n7664 & ~n7665;
  assign n7667 = n7544 & n7666;
  assign po0422 = n7662 | n7667;
  assign n7669 = ~pi0372 & ~n7544;
  assign n7670 = pi0372 & ~n7663;
  assign n7671 = n7560 & n7663;
  assign n7672 = ~n7670 & ~n7671;
  assign n7673 = n7544 & n7672;
  assign po0423 = n7669 | n7673;
  assign n7675 = ~pi0373 & ~n7544;
  assign n7676 = pi0373 & ~n7663;
  assign n7677 = ~n7580 & n7663;
  assign n7678 = ~n7676 & ~n7677;
  assign n7679 = n7544 & n7678;
  assign po0424 = n7675 | n7679;
  assign n7681 = ~pi0374 & ~n7544;
  assign n7682 = pi0374 & ~n7663;
  assign n7683 = ~n7587 & n7663;
  assign n7684 = ~n7682 & ~n7683;
  assign n7685 = n7544 & n7684;
  assign po0425 = n7681 | n7685;
  assign n7687 = ~pi0375 & ~n7544;
  assign n7688 = pi0375 & ~n7663;
  assign n7689 = ~n7594 & n7663;
  assign n7690 = ~n7688 & ~n7689;
  assign n7691 = n7544 & n7690;
  assign po0426 = n7687 | n7691;
  assign n7693 = ~pi0376 & ~n7544;
  assign n7694 = pi0376 & ~n7663;
  assign n7695 = ~n7601 & n7663;
  assign n7696 = ~n7694 & ~n7695;
  assign n7697 = n7544 & n7696;
  assign po0427 = n7693 | n7697;
  assign n7699 = ~pi0377 & ~n7544;
  assign n7700 = pi0377 & ~n7663;
  assign n7701 = ~n7608 & n7663;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = n7544 & n7702;
  assign po0428 = n7699 | n7703;
  assign n7705 = ~pi0378 & ~n7544;
  assign n7706 = pi0378 & ~n7663;
  assign n7707 = ~n7615 & n7663;
  assign n7708 = ~n7706 & ~n7707;
  assign n7709 = n7544 & n7708;
  assign po0429 = n7705 | n7709;
  assign n7711 = ~pi0379 & ~n7544;
  assign n7712 = pi0379 & ~n7663;
  assign n7713 = ~n7622 & n7663;
  assign n7714 = ~n7712 & ~n7713;
  assign n7715 = n7544 & n7714;
  assign po0430 = n7711 | n7715;
  assign n7717 = ~pi0380 & ~n7544;
  assign n7718 = pi0380 & ~n7663;
  assign n7719 = ~n7629 & n7663;
  assign n7720 = ~n7718 & ~n7719;
  assign n7721 = n7544 & n7720;
  assign po0431 = n7717 | n7721;
  assign n7723 = ~pi0381 & ~n7544;
  assign n7724 = pi0381 & ~n7663;
  assign n7725 = ~n7636 & n7663;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = n7544 & n7726;
  assign po0432 = n7723 | n7727;
  assign n7729 = ~pi0382 & ~n7544;
  assign n7730 = pi0382 & ~n7663;
  assign n7731 = ~n7643 & n7663;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 = n7544 & n7732;
  assign po0433 = n7729 | n7733;
  assign n7735 = ~pi0383 & ~n7544;
  assign n7736 = pi0383 & ~n7663;
  assign n7737 = ~n7650 & n7663;
  assign n7738 = ~n7736 & ~n7737;
  assign n7739 = n7544 & n7738;
  assign po0434 = n7735 | n7739;
  assign n7741 = ~pi0384 & ~n7544;
  assign n7742 = pi0384 & ~n7663;
  assign n7743 = ~n7657 & n7663;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = n7544 & n7744;
  assign po0435 = n7741 | n7745;
  assign n7747 = ~pi0385 & ~n7544;
  assign n7748 = n7454 & ~n7551;
  assign n7749 = ~pi0385 & ~n7454;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = n7544 & ~n7750;
  assign po0436 = n7747 | n7751;
  assign n7753 = ~pi0386 & ~n7544;
  assign n7754 = n7454 & ~n7560;
  assign n7755 = ~pi0386 & ~n7454;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = n7544 & ~n7756;
  assign po0437 = n7753 | n7757;
  assign n7759 = ~pi0387 & ~n7544;
  assign n7760 = n7454 & n7580;
  assign n7761 = ~pi0387 & ~n7454;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = n7544 & ~n7762;
  assign po0438 = n7759 | n7763;
  assign n7765 = ~pi0388 & ~n7544;
  assign n7766 = n7454 & n7587;
  assign n7767 = ~pi0388 & ~n7454;
  assign n7768 = ~n7766 & ~n7767;
  assign n7769 = n7544 & ~n7768;
  assign po0439 = n7765 | n7769;
  assign n7771 = ~pi0389 & ~n7544;
  assign n7772 = n7454 & n7594;
  assign n7773 = ~pi0389 & ~n7454;
  assign n7774 = ~n7772 & ~n7773;
  assign n7775 = n7544 & ~n7774;
  assign po0440 = n7771 | n7775;
  assign n7777 = ~pi0390 & ~n7544;
  assign n7778 = n7454 & n7601;
  assign n7779 = ~pi0390 & ~n7454;
  assign n7780 = ~n7778 & ~n7779;
  assign n7781 = n7544 & ~n7780;
  assign po0441 = n7777 | n7781;
  assign n7783 = ~pi0391 & ~n7544;
  assign n7784 = n7454 & n7608;
  assign n7785 = ~pi0391 & ~n7454;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = n7544 & ~n7786;
  assign po0442 = n7783 | n7787;
  assign n7789 = ~pi0392 & ~n7544;
  assign n7790 = n7454 & n7615;
  assign n7791 = ~pi0392 & ~n7454;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = n7544 & ~n7792;
  assign po0443 = n7789 | n7793;
  assign n7795 = ~pi0393 & ~n7544;
  assign n7796 = n7454 & n7622;
  assign n7797 = ~pi0393 & ~n7454;
  assign n7798 = ~n7796 & ~n7797;
  assign n7799 = n7544 & ~n7798;
  assign po0444 = n7795 | n7799;
  assign n7801 = ~pi0394 & ~n7544;
  assign n7802 = n7454 & n7629;
  assign n7803 = ~pi0394 & ~n7454;
  assign n7804 = ~n7802 & ~n7803;
  assign n7805 = n7544 & ~n7804;
  assign po0445 = n7801 | n7805;
  assign n7807 = ~pi0395 & ~n7544;
  assign n7808 = n7454 & n7636;
  assign n7809 = ~pi0395 & ~n7454;
  assign n7810 = ~n7808 & ~n7809;
  assign n7811 = n7544 & ~n7810;
  assign po0446 = n7807 | n7811;
  assign n7813 = ~pi0396 & ~n7544;
  assign n7814 = n7454 & n7643;
  assign n7815 = ~pi0396 & ~n7454;
  assign n7816 = ~n7814 & ~n7815;
  assign n7817 = n7544 & ~n7816;
  assign po0447 = n7813 | n7817;
  assign n7819 = ~pi0397 & ~n7544;
  assign n7820 = n7454 & n7650;
  assign n7821 = ~pi0397 & ~n7454;
  assign n7822 = ~n7820 & ~n7821;
  assign n7823 = n7544 & ~n7822;
  assign po0448 = n7819 | n7823;
  assign n7825 = ~pi0398 & ~n7544;
  assign n7826 = n7454 & n7657;
  assign n7827 = ~pi0398 & ~n7454;
  assign n7828 = ~n7826 & ~n7827;
  assign n7829 = n7544 & ~n7828;
  assign po0449 = n7825 | n7829;
  assign n7831 = pi0803 & n7453;
  assign n7832 = ~pi1138 & pi1152;
  assign n7833 = pi0923 & n7832;
  assign n7834 = ~n7831 & ~n7833;
  assign n7835 = pi1875 & n7548;
  assign n7836 = n7834 & ~n7835;
  assign n7837 = n7454 & ~n7836;
  assign n7838 = ~pi0399 & ~n7454;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = n7544 & ~n7839;
  assign n7841 = ~pi0399 & ~n7544;
  assign po0450 = n7840 | n7841;
  assign n7843 = ~pi0400 & ~n7566;
  assign n7844 = pi0794 & n7453;
  assign n7845 = pi0335 & n7832;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = pi0814 & n7548;
  assign n7848 = n7846 & ~n7847;
  assign n7849 = n7566 & ~n7848;
  assign n7850 = ~n7843 & ~n7849;
  assign n7851 = n7544 & ~n7850;
  assign n7852 = ~pi0400 & ~n7544;
  assign po0451 = n7851 | n7852;
  assign n7854 = ~pi0401 & ~n7566;
  assign n7855 = pi0795 & n7453;
  assign n7856 = pi0233 & n7832;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = pi0480 & n7548;
  assign n7859 = n7857 & ~n7858;
  assign n7860 = n7566 & ~n7859;
  assign n7861 = ~n7854 & ~n7860;
  assign n7862 = n7544 & ~n7861;
  assign n7863 = ~pi0401 & ~n7544;
  assign po0452 = n7862 | n7863;
  assign n7865 = ~pi0402 & ~n7566;
  assign n7866 = pi0197 & n7832;
  assign n7867 = pi0213 & n7548;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = pi1935 & n7453;
  assign n7870 = n7868 & ~n7869;
  assign n7871 = n7566 & ~n7870;
  assign n7872 = ~n7865 & ~n7871;
  assign n7873 = n7544 & ~n7872;
  assign n7874 = ~pi0402 & ~n7544;
  assign po0453 = n7873 | n7874;
  assign n7876 = ~pi0403 & ~n7663;
  assign n7877 = pi0193 & n7832;
  assign n7878 = pi0208 & n7548;
  assign n7879 = ~n7877 & ~n7878;
  assign n7880 = pi1926 & n7453;
  assign n7881 = n7879 & ~n7880;
  assign n7882 = n7663 & ~n7881;
  assign n7883 = ~n7876 & ~n7882;
  assign n7884 = n7544 & ~n7883;
  assign n7885 = ~pi0403 & ~n7544;
  assign po0454 = n7884 | n7885;
  assign n7887 = ~pi0404 & ~n7663;
  assign n7888 = pi0798 & n7453;
  assign n7889 = pi1978 & n7832;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = pi1961 & n7548;
  assign n7892 = n7890 & ~n7891;
  assign n7893 = n7663 & ~n7892;
  assign n7894 = ~n7887 & ~n7893;
  assign n7895 = n7544 & ~n7894;
  assign n7896 = ~pi0404 & ~n7544;
  assign po0455 = n7895 | n7896;
  assign n7898 = ~pi0405 & ~n7663;
  assign n7899 = n7663 & ~n7836;
  assign n7900 = ~n7898 & ~n7899;
  assign n7901 = n7544 & ~n7900;
  assign n7902 = ~pi0405 & ~n7544;
  assign po0456 = n7901 | n7902;
  assign n7904 = ~pi0406 & ~n7663;
  assign n7905 = pi0657 & n7453;
  assign n7906 = pi0877 & n7832;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = pi0947 & n7548;
  assign n7909 = n7907 & ~n7908;
  assign n7910 = n7663 & ~n7909;
  assign n7911 = ~n7904 & ~n7910;
  assign n7912 = n7544 & ~n7911;
  assign n7913 = ~pi0406 & ~n7544;
  assign po0457 = n7912 | n7913;
  assign n7915 = n7454 & ~n7870;
  assign n7916 = ~pi0407 & ~n7454;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = n7544 & ~n7917;
  assign n7919 = ~pi0407 & ~n7544;
  assign po0458 = n7918 | n7919;
  assign n7921 = n7454 & ~n7881;
  assign n7922 = ~pi0408 & ~n7454;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = n7544 & ~n7923;
  assign n7925 = ~pi0408 & ~n7544;
  assign po0459 = n7924 | n7925;
  assign n7927 = pi0801 & n7453;
  assign n7928 = pi1875 & n7832;
  assign n7929 = ~n7927 & ~n7928;
  assign n7930 = pi1926 & n7548;
  assign n7931 = n7929 & ~n7930;
  assign n7932 = n7454 & ~n7931;
  assign n7933 = ~pi0409 & ~n7454;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = n7544 & ~n7934;
  assign n7936 = ~pi0409 & ~n7544;
  assign po0460 = n7935 | n7936;
  assign n7938 = pi0802 & n7453;
  assign n7939 = pi0947 & n7832;
  assign n7940 = ~n7938 & ~n7939;
  assign n7941 = pi1901 & n7548;
  assign n7942 = n7940 & ~n7941;
  assign n7943 = n7454 & ~n7942;
  assign n7944 = ~pi0410 & ~n7454;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = n7544 & ~n7945;
  assign n7947 = ~pi0410 & ~n7544;
  assign po0461 = n7946 | n7947;
  assign n7949 = pi0411 & ~n7451;
  assign n7950 = ~pi0411 & pi0635;
  assign n7951 = pi0411 & ~pi0635;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = n7453 & ~n7952;
  assign n7954 = ~pi0411 & ~n7453;
  assign n7955 = ~n7953 & ~n7954;
  assign n7956 = n7451 & ~n7955;
  assign n7957 = ~n7949 & ~n7956;
  assign po0462 = pi1150 & ~n7957;
  assign n7959 = pi0412 & ~n7451;
  assign n7960 = ~n7566 & ~n7663;
  assign n7961 = ~n7453 & ~n7960;
  assign n7962 = ~pi0412 & n7459;
  assign n7963 = pi0412 & ~n7459;
  assign n7964 = ~n7962 & ~n7963;
  assign n7965 = n7453 & ~n7964;
  assign n7966 = ~n7961 & ~n7965;
  assign n7967 = n7451 & ~n7966;
  assign n7968 = ~n7959 & ~n7967;
  assign po0463 = pi1150 & ~n7968;
  assign n7970 = pi1382 & n5455;
  assign n7971 = pi1357 & n5200;
  assign n7972 = pi1792 & n7335;
  assign n7973 = pi1332 & n5199;
  assign n7974 = ~n7972 & ~n7973;
  assign n7975 = ~n7971 & n7974;
  assign n7976 = ~n7970 & n7975;
  assign n7977 = ~pi0353 & ~n7976;
  assign n7978 = pi1372 & n5455;
  assign n7979 = pi1347 & n5200;
  assign n7980 = ~n7978 & ~n7979;
  assign n7981 = pi1322 & n5199;
  assign n7982 = pi0956 & n7335;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = n7980 & n7983;
  assign n7985 = pi0353 & ~n7984;
  assign n7986 = ~n7977 & ~n7985;
  assign n7987 = n5197 & ~n7986;
  assign n7988 = pi1361 & n5455;
  assign n7989 = pi1336 & n5200;
  assign n7990 = pi1669 & n7335;
  assign n7991 = pi1311 & n5199;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = ~n7989 & n7992;
  assign n7994 = ~n7988 & n7993;
  assign n7995 = n7349 & ~n7994;
  assign n7996 = pi1384 & n5455;
  assign n7997 = pi1359 & n5200;
  assign n7998 = pi1683 & n7335;
  assign n7999 = pi1334 & n5199;
  assign n8000 = ~n7998 & ~n7999;
  assign n8001 = ~n7997 & n8000;
  assign n8002 = ~n7996 & n8001;
  assign n8003 = n7340 & ~n8002;
  assign n8004 = ~n7995 & ~n8003;
  assign n8005 = ~n7987 & n8004;
  assign n8006 = n5196 & ~n8005;
  assign n8007 = ~pi0413 & ~n5196;
  assign n8008 = ~n8006 & ~n8007;
  assign po0464 = pi1035 & ~n8008;
  assign n8010 = pi1027 & n5455;
  assign n8011 = pi1039 & n5200;
  assign n8012 = pi0961 & n7335;
  assign n8013 = pi1054 & n5199;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = ~n8011 & n8014;
  assign n8016 = ~n8010 & n8015;
  assign n8017 = ~pi0353 & ~n8016;
  assign n8018 = pi1374 & n5455;
  assign n8019 = pi1349 & n5200;
  assign n8020 = ~n8018 & ~n8019;
  assign n8021 = pi1324 & n5199;
  assign n8022 = pi1675 & n7335;
  assign n8023 = ~n8021 & ~n8022;
  assign n8024 = n8020 & n8023;
  assign n8025 = pi0353 & ~n8024;
  assign n8026 = ~n8017 & ~n8025;
  assign n8027 = n5197 & ~n8026;
  assign n8028 = pi1363 & n5455;
  assign n8029 = pi1338 & n5200;
  assign n8030 = pi0952 & n7335;
  assign n8031 = pi1313 & n5199;
  assign n8032 = ~n8030 & ~n8031;
  assign n8033 = ~n8029 & n8032;
  assign n8034 = ~n8028 & n8033;
  assign n8035 = n7349 & ~n8034;
  assign n8036 = pi1312 & n5199;
  assign n8037 = pi1337 & n5200;
  assign n8038 = pi1670 & n7335;
  assign n8039 = pi1362 & n5455;
  assign n8040 = ~n8038 & ~n8039;
  assign n8041 = ~n8037 & n8040;
  assign n8042 = ~n8036 & n8041;
  assign n8043 = n7340 & ~n8042;
  assign n8044 = ~n8035 & ~n8043;
  assign n8045 = ~n8027 & n8044;
  assign n8046 = n5196 & ~n8045;
  assign n8047 = ~pi0414 & ~n5196;
  assign n8048 = ~n8046 & ~n8047;
  assign po0465 = pi1035 & ~n8048;
  assign n8050 = ~pi0353 & ~n7994;
  assign n8051 = pi1375 & n5455;
  assign n8052 = pi1350 & n5200;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = pi1325 & n5199;
  assign n8055 = pi1678 & n7335;
  assign n8056 = ~n8054 & ~n8055;
  assign n8057 = n8053 & n8056;
  assign n8058 = pi0353 & ~n8057;
  assign n8059 = ~n8050 & ~n8058;
  assign n8060 = n5197 & ~n8059;
  assign n8061 = pi1314 & n5199;
  assign n8062 = pi1339 & n5200;
  assign n8063 = pi0953 & n7335;
  assign n8064 = pi1364 & n5455;
  assign n8065 = ~n8063 & ~n8064;
  assign n8066 = ~n8062 & n8065;
  assign n8067 = ~n8061 & n8066;
  assign n8068 = n7349 & ~n8067;
  assign n8069 = pi1041 & n5455;
  assign n8070 = pi1052 & n5200;
  assign n8071 = pi1818 & n7335;
  assign n8072 = pi1065 & n5199;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = ~n8070 & n8073;
  assign n8075 = ~n8069 & n8074;
  assign n8076 = n7340 & ~n8075;
  assign n8077 = ~n8068 & ~n8076;
  assign n8078 = ~n8060 & n8077;
  assign n8079 = n5196 & ~n8078;
  assign n8080 = ~pi0415 & ~n5196;
  assign n8081 = ~n8079 & ~n8080;
  assign po0466 = pi1035 & ~n8081;
  assign n8083 = ~pi0353 & ~n8042;
  assign n8084 = pi1056 & n5199;
  assign n8085 = pi1676 & n7335;
  assign n8086 = ~n8084 & ~n8085;
  assign n8087 = pi1033 & n5455;
  assign n8088 = pi1045 & n5200;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = n8086 & n8089;
  assign n8091 = pi0353 & ~n8090;
  assign n8092 = ~n8083 & ~n8091;
  assign n8093 = n5197 & ~n8092;
  assign n8094 = pi1365 & n5455;
  assign n8095 = pi1315 & n5199;
  assign n8096 = ~n8094 & ~n8095;
  assign n8097 = pi1340 & n5200;
  assign n8098 = pi1671 & n7335;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = n8096 & n8099;
  assign n8101 = n7349 & ~n8100;
  assign n8102 = n7340 & ~n8034;
  assign n8103 = ~n8101 & ~n8102;
  assign n8104 = ~n8093 & n8103;
  assign n8105 = n5196 & ~n8104;
  assign n8106 = ~pi0416 & ~n5196;
  assign n8107 = ~n8105 & ~n8106;
  assign po0467 = pi1035 & ~n8107;
  assign n8109 = ~pi0353 & ~n8075;
  assign n8110 = pi1326 & n5199;
  assign n8111 = pi1677 & n7335;
  assign n8112 = ~n8110 & ~n8111;
  assign n8113 = pi1376 & n5455;
  assign n8114 = pi1351 & n5200;
  assign n8115 = ~n8113 & ~n8114;
  assign n8116 = n8112 & n8115;
  assign n8117 = pi0353 & ~n8116;
  assign n8118 = ~n8109 & ~n8117;
  assign n8119 = n5197 & ~n8118;
  assign n8120 = n7349 & ~n7431;
  assign n8121 = n7340 & ~n8067;
  assign n8122 = ~n8120 & ~n8121;
  assign n8123 = ~n8119 & n8122;
  assign n8124 = n5196 & ~n8123;
  assign n8125 = ~pi0417 & ~n5196;
  assign n8126 = ~n8124 & ~n8125;
  assign po0468 = pi1035 & ~n8126;
  assign n8128 = pi1383 & n5455;
  assign n8129 = pi1333 & n5199;
  assign n8130 = pi1358 & n5200;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = pi0960 & n7335;
  assign n8133 = n8131 & ~n8132;
  assign n8134 = ~n8128 & n8133;
  assign n8135 = ~pi0353 & ~n8134;
  assign n8136 = pi1032 & n5455;
  assign n8137 = pi1046 & n5200;
  assign n8138 = ~n8136 & ~n8137;
  assign n8139 = pi1060 & n5199;
  assign n8140 = pi1806 & n7335;
  assign n8141 = ~n8139 & ~n8140;
  assign n8142 = n8138 & n8141;
  assign n8143 = pi0353 & ~n8142;
  assign n8144 = ~n8135 & ~n8143;
  assign n8145 = n5197 & ~n8144;
  assign n8146 = n7349 & ~n8042;
  assign n8147 = n7340 & ~n8016;
  assign n8148 = ~n8146 & ~n8147;
  assign n8149 = ~n8145 & n8148;
  assign n8150 = n5196 & ~n8149;
  assign n8151 = ~pi0418 & ~n5196;
  assign n8152 = ~n8150 & ~n8151;
  assign po0469 = pi1035 & ~n8152;
  assign n8154 = ~pi0353 & ~n8067;
  assign n8155 = pi1029 & n5455;
  assign n8156 = pi1044 & n5200;
  assign n8157 = ~n8155 & ~n8156;
  assign n8158 = pi1053 & n5199;
  assign n8159 = pi1799 & n7335;
  assign n8160 = ~n8158 & ~n8159;
  assign n8161 = n8157 & n8160;
  assign n8162 = pi0353 & ~n8161;
  assign n8163 = ~n8154 & ~n8162;
  assign n8164 = n5197 & ~n8163;
  assign n8165 = pi1367 & n5455;
  assign n8166 = pi1342 & n5200;
  assign n8167 = pi1317 & n5199;
  assign n8168 = pi1672 & n7335;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = ~n8166 & n8169;
  assign n8171 = ~n8165 & n8170;
  assign n8172 = n7349 & ~n8171;
  assign n8173 = n7340 & ~n7431;
  assign n8174 = ~n8172 & ~n8173;
  assign n8175 = ~n8164 & n8174;
  assign n8176 = n5196 & ~n8175;
  assign n8177 = ~pi0419 & ~n5196;
  assign n8178 = ~n8176 & ~n8177;
  assign po0470 = pi1035 & ~n8178;
  assign n8180 = ~pi0353 & ~n8002;
  assign n8181 = pi1373 & n5455;
  assign n8182 = pi1348 & n5200;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = pi1323 & n5199;
  assign n8185 = pi0957 & n7335;
  assign n8186 = ~n8184 & ~n8185;
  assign n8187 = n8183 & n8186;
  assign n8188 = pi0353 & ~n8187;
  assign n8189 = ~n8180 & ~n8188;
  assign n8190 = n5197 & ~n8189;
  assign n8191 = n7349 & ~n8075;
  assign n8192 = n7340 & ~n7994;
  assign n8193 = ~n8191 & ~n8192;
  assign n8194 = ~n8190 & n8193;
  assign n8195 = n5196 & ~n8194;
  assign n8196 = ~pi0420 & ~n5196;
  assign n8197 = ~n8195 & ~n8196;
  assign po0471 = pi1035 & ~n8197;
  assign n8199 = ~pi0353 & ~n8100;
  assign n8200 = pi1379 & n5455;
  assign n8201 = pi1354 & n5200;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = pi1329 & n5199;
  assign n8204 = pi0958 & n7335;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = n8202 & n8205;
  assign n8207 = pi0353 & ~n8206;
  assign n8208 = ~n8199 & ~n8207;
  assign n8209 = n5197 & ~n8208;
  assign n8210 = pi1368 & n5455;
  assign n8211 = pi1343 & n5200;
  assign n8212 = pi1318 & n5199;
  assign n8213 = pi0955 & n7335;
  assign n8214 = ~n8212 & ~n8213;
  assign n8215 = ~n8211 & n8214;
  assign n8216 = ~n8210 & n8215;
  assign n8217 = n7349 & ~n8216;
  assign n8218 = pi1366 & n5455;
  assign n8219 = pi1341 & n5200;
  assign n8220 = pi1316 & n5199;
  assign n8221 = pi1808 & n7335;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = ~n8219 & n8222;
  assign n8224 = ~n8218 & n8223;
  assign n8225 = n7340 & ~n8224;
  assign n8226 = ~n8217 & ~n8225;
  assign n8227 = ~n8209 & n8226;
  assign n8228 = n5196 & ~n8227;
  assign n8229 = ~pi0421 & ~n5196;
  assign n8230 = ~n8228 & ~n8229;
  assign po0472 = pi1035 & ~n8230;
  assign n8232 = ~pi0353 & ~n8034;
  assign n8233 = pi1377 & n5455;
  assign n8234 = pi1352 & n5200;
  assign n8235 = ~n8233 & ~n8234;
  assign n8236 = pi1327 & n5199;
  assign n8237 = pi1680 & n7335;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = n8235 & n8238;
  assign n8240 = pi0353 & ~n8239;
  assign n8241 = ~n8232 & ~n8240;
  assign n8242 = n5197 & ~n8241;
  assign n8243 = n7349 & ~n8224;
  assign n8244 = n7340 & ~n8100;
  assign n8245 = ~n8243 & ~n8244;
  assign n8246 = ~n8242 & n8245;
  assign n8247 = n5196 & ~n8246;
  assign n8248 = ~pi0422 & ~n5196;
  assign n8249 = ~n8247 & ~n8248;
  assign po0473 = pi1035 & ~n8249;
  assign n8251 = pi0353 & ~n8224;
  assign n8252 = ~pi0353 & ~n7339;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = n5197 & ~n8253;
  assign n8255 = pi1028 & n5455;
  assign n8256 = pi1042 & n5200;
  assign n8257 = pi1682 & n7335;
  assign n8258 = pi1055 & n5199;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = ~n8256 & n8259;
  assign n8261 = ~n8255 & n8260;
  assign n8262 = n7349 & ~n8261;
  assign n8263 = n7340 & ~n7348;
  assign n8264 = ~n8262 & ~n8263;
  assign n8265 = ~n8254 & n8264;
  assign n8266 = n5196 & ~n8265;
  assign n8267 = ~pi0423 & ~n5196;
  assign n8268 = ~n8266 & ~n8267;
  assign po0474 = pi1035 & ~n8268;
  assign n8270 = ~pi0353 & ~n7409;
  assign n8271 = pi0353 & ~n8171;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = n5197 & ~n8272;
  assign n8274 = n7349 & ~n7976;
  assign n8275 = n7340 & ~n7441;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n8273 & n8276;
  assign n8278 = n5196 & ~n8277;
  assign n8279 = ~pi0424 & ~n5196;
  assign n8280 = ~n8278 & ~n8279;
  assign po0475 = pi1035 & ~n8280;
  assign n8282 = ~pi0353 & ~n7348;
  assign n8283 = pi0353 & ~n8216;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = n5197 & ~n8284;
  assign n8286 = n7349 & ~n8134;
  assign n8287 = n7340 & ~n8261;
  assign n8288 = ~n8286 & ~n8287;
  assign n8289 = ~n8285 & n8288;
  assign n8290 = n5196 & ~n8289;
  assign n8291 = ~pi0425 & ~n5196;
  assign n8292 = ~n8290 & ~n8291;
  assign po0476 = pi1035 & ~n8292;
  assign n8294 = ~pi0353 & ~n7441;
  assign n8295 = pi1370 & n5455;
  assign n8296 = pi1345 & n5200;
  assign n8297 = ~n8295 & ~n8296;
  assign n8298 = pi1320 & n5199;
  assign n8299 = pi1815 & n7335;
  assign n8300 = ~n8298 & ~n8299;
  assign n8301 = n8297 & n8300;
  assign n8302 = pi0353 & ~n8301;
  assign n8303 = ~n8294 & ~n8302;
  assign n8304 = n5197 & ~n8303;
  assign n8305 = n7349 & ~n8002;
  assign n8306 = n7340 & ~n7976;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = ~n8304 & n8307;
  assign n8309 = n5196 & ~n8308;
  assign n8310 = ~pi0426 & ~n5196;
  assign n8311 = ~n8309 & ~n8310;
  assign po0477 = pi1035 & ~n8311;
  assign n8313 = ~pi0353 & ~n8261;
  assign n8314 = pi1371 & n5455;
  assign n8315 = pi1346 & n5200;
  assign n8316 = ~n8314 & ~n8315;
  assign n8317 = pi1321 & n5199;
  assign n8318 = pi1674 & n7335;
  assign n8319 = ~n8317 & ~n8318;
  assign n8320 = n8316 & n8319;
  assign n8321 = pi0353 & ~n8320;
  assign n8322 = ~n8313 & ~n8321;
  assign n8323 = n5197 & ~n8322;
  assign n8324 = n7349 & ~n8016;
  assign n8325 = n7340 & ~n8134;
  assign n8326 = ~n8324 & ~n8325;
  assign n8327 = ~n8323 & n8326;
  assign n8328 = n5196 & ~n8327;
  assign n8329 = ~pi0427 & ~n5196;
  assign n8330 = ~n8328 & ~n8329;
  assign po0478 = pi1035 & ~n8330;
  assign n8332 = ~pi0428 & ~n5215;
  assign n8333 = pi1458 & n5481;
  assign n8334 = pi1766 & n7359;
  assign n8335 = pi1408 & n5218;
  assign n8336 = pi1433 & n5219;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = ~n8334 & n8337;
  assign n8339 = ~n8333 & n8338;
  assign n8340 = ~pi0354 & ~n8339;
  assign n8341 = pi1812 & n5481;
  assign n8342 = pi1826 & n5219;
  assign n8343 = ~n8341 & ~n8342;
  assign n8344 = pi1021 & n5218;
  assign n8345 = pi0966 & n7359;
  assign n8346 = ~n8344 & ~n8345;
  assign n8347 = n8343 & n8346;
  assign n8348 = pi0354 & ~n8347;
  assign n8349 = ~n8340 & ~n8348;
  assign n8350 = n5216 & ~n8349;
  assign n8351 = pi1437 & n5481;
  assign n8352 = pi1412 & n5219;
  assign n8353 = pi1387 & n5218;
  assign n8354 = pi1684 & n7359;
  assign n8355 = ~n8353 & ~n8354;
  assign n8356 = ~n8352 & n8355;
  assign n8357 = ~n8351 & n8356;
  assign n8358 = n7364 & ~n8357;
  assign n8359 = pi1801 & n5481;
  assign n8360 = pi1805 & n5219;
  assign n8361 = pi1829 & n5218;
  assign n8362 = pi1698 & n7359;
  assign n8363 = ~n8361 & ~n8362;
  assign n8364 = ~n8360 & n8363;
  assign n8365 = ~n8359 & n8364;
  assign n8366 = n7373 & ~n8365;
  assign n8367 = ~n8358 & ~n8366;
  assign n8368 = ~n8350 & n8367;
  assign n8369 = n5215 & ~n8368;
  assign n8370 = ~n8332 & ~n8369;
  assign po0479 = pi1169 & ~n8370;
  assign n8372 = ~pi0429 & ~n5215;
  assign n8373 = pi1459 & n5481;
  assign n8374 = pi0970 & n7359;
  assign n8375 = pi1434 & n5219;
  assign n8376 = pi1409 & n5218;
  assign n8377 = ~n8375 & ~n8376;
  assign n8378 = ~n8374 & n8377;
  assign n8379 = ~n8373 & n8378;
  assign n8380 = ~pi0354 & ~n8379;
  assign n8381 = pi1448 & n5481;
  assign n8382 = pi1422 & n5219;
  assign n8383 = ~n8381 & ~n8382;
  assign n8384 = pi1398 & n5218;
  assign n8385 = pi1770 & n7359;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = n8383 & n8386;
  assign n8388 = pi0354 & ~n8387;
  assign n8389 = ~n8380 & ~n8388;
  assign n8390 = n5216 & ~n8389;
  assign n8391 = pi1816 & n5481;
  assign n8392 = pi1823 & n5219;
  assign n8393 = pi1024 & n5218;
  assign n8394 = pi1685 & n7359;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = ~n8392 & n8395;
  assign n8397 = ~n8391 & n8396;
  assign n8398 = n7364 & ~n8397;
  assign n8399 = pi1460 & n5481;
  assign n8400 = pi1410 & n5218;
  assign n8401 = pi1435 & n5219;
  assign n8402 = pi0971 & n7359;
  assign n8403 = ~n8401 & ~n8402;
  assign n8404 = ~n8400 & n8403;
  assign n8405 = ~n8399 & n8404;
  assign n8406 = n7373 & ~n8405;
  assign n8407 = ~n8398 & ~n8406;
  assign n8408 = ~n8390 & n8407;
  assign n8409 = n5215 & ~n8408;
  assign n8410 = ~n8372 & ~n8409;
  assign po0480 = pi1169 & ~n8410;
  assign n8412 = ~pi0430 & ~n5215;
  assign n8413 = ~pi0354 & ~n8365;
  assign n8414 = pi1449 & n5481;
  assign n8415 = pi1423 & n5219;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = pi1399 & n5218;
  assign n8418 = pi0967 & n7359;
  assign n8419 = ~n8417 & ~n8418;
  assign n8420 = n8416 & n8419;
  assign n8421 = pi0354 & ~n8420;
  assign n8422 = ~n8413 & ~n8421;
  assign n8423 = n5216 & ~n8422;
  assign n8424 = pi1438 & n5481;
  assign n8425 = pi1388 & n5218;
  assign n8426 = pi1790 & n7359;
  assign n8427 = pi1413 & n5219;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = ~n8425 & n8428;
  assign n8430 = ~n8424 & n8429;
  assign n8431 = n7364 & ~n8430;
  assign n8432 = n7373 & ~n8357;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = ~n8423 & n8433;
  assign n8435 = n5215 & ~n8434;
  assign n8436 = ~n8412 & ~n8435;
  assign po0481 = pi1169 & ~n8436;
  assign n8438 = ~pi0431 & ~n5215;
  assign n8439 = ~pi0354 & ~n8357;
  assign n8440 = pi1810 & n5481;
  assign n8441 = pi1819 & n5219;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = pi1019 & n5218;
  assign n8444 = pi1691 & n7359;
  assign n8445 = ~n8443 & ~n8444;
  assign n8446 = n8442 & n8445;
  assign n8447 = pi0354 & ~n8446;
  assign n8448 = ~n8439 & ~n8447;
  assign n8449 = n5216 & ~n8448;
  assign n8450 = n7373 & ~n8430;
  assign n8451 = pi1440 & n5481;
  assign n8452 = pi0963 & n7359;
  assign n8453 = pi1390 & n5218;
  assign n8454 = pi1415 & n5219;
  assign n8455 = ~n8453 & ~n8454;
  assign n8456 = ~n8452 & n8455;
  assign n8457 = ~n8451 & n8456;
  assign n8458 = n7364 & ~n8457;
  assign n8459 = ~n8450 & ~n8458;
  assign n8460 = ~n8449 & n8459;
  assign n8461 = n5215 & ~n8460;
  assign n8462 = ~n8438 & ~n8461;
  assign po0482 = pi1169 & ~n8462;
  assign n8464 = ~pi0432 & ~n5215;
  assign n8465 = ~pi0354 & ~n8397;
  assign n8466 = pi1451 & n5481;
  assign n8467 = pi1425 & n5219;
  assign n8468 = ~n8466 & ~n8467;
  assign n8469 = pi1401 & n5218;
  assign n8470 = pi1692 & n7359;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = n8468 & n8471;
  assign n8473 = pi0354 & ~n8472;
  assign n8474 = ~n8465 & ~n8473;
  assign n8475 = n5216 & ~n8474;
  assign n8476 = pi1439 & n5481;
  assign n8477 = pi1389 & n5218;
  assign n8478 = pi0962 & n7359;
  assign n8479 = pi1414 & n5219;
  assign n8480 = ~n8478 & ~n8479;
  assign n8481 = ~n8477 & n8480;
  assign n8482 = ~n8476 & n8481;
  assign n8483 = n7373 & ~n8482;
  assign n8484 = pi1813 & n5481;
  assign n8485 = pi1827 & n5219;
  assign n8486 = pi1686 & n7359;
  assign n8487 = pi1022 & n5218;
  assign n8488 = ~n8486 & ~n8487;
  assign n8489 = ~n8485 & n8488;
  assign n8490 = ~n8484 & n8489;
  assign n8491 = n7364 & ~n8490;
  assign n8492 = ~n8483 & ~n8491;
  assign n8493 = ~n8475 & n8492;
  assign n8494 = n5215 & ~n8493;
  assign n8495 = ~n8464 & ~n8494;
  assign po0483 = pi1169 & ~n8495;
  assign n8497 = ~pi0433 & ~n5215;
  assign n8498 = ~pi0354 & ~n8430;
  assign n8499 = pi1452 & n5481;
  assign n8500 = pi1426 & n5219;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = pi1402 & n5218;
  assign n8503 = pi1778 & n7359;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = n8501 & n8504;
  assign n8506 = pi0354 & ~n8505;
  assign n8507 = ~n8498 & ~n8506;
  assign n8508 = n5216 & ~n8507;
  assign n8509 = pi1441 & n5481;
  assign n8510 = pi1416 & n5219;
  assign n8511 = pi0964 & n7359;
  assign n8512 = pi1392 & n5218;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = ~n8510 & n8513;
  assign n8515 = ~n8509 & n8514;
  assign n8516 = n7364 & ~n8515;
  assign n8517 = n7373 & ~n8457;
  assign n8518 = ~n8516 & ~n8517;
  assign n8519 = ~n8508 & n8518;
  assign n8520 = n5215 & ~n8519;
  assign n8521 = ~n8497 & ~n8520;
  assign po0484 = pi1169 & ~n8521;
  assign n8523 = ~pi0354 & ~n8457;
  assign n8524 = pi1428 & n5219;
  assign n8525 = pi1404 & n5218;
  assign n8526 = pi1454 & n5481;
  assign n8527 = pi1769 & n7359;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = ~n8525 & n8528;
  assign n8530 = ~n8524 & n8529;
  assign n8531 = pi0354 & ~n8530;
  assign n8532 = ~n8523 & ~n8531;
  assign n8533 = n5216 & ~n8532;
  assign n8534 = pi1687 & n7359;
  assign n8535 = pi1443 & n5481;
  assign n8536 = pi1394 & n5218;
  assign n8537 = pi1418 & n5219;
  assign n8538 = ~n8536 & ~n8537;
  assign n8539 = ~n8535 & n8538;
  assign n8540 = ~n8534 & n8539;
  assign n8541 = n7364 & ~n8540;
  assign n8542 = n7373 & ~n8515;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = ~n8533 & n8543;
  assign n8545 = n5215 & ~n8544;
  assign n8546 = ~pi0434 & ~n5215;
  assign n8547 = ~n8545 & ~n8546;
  assign po0485 = pi1169 & ~n8547;
  assign n8549 = ~pi0435 & ~n5215;
  assign n8550 = ~pi0354 & ~n8490;
  assign n8551 = pi1429 & n5219;
  assign n8552 = pi0968 & n7359;
  assign n8553 = pi1455 & n5481;
  assign n8554 = pi1405 & n5218;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = ~n8552 & n8555;
  assign n8557 = ~n8551 & n8556;
  assign n8558 = pi0354 & ~n8557;
  assign n8559 = ~n8550 & ~n8558;
  assign n8560 = n5216 & ~n8559;
  assign n8561 = pi1442 & n5481;
  assign n8562 = pi1393 & n5218;
  assign n8563 = pi1788 & n7359;
  assign n8564 = pi1417 & n5219;
  assign n8565 = ~n8563 & ~n8564;
  assign n8566 = ~n8562 & n8565;
  assign n8567 = ~n8561 & n8566;
  assign n8568 = n7373 & ~n8567;
  assign n8569 = pi1809 & n5481;
  assign n8570 = pi0965 & n7359;
  assign n8571 = pi1825 & n5219;
  assign n8572 = pi1023 & n5218;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = ~n8570 & n8573;
  assign n8575 = ~n8569 & n8574;
  assign n8576 = n7364 & ~n8575;
  assign n8577 = ~n8568 & ~n8576;
  assign n8578 = ~n8560 & n8577;
  assign n8579 = n5215 & ~n8578;
  assign n8580 = ~n8549 & ~n8579;
  assign po0486 = pi1169 & ~n8580;
  assign n8582 = ~pi0354 & ~n7395;
  assign n8583 = pi0354 & ~n8515;
  assign n8584 = ~n8582 & ~n8583;
  assign n8585 = n5216 & ~n8584;
  assign n8586 = n7373 & ~n7387;
  assign n8587 = pi1803 & n5481;
  assign n8588 = pi1830 & n5218;
  assign n8589 = pi1431 & n5219;
  assign n8590 = pi0969 & n7359;
  assign n8591 = ~n8589 & ~n8590;
  assign n8592 = ~n8588 & n8591;
  assign n8593 = ~n8587 & n8592;
  assign n8594 = n7364 & ~n8593;
  assign n8595 = ~n8586 & ~n8594;
  assign n8596 = ~n8585 & n8595;
  assign n8597 = n5215 & ~n8596;
  assign n8598 = ~pi0436 & ~n5215;
  assign n8599 = ~n8597 & ~n8598;
  assign po0487 = pi1169 & ~n8599;
  assign n8601 = pi0354 & ~n8567;
  assign n8602 = ~pi0354 & ~n7372;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = n5216 & ~n8603;
  assign n8605 = ~n7363 & n7373;
  assign n8606 = pi1457 & n5481;
  assign n8607 = pi1697 & n7359;
  assign n8608 = pi1407 & n5218;
  assign n8609 = pi1432 & n5219;
  assign n8610 = ~n8608 & ~n8609;
  assign n8611 = ~n8607 & n8610;
  assign n8612 = ~n8606 & n8611;
  assign n8613 = n7364 & ~n8612;
  assign n8614 = ~n8605 & ~n8613;
  assign n8615 = ~n8604 & n8614;
  assign n8616 = n5215 & ~n8615;
  assign n8617 = ~pi0437 & ~n5215;
  assign n8618 = ~n8616 & ~n8617;
  assign po0488 = pi1169 & ~n8618;
  assign n8620 = pi0354 & ~n8540;
  assign n8621 = ~pi0354 & ~n7387;
  assign n8622 = ~n8620 & ~n8621;
  assign n8623 = n5216 & ~n8622;
  assign n8624 = n7373 & ~n8593;
  assign n8625 = n7364 & ~n8339;
  assign n8626 = ~n8624 & ~n8625;
  assign n8627 = ~n8623 & n8626;
  assign n8628 = n5215 & ~n8627;
  assign n8629 = ~pi0438 & ~n5215;
  assign n8630 = ~n8628 & ~n8629;
  assign po0489 = pi1169 & ~n8630;
  assign n8632 = ~pi0439 & ~n5215;
  assign n8633 = ~pi0354 & ~n8593;
  assign n8634 = pi1420 & n5219;
  assign n8635 = pi1396 & n5218;
  assign n8636 = pi1445 & n5481;
  assign n8637 = pi1782 & n7359;
  assign n8638 = ~n8636 & ~n8637;
  assign n8639 = ~n8635 & n8638;
  assign n8640 = ~n8634 & n8639;
  assign n8641 = pi0354 & ~n8640;
  assign n8642 = ~n8633 & ~n8641;
  assign n8643 = n5216 & ~n8642;
  assign n8644 = n7364 & ~n8365;
  assign n8645 = n7373 & ~n8339;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = ~n8643 & n8646;
  assign n8648 = n5215 & ~n8647;
  assign n8649 = ~n8632 & ~n8648;
  assign po0490 = pi1169 & ~n8649;
  assign n8651 = ~pi0440 & ~n5215;
  assign n8652 = ~pi0354 & ~n8612;
  assign n8653 = pi1446 & n5481;
  assign n8654 = pi1421 & n5219;
  assign n8655 = ~n8653 & ~n8654;
  assign n8656 = pi1397 & n5218;
  assign n8657 = pi1689 & n7359;
  assign n8658 = ~n8656 & ~n8657;
  assign n8659 = n8655 & n8658;
  assign n8660 = pi0354 & ~n8659;
  assign n8661 = ~n8652 & ~n8660;
  assign n8662 = n5216 & ~n8661;
  assign n8663 = n7364 & ~n8405;
  assign n8664 = n7373 & ~n8379;
  assign n8665 = ~n8663 & ~n8664;
  assign n8666 = ~n8662 & n8665;
  assign n8667 = n5215 & ~n8666;
  assign n8668 = ~n8651 & ~n8667;
  assign po0491 = pi1169 & ~n8668;
  assign n8670 = ~pi0441 & ~n7546;
  assign n8671 = pi0791 & n7453;
  assign n8672 = pi1962 & n7832;
  assign n8673 = ~n8671 & ~n8672;
  assign n8674 = pi1979 & n7548;
  assign n8675 = n8673 & ~n8674;
  assign n8676 = n7546 & ~n8675;
  assign n8677 = ~n8670 & ~n8676;
  assign n8678 = n7544 & ~n8677;
  assign n8679 = ~pi0441 & ~n7544;
  assign po0492 = n8678 | n8679;
  assign n8681 = ~pi0442 & ~n7546;
  assign n8682 = pi0792 & n7453;
  assign n8683 = pi0814 & n7832;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = pi0877 & n7548;
  assign n8686 = n8684 & ~n8685;
  assign n8687 = n7546 & ~n8686;
  assign n8688 = ~n8681 & ~n8687;
  assign n8689 = n7544 & ~n8688;
  assign n8690 = ~pi0442 & ~n7544;
  assign po0493 = n8689 | n8690;
  assign n8692 = ~pi0443 & ~n7546;
  assign n8693 = pi0793 & n7453;
  assign n8694 = pi0480 & n7832;
  assign n8695 = ~n8693 & ~n8694;
  assign n8696 = pi0871 & n7548;
  assign n8697 = n8695 & ~n8696;
  assign n8698 = n7546 & ~n8697;
  assign n8699 = ~n8692 & ~n8698;
  assign n8700 = n7544 & ~n8699;
  assign n8701 = ~pi0443 & ~n7544;
  assign po0494 = n8700 | n8701;
  assign n8703 = ~pi0444 & ~n7546;
  assign n8704 = n7546 & ~n7848;
  assign n8705 = ~n8703 & ~n8704;
  assign n8706 = n7544 & ~n8705;
  assign n8707 = ~pi0444 & ~n7544;
  assign po0495 = n8706 | n8707;
  assign n8709 = ~pi0445 & ~n7546;
  assign n8710 = n7546 & ~n7859;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = n7544 & ~n8711;
  assign n8713 = ~pi0445 & ~n7544;
  assign po0496 = n8712 | n8713;
  assign n8715 = ~pi0446 & ~n7546;
  assign n8716 = pi0796 & n7453;
  assign n8717 = pi0213 & n7832;
  assign n8718 = ~n8716 & ~n8717;
  assign n8719 = pi0335 & n7548;
  assign n8720 = n8718 & ~n8719;
  assign n8721 = n7546 & ~n8720;
  assign n8722 = ~n8715 & ~n8721;
  assign n8723 = n7544 & ~n8722;
  assign n8724 = ~pi0446 & ~n7544;
  assign po0497 = n8723 | n8724;
  assign n8726 = ~pi0447 & ~n7546;
  assign n8727 = pi0797 & n7453;
  assign n8728 = pi0208 & n7832;
  assign n8729 = ~n8727 & ~n8728;
  assign n8730 = pi0233 & n7548;
  assign n8731 = n8729 & ~n8730;
  assign n8732 = n7546 & ~n8731;
  assign n8733 = ~n8726 & ~n8732;
  assign n8734 = n7544 & ~n8733;
  assign n8735 = ~pi0447 & ~n7544;
  assign po0498 = n8734 | n8735;
  assign n8737 = ~pi0448 & ~n7546;
  assign n8738 = n7546 & ~n7892;
  assign n8739 = ~n8737 & ~n8738;
  assign n8740 = n7544 & ~n8739;
  assign n8741 = ~pi0448 & ~n7544;
  assign po0499 = n8740 | n8741;
  assign n8743 = ~pi0946 & pi1930;
  assign n8744 = pi0836 & n8743;
  assign n8745 = pi0449 & ~n8744;
  assign n8746 = pi1144 & pi1905;
  assign po0500 = n8745 | n8746;
  assign n8748 = ~pi1907 & n5253;
  assign po0501 = ~pi0450 | n8748;
  assign n8750 = ~pi1904 & n5272;
  assign po0502 = ~pi0451 | n8750;
  assign n8752 = ~pi1909 & n5291;
  assign po0503 = ~pi0452 | n8752;
  assign n8754 = ~pi1910 & n5234;
  assign po0504 = ~pi0453 | n8754;
  assign n8756 = pi0354 & ~n8575;
  assign n8757 = ~pi0354 & ~n7363;
  assign n8758 = ~n8756 & ~n8757;
  assign n8759 = n5216 & ~n8758;
  assign n8760 = n7364 & ~n8379;
  assign n8761 = n7373 & ~n8612;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = ~n8759 & n8762;
  assign n8764 = n5215 & ~n8763;
  assign n8765 = ~pi0454 & ~n5215;
  assign n8766 = ~n8764 & ~n8765;
  assign po0505 = pi1169 & ~n8766;
  assign n8768 = ~pi0455 & ~n5215;
  assign n8769 = ~pi0354 & ~n8482;
  assign n8770 = pi1453 & n5481;
  assign n8771 = pi1427 & n5219;
  assign n8772 = ~n8770 & ~n8771;
  assign n8773 = pi1403 & n5218;
  assign n8774 = pi1695 & n7359;
  assign n8775 = ~n8773 & ~n8774;
  assign n8776 = n8772 & n8775;
  assign n8777 = pi0354 & ~n8776;
  assign n8778 = ~n8769 & ~n8777;
  assign n8779 = n5216 & ~n8778;
  assign n8780 = n7364 & ~n8567;
  assign n8781 = n7373 & ~n8490;
  assign n8782 = ~n8780 & ~n8781;
  assign n8783 = ~n8779 & n8782;
  assign n8784 = n5215 & ~n8783;
  assign n8785 = ~n8768 & ~n8784;
  assign po0506 = pi1169 & ~n8785;
  assign n8787 = ~pi0457 & ~n5215;
  assign n8788 = ~pi0354 & ~n8405;
  assign n8789 = pi1450 & n5481;
  assign n8790 = pi1424 & n5219;
  assign n8791 = ~n8789 & ~n8790;
  assign n8792 = pi1400 & n5218;
  assign n8793 = pi1693 & n7359;
  assign n8794 = ~n8792 & ~n8793;
  assign n8795 = n8791 & n8794;
  assign n8796 = pi0354 & ~n8795;
  assign n8797 = ~n8788 & ~n8796;
  assign n8798 = n5216 & ~n8797;
  assign n8799 = n7364 & ~n8482;
  assign n8800 = n7373 & ~n8397;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8798 & n8801;
  assign n8803 = n5215 & ~n8802;
  assign n8804 = ~n8787 & ~n8803;
  assign po0508 = pi1169 & ~n8804;
  assign n8806 = ~pi1134 & ~pi1146;
  assign n8807 = ~pi0790 & n8806;
  assign po1927 = pi0939 & pi1952;
  assign n8809 = ~pi1876 & po1927;
  assign n8810 = ~n8807 & n8809;
  assign n8811 = ~pi0458 & ~n8810;
  assign n8812 = ~pi0601 & ~pi0602;
  assign n8813 = pi0458 & ~n8812;
  assign n8814 = pi1134 & ~pi1146;
  assign n8815 = pi0196 & n8814;
  assign n8816 = pi1886 & n8806;
  assign n8817 = ~n8815 & ~n8816;
  assign n8818 = n8812 & n8817;
  assign n8819 = ~n8813 & ~n8818;
  assign n8820 = n8810 & n8819;
  assign po0509 = n8811 | n8820;
  assign n8822 = ~pi0459 & ~n8810;
  assign n8823 = pi0601 & pi0602;
  assign n8824 = pi0212 & n8806;
  assign n8825 = n8823 & n8824;
  assign n8826 = ~pi0459 & ~n8823;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = n8810 & ~n8827;
  assign po0510 = n8822 | n8828;
  assign n8830 = ~pi0460 & ~n8810;
  assign n8831 = pi0819 & n8806;
  assign n8832 = n8823 & n8831;
  assign n8833 = ~pi0460 & ~n8823;
  assign n8834 = ~n8832 & ~n8833;
  assign n8835 = n8810 & ~n8834;
  assign po0511 = n8830 | n8835;
  assign n8837 = ~pi1157 & ~pi1158;
  assign n8838 = ~pi0821 & n8837;
  assign po1932 = pi0938 & ~pi1931;
  assign n8840 = pi1881 & po1932;
  assign n8841 = ~n8838 & n8840;
  assign n8842 = ~pi0461 & ~n8841;
  assign n8843 = pi0746 & pi0843;
  assign n8844 = pi0195 & n8837;
  assign n8845 = n8843 & n8844;
  assign n8846 = ~pi0461 & ~n8843;
  assign n8847 = ~n8845 & ~n8846;
  assign n8848 = n8841 & ~n8847;
  assign po0512 = n8842 | n8848;
  assign n8850 = ~pi0462 & ~n8841;
  assign n8851 = pi0333 & n8837;
  assign n8852 = n8843 & n8851;
  assign n8853 = ~pi0462 & ~n8843;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = n8841 & ~n8854;
  assign po0513 = n8850 | n8855;
  assign n8857 = pi0463 & ~n8809;
  assign n8858 = pi0463 & n8823;
  assign n8859 = ~pi0463 & ~n8823;
  assign n8860 = ~n8858 & ~n8859;
  assign n8861 = ~n8806 & n8860;
  assign n8862 = pi0601 & pi0790;
  assign n8863 = pi0602 & n8862;
  assign n8864 = pi0463 & ~n8863;
  assign n8865 = ~pi0463 & n8863;
  assign n8866 = ~n8864 & ~n8865;
  assign n8867 = n8806 & ~n8866;
  assign n8868 = ~n8861 & ~n8867;
  assign n8869 = n8809 & ~n8868;
  assign n8870 = ~n8857 & ~n8869;
  assign po0514 = pi1036 & ~n8870;
  assign n8872 = ~pi0464 & ~n8841;
  assign n8873 = pi0883 & n8837;
  assign n8874 = n8843 & n8873;
  assign n8875 = ~pi0464 & ~n8843;
  assign n8876 = ~n8874 & ~n8875;
  assign n8877 = n8841 & ~n8876;
  assign po0515 = n8872 | n8877;
  assign n8879 = ~pi0465 & ~n8841;
  assign n8880 = pi0746 & ~pi0843;
  assign n8881 = pi0465 & ~n8880;
  assign n8882 = pi0211 & n8837;
  assign n8883 = n8880 & ~n8882;
  assign n8884 = ~n8881 & ~n8883;
  assign n8885 = n8841 & n8884;
  assign po0516 = n8879 | n8885;
  assign n8887 = ~pi0466 & ~n8841;
  assign n8888 = pi0466 & ~n8880;
  assign n8889 = pi0818 & n8837;
  assign n8890 = n8880 & ~n8889;
  assign n8891 = ~n8888 & ~n8890;
  assign n8892 = n8841 & n8891;
  assign po0517 = n8887 | n8892;
  assign n8894 = ~pi0467 & ~n8841;
  assign n8895 = pi0467 & ~n8880;
  assign n8896 = pi0951 & n8837;
  assign n8897 = n8880 & ~n8896;
  assign n8898 = ~n8895 & ~n8897;
  assign n8899 = n8841 & n8898;
  assign po0518 = n8894 | n8899;
  assign n8901 = ~pi0468 & ~n8841;
  assign n8902 = ~pi0746 & pi0843;
  assign n8903 = pi0468 & ~n8902;
  assign n8904 = ~n8882 & n8902;
  assign n8905 = ~n8903 & ~n8904;
  assign n8906 = n8841 & n8905;
  assign po0519 = n8901 | n8906;
  assign n8908 = ~pi0469 & ~n8841;
  assign n8909 = pi0469 & ~n8902;
  assign n8910 = pi0481 & n8837;
  assign n8911 = n8902 & ~n8910;
  assign n8912 = ~n8909 & ~n8911;
  assign n8913 = n8841 & n8912;
  assign po0520 = n8908 | n8913;
  assign n8915 = ~pi0470 & ~n8841;
  assign n8916 = pi0470 & ~n8902;
  assign n8917 = ~n8873 & n8902;
  assign n8918 = ~n8916 & ~n8917;
  assign n8919 = n8841 & n8918;
  assign po0521 = n8915 | n8919;
  assign n8921 = ~pi0471 & ~n8810;
  assign n8922 = ~pi0601 & pi0602;
  assign n8923 = pi0471 & ~n8922;
  assign n8924 = ~n8831 & n8922;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = n8810 & n8925;
  assign po0522 = n8921 | n8926;
  assign n8928 = n7454 & ~n8720;
  assign n8929 = ~pi0472 & ~n7454;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = n7544 & ~n8930;
  assign n8932 = ~pi0472 & ~n7544;
  assign po0523 = n8931 | n8932;
  assign n8934 = n7454 & ~n8675;
  assign n8935 = ~pi0473 & ~n7454;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = n7544 & ~n8936;
  assign n8938 = ~pi0473 & ~n7544;
  assign po0524 = n8937 | n8938;
  assign n8940 = n7454 & ~n7859;
  assign n8941 = ~pi0474 & ~n7454;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = n7544 & ~n8942;
  assign n8944 = ~pi0474 & ~n7544;
  assign po0525 = n8943 | n8944;
  assign n8946 = pi0601 & ~pi0602;
  assign n8947 = ~pi0475 & ~n8946;
  assign n8948 = pi0831 & n8806;
  assign n8949 = ~pi1134 & pi1146;
  assign n8950 = pi1983 & n8949;
  assign n8951 = ~n8948 & ~n8950;
  assign n8952 = pi1984 & n8814;
  assign n8953 = n8951 & ~n8952;
  assign n8954 = n8946 & ~n8953;
  assign n8955 = ~n8947 & ~n8954;
  assign n8956 = n8810 & ~n8955;
  assign n8957 = ~pi0475 & ~n8810;
  assign po0526 = n8956 | n8957;
  assign n8959 = ~pi0476 & ~n7566;
  assign n8960 = n7566 & ~n8731;
  assign n8961 = ~n8959 & ~n8960;
  assign n8962 = n7544 & ~n8961;
  assign n8963 = ~pi0476 & ~n7544;
  assign po0527 = n8962 | n8963;
  assign n8965 = ~pi0477 & ~n7566;
  assign n8966 = n7566 & ~n7942;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = n7544 & ~n8967;
  assign n8969 = ~pi0477 & ~n7544;
  assign po0528 = n8968 | n8969;
  assign n8971 = pi0876 & ~pi2056;
  assign n8972 = pi0478 & pi2056;
  assign po0529 = n8971 | n8972;
  assign n8974 = pi0876 & ~pi2057;
  assign n8975 = pi0479 & pi2057;
  assign po0530 = n8974 | n8975;
  assign n8977 = pi0876 & ~pi2058;
  assign n8978 = pi0480 & pi2058;
  assign po0531 = n8977 | n8978;
  assign n8980 = pi0876 & ~pi2059;
  assign n8981 = pi0481 & pi2059;
  assign po0532 = n8980 | n8981;
  assign n8983 = ~pi0482 & ~n8810;
  assign n8984 = pi0482 & ~n8922;
  assign n8985 = n8817 & n8922;
  assign n8986 = ~n8984 & ~n8985;
  assign n8987 = n8810 & n8986;
  assign po0533 = n8983 | n8987;
  assign n8989 = ~pi0483 & ~n8810;
  assign n8990 = pi0483 & ~n8922;
  assign n8991 = pi0192 & n8814;
  assign n8992 = pi1852 & n8806;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = n8922 & n8993;
  assign n8995 = ~n8990 & ~n8994;
  assign n8996 = n8810 & n8995;
  assign po0534 = n8989 | n8996;
  assign n8998 = ~pi0484 & ~n8810;
  assign n8999 = pi0484 & ~n8922;
  assign n9000 = pi0950 & n8806;
  assign n9001 = n8922 & ~n9000;
  assign n9002 = ~n8999 & ~n9001;
  assign n9003 = n8810 & n9002;
  assign po0535 = n8998 | n9003;
  assign n9005 = ~pi0485 & ~n8810;
  assign n9006 = pi0485 & ~n8922;
  assign n9007 = pi0915 & n8806;
  assign n9008 = n8922 & ~n9007;
  assign n9009 = ~n9006 & ~n9008;
  assign n9010 = n8810 & n9009;
  assign po0536 = n9005 | n9010;
  assign n9012 = ~pi0486 & ~n8810;
  assign n9013 = pi0486 & ~n8922;
  assign n9014 = pi0882 & n8806;
  assign n9015 = n8922 & ~n9014;
  assign n9016 = ~n9013 & ~n9015;
  assign n9017 = n8810 & n9016;
  assign po0537 = n9012 | n9017;
  assign n9019 = ~pi0487 & ~n8841;
  assign n9020 = ~pi0746 & ~pi0843;
  assign n9021 = pi0487 & ~n9020;
  assign n9022 = ~pi1157 & pi1158;
  assign n9023 = pi0195 & n9022;
  assign n9024 = pi1883 & n8837;
  assign n9025 = ~n9023 & ~n9024;
  assign n9026 = n9020 & n9025;
  assign n9027 = ~n9021 & ~n9026;
  assign n9028 = n8841 & n9027;
  assign po0538 = n9019 | n9028;
  assign n9030 = ~pi0488 & ~n8841;
  assign n9031 = pi0488 & ~n9020;
  assign n9032 = pi0191 & n9022;
  assign n9033 = pi1853 & n8837;
  assign n9034 = ~n9032 & ~n9033;
  assign n9035 = n9020 & n9034;
  assign n9036 = ~n9031 & ~n9035;
  assign n9037 = n8841 & n9036;
  assign po0539 = n9030 | n9037;
  assign n9039 = ~pi0489 & ~n8810;
  assign n9040 = pi0489 & ~n8922;
  assign n9041 = pi0866 & n8806;
  assign n9042 = n8922 & ~n9041;
  assign n9043 = ~n9040 & ~n9042;
  assign n9044 = n8810 & n9043;
  assign po0540 = n9039 | n9044;
  assign n9046 = ~pi0490 & ~n8810;
  assign n9047 = pi0490 & ~n8922;
  assign n9048 = pi0479 & n8806;
  assign n9049 = n8922 & ~n9048;
  assign n9050 = ~n9047 & ~n9049;
  assign n9051 = n8810 & n9050;
  assign po0541 = n9046 | n9051;
  assign n9053 = ~pi0491 & ~n8810;
  assign n9054 = pi0491 & ~n8922;
  assign n9055 = pi0334 & n8806;
  assign n9056 = n8922 & ~n9055;
  assign n9057 = ~n9054 & ~n9056;
  assign n9058 = n8810 & n9057;
  assign po0542 = n9053 | n9058;
  assign n9060 = ~pi0492 & ~n8810;
  assign n9061 = pi0492 & ~n8922;
  assign n9062 = pi0235 & n8806;
  assign n9063 = n8922 & ~n9062;
  assign n9064 = ~n9061 & ~n9063;
  assign n9065 = n8810 & n9064;
  assign po0543 = n9060 | n9065;
  assign n9067 = ~pi0493 & ~n8841;
  assign n9068 = pi0493 & ~n8902;
  assign n9069 = n8902 & n9025;
  assign n9070 = ~n9068 & ~n9069;
  assign n9071 = n8841 & n9070;
  assign po0544 = n9067 | n9071;
  assign n9073 = ~pi0494 & ~n8841;
  assign n9074 = pi0494 & ~n8902;
  assign n9075 = n8902 & n9034;
  assign n9076 = ~n9074 & ~n9075;
  assign n9077 = n8841 & n9076;
  assign po0545 = n9073 | n9077;
  assign n9079 = ~pi0495 & ~n8841;
  assign n9080 = pi0495 & ~n8902;
  assign n9081 = ~n8896 & n8902;
  assign n9082 = ~n9080 & ~n9081;
  assign n9083 = n8841 & n9082;
  assign po0546 = n9079 | n9083;
  assign n9085 = ~pi0496 & ~n8841;
  assign n9086 = pi0496 & ~n8902;
  assign n9087 = pi0916 & n8837;
  assign n9088 = n8902 & ~n9087;
  assign n9089 = ~n9086 & ~n9088;
  assign n9090 = n8841 & n9089;
  assign po0547 = n9085 | n9090;
  assign n9092 = ~pi0497 & ~n8810;
  assign n9093 = pi0497 & ~n8922;
  assign n9094 = ~n8824 & n8922;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = n8810 & n9095;
  assign po0548 = n9092 | n9096;
  assign n9098 = ~pi0498 & ~n8841;
  assign n9099 = pi0498 & ~n8902;
  assign n9100 = pi0870 & n8837;
  assign n9101 = n8902 & ~n9100;
  assign n9102 = ~n9099 & ~n9101;
  assign n9103 = n8841 & n9102;
  assign po0549 = n9098 | n9103;
  assign n9105 = ~pi0499 & ~n8841;
  assign n9106 = pi0499 & ~n8902;
  assign n9107 = ~n8889 & n8902;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = n8841 & n9108;
  assign po0550 = n9105 | n9109;
  assign n9111 = ~pi0500 & ~n8841;
  assign n9112 = pi0500 & ~n8902;
  assign n9113 = ~n8851 & n8902;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = n8841 & n9114;
  assign po0551 = n9111 | n9115;
  assign n9117 = ~pi0501 & ~n8810;
  assign n9118 = pi0501 & ~n8922;
  assign n9119 = pi0207 & n8806;
  assign n9120 = n8922 & ~n9119;
  assign n9121 = ~n9118 & ~n9120;
  assign n9122 = n8810 & n9121;
  assign po0552 = n9117 | n9122;
  assign n9124 = ~pi0502 & ~n8841;
  assign n9125 = pi0502 & ~n8902;
  assign n9126 = pi0231 & n8837;
  assign n9127 = n8902 & ~n9126;
  assign n9128 = ~n9125 & ~n9127;
  assign n9129 = n8841 & n9128;
  assign po0553 = n9124 | n9129;
  assign n9131 = ~pi0503 & ~n8841;
  assign n9132 = pi0503 & ~n8902;
  assign n9133 = pi0206 & n8837;
  assign n9134 = n8902 & ~n9133;
  assign n9135 = ~n9132 & ~n9134;
  assign n9136 = n8841 & n9135;
  assign po0554 = n9131 | n9136;
  assign n9138 = ~pi0504 & ~n8841;
  assign n9139 = pi0504 & ~n8902;
  assign n9140 = ~n8844 & n8902;
  assign n9141 = ~n9139 & ~n9140;
  assign n9142 = n8841 & n9141;
  assign po0555 = n9138 | n9142;
  assign n9144 = ~pi0505 & ~n8841;
  assign n9145 = pi0505 & ~n8902;
  assign n9146 = pi0191 & n8837;
  assign n9147 = n8902 & ~n9146;
  assign n9148 = ~n9145 & ~n9147;
  assign n9149 = n8841 & n9148;
  assign po0556 = n9144 | n9149;
  assign n9151 = ~pi0506 & ~n8810;
  assign n9152 = pi0506 & ~n8922;
  assign n9153 = pi0196 & n8806;
  assign n9154 = n8922 & ~n9153;
  assign n9155 = ~n9152 & ~n9154;
  assign n9156 = n8810 & n9155;
  assign po0557 = n9151 | n9156;
  assign n9158 = ~pi0507 & ~n8841;
  assign n9159 = pi0507 & ~n8880;
  assign n9160 = n8880 & n9025;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = n8841 & n9161;
  assign po0558 = n9158 | n9162;
  assign n9164 = ~pi0508 & ~n8841;
  assign n9165 = pi0508 & ~n8880;
  assign n9166 = n8880 & n9034;
  assign n9167 = ~n9165 & ~n9166;
  assign n9168 = n8841 & n9167;
  assign po0559 = n9164 | n9168;
  assign n9170 = ~pi0509 & ~n8810;
  assign n9171 = pi0509 & ~n8922;
  assign n9172 = pi0192 & n8806;
  assign n9173 = n8922 & ~n9172;
  assign n9174 = ~n9171 & ~n9173;
  assign n9175 = n8810 & n9174;
  assign po0560 = n9170 | n9175;
  assign n9177 = ~pi0510 & ~n8841;
  assign n9178 = pi0510 & ~n8880;
  assign n9179 = n8880 & ~n9087;
  assign n9180 = ~n9178 & ~n9179;
  assign n9181 = n8841 & n9180;
  assign po0561 = n9177 | n9181;
  assign n9183 = ~pi0511 & ~n8841;
  assign n9184 = pi0511 & ~n8880;
  assign n9185 = ~n8873 & n8880;
  assign n9186 = ~n9184 & ~n9185;
  assign n9187 = n8841 & n9186;
  assign po0562 = n9183 | n9187;
  assign n9189 = ~pi0512 & ~n8841;
  assign n9190 = pi0512 & ~n8880;
  assign n9191 = n8880 & ~n9100;
  assign n9192 = ~n9190 & ~n9191;
  assign n9193 = n8841 & n9192;
  assign po0563 = n9189 | n9193;
  assign n9195 = ~pi0513 & ~n8841;
  assign n9196 = pi0513 & ~n8880;
  assign n9197 = n8880 & ~n8910;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = n8841 & n9198;
  assign po0564 = n9195 | n9199;
  assign n9201 = ~pi0514 & ~n8841;
  assign n9202 = pi0514 & ~n8880;
  assign n9203 = ~n8851 & n8880;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = n8841 & n9204;
  assign po0565 = n9201 | n9205;
  assign n9207 = ~pi0515 & ~n8841;
  assign n9208 = pi0515 & ~n8880;
  assign n9209 = n8880 & ~n9126;
  assign n9210 = ~n9208 & ~n9209;
  assign n9211 = n8841 & n9210;
  assign po0566 = n9207 | n9211;
  assign n9213 = ~pi0516 & ~n8841;
  assign n9214 = pi0516 & ~n8880;
  assign n9215 = n8880 & ~n9133;
  assign n9216 = ~n9214 & ~n9215;
  assign n9217 = n8841 & n9216;
  assign po0567 = n9213 | n9217;
  assign n9219 = ~pi0517 & ~n8841;
  assign n9220 = pi0517 & ~n8880;
  assign n9221 = ~n8844 & n8880;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = n8841 & n9222;
  assign po0568 = n9219 | n9223;
  assign n9225 = ~pi0518 & ~n8841;
  assign n9226 = pi0518 & ~n8880;
  assign n9227 = n8880 & ~n9146;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = n8841 & n9228;
  assign po0569 = n9225 | n9229;
  assign n9231 = ~pi0519 & ~n8841;
  assign n9232 = n8843 & ~n9025;
  assign n9233 = ~pi0519 & ~n8843;
  assign n9234 = ~n9232 & ~n9233;
  assign n9235 = n8841 & ~n9234;
  assign po0570 = n9231 | n9235;
  assign n9237 = ~pi0520 & ~n8841;
  assign n9238 = n8843 & ~n9034;
  assign n9239 = ~pi0520 & ~n8843;
  assign n9240 = ~n9238 & ~n9239;
  assign n9241 = n8841 & ~n9240;
  assign po0571 = n9237 | n9241;
  assign n9243 = ~pi0521 & ~n8841;
  assign n9244 = n8843 & n8896;
  assign n9245 = ~pi0521 & ~n8843;
  assign n9246 = ~n9244 & ~n9245;
  assign n9247 = n8841 & ~n9246;
  assign po0572 = n9243 | n9247;
  assign n9249 = ~pi0522 & ~n8841;
  assign n9250 = n8843 & n9087;
  assign n9251 = ~pi0522 & ~n8843;
  assign n9252 = ~n9250 & ~n9251;
  assign n9253 = n8841 & ~n9252;
  assign po0573 = n9249 | n9253;
  assign n9255 = ~pi0523 & ~n8841;
  assign n9256 = n8843 & n9100;
  assign n9257 = ~pi0523 & ~n8843;
  assign n9258 = ~n9256 & ~n9257;
  assign n9259 = n8841 & ~n9258;
  assign po0574 = n9255 | n9259;
  assign n9261 = ~pi0524 & ~n8841;
  assign n9262 = n8843 & n8889;
  assign n9263 = ~pi0524 & ~n8843;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = n8841 & ~n9264;
  assign po0575 = n9261 | n9265;
  assign n9267 = ~pi0525 & ~n8841;
  assign n9268 = n8843 & n8910;
  assign n9269 = ~pi0525 & ~n8843;
  assign n9270 = ~n9268 & ~n9269;
  assign n9271 = n8841 & ~n9270;
  assign po0576 = n9267 | n9271;
  assign n9273 = ~pi0526 & ~n8841;
  assign n9274 = n8843 & n9126;
  assign n9275 = ~pi0526 & ~n8843;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = n8841 & ~n9276;
  assign po0577 = n9273 | n9277;
  assign n9279 = ~pi0527 & ~n8841;
  assign n9280 = n8843 & n8882;
  assign n9281 = ~pi0527 & ~n8843;
  assign n9282 = ~n9280 & ~n9281;
  assign n9283 = n8841 & ~n9282;
  assign po0578 = n9279 | n9283;
  assign n9285 = ~pi0528 & ~n8841;
  assign n9286 = n8843 & n9133;
  assign n9287 = ~pi0528 & ~n8843;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = n8841 & ~n9288;
  assign po0579 = n9285 | n9289;
  assign n9291 = ~pi0529 & ~n8841;
  assign n9292 = n8843 & n9146;
  assign n9293 = ~pi0529 & ~n8843;
  assign n9294 = ~n9292 & ~n9293;
  assign n9295 = n8841 & ~n9294;
  assign po0580 = n9291 | n9295;
  assign n9297 = ~pi0530 & ~n8810;
  assign n9298 = ~n8817 & n8823;
  assign n9299 = ~pi0530 & ~n8823;
  assign n9300 = ~n9298 & ~n9299;
  assign n9301 = n8810 & ~n9300;
  assign po0581 = n9297 | n9301;
  assign n9303 = ~pi0531 & ~n8810;
  assign n9304 = n8823 & ~n8993;
  assign n9305 = ~pi0531 & ~n8823;
  assign n9306 = ~n9304 & ~n9305;
  assign n9307 = n8810 & ~n9306;
  assign po0582 = n9303 | n9307;
  assign n9309 = ~pi0532 & ~n8810;
  assign n9310 = n8823 & n9000;
  assign n9311 = ~pi0532 & ~n8823;
  assign n9312 = ~n9310 & ~n9311;
  assign n9313 = n8810 & ~n9312;
  assign po0583 = n9309 | n9313;
  assign n9315 = ~pi0533 & ~n8810;
  assign n9316 = n8823 & n9007;
  assign n9317 = ~pi0533 & ~n8823;
  assign n9318 = ~n9316 & ~n9317;
  assign n9319 = n8810 & ~n9318;
  assign po0584 = n9315 | n9319;
  assign n9321 = ~pi0534 & ~n8810;
  assign n9322 = n8823 & n9014;
  assign n9323 = ~pi0534 & ~n8823;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = n8810 & ~n9324;
  assign po0585 = n9321 | n9325;
  assign n9327 = ~pi0535 & ~n8810;
  assign n9328 = n8823 & n9041;
  assign n9329 = ~pi0535 & ~n8823;
  assign n9330 = ~n9328 & ~n9329;
  assign n9331 = n8810 & ~n9330;
  assign po0586 = n9327 | n9331;
  assign n9333 = ~pi0536 & ~n8810;
  assign n9334 = n8823 & n9048;
  assign n9335 = ~pi0536 & ~n8823;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = n8810 & ~n9336;
  assign po0587 = n9333 | n9337;
  assign n9339 = ~pi0537 & ~n8810;
  assign n9340 = n8823 & n9055;
  assign n9341 = ~pi0537 & ~n8823;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = n8810 & ~n9342;
  assign po0588 = n9339 | n9343;
  assign n9345 = ~pi0538 & ~n8810;
  assign n9346 = n8823 & n9062;
  assign n9347 = ~pi0538 & ~n8823;
  assign n9348 = ~n9346 & ~n9347;
  assign n9349 = n8810 & ~n9348;
  assign po0589 = n9345 | n9349;
  assign n9351 = ~pi0539 & ~n8810;
  assign n9352 = n8823 & n9119;
  assign n9353 = ~pi0539 & ~n8823;
  assign n9354 = ~n9352 & ~n9353;
  assign n9355 = n8810 & ~n9354;
  assign po0590 = n9351 | n9355;
  assign n9357 = ~pi0540 & ~n8810;
  assign n9358 = n8823 & n9153;
  assign n9359 = ~pi0540 & ~n8823;
  assign n9360 = ~n9358 & ~n9359;
  assign n9361 = n8810 & ~n9360;
  assign po0591 = n9357 | n9361;
  assign n9363 = ~pi0541 & ~n8810;
  assign n9364 = n8823 & n9172;
  assign n9365 = ~pi0541 & ~n8823;
  assign n9366 = ~n9364 & ~n9365;
  assign n9367 = n8810 & ~n9366;
  assign po0592 = n9363 | n9367;
  assign n9369 = ~pi0542 & ~n8810;
  assign n9370 = pi0542 & ~n8812;
  assign n9371 = n8812 & n8993;
  assign n9372 = ~n9370 & ~n9371;
  assign n9373 = n8810 & n9372;
  assign po0593 = n9369 | n9373;
  assign n9375 = ~pi0543 & ~n8810;
  assign n9376 = pi0543 & ~n8946;
  assign n9377 = n8817 & n8946;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = n8810 & n9378;
  assign po0594 = n9375 | n9379;
  assign n9381 = ~pi0544 & ~n8810;
  assign n9382 = pi0544 & ~n8946;
  assign n9383 = n8946 & n8993;
  assign n9384 = ~n9382 & ~n9383;
  assign n9385 = n8810 & n9384;
  assign po0595 = n9381 | n9385;
  assign n9387 = ~pi0545 & ~n8810;
  assign n9388 = pi0545 & ~n8946;
  assign n9389 = n8946 & ~n9007;
  assign n9390 = ~n9388 & ~n9389;
  assign n9391 = n8810 & n9390;
  assign po0596 = n9387 | n9391;
  assign n9393 = ~pi0546 & ~n8810;
  assign n9394 = pi0546 & ~n8946;
  assign n9395 = n8946 & ~n9014;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = n8810 & n9396;
  assign po0597 = n9393 | n9397;
  assign n9399 = ~pi0547 & ~n8810;
  assign n9400 = pi0547 & ~n8946;
  assign n9401 = n8946 & ~n9041;
  assign n9402 = ~n9400 & ~n9401;
  assign n9403 = n8810 & n9402;
  assign po0598 = n9399 | n9403;
  assign n9405 = ~pi0548 & ~n8810;
  assign n9406 = pi0548 & ~n8946;
  assign n9407 = ~n8831 & n8946;
  assign n9408 = ~n9406 & ~n9407;
  assign n9409 = n8810 & n9408;
  assign po0599 = n9405 | n9409;
  assign n9411 = ~pi0549 & ~n8810;
  assign n9412 = pi0549 & ~n8946;
  assign n9413 = n8946 & ~n9048;
  assign n9414 = ~n9412 & ~n9413;
  assign n9415 = n8810 & n9414;
  assign po0600 = n9411 | n9415;
  assign n9417 = ~pi0550 & ~n8810;
  assign n9418 = pi0550 & ~n8946;
  assign n9419 = n8946 & ~n9055;
  assign n9420 = ~n9418 & ~n9419;
  assign n9421 = n8810 & n9420;
  assign po0601 = n9417 | n9421;
  assign n9423 = ~pi0551 & ~n8810;
  assign n9424 = pi0551 & ~n8946;
  assign n9425 = n8946 & ~n9062;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = n8810 & n9426;
  assign po0602 = n9423 | n9427;
  assign n9429 = ~pi0552 & ~n8810;
  assign n9430 = pi0552 & ~n8946;
  assign n9431 = ~n8824 & n8946;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = n8810 & n9432;
  assign po0603 = n9429 | n9433;
  assign n9435 = ~pi0553 & ~n8810;
  assign n9436 = pi0553 & ~n8946;
  assign n9437 = n8946 & ~n9119;
  assign n9438 = ~n9436 & ~n9437;
  assign n9439 = n8810 & n9438;
  assign po0604 = n9435 | n9439;
  assign n9441 = ~pi0554 & ~n8810;
  assign n9442 = pi0554 & ~n8946;
  assign n9443 = n8946 & ~n9000;
  assign n9444 = ~n9442 & ~n9443;
  assign n9445 = n8810 & n9444;
  assign po0605 = n9441 | n9445;
  assign n9447 = ~pi0555 & ~n8810;
  assign n9448 = pi0555 & ~n8946;
  assign n9449 = n8946 & ~n9153;
  assign n9450 = ~n9448 & ~n9449;
  assign n9451 = n8810 & n9450;
  assign po0606 = n9447 | n9451;
  assign n9453 = ~pi0556 & ~n8810;
  assign n9454 = pi0556 & ~n8946;
  assign n9455 = n8946 & ~n9172;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = n8810 & n9456;
  assign po0607 = n9453 | n9457;
  assign n9459 = n7454 & ~n7909;
  assign n9460 = ~pi0557 & ~n7454;
  assign n9461 = ~n9459 & ~n9460;
  assign n9462 = n7544 & ~n9461;
  assign n9463 = ~pi0557 & ~n7544;
  assign po0608 = n9462 | n9463;
  assign n9465 = pi0871 & n7832;
  assign n9466 = pi0923 & n7548;
  assign n9467 = ~n9465 & ~n9466;
  assign n9468 = pi0804 & n7453;
  assign n9469 = n9467 & ~n9468;
  assign n9470 = n7454 & ~n9469;
  assign n9471 = ~pi0558 & ~n7454;
  assign n9472 = ~n9470 & ~n9471;
  assign n9473 = n7544 & ~n9472;
  assign n9474 = ~pi0558 & ~n7544;
  assign po0609 = n9473 | n9474;
  assign n9476 = ~pi0559 & ~n8922;
  assign n9477 = pi0824 & n8806;
  assign n9478 = pi1980 & n8949;
  assign n9479 = ~n9477 & ~n9478;
  assign n9480 = pi1960 & n8814;
  assign n9481 = n9479 & ~n9480;
  assign n9482 = n8922 & ~n9481;
  assign n9483 = ~n9476 & ~n9482;
  assign n9484 = n8810 & ~n9483;
  assign n9485 = ~pi0559 & ~n8810;
  assign po0610 = n9484 | n9485;
  assign n9487 = ~pi0560 & ~n8922;
  assign n9488 = pi0822 & n8806;
  assign n9489 = pi1852 & n8949;
  assign n9490 = ~n9488 & ~n9489;
  assign n9491 = pi1924 & n8814;
  assign n9492 = n9490 & ~n9491;
  assign n9493 = n8922 & ~n9492;
  assign n9494 = ~n9487 & ~n9493;
  assign n9495 = n8810 & ~n9494;
  assign n9496 = ~pi0560 & ~n8810;
  assign po0611 = n9495 | n9496;
  assign n9498 = ~pi0561 & ~n8922;
  assign n9499 = pi0827 & n8806;
  assign n9500 = pi0950 & n8949;
  assign n9501 = ~n9499 & ~n9500;
  assign n9502 = pi1886 & n8814;
  assign n9503 = n9501 & ~n9502;
  assign n9504 = n8922 & ~n9503;
  assign n9505 = ~n9498 & ~n9504;
  assign n9506 = n8810 & ~n9505;
  assign n9507 = ~pi0561 & ~n8810;
  assign po0612 = n9506 | n9507;
  assign n9509 = pi0823 & n8806;
  assign n9510 = pi1924 & n8949;
  assign n9511 = ~n9509 & ~n9510;
  assign n9512 = pi1980 & n8814;
  assign n9513 = n9511 & ~n9512;
  assign n9514 = n8823 & ~n9513;
  assign n9515 = ~pi0562 & ~n8823;
  assign n9516 = ~n9514 & ~n9515;
  assign n9517 = n8810 & ~n9516;
  assign n9518 = ~pi0562 & ~n8810;
  assign po0613 = n9517 | n9518;
  assign n9520 = ~pi0563 & ~n8922;
  assign n9521 = pi0866 & n8949;
  assign n9522 = pi0915 & n8814;
  assign n9523 = ~n9521 & ~n9522;
  assign n9524 = pi0829 & n8806;
  assign n9525 = n9523 & ~n9524;
  assign n9526 = n8922 & ~n9525;
  assign n9527 = ~n9520 & ~n9526;
  assign n9528 = n8810 & ~n9527;
  assign n9529 = ~pi0563 & ~n8810;
  assign po0614 = n9528 | n9529;
  assign n9531 = ~pi0564 & ~n7566;
  assign n9532 = n7566 & ~n8675;
  assign n9533 = ~n9531 & ~n9532;
  assign n9534 = n7544 & ~n9533;
  assign n9535 = ~pi0564 & ~n7544;
  assign po0615 = n9534 | n9535;
  assign n9537 = ~pi0565 & ~n7566;
  assign n9538 = n7566 & ~n8686;
  assign n9539 = ~n9537 & ~n9538;
  assign n9540 = n7544 & ~n9539;
  assign n9541 = ~pi0565 & ~n7544;
  assign po0616 = n9540 | n9541;
  assign n9543 = ~pi0566 & ~n7566;
  assign n9544 = n7566 & ~n8697;
  assign n9545 = ~n9543 & ~n9544;
  assign n9546 = n7544 & ~n9545;
  assign n9547 = ~pi0566 & ~n7544;
  assign po0617 = n9546 | n9547;
  assign n9549 = pi0825 & n8806;
  assign n9550 = pi1934 & n8949;
  assign n9551 = ~n9549 & ~n9550;
  assign n9552 = pi1983 & n8814;
  assign n9553 = n9551 & ~n9552;
  assign n9554 = n8823 & ~n9553;
  assign n9555 = ~pi0567 & ~n8823;
  assign n9556 = ~n9554 & ~n9555;
  assign n9557 = n8810 & ~n9556;
  assign n9558 = ~pi0567 & ~n8810;
  assign po0618 = n9557 | n9558;
  assign n9560 = n8823 & ~n9525;
  assign n9561 = ~pi0568 & ~n8823;
  assign n9562 = ~n9560 & ~n9561;
  assign n9563 = n8810 & ~n9562;
  assign n9564 = ~pi0568 & ~n8810;
  assign po0619 = n9563 | n9564;
  assign n9566 = ~pi0569 & ~n7566;
  assign n9567 = n7566 & ~n8720;
  assign n9568 = ~n9566 & ~n9567;
  assign n9569 = n7544 & ~n9568;
  assign n9570 = ~pi0569 & ~n7544;
  assign po0620 = n9569 | n9570;
  assign n9572 = ~pi0570 & ~n7566;
  assign n9573 = n7566 & ~n7892;
  assign n9574 = ~n9572 & ~n9573;
  assign n9575 = n7544 & ~n9574;
  assign n9576 = ~pi0570 & ~n7544;
  assign po0621 = n9575 | n9576;
  assign n9578 = ~pi0571 & ~n7566;
  assign n9579 = pi0799 & n7453;
  assign n9580 = pi1935 & n7832;
  assign n9581 = ~n9579 & ~n9580;
  assign n9582 = pi1962 & n7548;
  assign n9583 = n9581 & ~n9582;
  assign n9584 = n7566 & ~n9583;
  assign n9585 = ~n9578 & ~n9584;
  assign n9586 = n7544 & ~n9585;
  assign n9587 = ~pi0571 & ~n7544;
  assign po0622 = n9586 | n9587;
  assign n9589 = ~pi0572 & ~n7566;
  assign n9590 = pi0800 & n7453;
  assign n9591 = pi1926 & n7832;
  assign n9592 = ~n9590 & ~n9591;
  assign n9593 = pi1978 & n7548;
  assign n9594 = n9592 & ~n9593;
  assign n9595 = n7566 & ~n9594;
  assign n9596 = ~n9589 & ~n9595;
  assign n9597 = n7544 & ~n9596;
  assign n9598 = ~pi0572 & ~n7544;
  assign po0623 = n9597 | n9598;
  assign n9600 = ~pi0573 & ~n7566;
  assign n9601 = pi0751 & n7453;
  assign n9602 = pi1901 & n7832;
  assign n9603 = ~n9601 & ~n9602;
  assign n9604 = pi1935 & n7548;
  assign n9605 = n9603 & ~n9604;
  assign n9606 = n7566 & ~n9605;
  assign n9607 = ~n9600 & ~n9606;
  assign n9608 = n7544 & ~n9607;
  assign n9609 = ~pi0573 & ~n7544;
  assign po0624 = n9608 | n9609;
  assign n9611 = ~pi0574 & ~n7566;
  assign n9612 = n7566 & ~n7931;
  assign n9613 = ~n9611 & ~n9612;
  assign n9614 = n7544 & ~n9613;
  assign n9615 = ~pi0574 & ~n7544;
  assign po0625 = n9614 | n9615;
  assign n9617 = ~pi0575 & ~n7566;
  assign n9618 = n7566 & ~n7836;
  assign n9619 = ~n9617 & ~n9618;
  assign n9620 = n7544 & ~n9619;
  assign n9621 = ~pi0575 & ~n7544;
  assign po0626 = n9620 | n9621;
  assign n9623 = ~pi0576 & ~n7566;
  assign n9624 = n7566 & ~n7909;
  assign n9625 = ~n9623 & ~n9624;
  assign n9626 = n7544 & ~n9625;
  assign n9627 = ~pi0576 & ~n7544;
  assign po0627 = n9626 | n9627;
  assign n9629 = ~pi0577 & ~n7566;
  assign n9630 = n7566 & ~n9469;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = n7544 & ~n9631;
  assign n9633 = ~pi0577 & ~n7544;
  assign po0628 = n9632 | n9633;
  assign n9635 = ~pi0578 & ~n7663;
  assign n9636 = n7663 & ~n8675;
  assign n9637 = ~n9635 & ~n9636;
  assign n9638 = n7544 & ~n9637;
  assign n9639 = ~pi0578 & ~n7544;
  assign po0629 = n9638 | n9639;
  assign n9641 = ~pi0579 & ~n7663;
  assign n9642 = n7663 & ~n8686;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = n7544 & ~n9643;
  assign n9645 = ~pi0579 & ~n7544;
  assign po0630 = n9644 | n9645;
  assign n9647 = ~pi0580 & ~n7663;
  assign n9648 = n7663 & ~n8697;
  assign n9649 = ~n9647 & ~n9648;
  assign n9650 = n7544 & ~n9649;
  assign n9651 = ~pi0580 & ~n7544;
  assign po0631 = n9650 | n9651;
  assign n9653 = ~pi0581 & ~n7663;
  assign n9654 = n7663 & ~n7859;
  assign n9655 = ~n9653 & ~n9654;
  assign n9656 = n7544 & ~n9655;
  assign n9657 = ~pi0581 & ~n7544;
  assign po0632 = n9656 | n9657;
  assign n9659 = ~pi0582 & ~n7663;
  assign n9660 = n7663 & ~n8720;
  assign n9661 = ~n9659 & ~n9660;
  assign n9662 = n7544 & ~n9661;
  assign n9663 = ~pi0582 & ~n7544;
  assign po0633 = n9662 | n9663;
  assign n9665 = ~pi0583 & ~n7663;
  assign n9666 = n7663 & ~n8731;
  assign n9667 = ~n9665 & ~n9666;
  assign n9668 = n7544 & ~n9667;
  assign n9669 = ~pi0583 & ~n7544;
  assign po0634 = n9668 | n9669;
  assign n9671 = ~pi0584 & ~n7663;
  assign n9672 = n7663 & ~n7870;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = n7544 & ~n9673;
  assign n9675 = ~pi0584 & ~n7544;
  assign po0635 = n9674 | n9675;
  assign n9677 = ~pi0585 & ~n7566;
  assign n9678 = n7566 & ~n7881;
  assign n9679 = ~n9677 & ~n9678;
  assign n9680 = n7544 & ~n9679;
  assign n9681 = ~pi0585 & ~n7544;
  assign po0636 = n9680 | n9681;
  assign n9683 = ~pi0586 & ~n7663;
  assign n9684 = n7663 & ~n7848;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = n7544 & ~n9685;
  assign n9687 = ~pi0586 & ~n7544;
  assign po0637 = n9686 | n9687;
  assign n9689 = ~pi0587 & ~n7663;
  assign n9690 = n7663 & ~n9583;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = n7544 & ~n9691;
  assign n9693 = ~pi0587 & ~n7544;
  assign po0638 = n9692 | n9693;
  assign n9695 = ~pi0588 & ~n7663;
  assign n9696 = n7663 & ~n9594;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = n7544 & ~n9697;
  assign n9699 = ~pi0588 & ~n7544;
  assign po0639 = n9698 | n9699;
  assign n9701 = ~pi0589 & ~n7663;
  assign n9702 = n7663 & ~n7942;
  assign n9703 = ~n9701 & ~n9702;
  assign n9704 = n7544 & ~n9703;
  assign n9705 = ~pi0589 & ~n7544;
  assign po0640 = n9704 | n9705;
  assign n9707 = ~pi0590 & ~n7663;
  assign n9708 = n7663 & ~n9605;
  assign n9709 = ~n9707 & ~n9708;
  assign n9710 = n7544 & ~n9709;
  assign n9711 = ~pi0590 & ~n7544;
  assign po0641 = n9710 | n9711;
  assign n9713 = ~pi0591 & ~n7663;
  assign n9714 = n7663 & ~n7931;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = n7544 & ~n9715;
  assign n9717 = ~pi0591 & ~n7544;
  assign po0642 = n9716 | n9717;
  assign n9719 = ~pi0592 & ~n7663;
  assign n9720 = n7663 & ~n9469;
  assign n9721 = ~n9719 & ~n9720;
  assign n9722 = n7544 & ~n9721;
  assign n9723 = ~pi0592 & ~n7544;
  assign po0643 = n9722 | n9723;
  assign n9725 = n7454 & ~n8697;
  assign n9726 = ~pi0593 & ~n7454;
  assign n9727 = ~n9725 & ~n9726;
  assign n9728 = n7544 & ~n9727;
  assign n9729 = ~pi0593 & ~n7544;
  assign po0644 = n9728 | n9729;
  assign n9731 = n7454 & ~n7848;
  assign n9732 = ~pi0594 & ~n7454;
  assign n9733 = ~n9731 & ~n9732;
  assign n9734 = n7544 & ~n9733;
  assign n9735 = ~pi0594 & ~n7544;
  assign po0645 = n9734 | n9735;
  assign n9737 = n7454 & ~n8731;
  assign n9738 = ~pi0595 & ~n7454;
  assign n9739 = ~n9737 & ~n9738;
  assign n9740 = n7544 & ~n9739;
  assign n9741 = ~pi0595 & ~n7544;
  assign po0646 = n9740 | n9741;
  assign n9743 = n7454 & ~n8686;
  assign n9744 = ~pi0596 & ~n7454;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = n7544 & ~n9745;
  assign n9747 = ~pi0596 & ~n7544;
  assign po0647 = n9746 | n9747;
  assign n9749 = n7454 & ~n9583;
  assign n9750 = ~pi0597 & ~n7454;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = n7544 & ~n9751;
  assign n9753 = ~pi0597 & ~n7544;
  assign po0648 = n9752 | n9753;
  assign n9755 = n7454 & ~n9594;
  assign n9756 = ~pi0598 & ~n7454;
  assign n9757 = ~n9755 & ~n9756;
  assign n9758 = n7544 & ~n9757;
  assign n9759 = ~pi0598 & ~n7544;
  assign po0649 = n9758 | n9759;
  assign n9761 = n7454 & ~n9605;
  assign n9762 = ~pi0599 & ~n7454;
  assign n9763 = ~n9761 & ~n9762;
  assign n9764 = n7544 & ~n9763;
  assign n9765 = ~pi0599 & ~n7544;
  assign po0650 = n9764 | n9765;
  assign n9767 = n7454 & ~n7892;
  assign n9768 = ~pi0600 & ~n7454;
  assign n9769 = ~n9767 & ~n9768;
  assign n9770 = n7544 & ~n9769;
  assign n9771 = ~pi0600 & ~n7544;
  assign po0651 = n9770 | n9771;
  assign n9773 = pi0601 & ~n8809;
  assign n9774 = ~pi0601 & pi0790;
  assign n9775 = pi0601 & ~pi0790;
  assign n9776 = ~n9774 & ~n9775;
  assign n9777 = n8806 & ~n9776;
  assign n9778 = ~pi0601 & ~n8806;
  assign n9779 = ~n9777 & ~n9778;
  assign n9780 = n8809 & ~n9779;
  assign n9781 = ~n9773 & ~n9780;
  assign po0652 = pi1036 & ~n9781;
  assign n9783 = pi0602 & ~n8809;
  assign n9784 = ~n8922 & ~n8946;
  assign n9785 = ~n8806 & ~n9784;
  assign n9786 = ~pi0602 & n8862;
  assign n9787 = pi0602 & ~n8862;
  assign n9788 = ~n9786 & ~n9787;
  assign n9789 = n8806 & ~n9788;
  assign n9790 = ~n9785 & ~n9789;
  assign n9791 = n8809 & ~n9790;
  assign n9792 = ~n9783 & ~n9791;
  assign po0653 = pi1036 & ~n9792;
  assign n9794 = ~pi0603 & ~n8812;
  assign n9795 = n8812 & ~n9553;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = n8810 & ~n9796;
  assign n9798 = ~pi0603 & ~n8810;
  assign po0654 = n9797 | n9798;
  assign n9800 = ~pi0604 & ~n7546;
  assign n9801 = n7546 & ~n7931;
  assign n9802 = ~n9800 & ~n9801;
  assign n9803 = n7544 & ~n9802;
  assign n9804 = ~pi0604 & ~n7544;
  assign po0655 = n9803 | n9804;
  assign n9806 = ~pi0605 & ~n8812;
  assign n9807 = pi0813 & n8806;
  assign n9808 = pi0235 & n8949;
  assign n9809 = ~n9807 & ~n9808;
  assign n9810 = pi0479 & n8814;
  assign n9811 = n9809 & ~n9810;
  assign n9812 = n8812 & ~n9811;
  assign n9813 = ~n9806 & ~n9812;
  assign n9814 = n8810 & ~n9813;
  assign n9815 = ~pi0605 & ~n8810;
  assign po0656 = n9814 | n9815;
  assign n9817 = ~pi0606 & ~n8812;
  assign n9818 = pi0835 & n8806;
  assign n9819 = pi0334 & n8949;
  assign n9820 = ~n9818 & ~n9819;
  assign n9821 = pi0819 & n8814;
  assign n9822 = n9820 & ~n9821;
  assign n9823 = n8812 & ~n9822;
  assign n9824 = ~n9817 & ~n9823;
  assign n9825 = n8810 & ~n9824;
  assign n9826 = ~pi0606 & ~n8810;
  assign po0657 = n9825 | n9826;
  assign n9828 = ~pi0607 & ~n7546;
  assign n9829 = n7546 & ~n7870;
  assign n9830 = ~n9828 & ~n9829;
  assign n9831 = n7544 & ~n9830;
  assign n9832 = ~pi0607 & ~n7544;
  assign po0658 = n9831 | n9832;
  assign n9834 = n7546 & n7580;
  assign n9835 = ~pi0608 & ~n7546;
  assign n9836 = ~n9834 & ~n9835;
  assign n9837 = n7544 & ~n9836;
  assign n9838 = ~pi0608 & ~n7544;
  assign po0659 = n9837 | n9838;
  assign n9840 = n7546 & n7587;
  assign n9841 = ~pi0609 & ~n7546;
  assign n9842 = ~n9840 & ~n9841;
  assign n9843 = n7544 & ~n9842;
  assign n9844 = ~pi0609 & ~n7544;
  assign po0660 = n9843 | n9844;
  assign n9846 = n7546 & n7594;
  assign n9847 = ~pi0610 & ~n7546;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = n7544 & ~n9848;
  assign n9850 = ~pi0610 & ~n7544;
  assign po0661 = n9849 | n9850;
  assign n9852 = n7546 & n7601;
  assign n9853 = ~pi0611 & ~n7546;
  assign n9854 = ~n9852 & ~n9853;
  assign n9855 = n7544 & ~n9854;
  assign n9856 = ~pi0611 & ~n7544;
  assign po0662 = n9855 | n9856;
  assign n9858 = n7546 & n7608;
  assign n9859 = ~pi0612 & ~n7546;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = n7544 & ~n9860;
  assign n9862 = ~pi0612 & ~n7544;
  assign po0663 = n9861 | n9862;
  assign n9864 = n7546 & n7615;
  assign n9865 = ~pi0613 & ~n7546;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = n7544 & ~n9866;
  assign n9868 = ~pi0613 & ~n7544;
  assign po0664 = n9867 | n9868;
  assign n9870 = n8812 & n9007;
  assign n9871 = ~pi0614 & ~n8812;
  assign n9872 = ~n9870 & ~n9871;
  assign n9873 = n8810 & ~n9872;
  assign n9874 = ~pi0614 & ~n8810;
  assign po0665 = n9873 | n9874;
  assign n9876 = n7546 & n7622;
  assign n9877 = ~pi0615 & ~n7546;
  assign n9878 = ~n9876 & ~n9877;
  assign n9879 = n7544 & ~n9878;
  assign n9880 = ~pi0615 & ~n7544;
  assign po0666 = n9879 | n9880;
  assign n9882 = n7546 & n7629;
  assign n9883 = ~pi0616 & ~n7546;
  assign n9884 = ~n9882 & ~n9883;
  assign n9885 = n7544 & ~n9884;
  assign n9886 = ~pi0616 & ~n7544;
  assign po0667 = n9885 | n9886;
  assign n9888 = n8812 & n9014;
  assign n9889 = ~pi0617 & ~n8812;
  assign n9890 = ~n9888 & ~n9889;
  assign n9891 = n8810 & ~n9890;
  assign n9892 = ~pi0617 & ~n8810;
  assign po0668 = n9891 | n9892;
  assign n9894 = n7546 & n7636;
  assign n9895 = ~pi0618 & ~n7546;
  assign n9896 = ~n9894 & ~n9895;
  assign n9897 = n7544 & ~n9896;
  assign n9898 = ~pi0618 & ~n7544;
  assign po0669 = n9897 | n9898;
  assign n9900 = n7546 & n7643;
  assign n9901 = ~pi0619 & ~n7546;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = n7544 & ~n9902;
  assign n9904 = ~pi0619 & ~n7544;
  assign po0670 = n9903 | n9904;
  assign n9906 = ~pi0620 & ~n7546;
  assign n9907 = n7546 & ~n9583;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = n7544 & ~n9908;
  assign n9910 = ~pi0620 & ~n7544;
  assign po0671 = n9909 | n9910;
  assign n9912 = n7546 & n7650;
  assign n9913 = ~pi0621 & ~n7546;
  assign n9914 = ~n9912 & ~n9913;
  assign n9915 = n7544 & ~n9914;
  assign n9916 = ~pi0621 & ~n7544;
  assign po0672 = n9915 | n9916;
  assign n9918 = n7546 & n7657;
  assign n9919 = ~pi0622 & ~n7546;
  assign n9920 = ~n9918 & ~n9919;
  assign n9921 = n7544 & ~n9920;
  assign n9922 = ~pi0622 & ~n7544;
  assign po0673 = n9921 | n9922;
  assign n9924 = ~pi0623 & ~n7546;
  assign n9925 = n7546 & ~n9594;
  assign n9926 = ~n9924 & ~n9925;
  assign n9927 = n7544 & ~n9926;
  assign n9928 = ~pi0623 & ~n7544;
  assign po0674 = n9927 | n9928;
  assign n9930 = n8812 & n9048;
  assign n9931 = ~pi0624 & ~n8812;
  assign n9932 = ~n9930 & ~n9931;
  assign n9933 = n8810 & ~n9932;
  assign n9934 = ~pi0624 & ~n8810;
  assign po0675 = n9933 | n9934;
  assign n9936 = ~pi0625 & ~n7546;
  assign n9937 = n7546 & ~n9605;
  assign n9938 = ~n9936 & ~n9937;
  assign n9939 = n7544 & ~n9938;
  assign n9940 = ~pi0625 & ~n7544;
  assign po0676 = n9939 | n9940;
  assign n9942 = n8812 & n9055;
  assign n9943 = ~pi0626 & ~n8812;
  assign n9944 = ~n9942 & ~n9943;
  assign n9945 = n8810 & ~n9944;
  assign n9946 = ~pi0626 & ~n8810;
  assign po0677 = n9945 | n9946;
  assign n9948 = n8812 & n9062;
  assign n9949 = ~pi0627 & ~n8812;
  assign n9950 = ~n9948 & ~n9949;
  assign n9951 = n8810 & ~n9950;
  assign n9952 = ~pi0627 & ~n8810;
  assign po0678 = n9951 | n9952;
  assign n9954 = ~pi0628 & ~n7546;
  assign n9955 = n7546 & ~n7942;
  assign n9956 = ~n9954 & ~n9955;
  assign n9957 = n7544 & ~n9956;
  assign n9958 = ~pi0628 & ~n7544;
  assign po0679 = n9957 | n9958;
  assign n9960 = n8812 & n8824;
  assign n9961 = ~pi0629 & ~n8812;
  assign n9962 = ~n9960 & ~n9961;
  assign n9963 = n8810 & ~n9962;
  assign n9964 = ~pi0629 & ~n8810;
  assign po0680 = n9963 | n9964;
  assign n9966 = ~pi0630 & ~n7546;
  assign n9967 = n7546 & ~n7836;
  assign n9968 = ~n9966 & ~n9967;
  assign n9969 = n7544 & ~n9968;
  assign n9970 = ~pi0630 & ~n7544;
  assign po0681 = n9969 | n9970;
  assign n9972 = ~pi0631 & ~n7546;
  assign n9973 = n7546 & ~n7909;
  assign n9974 = ~n9972 & ~n9973;
  assign n9975 = n7544 & ~n9974;
  assign n9976 = ~pi0631 & ~n7544;
  assign po0682 = n9975 | n9976;
  assign n9978 = n8812 & n9119;
  assign n9979 = ~pi0632 & ~n8812;
  assign n9980 = ~n9978 & ~n9979;
  assign n9981 = n8810 & ~n9980;
  assign n9982 = ~pi0632 & ~n8810;
  assign po0683 = n9981 | n9982;
  assign n9984 = ~pi0633 & ~n7546;
  assign n9985 = n7546 & ~n9469;
  assign n9986 = ~n9984 & ~n9985;
  assign n9987 = n7544 & ~n9986;
  assign n9988 = ~pi0633 & ~n7544;
  assign po0684 = n9987 | n9988;
  assign n9990 = ~pi0634 & ~n8812;
  assign n9991 = n8812 & ~n9492;
  assign n9992 = ~n9990 & ~n9991;
  assign n9993 = n8810 & ~n9992;
  assign n9994 = ~pi0634 & ~n8810;
  assign po0685 = n9993 | n9994;
  assign n9996 = pi0635 & pi1150;
  assign n9997 = ~n7451 & n9996;
  assign n9998 = pi0635 & ~n7453;
  assign n9999 = ~n7543 & ~n9998;
  assign n10000 = n7451 & ~n9999;
  assign n10001 = pi1150 & n10000;
  assign po0686 = n9997 | n10001;
  assign n10003 = pi2020 & n7451;
  assign po0687 = ~pi0636 | n10003;
  assign n10005 = ~pi0637 & ~n8812;
  assign n10006 = n8812 & ~n9481;
  assign n10007 = ~n10005 & ~n10006;
  assign n10008 = n8810 & ~n10007;
  assign n10009 = ~pi0637 & ~n8810;
  assign po0688 = n10008 | n10009;
  assign n10011 = ~pi0638 & ~n7546;
  assign n10012 = n7546 & ~n7881;
  assign n10013 = ~n10011 & ~n10012;
  assign n10014 = n7544 & ~n10013;
  assign n10015 = ~pi0638 & ~n7544;
  assign po0689 = n10014 | n10015;
  assign n10017 = pi0192 & n8949;
  assign n10018 = pi0207 & n8814;
  assign n10019 = ~n10017 & ~n10018;
  assign n10020 = pi1924 & n8806;
  assign n10021 = n10019 & ~n10020;
  assign n10022 = n8823 & ~n10021;
  assign n10023 = ~pi0639 & ~n8823;
  assign n10024 = ~n10022 & ~n10023;
  assign n10025 = n8810 & ~n10024;
  assign n10026 = ~pi0639 & ~n8810;
  assign po0690 = n10025 | n10026;
  assign n10028 = ~pi0641 & ~n8812;
  assign n10029 = pi0820 & n8806;
  assign n10030 = pi0479 & n8949;
  assign n10031 = ~n10029 & ~n10030;
  assign n10032 = pi0866 & n8814;
  assign n10033 = n10031 & ~n10032;
  assign n10034 = n8812 & ~n10033;
  assign n10035 = ~n10028 & ~n10034;
  assign n10036 = n8810 & ~n10035;
  assign n10037 = ~pi0641 & ~n8810;
  assign po0692 = n10036 | n10037;
  assign n10039 = ~pi0642 & ~n9020;
  assign n10040 = pi1933 & n9022;
  assign n10041 = pi0857 & n8837;
  assign n10042 = ~n10040 & ~n10041;
  assign n10043 = pi1157 & ~pi1158;
  assign n10044 = pi1883 & n10043;
  assign n10045 = n10042 & ~n10044;
  assign n10046 = n9020 & ~n10045;
  assign n10047 = ~n10039 & ~n10046;
  assign n10048 = n8841 & ~n10047;
  assign n10049 = ~pi0642 & ~n8841;
  assign po0693 = n10048 | n10049;
  assign n10051 = pi0643 & ~n8840;
  assign n10052 = pi0643 & n8843;
  assign n10053 = ~pi0643 & ~n8843;
  assign n10054 = ~n10052 & ~n10053;
  assign n10055 = ~n8837 & n10054;
  assign n10056 = pi0821 & pi0843;
  assign n10057 = pi0746 & n10056;
  assign n10058 = pi0643 & ~n10057;
  assign n10059 = ~pi0643 & n10057;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = n8837 & ~n10060;
  assign n10062 = ~n10055 & ~n10061;
  assign n10063 = n8840 & ~n10062;
  assign n10064 = ~n10051 & ~n10063;
  assign po0694 = pi1145 & ~n10064;
  assign n10066 = ~pi0644 & ~n9020;
  assign n10067 = pi0883 & n10043;
  assign n10068 = pi0951 & n9022;
  assign n10069 = ~n10067 & ~n10068;
  assign n10070 = pi0858 & n8837;
  assign n10071 = n10069 & ~n10070;
  assign n10072 = n9020 & ~n10071;
  assign n10073 = ~n10066 & ~n10072;
  assign n10074 = n8841 & ~n10073;
  assign n10075 = ~pi0644 & ~n8841;
  assign po0695 = n10074 | n10075;
  assign n10077 = ~pi0645 & ~n8946;
  assign n10078 = pi0828 & n8806;
  assign n10079 = pi0882 & n8949;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = pi0950 & n8814;
  assign n10082 = n10080 & ~n10081;
  assign n10083 = n8946 & ~n10082;
  assign n10084 = ~n10077 & ~n10083;
  assign n10085 = n8810 & ~n10084;
  assign n10086 = ~pi0645 & ~n8810;
  assign po0696 = n10085 | n10086;
  assign n10088 = ~pi0646 & ~n9020;
  assign n10089 = pi1958 & n9022;
  assign n10090 = pi0854 & n8837;
  assign n10091 = ~n10089 & ~n10090;
  assign n10092 = pi1933 & n10043;
  assign n10093 = n10091 & ~n10092;
  assign n10094 = n9020 & ~n10093;
  assign n10095 = ~n10088 & ~n10094;
  assign n10096 = n8841 & ~n10095;
  assign n10097 = ~pi0646 & ~n8841;
  assign po0697 = n10096 | n10097;
  assign n10099 = n8851 & n9020;
  assign n10100 = ~pi0647 & ~n9020;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = n8841 & ~n10101;
  assign n10103 = ~pi0647 & ~n8841;
  assign po0698 = n10102 | n10103;
  assign n10105 = ~pi0648 & ~n8946;
  assign n10106 = n8946 & ~n9503;
  assign n10107 = ~n10105 & ~n10106;
  assign n10108 = n8810 & ~n10107;
  assign n10109 = ~pi0648 & ~n8810;
  assign po0699 = n10108 | n10109;
  assign n10111 = ~pi0649 & ~n9020;
  assign n10112 = pi0206 & n9022;
  assign n10113 = pi0191 & n10043;
  assign n10114 = ~n10112 & ~n10113;
  assign n10115 = pi1925 & n8837;
  assign n10116 = n10114 & ~n10115;
  assign n10117 = n9020 & ~n10116;
  assign n10118 = ~n10111 & ~n10117;
  assign n10119 = n8841 & ~n10118;
  assign n10120 = ~pi0649 & ~n8841;
  assign po0700 = n10119 | n10120;
  assign n10122 = ~pi0650 & ~n9020;
  assign n10123 = pi0851 & n8837;
  assign n10124 = pi0481 & n9022;
  assign n10125 = ~n10123 & ~n10124;
  assign n10126 = pi0231 & n10043;
  assign n10127 = n10125 & ~n10126;
  assign n10128 = n9020 & ~n10127;
  assign n10129 = ~n10122 & ~n10128;
  assign n10130 = n8841 & ~n10129;
  assign n10131 = ~pi0650 & ~n8841;
  assign po0701 = n10130 | n10131;
  assign n10133 = ~pi0651 & ~n8946;
  assign n10134 = n8946 & ~n9481;
  assign n10135 = ~n10133 & ~n10134;
  assign n10136 = n8810 & ~n10135;
  assign n10137 = ~pi0651 & ~n8810;
  assign po0702 = n10136 | n10137;
  assign n10139 = ~pi0652 & ~n8946;
  assign n10140 = pi0833 & n8806;
  assign n10141 = pi0207 & n8949;
  assign n10142 = ~n10140 & ~n10141;
  assign n10143 = pi0235 & n8814;
  assign n10144 = n10142 & ~n10143;
  assign n10145 = n8946 & ~n10144;
  assign n10146 = ~n10139 & ~n10145;
  assign n10147 = n8810 & ~n10146;
  assign n10148 = ~pi0652 & ~n8810;
  assign po0703 = n10147 | n10148;
  assign n10150 = ~pi0653 & ~n8946;
  assign n10151 = n8946 & ~n9811;
  assign n10152 = ~n10150 & ~n10151;
  assign n10153 = n8810 & ~n10152;
  assign n10154 = ~pi0653 & ~n8810;
  assign po0704 = n10153 | n10154;
  assign n10156 = ~pi0654 & ~n8946;
  assign n10157 = pi0832 & n8806;
  assign n10158 = pi0819 & n8949;
  assign n10159 = ~n10157 & ~n10158;
  assign n10160 = pi0882 & n8814;
  assign n10161 = n10159 & ~n10160;
  assign n10162 = n8946 & ~n10161;
  assign n10163 = ~n10156 & ~n10162;
  assign n10164 = n8810 & ~n10163;
  assign n10165 = ~pi0654 & ~n8810;
  assign po0705 = n10164 | n10165;
  assign n10167 = n8823 & ~n10082;
  assign n10168 = ~pi0655 & ~n8823;
  assign n10169 = ~n10167 & ~n10168;
  assign n10170 = n8810 & ~n10169;
  assign n10171 = ~pi0655 & ~n8810;
  assign po0706 = n10170 | n10171;
  assign n10173 = n8812 & n9041;
  assign n10174 = ~pi0656 & ~n8812;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = n8810 & ~n10175;
  assign n10177 = ~pi0656 & ~n8810;
  assign po0707 = n10176 | n10177;
  assign n10179 = ~pi0635 & n7451;
  assign n10180 = pi0657 & ~n10179;
  assign n10181 = pi0814 & n10179;
  assign po0708 = n10180 | n10181;
  assign n10183 = ~pi0658 & ~n8880;
  assign n10184 = pi0850 & n8837;
  assign n10185 = pi0818 & n9022;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = pi0333 & n10043;
  assign n10188 = n10186 & ~n10187;
  assign n10189 = n8880 & ~n10188;
  assign n10190 = ~n10183 & ~n10189;
  assign n10191 = n8841 & ~n10190;
  assign n10192 = ~pi0658 & ~n8841;
  assign po0709 = n10191 | n10192;
  assign n10194 = n8823 & ~n9811;
  assign n10195 = ~pi0659 & ~n8823;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = n8810 & ~n10196;
  assign n10198 = ~pi0659 & ~n8810;
  assign po0710 = n10197 | n10198;
  assign n10200 = n8823 & ~n8953;
  assign n10201 = ~pi0660 & ~n8823;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = n8810 & ~n10202;
  assign n10204 = ~pi0660 & ~n8810;
  assign po0711 = n10203 | n10204;
  assign n10206 = n8843 & ~n10045;
  assign n10207 = ~pi0661 & ~n8843;
  assign n10208 = ~n10206 & ~n10207;
  assign n10209 = n8841 & ~n10208;
  assign n10210 = ~pi0661 & ~n8841;
  assign po0712 = n10209 | n10210;
  assign n10212 = pi1959 & n9022;
  assign n10213 = pi0853 & n8837;
  assign n10214 = ~n10212 & ~n10213;
  assign n10215 = pi1981 & n10043;
  assign n10216 = n10214 & ~n10215;
  assign n10217 = n8843 & ~n10216;
  assign n10218 = ~pi0662 & ~n8843;
  assign n10219 = ~n10217 & ~n10218;
  assign n10220 = n8841 & ~n10219;
  assign n10221 = ~pi0662 & ~n8841;
  assign po0713 = n10220 | n10221;
  assign n10223 = pi0852 & n8837;
  assign n10224 = pi0231 & n9022;
  assign n10225 = ~n10223 & ~n10224;
  assign n10226 = pi0206 & n10043;
  assign n10227 = n10225 & ~n10226;
  assign n10228 = n8843 & ~n10227;
  assign n10229 = ~pi0663 & ~n8843;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = n8841 & ~n10230;
  assign n10232 = ~pi0663 & ~n8841;
  assign po0714 = n10231 | n10232;
  assign n10234 = ~pi0664 & ~n8880;
  assign n10235 = pi1925 & n9022;
  assign n10236 = pi0855 & n8837;
  assign n10237 = ~n10235 & ~n10236;
  assign n10238 = pi1853 & n10043;
  assign n10239 = n10237 & ~n10238;
  assign n10240 = n8880 & ~n10239;
  assign n10241 = ~n10234 & ~n10240;
  assign n10242 = n8841 & ~n10241;
  assign n10243 = ~pi0664 & ~n8841;
  assign po0715 = n10242 | n10243;
  assign n10245 = ~pi0665 & ~n8880;
  assign n10246 = n8880 & ~n10093;
  assign n10247 = ~n10245 & ~n10246;
  assign n10248 = n8841 & ~n10247;
  assign n10249 = ~pi0665 & ~n8841;
  assign po0716 = n10248 | n10249;
  assign n10251 = ~pi0666 & ~n8946;
  assign n10252 = n8946 & ~n9525;
  assign n10253 = ~n10251 & ~n10252;
  assign n10254 = n8810 & ~n10253;
  assign n10255 = ~pi0666 & ~n8810;
  assign po0717 = n10254 | n10255;
  assign n10257 = ~pi0667 & ~n8922;
  assign n10258 = n8922 & ~n8953;
  assign n10259 = ~n10257 & ~n10258;
  assign n10260 = n8810 & ~n10259;
  assign n10261 = ~pi0667 & ~n8810;
  assign po0718 = n10260 | n10261;
  assign n10263 = ~pi0668 & ~n8922;
  assign n10264 = n8922 & ~n10033;
  assign n10265 = ~n10263 & ~n10264;
  assign n10266 = n8810 & ~n10265;
  assign n10267 = ~pi0668 & ~n8810;
  assign po0719 = n10266 | n10267;
  assign n10269 = ~pi0669 & ~n8922;
  assign n10270 = n8922 & ~n9822;
  assign n10271 = ~n10269 & ~n10270;
  assign n10272 = n8810 & ~n10271;
  assign n10273 = ~pi0669 & ~n8810;
  assign po0720 = n10272 | n10273;
  assign n10275 = ~pi0670 & ~n8922;
  assign n10276 = n8922 & ~n9811;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = n8810 & ~n10277;
  assign n10279 = ~pi0670 & ~n8810;
  assign po0721 = n10278 | n10279;
  assign n10281 = ~pi0671 & ~n8922;
  assign n10282 = pi0834 & n8806;
  assign n10283 = pi0212 & n8949;
  assign n10284 = ~n10282 & ~n10283;
  assign n10285 = pi0334 & n8814;
  assign n10286 = n10284 & ~n10285;
  assign n10287 = n8922 & ~n10286;
  assign n10288 = ~n10281 & ~n10287;
  assign n10289 = n8810 & ~n10288;
  assign n10290 = ~pi0671 & ~n8810;
  assign po0722 = n10289 | n10290;
  assign n10292 = ~pi0672 & ~n8922;
  assign n10293 = n8922 & ~n10144;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = n8810 & ~n10294;
  assign n10296 = ~pi0672 & ~n8810;
  assign po0723 = n10295 | n10296;
  assign n10298 = ~pi0673 & ~n8922;
  assign n10299 = pi0196 & n8949;
  assign n10300 = pi0212 & n8814;
  assign n10301 = ~n10299 & ~n10300;
  assign n10302 = pi1934 & n8806;
  assign n10303 = n10301 & ~n10302;
  assign n10304 = n8922 & ~n10303;
  assign n10305 = ~n10298 & ~n10304;
  assign n10306 = n8810 & ~n10305;
  assign n10307 = ~pi0673 & ~n8810;
  assign po0724 = n10306 | n10307;
  assign n10309 = ~pi0674 & ~n8922;
  assign n10310 = n8922 & ~n10161;
  assign n10311 = ~n10309 & ~n10310;
  assign n10312 = n8810 & ~n10311;
  assign n10313 = ~pi0674 & ~n8810;
  assign po0725 = n10312 | n10313;
  assign n10315 = ~pi0675 & ~n8902;
  assign n10316 = pi1947 & n9022;
  assign n10317 = pi0848 & n8837;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = pi1958 & n10043;
  assign n10320 = n10318 & ~n10319;
  assign n10321 = n8902 & ~n10320;
  assign n10322 = ~n10315 & ~n10321;
  assign n10323 = n8841 & ~n10322;
  assign n10324 = ~pi0675 & ~n8841;
  assign po0726 = n10323 | n10324;
  assign n10326 = ~pi0676 & ~n8902;
  assign n10327 = pi0846 & n8837;
  assign n10328 = pi0818 & n10043;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = pi0883 & n9022;
  assign n10331 = n10329 & ~n10330;
  assign n10332 = n8902 & ~n10331;
  assign n10333 = ~n10326 & ~n10332;
  assign n10334 = n8841 & ~n10333;
  assign n10335 = ~pi0676 & ~n8841;
  assign po0727 = n10334 | n10335;
  assign n10337 = ~pi0677 & ~n8902;
  assign n10338 = n8902 & ~n10188;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = n8841 & ~n10339;
  assign n10341 = ~pi0677 & ~n8841;
  assign po0728 = n10340 | n10341;
  assign n10343 = ~pi0678 & ~n8902;
  assign n10344 = n8902 & ~n10127;
  assign n10345 = ~n10343 & ~n10344;
  assign n10346 = n8841 & ~n10345;
  assign n10347 = ~pi0678 & ~n8841;
  assign po0729 = n10346 | n10347;
  assign n10349 = ~pi0679 & ~n8902;
  assign n10350 = pi0847 & n8837;
  assign n10351 = pi0333 & n9022;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = pi0211 & n10043;
  assign n10354 = n10352 & ~n10353;
  assign n10355 = n8902 & ~n10354;
  assign n10356 = ~n10349 & ~n10355;
  assign n10357 = n8841 & ~n10356;
  assign n10358 = ~pi0679 & ~n8841;
  assign po0730 = n10357 | n10358;
  assign n10360 = ~pi0680 & ~n8902;
  assign n10361 = pi0211 & n9022;
  assign n10362 = pi0195 & n10043;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = pi1933 & n8837;
  assign n10365 = n10363 & ~n10364;
  assign n10366 = n8902 & ~n10365;
  assign n10367 = ~n10360 & ~n10366;
  assign n10368 = n8841 & ~n10367;
  assign n10369 = ~pi0680 & ~n8841;
  assign po0731 = n10368 | n10369;
  assign n10371 = ~pi0681 & ~n8902;
  assign n10372 = n8902 & ~n10116;
  assign n10373 = ~n10371 & ~n10372;
  assign n10374 = n8841 & ~n10373;
  assign n10375 = ~pi0681 & ~n8841;
  assign po0732 = n10374 | n10375;
  assign n10377 = ~pi0682 & ~n8902;
  assign n10378 = n8902 & ~n10216;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = n8841 & ~n10379;
  assign n10381 = ~pi0682 & ~n8841;
  assign po0733 = n10380 | n10381;
  assign n10383 = ~pi0683 & ~n8902;
  assign n10384 = n8902 & ~n10093;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = n8841 & ~n10385;
  assign n10387 = ~pi0683 & ~n8841;
  assign po0734 = n10386 | n10387;
  assign n10389 = ~pi0684 & ~n8902;
  assign n10390 = pi1981 & n9022;
  assign n10391 = pi0845 & n8837;
  assign n10392 = ~n10390 & ~n10391;
  assign n10393 = pi1925 & n10043;
  assign n10394 = n10392 & ~n10393;
  assign n10395 = n8902 & ~n10394;
  assign n10396 = ~n10389 & ~n10395;
  assign n10397 = n8841 & ~n10396;
  assign n10398 = ~pi0684 & ~n8841;
  assign po0735 = n10397 | n10398;
  assign n10400 = ~pi0685 & ~n8902;
  assign n10401 = n8902 & ~n10045;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = n8841 & ~n10402;
  assign n10404 = ~pi0685 & ~n8841;
  assign po0736 = n10403 | n10404;
  assign n10406 = ~pi0686 & ~n8902;
  assign n10407 = n8902 & ~n10239;
  assign n10408 = ~n10406 & ~n10407;
  assign n10409 = n8841 & ~n10408;
  assign n10410 = ~pi0686 & ~n8841;
  assign po0737 = n10409 | n10410;
  assign n10412 = ~pi0687 & ~n8902;
  assign n10413 = pi1883 & n9022;
  assign n10414 = pi0856 & n8837;
  assign n10415 = ~n10413 & ~n10414;
  assign n10416 = pi0951 & n10043;
  assign n10417 = n10415 & ~n10416;
  assign n10418 = n8902 & ~n10417;
  assign n10419 = ~n10412 & ~n10418;
  assign n10420 = n8841 & ~n10419;
  assign n10421 = ~pi0687 & ~n8841;
  assign po0738 = n10420 | n10421;
  assign n10423 = ~pi0688 & ~n8902;
  assign n10424 = pi1853 & n9022;
  assign n10425 = pi0859 & n8837;
  assign n10426 = ~n10424 & ~n10425;
  assign n10427 = pi0916 & n10043;
  assign n10428 = n10426 & ~n10427;
  assign n10429 = n8902 & ~n10428;
  assign n10430 = ~n10423 & ~n10429;
  assign n10431 = n8841 & ~n10430;
  assign n10432 = ~pi0688 & ~n8841;
  assign po0739 = n10431 | n10432;
  assign n10434 = ~pi0689 & ~n8902;
  assign n10435 = n8902 & ~n10071;
  assign n10436 = ~n10434 & ~n10435;
  assign n10437 = n8841 & ~n10436;
  assign n10438 = ~pi0689 & ~n8841;
  assign po0740 = n10437 | n10438;
  assign n10440 = ~pi0690 & ~n8880;
  assign n10441 = n8880 & ~n10320;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = n8841 & ~n10442;
  assign n10444 = ~pi0690 & ~n8841;
  assign po0741 = n10443 | n10444;
  assign n10446 = ~pi0691 & ~n8880;
  assign n10447 = n8880 & ~n10331;
  assign n10448 = ~n10446 & ~n10447;
  assign n10449 = n8841 & ~n10448;
  assign n10450 = ~pi0691 & ~n8841;
  assign po0742 = n10449 | n10450;
  assign n10452 = ~pi0692 & ~n8880;
  assign n10453 = pi0849 & n8837;
  assign n10454 = pi0481 & n10043;
  assign n10455 = ~n10453 & ~n10454;
  assign n10456 = pi0870 & n9022;
  assign n10457 = n10455 & ~n10456;
  assign n10458 = n8880 & ~n10457;
  assign n10459 = ~n10452 & ~n10458;
  assign n10460 = n8841 & ~n10459;
  assign n10461 = ~pi0692 & ~n8841;
  assign po0743 = n10460 | n10461;
  assign n10463 = ~pi0693 & ~n8880;
  assign n10464 = n8880 & ~n10354;
  assign n10465 = ~n10463 & ~n10464;
  assign n10466 = n8841 & ~n10465;
  assign n10467 = ~pi0693 & ~n8841;
  assign po0744 = n10466 | n10467;
  assign n10469 = ~pi0694 & ~n8880;
  assign n10470 = n8880 & ~n10227;
  assign n10471 = ~n10469 & ~n10470;
  assign n10472 = n8841 & ~n10471;
  assign n10473 = ~pi0694 & ~n8841;
  assign po0745 = n10472 | n10473;
  assign n10475 = ~pi0695 & ~n8880;
  assign n10476 = n8880 & ~n10365;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = n8841 & ~n10477;
  assign n10479 = ~pi0695 & ~n8841;
  assign po0746 = n10478 | n10479;
  assign n10481 = ~pi0696 & ~n8880;
  assign n10482 = n8880 & ~n10116;
  assign n10483 = ~n10481 & ~n10482;
  assign n10484 = n8841 & ~n10483;
  assign n10485 = ~pi0696 & ~n8841;
  assign po0747 = n10484 | n10485;
  assign n10487 = ~pi0697 & ~n8880;
  assign n10488 = n8880 & ~n10216;
  assign n10489 = ~n10487 & ~n10488;
  assign n10490 = n8841 & ~n10489;
  assign n10491 = ~pi0697 & ~n8841;
  assign po0748 = n10490 | n10491;
  assign n10493 = ~pi0698 & ~n8922;
  assign n10494 = n8922 & ~n9513;
  assign n10495 = ~n10493 & ~n10494;
  assign n10496 = n8810 & ~n10495;
  assign n10497 = ~pi0698 & ~n8810;
  assign po0749 = n10496 | n10497;
  assign n10499 = ~pi0699 & ~n8880;
  assign n10500 = n8880 & ~n10394;
  assign n10501 = ~n10499 & ~n10500;
  assign n10502 = n8841 & ~n10501;
  assign n10503 = ~pi0699 & ~n8841;
  assign po0750 = n10502 | n10503;
  assign n10505 = ~pi0700 & ~n8922;
  assign n10506 = pi0826 & n8806;
  assign n10507 = pi1886 & n8949;
  assign n10508 = ~n10506 & ~n10507;
  assign n10509 = pi1934 & n8814;
  assign n10510 = n10508 & ~n10509;
  assign n10511 = n8922 & ~n10510;
  assign n10512 = ~n10505 & ~n10511;
  assign n10513 = n8810 & ~n10512;
  assign n10514 = ~pi0700 & ~n8810;
  assign po0751 = n10513 | n10514;
  assign n10516 = ~pi0701 & ~n8880;
  assign n10517 = n8880 & ~n10045;
  assign n10518 = ~n10516 & ~n10517;
  assign n10519 = n8841 & ~n10518;
  assign n10520 = ~pi0701 & ~n8841;
  assign po0752 = n10519 | n10520;
  assign n10522 = ~pi0702 & ~n8880;
  assign n10523 = n8880 & ~n10417;
  assign n10524 = ~n10522 & ~n10523;
  assign n10525 = n8841 & ~n10524;
  assign n10526 = ~pi0702 & ~n8841;
  assign po0753 = n10525 | n10526;
  assign n10528 = ~pi0703 & ~n8880;
  assign n10529 = n8880 & ~n10428;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = n8841 & ~n10530;
  assign n10532 = ~pi0703 & ~n8841;
  assign po0754 = n10531 | n10532;
  assign n10534 = ~pi0704 & ~n8880;
  assign n10535 = n8880 & ~n10071;
  assign n10536 = ~n10534 & ~n10535;
  assign n10537 = n8841 & ~n10536;
  assign n10538 = ~pi0704 & ~n8841;
  assign po0755 = n10537 | n10538;
  assign n10540 = n8843 & ~n10320;
  assign n10541 = ~pi0705 & ~n8843;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = n8841 & ~n10542;
  assign n10544 = ~pi0705 & ~n8841;
  assign po0756 = n10543 | n10544;
  assign n10546 = n8843 & ~n10331;
  assign n10547 = ~pi0706 & ~n8843;
  assign n10548 = ~n10546 & ~n10547;
  assign n10549 = n8841 & ~n10548;
  assign n10550 = ~pi0706 & ~n8841;
  assign po0757 = n10549 | n10550;
  assign n10552 = n8843 & ~n10457;
  assign n10553 = ~pi0707 & ~n8843;
  assign n10554 = ~n10552 & ~n10553;
  assign n10555 = n8841 & ~n10554;
  assign n10556 = ~pi0707 & ~n8841;
  assign po0758 = n10555 | n10556;
  assign n10558 = n8843 & ~n10188;
  assign n10559 = ~pi0708 & ~n8843;
  assign n10560 = ~n10558 & ~n10559;
  assign n10561 = n8841 & ~n10560;
  assign n10562 = ~pi0708 & ~n8841;
  assign po0759 = n10561 | n10562;
  assign n10564 = n8843 & ~n10127;
  assign n10565 = ~pi0709 & ~n8843;
  assign n10566 = ~n10564 & ~n10565;
  assign n10567 = n8841 & ~n10566;
  assign n10568 = ~pi0709 & ~n8841;
  assign po0760 = n10567 | n10568;
  assign n10570 = n8843 & ~n10354;
  assign n10571 = ~pi0710 & ~n8843;
  assign n10572 = ~n10570 & ~n10571;
  assign n10573 = n8841 & ~n10572;
  assign n10574 = ~pi0710 & ~n8841;
  assign po0761 = n10573 | n10574;
  assign n10576 = ~pi0711 & ~n8880;
  assign n10577 = n8880 & ~n10127;
  assign n10578 = ~n10576 & ~n10577;
  assign n10579 = n8841 & ~n10578;
  assign n10580 = ~pi0711 & ~n8841;
  assign po0762 = n10579 | n10580;
  assign n10582 = n8843 & ~n10365;
  assign n10583 = ~pi0712 & ~n8843;
  assign n10584 = ~n10582 & ~n10583;
  assign n10585 = n8841 & ~n10584;
  assign n10586 = ~pi0712 & ~n8841;
  assign po0763 = n10585 | n10586;
  assign n10588 = n8843 & ~n10116;
  assign n10589 = ~pi0713 & ~n8843;
  assign n10590 = ~n10588 & ~n10589;
  assign n10591 = n8841 & ~n10590;
  assign n10592 = ~pi0713 & ~n8841;
  assign po0764 = n10591 | n10592;
  assign n10594 = ~pi0714 & ~n8922;
  assign n10595 = pi0830 & n8806;
  assign n10596 = pi0915 & n8949;
  assign n10597 = ~n10595 & ~n10596;
  assign n10598 = pi1852 & n8814;
  assign n10599 = n10597 & ~n10598;
  assign n10600 = n8922 & ~n10599;
  assign n10601 = ~n10594 & ~n10600;
  assign n10602 = n8810 & ~n10601;
  assign n10603 = ~pi0714 & ~n8810;
  assign po0765 = n10602 | n10603;
  assign n10605 = n8843 & ~n10093;
  assign n10606 = ~pi0715 & ~n8843;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = n8841 & ~n10607;
  assign n10609 = ~pi0715 & ~n8841;
  assign po0766 = n10608 | n10609;
  assign n10611 = n8843 & ~n10394;
  assign n10612 = ~pi0716 & ~n8843;
  assign n10613 = ~n10611 & ~n10612;
  assign n10614 = n8841 & ~n10613;
  assign n10615 = ~pi0716 & ~n8841;
  assign po0767 = n10614 | n10615;
  assign n10617 = n8843 & ~n10239;
  assign n10618 = ~pi0717 & ~n8843;
  assign n10619 = ~n10617 & ~n10618;
  assign n10620 = n8841 & ~n10619;
  assign n10621 = ~pi0717 & ~n8841;
  assign po0768 = n10620 | n10621;
  assign n10623 = n8843 & ~n10417;
  assign n10624 = ~pi0718 & ~n8843;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = n8841 & ~n10625;
  assign n10627 = ~pi0718 & ~n8841;
  assign po0769 = n10626 | n10627;
  assign n10629 = n8843 & ~n10428;
  assign n10630 = ~pi0719 & ~n8843;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = n8841 & ~n10631;
  assign n10633 = ~pi0719 & ~n8841;
  assign po0770 = n10632 | n10633;
  assign n10635 = ~pi0720 & ~n8922;
  assign n10636 = n8922 & ~n10082;
  assign n10637 = ~n10635 & ~n10636;
  assign n10638 = n8810 & ~n10637;
  assign n10639 = ~pi0720 & ~n8810;
  assign po0771 = n10638 | n10639;
  assign n10641 = pi0870 & n10043;
  assign n10642 = pi0916 & n9022;
  assign n10643 = ~n10641 & ~n10642;
  assign n10644 = pi0844 & n8837;
  assign n10645 = n10643 & ~n10644;
  assign n10646 = n8843 & ~n10645;
  assign n10647 = ~pi0721 & ~n8843;
  assign n10648 = ~n10646 & ~n10647;
  assign n10649 = n8841 & ~n10648;
  assign n10650 = ~pi0721 & ~n8841;
  assign po0772 = n10649 | n10650;
  assign n10652 = n8843 & ~n10071;
  assign n10653 = ~pi0722 & ~n8843;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 = n8841 & ~n10654;
  assign n10656 = ~pi0722 & ~n8841;
  assign po0773 = n10655 | n10656;
  assign n10658 = n8823 & ~n10161;
  assign n10659 = ~pi0723 & ~n8823;
  assign n10660 = ~n10658 & ~n10659;
  assign n10661 = n8810 & ~n10660;
  assign n10662 = ~pi0723 & ~n8810;
  assign po0774 = n10661 | n10662;
  assign n10664 = n8823 & ~n10033;
  assign n10665 = ~pi0724 & ~n8823;
  assign n10666 = ~n10664 & ~n10665;
  assign n10667 = n8810 & ~n10666;
  assign n10668 = ~pi0724 & ~n8810;
  assign po0775 = n10667 | n10668;
  assign n10670 = n8823 & ~n9822;
  assign n10671 = ~pi0725 & ~n8823;
  assign n10672 = ~n10670 & ~n10671;
  assign n10673 = n8810 & ~n10672;
  assign n10674 = ~pi0725 & ~n8810;
  assign po0776 = n10673 | n10674;
  assign n10676 = n8823 & ~n10286;
  assign n10677 = ~pi0726 & ~n8823;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = n8810 & ~n10678;
  assign n10680 = ~pi0726 & ~n8810;
  assign po0777 = n10679 | n10680;
  assign n10682 = n8823 & ~n10144;
  assign n10683 = ~pi0727 & ~n8823;
  assign n10684 = ~n10682 & ~n10683;
  assign n10685 = n8810 & ~n10684;
  assign n10686 = ~pi0727 & ~n8810;
  assign po0778 = n10685 | n10686;
  assign n10688 = n8823 & ~n10303;
  assign n10689 = ~pi0728 & ~n8823;
  assign n10690 = ~n10688 & ~n10689;
  assign n10691 = n8810 & ~n10690;
  assign n10692 = ~pi0728 & ~n8810;
  assign po0779 = n10691 | n10692;
  assign n10694 = n8823 & ~n9481;
  assign n10695 = ~pi0729 & ~n8823;
  assign n10696 = ~n10694 & ~n10695;
  assign n10697 = n8810 & ~n10696;
  assign n10698 = ~pi0729 & ~n8810;
  assign po0780 = n10697 | n10698;
  assign n10700 = n8823 & ~n10510;
  assign n10701 = ~pi0730 & ~n8823;
  assign n10702 = ~n10700 & ~n10701;
  assign n10703 = n8810 & ~n10702;
  assign n10704 = ~pi0730 & ~n8810;
  assign po0781 = n10703 | n10704;
  assign n10706 = n8823 & ~n9492;
  assign n10707 = ~pi0731 & ~n8823;
  assign n10708 = ~n10706 & ~n10707;
  assign n10709 = n8810 & ~n10708;
  assign n10710 = ~pi0731 & ~n8810;
  assign po0782 = n10709 | n10710;
  assign n10712 = n8823 & ~n9503;
  assign n10713 = ~pi0732 & ~n8823;
  assign n10714 = ~n10712 & ~n10713;
  assign n10715 = n8810 & ~n10714;
  assign n10716 = ~pi0732 & ~n8810;
  assign po0783 = n10715 | n10716;
  assign n10718 = n8823 & ~n10599;
  assign n10719 = ~pi0733 & ~n8823;
  assign n10720 = ~n10718 & ~n10719;
  assign n10721 = n8810 & ~n10720;
  assign n10722 = ~pi0733 & ~n8810;
  assign po0784 = n10721 | n10722;
  assign n10724 = ~pi0734 & ~n8946;
  assign n10725 = n8946 & ~n10033;
  assign n10726 = ~n10724 & ~n10725;
  assign n10727 = n8810 & ~n10726;
  assign n10728 = ~pi0734 & ~n8810;
  assign po0785 = n10727 | n10728;
  assign n10730 = ~pi0735 & ~n8946;
  assign n10731 = n8946 & ~n9822;
  assign n10732 = ~n10730 & ~n10731;
  assign n10733 = n8810 & ~n10732;
  assign n10734 = ~pi0735 & ~n8810;
  assign po0786 = n10733 | n10734;
  assign n10736 = ~pi0736 & ~n8946;
  assign n10737 = n8946 & ~n10286;
  assign n10738 = ~n10736 & ~n10737;
  assign n10739 = n8810 & ~n10738;
  assign n10740 = ~pi0736 & ~n8810;
  assign po0787 = n10739 | n10740;
  assign n10742 = ~pi0737 & ~n8946;
  assign n10743 = n8946 & ~n10021;
  assign n10744 = ~n10742 & ~n10743;
  assign n10745 = n8810 & ~n10744;
  assign n10746 = ~pi0737 & ~n8810;
  assign po0788 = n10745 | n10746;
  assign n10748 = ~pi0738 & ~n8946;
  assign n10749 = n8946 & ~n10303;
  assign n10750 = ~n10748 & ~n10749;
  assign n10751 = n8810 & ~n10750;
  assign n10752 = ~pi0738 & ~n8810;
  assign po0789 = n10751 | n10752;
  assign n10754 = ~pi0739 & ~n8902;
  assign n10755 = n8902 & ~n10645;
  assign n10756 = ~n10754 & ~n10755;
  assign n10757 = n8841 & ~n10756;
  assign n10758 = ~pi0739 & ~n8841;
  assign po0790 = n10757 | n10758;
  assign n10760 = ~pi0740 & ~n8946;
  assign n10761 = n8946 & ~n9513;
  assign n10762 = ~n10760 & ~n10761;
  assign n10763 = n8810 & ~n10762;
  assign n10764 = ~pi0740 & ~n8810;
  assign po0791 = n10763 | n10764;
  assign n10766 = ~pi0741 & ~n8946;
  assign n10767 = n8946 & ~n10510;
  assign n10768 = ~n10766 & ~n10767;
  assign n10769 = n8810 & ~n10768;
  assign n10770 = ~pi0741 & ~n8810;
  assign po0792 = n10769 | n10770;
  assign n10772 = ~pi0742 & ~n8946;
  assign n10773 = n8946 & ~n9492;
  assign n10774 = ~n10772 & ~n10773;
  assign n10775 = n8810 & ~n10774;
  assign n10776 = ~pi0742 & ~n8810;
  assign po0793 = n10775 | n10776;
  assign n10778 = ~pi0743 & ~n8946;
  assign n10779 = n8946 & ~n9553;
  assign n10780 = ~n10778 & ~n10779;
  assign n10781 = n8810 & ~n10780;
  assign n10782 = ~pi0743 & ~n8810;
  assign po0794 = n10781 | n10782;
  assign n10784 = ~pi0744 & ~n8922;
  assign n10785 = n8922 & ~n9553;
  assign n10786 = ~n10784 & ~n10785;
  assign n10787 = n8810 & ~n10786;
  assign n10788 = ~pi0744 & ~n8810;
  assign po0795 = n10787 | n10788;
  assign n10790 = ~pi0745 & ~n8946;
  assign n10791 = n8946 & ~n10599;
  assign n10792 = ~n10790 & ~n10791;
  assign n10793 = n8810 & ~n10792;
  assign n10794 = ~pi0745 & ~n8810;
  assign po0796 = n10793 | n10794;
  assign n10796 = pi0746 & ~n8840;
  assign n10797 = ~n8880 & ~n8902;
  assign n10798 = ~n8837 & ~n10797;
  assign n10799 = ~pi0746 & n10056;
  assign n10800 = pi0746 & ~n10056;
  assign n10801 = ~n10799 & ~n10800;
  assign n10802 = n8837 & ~n10801;
  assign n10803 = ~n10798 & ~n10802;
  assign n10804 = n8840 & ~n10803;
  assign n10805 = ~n10796 & ~n10804;
  assign po0797 = pi1145 & ~n10805;
  assign n10807 = ~pi0747 & ~n8902;
  assign n10808 = n8902 & ~n10227;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = n8841 & ~n10809;
  assign n10811 = ~pi0747 & ~n8841;
  assign po0798 = n10810 | n10811;
  assign n10813 = ~pi0748 & ~n8902;
  assign n10814 = n8902 & ~n10457;
  assign n10815 = ~n10813 & ~n10814;
  assign n10816 = n8841 & ~n10815;
  assign n10817 = ~pi0748 & ~n8841;
  assign po0799 = n10816 | n10817;
  assign n10819 = ~pi0749 & ~n8922;
  assign n10820 = n8922 & ~n10021;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = n8810 & ~n10821;
  assign n10823 = ~pi0749 & ~n8810;
  assign po0800 = n10822 | n10823;
  assign n10825 = n8812 & n8831;
  assign n10826 = ~pi0750 & ~n8812;
  assign n10827 = ~n10825 & ~n10826;
  assign n10828 = n8810 & ~n10827;
  assign n10829 = ~pi0750 & ~n8810;
  assign po0801 = n10828 | n10829;
  assign n10831 = pi0751 & ~n10179;
  assign n10832 = pi0947 & n10179;
  assign po0802 = n10831 | n10832;
  assign n10834 = ~pi0752 & ~n8812;
  assign n10835 = n8812 & ~n10082;
  assign n10836 = ~n10834 & ~n10835;
  assign n10837 = n8810 & ~n10836;
  assign n10838 = ~pi0752 & ~n8810;
  assign po0803 = n10837 | n10838;
  assign n10840 = ~pi0753 & ~n8812;
  assign n10841 = n8812 & ~n10510;
  assign n10842 = ~n10840 & ~n10841;
  assign n10843 = n8810 & ~n10842;
  assign n10844 = ~pi0753 & ~n8810;
  assign po0804 = n10843 | n10844;
  assign n10846 = ~pi0754 & ~n9020;
  assign n10847 = n9020 & ~n10320;
  assign n10848 = ~n10846 & ~n10847;
  assign n10849 = n8841 & ~n10848;
  assign n10850 = ~pi0754 & ~n8841;
  assign po0805 = n10849 | n10850;
  assign n10852 = ~pi0755 & ~n9020;
  assign n10853 = n9020 & ~n10331;
  assign n10854 = ~n10852 & ~n10853;
  assign n10855 = n8841 & ~n10854;
  assign n10856 = ~pi0755 & ~n8841;
  assign po0806 = n10855 | n10856;
  assign n10858 = ~pi0756 & ~n9020;
  assign n10859 = n9020 & ~n10457;
  assign n10860 = ~n10858 & ~n10859;
  assign n10861 = n8841 & ~n10860;
  assign n10862 = ~pi0756 & ~n8841;
  assign po0807 = n10861 | n10862;
  assign n10864 = ~pi0757 & ~n9020;
  assign n10865 = n9020 & ~n10188;
  assign n10866 = ~n10864 & ~n10865;
  assign n10867 = n8841 & ~n10866;
  assign n10868 = ~pi0757 & ~n8841;
  assign po0808 = n10867 | n10868;
  assign n10870 = ~pi0758 & ~n9020;
  assign n10871 = n9020 & ~n10354;
  assign n10872 = ~n10870 & ~n10871;
  assign n10873 = n8841 & ~n10872;
  assign n10874 = ~pi0758 & ~n8841;
  assign po0809 = n10873 | n10874;
  assign n10876 = ~pi0759 & ~n9020;
  assign n10877 = n9020 & ~n10227;
  assign n10878 = ~n10876 & ~n10877;
  assign n10879 = n8841 & ~n10878;
  assign n10880 = ~pi0759 & ~n8841;
  assign po0810 = n10879 | n10880;
  assign n10882 = ~pi0760 & ~n9020;
  assign n10883 = n9020 & ~n10365;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = n8841 & ~n10884;
  assign n10886 = ~pi0760 & ~n8841;
  assign po0811 = n10885 | n10886;
  assign n10888 = ~pi0761 & ~n9020;
  assign n10889 = n9020 & ~n10216;
  assign n10890 = ~n10888 & ~n10889;
  assign n10891 = n8841 & ~n10890;
  assign n10892 = ~pi0761 & ~n8841;
  assign po0812 = n10891 | n10892;
  assign n10894 = n8896 & n9020;
  assign n10895 = ~pi0762 & ~n9020;
  assign n10896 = ~n10894 & ~n10895;
  assign n10897 = n8841 & ~n10896;
  assign n10898 = ~pi0762 & ~n8841;
  assign po0813 = n10897 | n10898;
  assign n10900 = n9020 & n9087;
  assign n10901 = ~pi0763 & ~n9020;
  assign n10902 = ~n10900 & ~n10901;
  assign n10903 = n8841 & ~n10902;
  assign n10904 = ~pi0763 & ~n8841;
  assign po0814 = n10903 | n10904;
  assign n10906 = n8873 & n9020;
  assign n10907 = ~pi0764 & ~n9020;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = n8841 & ~n10908;
  assign n10910 = ~pi0764 & ~n8841;
  assign po0815 = n10909 | n10910;
  assign n10912 = n9020 & n9100;
  assign n10913 = ~pi0765 & ~n9020;
  assign n10914 = ~n10912 & ~n10913;
  assign n10915 = n8841 & ~n10914;
  assign n10916 = ~pi0765 & ~n8841;
  assign po0816 = n10915 | n10916;
  assign n10918 = n8889 & n9020;
  assign n10919 = ~pi0766 & ~n9020;
  assign n10920 = ~n10918 & ~n10919;
  assign n10921 = n8841 & ~n10920;
  assign n10922 = ~pi0766 & ~n8841;
  assign po0817 = n10921 | n10922;
  assign n10924 = n8910 & n9020;
  assign n10925 = ~pi0767 & ~n9020;
  assign n10926 = ~n10924 & ~n10925;
  assign n10927 = n8841 & ~n10926;
  assign n10928 = ~pi0767 & ~n8841;
  assign po0818 = n10927 | n10928;
  assign n10930 = n9020 & n9126;
  assign n10931 = ~pi0768 & ~n9020;
  assign n10932 = ~n10930 & ~n10931;
  assign n10933 = n8841 & ~n10932;
  assign n10934 = ~pi0768 & ~n8841;
  assign po0819 = n10933 | n10934;
  assign n10936 = n8882 & n9020;
  assign n10937 = ~pi0769 & ~n9020;
  assign n10938 = ~n10936 & ~n10937;
  assign n10939 = n8841 & ~n10938;
  assign n10940 = ~pi0769 & ~n8841;
  assign po0820 = n10939 | n10940;
  assign n10942 = n9020 & n9133;
  assign n10943 = ~pi0770 & ~n9020;
  assign n10944 = ~n10942 & ~n10943;
  assign n10945 = n8841 & ~n10944;
  assign n10946 = ~pi0770 & ~n8841;
  assign po0821 = n10945 | n10946;
  assign n10948 = n8844 & n9020;
  assign n10949 = ~pi0771 & ~n9020;
  assign n10950 = ~n10948 & ~n10949;
  assign n10951 = n8841 & ~n10950;
  assign n10952 = ~pi0771 & ~n8841;
  assign po0822 = n10951 | n10952;
  assign n10954 = n9020 & n9146;
  assign n10955 = ~pi0772 & ~n9020;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = n8841 & ~n10956;
  assign n10958 = ~pi0772 & ~n8841;
  assign po0823 = n10957 | n10958;
  assign n10960 = ~pi0773 & ~n9020;
  assign n10961 = n9020 & ~n10394;
  assign n10962 = ~n10960 & ~n10961;
  assign n10963 = n8841 & ~n10962;
  assign n10964 = ~pi0773 & ~n8841;
  assign po0824 = n10963 | n10964;
  assign n10966 = ~pi0774 & ~n9020;
  assign n10967 = n9020 & ~n10239;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = n8841 & ~n10968;
  assign n10970 = ~pi0774 & ~n8841;
  assign po0825 = n10969 | n10970;
  assign n10972 = ~pi0775 & ~n9020;
  assign n10973 = n9020 & ~n10417;
  assign n10974 = ~n10972 & ~n10973;
  assign n10975 = n8841 & ~n10974;
  assign n10976 = ~pi0775 & ~n8841;
  assign po0826 = n10975 | n10976;
  assign n10978 = ~pi0776 & ~n9020;
  assign n10979 = n9020 & ~n10428;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = n8841 & ~n10980;
  assign n10982 = ~pi0776 & ~n8841;
  assign po0827 = n10981 | n10982;
  assign n10984 = ~pi0777 & ~n9020;
  assign n10985 = n9020 & ~n10645;
  assign n10986 = ~n10984 & ~n10985;
  assign n10987 = n8841 & ~n10986;
  assign n10988 = ~pi0777 & ~n8841;
  assign po0828 = n10987 | n10988;
  assign n10990 = ~pi0778 & ~n8812;
  assign n10991 = n8812 & ~n8953;
  assign n10992 = ~n10990 & ~n10991;
  assign n10993 = n8810 & ~n10992;
  assign n10994 = ~pi0778 & ~n8810;
  assign po0829 = n10993 | n10994;
  assign n10996 = ~pi0779 & ~n8812;
  assign n10997 = n8812 & ~n10161;
  assign n10998 = ~n10996 & ~n10997;
  assign n10999 = n8810 & ~n10998;
  assign n11000 = ~pi0779 & ~n8810;
  assign po0830 = n10999 | n11000;
  assign n11002 = ~pi0780 & ~n8812;
  assign n11003 = n8812 & ~n10286;
  assign n11004 = ~n11002 & ~n11003;
  assign n11005 = n8810 & ~n11004;
  assign n11006 = ~pi0780 & ~n8810;
  assign po0831 = n11005 | n11006;
  assign n11008 = ~pi0781 & ~n8812;
  assign n11009 = n8812 & ~n10144;
  assign n11010 = ~n11008 & ~n11009;
  assign n11011 = n8810 & ~n11010;
  assign n11012 = ~pi0781 & ~n8810;
  assign po0832 = n11011 | n11012;
  assign n11014 = ~pi0782 & ~n8812;
  assign n11015 = n8812 & ~n10303;
  assign n11016 = ~n11014 & ~n11015;
  assign n11017 = n8810 & ~n11016;
  assign n11018 = ~pi0782 & ~n8810;
  assign po0833 = n11017 | n11018;
  assign n11020 = ~pi0783 & ~n8812;
  assign n11021 = n8812 & ~n10021;
  assign n11022 = ~n11020 & ~n11021;
  assign n11023 = n8810 & ~n11022;
  assign n11024 = ~pi0783 & ~n8810;
  assign po0834 = n11023 | n11024;
  assign n11026 = n8812 & n9172;
  assign n11027 = ~pi0784 & ~n8812;
  assign n11028 = ~n11026 & ~n11027;
  assign n11029 = n8810 & ~n11028;
  assign n11030 = ~pi0784 & ~n8810;
  assign po0835 = n11029 | n11030;
  assign n11032 = ~pi0785 & ~n8812;
  assign n11033 = n8812 & ~n9513;
  assign n11034 = ~n11032 & ~n11033;
  assign n11035 = n8810 & ~n11034;
  assign n11036 = ~pi0785 & ~n8810;
  assign po0836 = n11035 | n11036;
  assign n11038 = n8812 & n9153;
  assign n11039 = ~pi0786 & ~n8812;
  assign n11040 = ~n11038 & ~n11039;
  assign n11041 = n8810 & ~n11040;
  assign n11042 = ~pi0786 & ~n8810;
  assign po0837 = n11041 | n11042;
  assign n11044 = ~pi0787 & ~n8812;
  assign n11045 = n8812 & ~n9503;
  assign n11046 = ~n11044 & ~n11045;
  assign n11047 = n8810 & ~n11046;
  assign n11048 = ~pi0787 & ~n8810;
  assign po0838 = n11047 | n11048;
  assign n11050 = ~pi0788 & ~n8812;
  assign n11051 = n8812 & ~n10599;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = n8810 & ~n11052;
  assign n11054 = ~pi0788 & ~n8810;
  assign po0839 = n11053 | n11054;
  assign n11056 = ~pi0789 & ~n8812;
  assign n11057 = n8812 & ~n9525;
  assign n11058 = ~n11056 & ~n11057;
  assign n11059 = n8810 & ~n11058;
  assign n11060 = ~pi0789 & ~n8810;
  assign po0840 = n11059 | n11060;
  assign n11062 = pi0790 & pi1036;
  assign n11063 = ~n8809 & n11062;
  assign n11064 = pi0790 & ~n8806;
  assign n11065 = ~n8807 & ~n11064;
  assign n11066 = n8809 & ~n11065;
  assign n11067 = pi1036 & n11066;
  assign po0841 = n11063 | n11067;
  assign n11069 = pi0791 & ~n10179;
  assign n11070 = pi1935 & n10179;
  assign po0842 = n11069 | n11070;
  assign n11072 = pi0792 & ~n10179;
  assign n11073 = pi0335 & n10179;
  assign po0843 = n11072 | n11073;
  assign n11075 = pi0793 & ~n10179;
  assign n11076 = pi0233 & n10179;
  assign po0844 = n11075 | n11076;
  assign n11078 = pi0794 & ~n10179;
  assign n11079 = pi0213 & n10179;
  assign po0845 = n11078 | n11079;
  assign n11081 = pi0795 & ~n10179;
  assign n11082 = pi0208 & n10179;
  assign po0846 = n11081 | n11082;
  assign n11084 = pi0796 & ~n10179;
  assign n11085 = pi0197 & n10179;
  assign po0847 = n11084 | n11085;
  assign n11087 = pi0797 & ~n10179;
  assign n11088 = pi0193 & n10179;
  assign po0848 = n11087 | n11088;
  assign n11090 = pi0798 & ~n10179;
  assign n11091 = pi1926 & n10179;
  assign po0849 = n11090 | n11091;
  assign n11093 = pi0799 & ~n10179;
  assign n11094 = pi1901 & n10179;
  assign po0850 = n11093 | n11094;
  assign n11096 = pi0800 & ~n10179;
  assign n11097 = pi1875 & n10179;
  assign po0851 = n11096 | n11097;
  assign n11099 = pi0801 & ~n10179;
  assign n11100 = pi0923 & n10179;
  assign po0852 = n11099 | n11100;
  assign n11102 = pi0802 & ~n10179;
  assign n11103 = pi0877 & n10179;
  assign po0853 = n11102 | n11103;
  assign n11105 = pi0803 & ~n10179;
  assign n11106 = pi0871 & n10179;
  assign po0854 = n11105 | n11106;
  assign n11108 = pi0804 & ~n10179;
  assign n11109 = pi0480 & n10179;
  assign po0855 = n11108 | n11109;
  assign n11111 = ~pi0805 & ~n8880;
  assign n11112 = n8880 & ~n10645;
  assign n11113 = ~n11111 & ~n11112;
  assign n11114 = n8841 & ~n11113;
  assign n11115 = ~pi0805 & ~n8841;
  assign po0856 = n11114 | n11115;
  assign n11117 = ~pi1903 & n5196;
  assign po0857 = ~pi0806 | n11117;
  assign n11119 = ~pi1908 & n5215;
  assign po0858 = ~pi0807 | n11119;
  assign n11121 = pi2055 & n8809;
  assign po0859 = ~pi0808 | n11121;
  assign n11123 = pi0946 & ~pi1930;
  assign n11124 = pi0809 & ~n11123;
  assign n11125 = ~pi1144 & pi1905;
  assign po0860 = n11124 | n11125;
  assign n11127 = pi0809 & n11123;
  assign n11128 = ~pi0810 & ~n11127;
  assign po0861 = ~n5425 & ~n11128;
  assign n11130 = n8812 & n9000;
  assign n11131 = ~pi0811 & ~n8812;
  assign n11132 = ~n11130 & ~n11131;
  assign n11133 = n8810 & ~n11132;
  assign n11134 = ~pi0811 & ~n8810;
  assign po0862 = n11133 | n11134;
  assign n11136 = ~pi0247 & ~pi2032;
  assign n11137 = pi0890 & pi2032;
  assign po0863 = n11136 | n11137;
  assign n11139 = ~pi0790 & n8809;
  assign n11140 = pi0813 & ~n11139;
  assign n11141 = pi0207 & n11139;
  assign po0864 = n11140 | n11141;
  assign n11143 = pi0891 & ~pi2058;
  assign n11144 = pi0814 & pi2058;
  assign po0865 = n11143 | n11144;
  assign n11146 = ~pi0815 & ~pi0908;
  assign po0866 = ~n5425 & ~n11146;
  assign n11148 = pi0816 & ~pi2060;
  assign n11149 = pi0891 & pi2060;
  assign po0867 = n11148 | n11149;
  assign n11151 = pi0891 & ~pi2056;
  assign n11152 = pi0817 & pi2056;
  assign po0868 = n11151 | n11152;
  assign n11154 = pi0891 & ~pi2059;
  assign n11155 = pi0818 & pi2059;
  assign po0869 = n11154 | n11155;
  assign n11157 = pi0891 & ~pi2057;
  assign n11158 = pi0819 & pi2057;
  assign po0870 = n11157 | n11158;
  assign n11160 = pi0820 & ~n11139;
  assign n11161 = pi0235 & n11139;
  assign po0871 = n11160 | n11161;
  assign n11163 = pi0821 & pi1145;
  assign n11164 = ~n8840 & n11163;
  assign n11165 = pi0821 & ~n8837;
  assign n11166 = ~n8838 & ~n11165;
  assign n11167 = n8840 & ~n11166;
  assign n11168 = pi1145 & n11167;
  assign po0872 = n11164 | n11168;
  assign n11170 = pi0822 & ~n11139;
  assign n11171 = pi0915 & n11139;
  assign po0873 = n11170 | n11171;
  assign n11173 = pi0823 & ~n11139;
  assign n11174 = pi1852 & n11139;
  assign po0874 = n11173 | n11174;
  assign n11176 = pi0824 & ~n11139;
  assign n11177 = pi1924 & n11139;
  assign po0875 = n11176 | n11177;
  assign n11179 = pi0825 & ~n11139;
  assign n11180 = pi1886 & n11139;
  assign po0876 = n11179 | n11180;
  assign n11182 = pi0826 & ~n11139;
  assign n11183 = pi0950 & n11139;
  assign po0877 = n11182 | n11183;
  assign n11185 = pi0827 & ~n11139;
  assign n11186 = pi0882 & n11139;
  assign po0878 = n11185 | n11186;
  assign n11188 = pi0828 & ~n11139;
  assign n11189 = pi0819 & n11139;
  assign po0879 = n11188 | n11189;
  assign n11191 = pi0829 & ~n11139;
  assign n11192 = pi0479 & n11139;
  assign po0880 = n11191 | n11192;
  assign n11194 = pi0830 & ~n11139;
  assign n11195 = pi0866 & n11139;
  assign po0881 = n11194 | n11195;
  assign n11197 = pi0831 & ~n11139;
  assign n11198 = pi1934 & n11139;
  assign po0882 = n11197 | n11198;
  assign n11200 = pi0832 & ~n11139;
  assign n11201 = pi0334 & n11139;
  assign po0883 = n11200 | n11201;
  assign n11203 = pi0833 & ~n11139;
  assign n11204 = pi0192 & n11139;
  assign po0884 = n11203 | n11204;
  assign n11206 = pi0834 & ~n11139;
  assign n11207 = pi0196 & n11139;
  assign po0885 = n11206 | n11207;
  assign n11209 = pi0835 & ~n11139;
  assign n11210 = pi0212 & n11139;
  assign po0886 = n11209 | n11210;
  assign n11212 = pi0449 & pi0836;
  assign n11213 = pi0449 & n11123;
  assign po0887 = n11212 | n11213;
  assign n11215 = pi0860 & pi0873;
  assign n11216 = ~pi0837 & ~n11215;
  assign po0888 = n11213 | n11216;
  assign n11218 = pi1176 & ~pi1904;
  assign n11219 = pi1176 & ~pi2005;
  assign n11220 = ~n11218 & ~n11219;
  assign n11221 = pi1176 & ~pi2138;
  assign n11222 = n11220 & ~n11221;
  assign n11223 = n5054 & ~n11222;
  assign n11224 = ~pi2138 & n11219;
  assign n11225 = ~n11218 & ~n11224;
  assign n11226 = n5062 & ~n11225;
  assign n11227 = n5065 & ~n11220;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = n5056 & n11218;
  assign n11230 = n11228 & ~n11229;
  assign po0889 = n11223 | ~n11230;
  assign n11232 = pi1035 & ~pi1903;
  assign n11233 = pi1035 & ~pi1987;
  assign n11234 = ~n11232 & ~n11233;
  assign n11235 = pi1035 & ~pi2140;
  assign n11236 = n11234 & ~n11235;
  assign n11237 = n5030 & ~n11236;
  assign n11238 = ~pi2140 & n11233;
  assign n11239 = ~n11232 & ~n11238;
  assign n11240 = n5038 & ~n11239;
  assign n11241 = n5041 & ~n11234;
  assign n11242 = ~n11240 & ~n11241;
  assign n11243 = n5032 & n11232;
  assign n11244 = n11242 & ~n11243;
  assign po0890 = n11237 | ~n11244;
  assign n11246 = ~pi0841 & ~pi0928;
  assign po0892 = ~n5425 & ~n11246;
  assign n11248 = ~pi0842 & ~pi0927;
  assign po0893 = ~n5425 & ~n11248;
  assign n11250 = pi0843 & ~n8840;
  assign n11251 = pi0821 & ~pi0843;
  assign n11252 = ~pi0821 & pi0843;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = n8837 & ~n11253;
  assign n11255 = ~pi0843 & ~n8837;
  assign n11256 = ~n11254 & ~n11255;
  assign n11257 = n8840 & ~n11256;
  assign n11258 = ~n11250 & ~n11257;
  assign po0894 = pi1145 & ~n11258;
  assign n11260 = ~pi0821 & n8840;
  assign n11261 = pi0844 & ~n11260;
  assign n11262 = pi0481 & n11260;
  assign po0895 = n11261 | n11262;
  assign n11264 = pi0845 & ~n11260;
  assign n11265 = pi1853 & n11260;
  assign po0896 = n11264 | n11265;
  assign n11267 = pi0846 & ~n11260;
  assign n11268 = pi0333 & n11260;
  assign po0897 = n11267 | n11268;
  assign n11270 = pi0847 & ~n11260;
  assign n11271 = pi0195 & n11260;
  assign po0898 = n11270 | n11271;
  assign n11273 = pi0848 & ~n11260;
  assign n11274 = pi1933 & n11260;
  assign po0899 = n11273 | n11274;
  assign n11276 = pi0849 & ~n11260;
  assign n11277 = pi0231 & n11260;
  assign po0900 = n11276 | n11277;
  assign n11279 = pi0850 & ~n11260;
  assign n11280 = pi0211 & n11260;
  assign po0901 = n11279 | n11280;
  assign n11282 = pi0851 & ~n11260;
  assign n11283 = pi0206 & n11260;
  assign po0902 = n11282 | n11283;
  assign n11285 = pi0852 & ~n11260;
  assign n11286 = pi0191 & n11260;
  assign po0903 = n11285 | n11286;
  assign n11288 = pi0853 & ~n11260;
  assign n11289 = pi1925 & n11260;
  assign po0904 = n11288 | n11289;
  assign n11291 = pi0854 & ~n11260;
  assign n11292 = pi1883 & n11260;
  assign po0905 = n11291 | n11292;
  assign n11294 = pi0855 & ~n11260;
  assign n11295 = pi0916 & n11260;
  assign po0906 = n11294 | n11295;
  assign n11297 = pi0856 & ~n11260;
  assign n11298 = pi0883 & n11260;
  assign po0907 = n11297 | n11298;
  assign n11300 = pi0857 & ~n11260;
  assign n11301 = pi0951 & n11260;
  assign po0908 = n11300 | n11301;
  assign n11303 = pi0858 & ~n11260;
  assign n11304 = pi0818 & n11260;
  assign po0909 = n11303 | n11304;
  assign n11306 = pi0859 & ~n11260;
  assign n11307 = pi0870 & n11260;
  assign po0910 = n11306 | n11307;
  assign n11309 = pi0860 & ~pi0873;
  assign n11310 = ~pi0837 & n8743;
  assign po0911 = n11309 | n11310;
  assign n11312 = pi1839 & ~pi1909;
  assign n11313 = pi1839 & ~pi2006;
  assign n11314 = ~n11312 & ~n11313;
  assign n11315 = pi1839 & ~pi2141;
  assign n11316 = n11314 & ~n11315;
  assign n11317 = n5129 & ~n11316;
  assign n11318 = ~pi2141 & n11313;
  assign n11319 = ~n11312 & ~n11318;
  assign n11320 = n5137 & ~n11319;
  assign n11321 = n5140 & ~n11314;
  assign n11322 = ~n11320 & ~n11321;
  assign n11323 = n5131 & n11312;
  assign n11324 = n11322 & ~n11323;
  assign po0912 = n11317 | ~n11324;
  assign n11326 = pi1838 & ~pi1910;
  assign n11327 = pi1838 & ~pi2007;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = pi1838 & ~pi2159;
  assign n11330 = n11328 & ~n11329;
  assign n11331 = n5153 & ~n11330;
  assign n11332 = ~pi2159 & n11327;
  assign n11333 = ~n11326 & ~n11332;
  assign n11334 = n5161 & ~n11333;
  assign n11335 = n5164 & ~n11328;
  assign n11336 = ~n11334 & ~n11335;
  assign n11337 = n5155 & n11326;
  assign n11338 = n11336 & ~n11337;
  assign po0913 = n11331 | ~n11338;
  assign n11340 = pi1164 & ~pi1907;
  assign n11341 = pi1164 & ~pi2004;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = pi1164 & ~pi2139;
  assign n11344 = n11342 & ~n11343;
  assign n11345 = n5081 & ~n11344;
  assign n11346 = ~pi2139 & n11341;
  assign n11347 = ~n11340 & ~n11346;
  assign n11348 = n5089 & ~n11347;
  assign n11349 = n5092 & ~n11342;
  assign n11350 = ~n11348 & ~n11349;
  assign n11351 = n5083 & n11340;
  assign n11352 = n11350 & ~n11351;
  assign po0914 = n11345 | ~n11352;
  assign n11354 = pi1169 & ~pi1908;
  assign n11355 = pi1169 & ~pi1988;
  assign n11356 = ~n11354 & ~n11355;
  assign n11357 = pi1169 & ~pi2158;
  assign n11358 = n11356 & ~n11357;
  assign n11359 = n5105 & ~n11358;
  assign n11360 = ~pi2158 & n11355;
  assign n11361 = ~n11354 & ~n11360;
  assign n11362 = n5113 & ~n11361;
  assign n11363 = n5116 & ~n11356;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = n5107 & n11354;
  assign n11366 = n11364 & ~n11365;
  assign po0915 = n11359 | ~n11366;
  assign po0916 = ~pi2254 & ~n7317;
  assign n11369 = pi0925 & ~pi2057;
  assign n11370 = pi0866 & pi2057;
  assign po0917 = n11369 | n11370;
  assign n11372 = pi0867 & ~pi2060;
  assign n11373 = pi0925 & pi2060;
  assign po0918 = n11372 | n11373;
  assign n11375 = pi0925 & ~pi2035;
  assign n11376 = pi0868 & pi2035;
  assign po0919 = n11375 | n11376;
  assign n11378 = pi0925 & ~pi2056;
  assign n11379 = pi0869 & pi2056;
  assign po0920 = n11378 | n11379;
  assign n11381 = pi0925 & ~pi2059;
  assign n11382 = pi0870 & pi2059;
  assign po0921 = n11381 | n11382;
  assign n11384 = pi0925 & ~pi2058;
  assign n11385 = pi0871 & pi2058;
  assign po0922 = n11384 | n11385;
  assign n11387 = pi2033 & n8840;
  assign po0923 = ~pi0872 | n11387;
  assign po0924 = pi0860 & n8743;
  assign po0925 = ~pi2252 & ~n7490;
  assign po0926 = ~pi2253 & ~n7514;
  assign n11392 = pi1768 & ~pi2058;
  assign n11393 = pi0877 & pi2058;
  assign po0928 = n11392 | n11393;
  assign n11395 = pi1768 & ~pi2056;
  assign n11396 = pi0878 & pi2056;
  assign po0929 = n11395 | n11396;
  assign n11398 = pi1844 & pi1884;
  assign n11399 = ~pi0914 & ~n11398;
  assign n11400 = pi0232 & n11399;
  assign n11401 = pi1839 & pi1930;
  assign n11402 = pi0879 & pi1839;
  assign n11403 = ~n11401 & ~n11402;
  assign n11404 = n11400 & ~n11403;
  assign po0930 = po1130 | n11404;
  assign n11406 = pi1879 & pi2134;
  assign n11407 = ~pi0880 & ~n11406;
  assign n11408 = ~pi1956 & ~pi2003;
  assign n11409 = pi1990 & pi2001;
  assign n11410 = n11408 & n11409;
  assign po0931 = ~n11407 & ~n11410;
  assign n11412 = pi1768 & ~pi2035;
  assign n11413 = pi0881 & pi2035;
  assign po0932 = n11412 | n11413;
  assign n11415 = pi1768 & ~pi2057;
  assign n11416 = pi0882 & pi2057;
  assign po0933 = n11415 | n11416;
  assign n11418 = pi1768 & ~pi2059;
  assign n11419 = pi0883 & pi2059;
  assign po0934 = n11418 | n11419;
  assign n11421 = pi0868 & pi1172;
  assign n11422 = ~pi0909 & ~n11421;
  assign n11423 = pi0232 & n11422;
  assign n11424 = pi1164 & pi1930;
  assign n11425 = pi0884 & pi1164;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = n11423 & ~n11426;
  assign po1126 = pi0884 & pi1930;
  assign po0935 = n11427 | po1126;
  assign n11430 = pi0881 & pi1187;
  assign n11431 = ~pi0910 & ~n11430;
  assign n11432 = pi0232 & n11431;
  assign n11433 = pi1035 & pi1930;
  assign n11434 = pi0885 & pi1035;
  assign n11435 = ~n11433 & ~n11434;
  assign n11436 = n11432 & ~n11435;
  assign po0936 = po1127 | n11436;
  assign n11438 = pi0949 & pi1170;
  assign n11439 = ~pi0911 & ~n11438;
  assign n11440 = pi0232 & n11439;
  assign n11441 = pi1169 & pi1930;
  assign n11442 = pi0886 & pi1169;
  assign n11443 = ~n11441 & ~n11442;
  assign n11444 = n11440 & ~n11443;
  assign po0937 = po1128 | n11444;
  assign n11446 = pi1177 & pi1850;
  assign n11447 = ~pi0907 & ~n11446;
  assign n11448 = pi0232 & n11447;
  assign n11449 = pi1176 & pi1930;
  assign n11450 = pi0887 & pi1176;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = n11448 & ~n11451;
  assign po0938 = po1129 | n11452;
  assign n11454 = pi1870 & pi1922;
  assign n11455 = ~pi0912 & ~n11454;
  assign n11456 = pi0232 & n11455;
  assign n11457 = pi1838 & pi1930;
  assign n11458 = pi0888 & pi1838;
  assign n11459 = ~n11457 & ~n11458;
  assign n11460 = n11456 & ~n11459;
  assign po0939 = po1131 | n11460;
  assign n11462 = pi0889 & ~pi1930;
  assign n11463 = pi0809 & pi1930;
  assign n11464 = pi0449 & pi1930;
  assign n11465 = ~n11463 & ~n11464;
  assign po0940 = n11462 | ~n11465;
  assign n11467 = ~pi0246 & ~pi2032;
  assign n11468 = pi1874 & pi2032;
  assign po0941 = n11467 | n11468;
  assign n11470 = pi0893 & pi0896;
  assign n11471 = pi0895 & pi0897;
  assign n11472 = pi0894 & n11471;
  assign n11473 = n11470 & n11472;
  assign n11474 = pi0892 & n11473;
  assign n11475 = ~pi0892 & ~n11473;
  assign n11476 = ~n11474 & ~n11475;
  assign n11477 = pi0894 & ~pi0895;
  assign n11478 = ~pi0897 & n11477;
  assign n11479 = ~pi0893 & n11478;
  assign n11480 = pi0892 & n11479;
  assign n11481 = pi0896 & n11480;
  assign n11482 = pi1878 & ~n11481;
  assign po0943 = n11476 & n11482;
  assign n11484 = pi0894 & pi0895;
  assign n11485 = ~pi0893 & n11484;
  assign n11486 = pi0893 & ~n11484;
  assign n11487 = ~n11485 & ~n11486;
  assign po0944 = n11482 & ~n11487;
  assign po0945 = ~pi0894 & n11482;
  assign n11490 = ~pi0894 & pi0895;
  assign n11491 = ~n11477 & ~n11490;
  assign po0946 = n11482 & ~n11491;
  assign n11493 = pi0893 & pi0897;
  assign n11494 = n11484 & n11493;
  assign n11495 = pi0896 & n11494;
  assign n11496 = ~pi0896 & ~n11494;
  assign n11497 = ~n11495 & ~n11496;
  assign po0947 = n11482 & n11497;
  assign n11499 = pi0893 & n11484;
  assign n11500 = pi0897 & n11499;
  assign n11501 = ~pi0897 & ~n11499;
  assign n11502 = ~n11500 & ~n11501;
  assign po0948 = n11482 & n11502;
  assign n11504 = ~pi2238 & ~pi2239;
  assign n11505 = ~pi2240 & n11504;
  assign n11506 = pi2242 & n11505;
  assign n11507 = ~pi2241 & n11506;
  assign n11508 = pi2104 & n11507;
  assign n11509 = pi2241 & ~pi2242;
  assign n11510 = pi2239 & n11509;
  assign n11511 = pi2240 & n11510;
  assign n11512 = ~pi2238 & n11511;
  assign n11513 = pi2130 & n11512;
  assign n11514 = ~n11508 & ~n11513;
  assign n11515 = pi2238 & n11511;
  assign n11516 = ~n11512 & ~n11515;
  assign n11517 = ~n11507 & n11516;
  assign n11518 = pi2238 & ~pi2239;
  assign n11519 = pi2240 & n11518;
  assign n11520 = pi1198 & n11519;
  assign n11521 = pi2240 & n11504;
  assign n11522 = pi2146 & n11521;
  assign n11523 = ~n11520 & ~n11522;
  assign n11524 = pi2134 & ~pi2238;
  assign n11525 = n5418 & n11524;
  assign n11526 = pi0810 & n5423;
  assign n11527 = ~n11525 & ~n11526;
  assign n11528 = n11523 & n11527;
  assign n11529 = ~pi2240 & n11518;
  assign n11530 = pi1172 & n11529;
  assign n11531 = n11528 & ~n11530;
  assign n11532 = ~pi2240 & n5422;
  assign n11533 = pi1844 & n11532;
  assign n11534 = pi2238 & pi2239;
  assign n11535 = ~pi2240 & n11534;
  assign n11536 = pi1153 & n11535;
  assign n11537 = ~n11533 & ~n11536;
  assign n11538 = n11531 & n11537;
  assign n11539 = n11517 & ~n11538;
  assign n11540 = pi2026 & n11515;
  assign n11541 = ~n11539 & ~n11540;
  assign po0949 = ~n11514 | ~n11541;
  assign n11543 = ~pi0221 & ~pi0935;
  assign n11544 = pi0221 & pi0935;
  assign n11545 = ~n11543 & ~n11544;
  assign n11546 = pi0225 & pi0918;
  assign n11547 = ~pi0225 & ~pi0918;
  assign po2190 = n11546 | n11547;
  assign n11549 = pi0217 & pi0941;
  assign n11550 = ~pi0217 & ~pi0941;
  assign n11551 = ~n11549 & ~n11550;
  assign n11552 = po2190 & ~n11551;
  assign n11553 = pi1937 & n11552;
  assign n11554 = n11545 & n11553;
  assign po0950 = ~pi0899 | n11554;
  assign n11556 = ~pi0237 & ~pi0945;
  assign n11557 = pi0237 & pi0945;
  assign n11558 = ~n11556 & ~n11557;
  assign n11559 = pi0236 & pi0919;
  assign n11560 = ~pi0236 & ~pi0919;
  assign po2191 = n11559 | n11560;
  assign n11562 = pi0214 & pi0942;
  assign n11563 = ~pi0214 & ~pi0942;
  assign n11564 = ~n11562 & ~n11563;
  assign n11565 = po2191 & ~n11564;
  assign n11566 = pi1938 & n11565;
  assign n11567 = n11558 & n11566;
  assign po0951 = ~pi0900 | n11567;
  assign n11569 = ~pi0223 & ~pi0937;
  assign n11570 = pi0223 & pi0937;
  assign n11571 = ~n11569 & ~n11570;
  assign n11572 = pi0226 & pi0922;
  assign n11573 = ~pi0226 & ~pi0922;
  assign po2192 = n11572 | n11573;
  assign n11575 = pi0219 & pi0944;
  assign n11576 = ~pi0219 & ~pi0944;
  assign n11577 = ~n11575 & ~n11576;
  assign n11578 = po2192 & ~n11577;
  assign n11579 = pi1940 & n11578;
  assign n11580 = n11571 & n11579;
  assign po0952 = ~pi0901 | n11580;
  assign n11582 = ~pi0222 & ~pi0931;
  assign n11583 = pi0222 & pi0931;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = pi0227 & pi0921;
  assign n11586 = ~pi0227 & ~pi0921;
  assign po2189 = n11585 | n11586;
  assign n11588 = pi0218 & pi0943;
  assign n11589 = ~pi0218 & ~pi0943;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = po2189 & ~n11590;
  assign n11592 = pi1936 & n11591;
  assign n11593 = n11584 & n11592;
  assign po0953 = ~pi0902 | n11593;
  assign n11595 = pi0903 & ~pi1930;
  assign po0954 = n11463 | n11595;
  assign n11597 = ~pi0220 & ~pi0934;
  assign n11598 = pi0220 & pi0934;
  assign n11599 = ~n11597 & ~n11598;
  assign n11600 = ~pi0224 & ~pi0917;
  assign n11601 = pi0224 & pi0917;
  assign po2210 = n11600 | n11601;
  assign n11603 = pi0216 & pi0940;
  assign n11604 = ~pi0216 & ~pi0940;
  assign n11605 = ~n11603 & ~n11604;
  assign n11606 = po2210 & ~n11605;
  assign n11607 = pi1941 & n11606;
  assign n11608 = n11599 & n11607;
  assign po0955 = ~pi0904 | n11608;
  assign n11610 = ~pi0239 & ~pi0936;
  assign n11611 = pi0239 & pi0936;
  assign n11612 = ~n11610 & ~n11611;
  assign n11613 = pi0238 & pi0920;
  assign n11614 = ~pi0238 & ~pi0920;
  assign po2209 = n11613 | n11614;
  assign n11616 = ~pi0215 & ~pi0930;
  assign n11617 = pi0215 & pi0930;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = po2209 & ~n11618;
  assign n11620 = pi1939 & n11619;
  assign n11621 = n11612 & n11620;
  assign po0956 = ~pi0905 | n11621;
  assign n11623 = pi1880 & ~pi2056;
  assign n11624 = pi0906 & pi2056;
  assign po0957 = n11623 | n11624;
  assign n11626 = pi0907 & pi1930;
  assign n11627 = ~pi1904 & ~pi1930;
  assign po0958 = n11626 | n11627;
  assign n11629 = pi1150 & pi2020;
  assign n11630 = pi1150 & ~pi2008;
  assign n11631 = ~n11629 & ~n11630;
  assign n11632 = pi1150 & ~pi2137;
  assign n11633 = n11631 & ~n11632;
  assign n11634 = n7304 & ~n11633;
  assign n11635 = ~pi2137 & n11630;
  assign n11636 = ~n11629 & ~n11635;
  assign n11637 = n7312 & ~n11636;
  assign n11638 = n7315 & ~n11631;
  assign n11639 = ~n11637 & ~n11638;
  assign n11640 = n7306 & n11629;
  assign n11641 = n11639 & ~n11640;
  assign po0959 = n11634 | ~n11641;
  assign n11643 = pi0909 & pi1930;
  assign n11644 = ~pi1907 & ~pi1930;
  assign po0960 = n11643 | n11644;
  assign n11646 = pi0910 & pi1930;
  assign n11647 = ~pi1903 & ~pi1930;
  assign po0961 = n11646 | n11647;
  assign n11649 = pi0911 & pi1930;
  assign n11650 = ~pi1908 & ~pi1930;
  assign po0962 = n11649 | n11650;
  assign n11652 = pi0912 & pi1930;
  assign n11653 = ~pi1910 & ~pi1930;
  assign po0963 = n11652 | n11653;
  assign n11655 = pi0913 & ~pi2060;
  assign n11656 = pi1880 & pi2060;
  assign po0964 = n11655 | n11656;
  assign n11658 = pi0914 & pi1930;
  assign n11659 = ~pi1909 & ~pi1930;
  assign po0965 = n11658 | n11659;
  assign n11661 = pi1880 & ~pi2057;
  assign n11662 = pi0915 & pi2057;
  assign po0966 = n11661 | n11662;
  assign n11664 = pi1880 & ~pi2059;
  assign n11665 = pi0916 & pi2059;
  assign po0967 = n11664 | n11665;
  assign n11667 = ~pi0917 & pi1941;
  assign n11668 = pi0917 & ~pi1941;
  assign n11669 = ~n11667 & ~n11668;
  assign po0968 = pi1838 & ~n11669;
  assign n11671 = ~pi0918 & pi1937;
  assign n11672 = pi0918 & ~pi1937;
  assign n11673 = ~n11671 & ~n11672;
  assign po0969 = pi1164 & ~n11673;
  assign n11675 = ~pi0919 & pi1938;
  assign n11676 = pi0919 & ~pi1938;
  assign n11677 = ~n11675 & ~n11676;
  assign po0970 = pi1035 & ~n11677;
  assign n11679 = ~pi0920 & pi1939;
  assign n11680 = pi0920 & ~pi1939;
  assign n11681 = ~n11679 & ~n11680;
  assign po0971 = pi1169 & ~n11681;
  assign n11683 = ~pi0921 & pi1936;
  assign n11684 = pi0921 & ~pi1936;
  assign n11685 = ~n11683 & ~n11684;
  assign po0972 = pi1176 & ~n11685;
  assign n11687 = ~pi0922 & pi1940;
  assign n11688 = pi0922 & ~pi1940;
  assign n11689 = ~n11687 & ~n11688;
  assign po0973 = pi1839 & ~n11689;
  assign n11691 = pi1880 & ~pi2058;
  assign n11692 = pi0923 & pi2058;
  assign po0974 = n11691 | n11692;
  assign n11694 = pi0926 & ~pi0933;
  assign n11695 = ~pi0932 & n11694;
  assign n11696 = ~pi0924 & ~n11695;
  assign po0975 = pi1878 & ~n11696;
  assign n11698 = n11481 & ~n11695;
  assign n11699 = pi0926 & ~n11698;
  assign n11700 = pi0932 & pi0933;
  assign n11701 = pi0926 & ~n11700;
  assign n11702 = ~pi0926 & n11700;
  assign n11703 = ~n11701 & ~n11702;
  assign n11704 = n11698 & ~n11703;
  assign n11705 = ~n11699 & ~n11704;
  assign po0977 = pi1878 & ~n11705;
  assign n11707 = pi1145 & pi2033;
  assign n11708 = pi1145 & ~pi2017;
  assign n11709 = ~n11707 & ~n11708;
  assign n11710 = pi1145 & ~pi2136;
  assign n11711 = n11709 & ~n11710;
  assign n11712 = n7477 & ~n11711;
  assign n11713 = ~pi2136 & n11708;
  assign n11714 = ~n11707 & ~n11713;
  assign n11715 = n7485 & ~n11714;
  assign n11716 = n7488 & ~n11709;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = n7479 & n11707;
  assign n11719 = n11717 & ~n11718;
  assign po0978 = n11712 | ~n11719;
  assign n11721 = pi1036 & pi2055;
  assign n11722 = pi1036 & ~pi2016;
  assign n11723 = ~n11721 & ~n11722;
  assign n11724 = pi1036 & ~pi2135;
  assign n11725 = n11723 & ~n11724;
  assign n11726 = n7501 & ~n11725;
  assign n11727 = ~pi2135 & n11722;
  assign n11728 = ~n11721 & ~n11727;
  assign n11729 = n7509 & ~n11728;
  assign n11730 = n7512 & ~n11723;
  assign n11731 = ~n11729 & ~n11730;
  assign n11732 = n7503 & n11721;
  assign n11733 = n11731 & ~n11732;
  assign po0979 = n11726 | ~n11733;
  assign n11735 = ~pi0913 & pi1151;
  assign n11736 = ~pi1857 & ~n11735;
  assign n11737 = pi0232 & n11736;
  assign n11738 = pi0929 & pi1150;
  assign n11739 = pi1150 & pi1943;
  assign n11740 = ~n11738 & ~n11739;
  assign n11741 = n11737 & ~n11740;
  assign po0980 = po1885 | n11741;
  assign n11743 = pi0930 & pi1169;
  assign n11744 = ~pi1939 & n11743;
  assign n11745 = pi0920 & ~pi0930;
  assign n11746 = ~pi0920 & pi0930;
  assign n11747 = ~n11745 & ~n11746;
  assign n11748 = pi1939 & ~n11747;
  assign n11749 = pi1169 & n11748;
  assign po0981 = n11744 | n11749;
  assign n11751 = pi0921 & pi0943;
  assign n11752 = ~pi0931 & n11751;
  assign n11753 = pi0931 & ~n11751;
  assign n11754 = ~n11752 & ~n11753;
  assign n11755 = pi1936 & ~n11754;
  assign n11756 = pi0931 & ~pi1936;
  assign n11757 = ~n11755 & ~n11756;
  assign po0982 = pi1176 & ~n11757;
  assign n11759 = pi0932 & ~n11698;
  assign n11760 = ~pi0932 & n11698;
  assign n11761 = ~n11759 & ~n11760;
  assign po0983 = pi1878 & ~n11761;
  assign n11763 = pi0933 & ~n11698;
  assign n11764 = pi0932 & ~pi0933;
  assign n11765 = ~pi0932 & pi0933;
  assign n11766 = ~n11764 & ~n11765;
  assign n11767 = n11698 & ~n11766;
  assign n11768 = ~n11763 & ~n11767;
  assign po0984 = pi1878 & ~n11768;
  assign n11770 = pi0917 & pi0940;
  assign n11771 = ~pi0934 & n11770;
  assign n11772 = pi0934 & ~n11770;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = pi1941 & ~n11773;
  assign n11775 = pi0934 & ~pi1941;
  assign n11776 = ~n11774 & ~n11775;
  assign po0985 = pi1838 & ~n11776;
  assign n11778 = pi0918 & pi0941;
  assign n11779 = ~pi0935 & n11778;
  assign n11780 = pi0935 & ~n11778;
  assign n11781 = ~n11779 & ~n11780;
  assign n11782 = pi1937 & ~n11781;
  assign n11783 = pi0935 & ~pi1937;
  assign n11784 = ~n11782 & ~n11783;
  assign po0986 = pi1164 & ~n11784;
  assign n11786 = pi0920 & pi0930;
  assign n11787 = ~pi0936 & n11786;
  assign n11788 = pi0936 & ~n11786;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = pi1939 & ~n11789;
  assign n11791 = pi0936 & ~pi1939;
  assign n11792 = ~n11790 & ~n11791;
  assign po0987 = pi1169 & ~n11792;
  assign n11794 = pi0922 & pi0944;
  assign n11795 = ~pi0937 & n11794;
  assign n11796 = pi0937 & ~n11794;
  assign n11797 = ~n11795 & ~n11796;
  assign n11798 = pi1940 & ~n11797;
  assign n11799 = pi0937 & ~pi1940;
  assign n11800 = ~n11798 & ~n11799;
  assign po0988 = pi1839 & ~n11800;
  assign n11802 = ~pi0816 & pi1153;
  assign n11803 = ~pi1856 & ~n11802;
  assign n11804 = pi0232 & n11803;
  assign n11805 = pi0938 & pi1145;
  assign n11806 = pi1145 & ~pi1931;
  assign n11807 = ~n11805 & ~n11806;
  assign n11808 = n11804 & ~n11807;
  assign po0989 = po1932 | n11808;
  assign n11810 = ~pi0867 & pi1163;
  assign n11811 = ~pi1877 & ~n11810;
  assign n11812 = pi0232 & n11811;
  assign n11813 = pi0939 & pi1036;
  assign n11814 = pi1036 & pi1952;
  assign n11815 = ~n11813 & ~n11814;
  assign n11816 = n11812 & ~n11815;
  assign po0990 = po1927 | n11816;
  assign n11818 = pi0940 & pi1838;
  assign n11819 = ~pi1941 & n11818;
  assign n11820 = pi0917 & ~pi0940;
  assign n11821 = ~pi0917 & pi0940;
  assign n11822 = ~n11820 & ~n11821;
  assign n11823 = pi1941 & ~n11822;
  assign n11824 = pi1838 & n11823;
  assign po0991 = n11819 | n11824;
  assign n11826 = pi0941 & pi1164;
  assign n11827 = ~pi1937 & n11826;
  assign n11828 = pi0918 & ~pi0941;
  assign n11829 = ~pi0918 & pi0941;
  assign n11830 = ~n11828 & ~n11829;
  assign n11831 = pi1937 & ~n11830;
  assign n11832 = pi1164 & n11831;
  assign po0992 = n11827 | n11832;
  assign n11834 = pi0942 & pi1035;
  assign n11835 = ~pi1938 & n11834;
  assign n11836 = pi0919 & ~pi0942;
  assign n11837 = ~pi0919 & pi0942;
  assign n11838 = ~n11836 & ~n11837;
  assign n11839 = pi1938 & ~n11838;
  assign n11840 = pi1035 & n11839;
  assign po0993 = n11835 | n11840;
  assign n11842 = pi0943 & pi1176;
  assign n11843 = ~pi1936 & n11842;
  assign n11844 = pi0921 & ~pi0943;
  assign n11845 = ~pi0921 & pi0943;
  assign n11846 = ~n11844 & ~n11845;
  assign n11847 = pi1936 & ~n11846;
  assign n11848 = pi1176 & n11847;
  assign po0994 = n11843 | n11848;
  assign n11850 = pi0944 & pi1839;
  assign n11851 = ~pi1940 & n11850;
  assign n11852 = pi0922 & ~pi0944;
  assign n11853 = ~pi0922 & pi0944;
  assign n11854 = ~n11852 & ~n11853;
  assign n11855 = pi1940 & ~n11854;
  assign n11856 = pi1839 & n11855;
  assign po0995 = n11851 | n11856;
  assign n11858 = pi0919 & pi0942;
  assign n11859 = ~pi0945 & n11858;
  assign n11860 = pi0945 & ~n11858;
  assign n11861 = ~n11859 & ~n11860;
  assign n11862 = pi1938 & ~n11861;
  assign n11863 = pi0945 & ~pi1938;
  assign n11864 = ~n11862 & ~n11863;
  assign po0996 = pi1035 & ~n11864;
  assign n11866 = pi1906 & ~pi2058;
  assign n11867 = pi0947 & pi2058;
  assign po0998 = n11866 | n11867;
  assign n11869 = pi1906 & ~pi2056;
  assign n11870 = pi0948 & pi2056;
  assign po0999 = n11869 | n11870;
  assign n11872 = pi1906 & ~pi2035;
  assign n11873 = pi0949 & pi2035;
  assign po1000 = n11872 | n11873;
  assign n11875 = pi1906 & ~pi2057;
  assign n11876 = pi0950 & pi2057;
  assign po1001 = n11875 | n11876;
  assign n11878 = pi1906 & ~pi2059;
  assign n11879 = pi0951 & pi2059;
  assign po1002 = n11878 | n11879;
  assign n11881 = pi0952 & ~pi1938;
  assign n11882 = ~pi0919 & ~pi0942;
  assign n11883 = pi0952 & ~n11882;
  assign n11884 = pi2174 & n11882;
  assign n11885 = ~n11883 & ~n11884;
  assign n11886 = pi1938 & ~n11885;
  assign po1003 = n11881 | n11886;
  assign n11888 = pi0953 & ~pi1938;
  assign n11889 = pi0953 & ~n11882;
  assign n11890 = pi2197 & n11882;
  assign n11891 = ~n11889 & ~n11890;
  assign n11892 = pi1938 & ~n11891;
  assign po1004 = n11888 | n11892;
  assign n11894 = pi0954 & ~pi1938;
  assign n11895 = pi0954 & ~n11882;
  assign n11896 = pi2196 & n11882;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = pi1938 & ~n11897;
  assign po1005 = n11894 | n11898;
  assign n11900 = pi0955 & ~pi1938;
  assign n11901 = pi0955 & ~n11882;
  assign n11902 = pi2179 & n11882;
  assign n11903 = ~n11901 & ~n11902;
  assign n11904 = pi1938 & ~n11903;
  assign po1006 = n11900 | n11904;
  assign n11906 = pi0956 & ~pi1938;
  assign n11907 = pi0956 & ~n11882;
  assign n11908 = pi2176 & n11882;
  assign n11909 = ~n11907 & ~n11908;
  assign n11910 = pi1938 & ~n11909;
  assign po1007 = n11906 | n11910;
  assign n11912 = pi0957 & ~pi1938;
  assign n11913 = pi0957 & ~n11882;
  assign n11914 = pi2169 & n11882;
  assign n11915 = ~n11913 & ~n11914;
  assign n11916 = pi1938 & ~n11915;
  assign po1008 = n11912 | n11916;
  assign n11918 = pi0958 & ~pi1938;
  assign n11919 = pi0958 & ~n11882;
  assign n11920 = pi2173 & n11882;
  assign n11921 = ~n11919 & ~n11920;
  assign n11922 = pi1938 & ~n11921;
  assign po1009 = n11918 | n11922;
  assign n11924 = pi0959 & ~pi1938;
  assign n11925 = pi0959 & ~n11882;
  assign n11926 = pi2167 & n11882;
  assign n11927 = ~n11925 & ~n11926;
  assign n11928 = pi1938 & ~n11927;
  assign po1010 = n11924 | n11928;
  assign n11930 = pi0960 & ~pi1938;
  assign n11931 = pi0960 & ~n11882;
  assign n11932 = pi2166 & n11882;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = pi1938 & ~n11933;
  assign po1011 = n11930 | n11934;
  assign n11936 = pi0961 & ~pi1938;
  assign n11937 = pi0961 & ~n11882;
  assign n11938 = pi2192 & n11882;
  assign n11939 = ~n11937 & ~n11938;
  assign n11940 = pi1938 & ~n11939;
  assign po1012 = n11936 | n11940;
  assign n11942 = pi0962 & ~pi1939;
  assign n11943 = ~pi0920 & ~pi0930;
  assign n11944 = pi0962 & ~n11943;
  assign n11945 = pi2174 & n11943;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = pi1939 & ~n11946;
  assign po1013 = n11942 | n11947;
  assign n11949 = pi0963 & ~pi1939;
  assign n11950 = pi0963 & ~n11943;
  assign n11951 = pi2197 & n11943;
  assign n11952 = ~n11950 & ~n11951;
  assign n11953 = pi1939 & ~n11952;
  assign po1014 = n11949 | n11953;
  assign n11955 = pi0964 & ~pi1939;
  assign n11956 = pi0964 & ~n11943;
  assign n11957 = pi2196 & n11943;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = pi1939 & ~n11958;
  assign po1015 = n11955 | n11959;
  assign n11961 = pi0965 & ~pi1939;
  assign n11962 = pi0965 & ~n11943;
  assign n11963 = pi2179 & n11943;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = pi1939 & ~n11964;
  assign po1016 = n11961 | n11965;
  assign n11967 = pi0966 & ~pi1939;
  assign n11968 = pi0966 & ~n11943;
  assign n11969 = pi2176 & n11943;
  assign n11970 = ~n11968 & ~n11969;
  assign n11971 = pi1939 & ~n11970;
  assign po1017 = n11967 | n11971;
  assign n11973 = pi0967 & ~pi1939;
  assign n11974 = pi0967 & ~n11943;
  assign n11975 = pi2169 & n11943;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = pi1939 & ~n11976;
  assign po1018 = n11973 | n11977;
  assign n11979 = pi0968 & ~pi1939;
  assign n11980 = pi0968 & ~n11943;
  assign n11981 = pi2173 & n11943;
  assign n11982 = ~n11980 & ~n11981;
  assign n11983 = pi1939 & ~n11982;
  assign po1019 = n11979 | n11983;
  assign n11985 = pi0969 & ~pi1939;
  assign n11986 = pi0969 & ~n11943;
  assign n11987 = pi2167 & n11943;
  assign n11988 = ~n11986 & ~n11987;
  assign n11989 = pi1939 & ~n11988;
  assign po1020 = n11985 | n11989;
  assign n11991 = pi0970 & ~pi1939;
  assign n11992 = pi0970 & ~n11943;
  assign n11993 = pi2166 & n11943;
  assign n11994 = ~n11992 & ~n11993;
  assign n11995 = pi1939 & ~n11994;
  assign po1021 = n11991 | n11995;
  assign n11997 = pi0971 & ~pi1939;
  assign n11998 = pi0971 & ~n11943;
  assign n11999 = pi2192 & n11943;
  assign n12000 = ~n11998 & ~n11999;
  assign n12001 = pi1939 & ~n12000;
  assign po1022 = n11997 | n12001;
  assign n12003 = pi0972 & ~pi1936;
  assign n12004 = ~pi0921 & ~pi0943;
  assign n12005 = pi0972 & ~n12004;
  assign n12006 = pi2174 & n12004;
  assign n12007 = ~n12005 & ~n12006;
  assign n12008 = pi1936 & ~n12007;
  assign po1023 = n12003 | n12008;
  assign n12010 = pi0973 & ~pi1936;
  assign n12011 = pi0973 & ~n12004;
  assign n12012 = pi2197 & n12004;
  assign n12013 = ~n12011 & ~n12012;
  assign n12014 = pi1936 & ~n12013;
  assign po1024 = n12010 | n12014;
  assign n12016 = pi0974 & ~pi1936;
  assign n12017 = pi0974 & ~n12004;
  assign n12018 = pi2196 & n12004;
  assign n12019 = ~n12017 & ~n12018;
  assign n12020 = pi1936 & ~n12019;
  assign po1025 = n12016 | n12020;
  assign n12022 = pi0975 & ~pi1936;
  assign n12023 = pi0975 & ~n12004;
  assign n12024 = pi2179 & n12004;
  assign n12025 = ~n12023 & ~n12024;
  assign n12026 = pi1936 & ~n12025;
  assign po1026 = n12022 | n12026;
  assign n12028 = pi0976 & ~pi1936;
  assign n12029 = pi0976 & ~n12004;
  assign n12030 = pi2176 & n12004;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = pi1936 & ~n12031;
  assign po1027 = n12028 | n12032;
  assign n12034 = pi0977 & ~pi1936;
  assign n12035 = pi0977 & ~n12004;
  assign n12036 = pi2169 & n12004;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = pi1936 & ~n12037;
  assign po1028 = n12034 | n12038;
  assign n12040 = pi0978 & ~pi1936;
  assign n12041 = pi0978 & ~n12004;
  assign n12042 = pi2173 & n12004;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = pi1936 & ~n12043;
  assign po1029 = n12040 | n12044;
  assign n12046 = pi0979 & ~pi1936;
  assign n12047 = pi0979 & ~n12004;
  assign n12048 = pi2167 & n12004;
  assign n12049 = ~n12047 & ~n12048;
  assign n12050 = pi1936 & ~n12049;
  assign po1030 = n12046 | n12050;
  assign n12052 = pi0980 & ~pi1936;
  assign n12053 = pi0980 & ~n12004;
  assign n12054 = pi2166 & n12004;
  assign n12055 = ~n12053 & ~n12054;
  assign n12056 = pi1936 & ~n12055;
  assign po1031 = n12052 | n12056;
  assign n12058 = pi0981 & ~pi1936;
  assign n12059 = pi0981 & ~n12004;
  assign n12060 = pi2192 & n12004;
  assign n12061 = ~n12059 & ~n12060;
  assign n12062 = pi1936 & ~n12061;
  assign po1032 = n12058 | n12062;
  assign n12064 = pi0982 & ~pi1940;
  assign n12065 = ~pi0922 & ~pi0944;
  assign n12066 = pi0982 & ~n12065;
  assign n12067 = pi2174 & n12065;
  assign n12068 = ~n12066 & ~n12067;
  assign n12069 = pi1940 & ~n12068;
  assign po1033 = n12064 | n12069;
  assign n12071 = pi0983 & ~pi1940;
  assign n12072 = pi0983 & ~n12065;
  assign n12073 = pi2197 & n12065;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = pi1940 & ~n12074;
  assign po1034 = n12071 | n12075;
  assign n12077 = pi0984 & ~pi1940;
  assign n12078 = pi0984 & ~n12065;
  assign n12079 = pi2196 & n12065;
  assign n12080 = ~n12078 & ~n12079;
  assign n12081 = pi1940 & ~n12080;
  assign po1035 = n12077 | n12081;
  assign n12083 = pi0985 & ~pi1940;
  assign n12084 = pi0985 & ~n12065;
  assign n12085 = pi2179 & n12065;
  assign n12086 = ~n12084 & ~n12085;
  assign n12087 = pi1940 & ~n12086;
  assign po1036 = n12083 | n12087;
  assign n12089 = pi0986 & ~pi1940;
  assign n12090 = pi0986 & ~n12065;
  assign n12091 = pi2176 & n12065;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = pi1940 & ~n12092;
  assign po1037 = n12089 | n12093;
  assign n12095 = pi0987 & ~pi1940;
  assign n12096 = pi0987 & ~n12065;
  assign n12097 = pi2169 & n12065;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = pi1940 & ~n12098;
  assign po1038 = n12095 | n12099;
  assign n12101 = pi0988 & ~pi1940;
  assign n12102 = pi0988 & ~n12065;
  assign n12103 = pi2173 & n12065;
  assign n12104 = ~n12102 & ~n12103;
  assign n12105 = pi1940 & ~n12104;
  assign po1039 = n12101 | n12105;
  assign n12107 = pi0989 & ~pi1940;
  assign n12108 = pi0989 & ~n12065;
  assign n12109 = pi2167 & n12065;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = pi1940 & ~n12110;
  assign po1040 = n12107 | n12111;
  assign n12113 = pi0990 & ~pi1940;
  assign n12114 = pi0990 & ~n12065;
  assign n12115 = pi2166 & n12065;
  assign n12116 = ~n12114 & ~n12115;
  assign n12117 = pi1940 & ~n12116;
  assign po1041 = n12113 | n12117;
  assign n12119 = pi0991 & ~pi1940;
  assign n12120 = pi0991 & ~n12065;
  assign n12121 = pi2192 & n12065;
  assign n12122 = ~n12120 & ~n12121;
  assign n12123 = pi1940 & ~n12122;
  assign po1042 = n12119 | n12123;
  assign n12125 = pi0992 & ~pi1937;
  assign n12126 = ~pi0918 & ~pi0941;
  assign n12127 = pi0992 & ~n12126;
  assign n12128 = pi2172 & n12126;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = pi1937 & ~n12129;
  assign po1043 = n12125 | n12130;
  assign n12132 = pi0993 & ~pi1937;
  assign n12133 = pi0993 & ~n12126;
  assign n12134 = pi2168 & n12126;
  assign n12135 = ~n12133 & ~n12134;
  assign n12136 = pi1937 & ~n12135;
  assign po1044 = n12132 | n12136;
  assign n12138 = pi0994 & ~pi1937;
  assign n12139 = pi0994 & ~n12126;
  assign n12140 = pi2178 & n12126;
  assign n12141 = ~n12139 & ~n12140;
  assign n12142 = pi1937 & ~n12141;
  assign po1045 = n12138 | n12142;
  assign n12144 = pi0995 & ~pi1941;
  assign n12145 = ~pi0917 & ~pi0940;
  assign n12146 = pi0995 & ~n12145;
  assign n12147 = pi2186 & n12145;
  assign n12148 = ~n12146 & ~n12147;
  assign n12149 = pi1941 & ~n12148;
  assign po1046 = n12144 | n12149;
  assign n12151 = pi0996 & ~pi1941;
  assign n12152 = pi0996 & ~n12145;
  assign n12153 = pi2172 & n12145;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = pi1941 & ~n12154;
  assign po1047 = n12151 | n12155;
  assign n12157 = pi0997 & ~pi1941;
  assign n12158 = pi0997 & ~n12145;
  assign n12159 = pi2168 & n12145;
  assign n12160 = ~n12158 & ~n12159;
  assign n12161 = pi1941 & ~n12160;
  assign po1048 = n12157 | n12161;
  assign n12163 = pi0998 & ~pi1941;
  assign n12164 = pi0998 & ~n12145;
  assign n12165 = pi2193 & n12145;
  assign n12166 = ~n12164 & ~n12165;
  assign n12167 = pi1941 & ~n12166;
  assign po1049 = n12163 | n12167;
  assign n12169 = pi0999 & ~pi1937;
  assign n12170 = pi0999 & ~n12126;
  assign n12171 = pi2198 & n12126;
  assign n12172 = ~n12170 & ~n12171;
  assign n12173 = pi1937 & ~n12172;
  assign po1050 = n12169 | n12173;
  assign n12175 = pi1000 & ~pi1937;
  assign n12176 = pi1000 & ~n12126;
  assign n12177 = pi2187 & n12126;
  assign n12178 = ~n12176 & ~n12177;
  assign n12179 = pi1937 & ~n12178;
  assign po1051 = n12175 | n12179;
  assign n12181 = pi1001 & ~pi1941;
  assign n12182 = pi1001 & ~n12145;
  assign n12183 = pi2170 & n12145;
  assign n12184 = ~n12182 & ~n12183;
  assign n12185 = pi1941 & ~n12184;
  assign po1052 = n12181 | n12185;
  assign n12187 = pi1002 & ~pi1941;
  assign n12188 = pi1002 & ~n12145;
  assign n12189 = pi2182 & n12145;
  assign n12190 = ~n12188 & ~n12189;
  assign n12191 = pi1941 & ~n12190;
  assign po1053 = n12187 | n12191;
  assign n12193 = pi1003 & ~pi1941;
  assign n12194 = pi1003 & ~n12145;
  assign n12195 = pi2175 & n12145;
  assign n12196 = ~n12194 & ~n12195;
  assign n12197 = pi1941 & ~n12196;
  assign po1054 = n12193 | n12197;
  assign n12199 = pi1004 & ~pi1941;
  assign n12200 = pi1004 & ~n12145;
  assign n12201 = pi2177 & n12145;
  assign n12202 = ~n12200 & ~n12201;
  assign n12203 = pi1941 & ~n12202;
  assign po1055 = n12199 | n12203;
  assign n12205 = pi1005 & ~pi1937;
  assign n12206 = pi1005 & ~n12126;
  assign n12207 = pi2181 & n12126;
  assign n12208 = ~n12206 & ~n12207;
  assign n12209 = pi1937 & ~n12208;
  assign po1056 = n12205 | n12209;
  assign n12211 = pi1006 & ~pi1941;
  assign n12212 = pi1006 & ~n12145;
  assign n12213 = pi2167 & n12145;
  assign n12214 = ~n12212 & ~n12213;
  assign n12215 = pi1941 & ~n12214;
  assign po1057 = n12211 | n12215;
  assign n12217 = pi1007 & ~pi1941;
  assign n12218 = pi1007 & ~n12145;
  assign n12219 = pi2188 & n12145;
  assign n12220 = ~n12218 & ~n12219;
  assign n12221 = pi1941 & ~n12220;
  assign po1058 = n12217 | n12221;
  assign n12223 = pi1008 & ~pi1937;
  assign n12224 = pi1008 & ~n12126;
  assign n12225 = pi2191 & n12126;
  assign n12226 = ~n12224 & ~n12225;
  assign n12227 = pi1937 & ~n12226;
  assign po1059 = n12223 | n12227;
  assign n12229 = pi1009 & ~pi1937;
  assign n12230 = pi1009 & ~n12126;
  assign n12231 = pi2175 & n12126;
  assign n12232 = ~n12230 & ~n12231;
  assign n12233 = pi1937 & ~n12232;
  assign po1060 = n12229 | n12233;
  assign n12235 = pi1010 & ~pi1937;
  assign n12236 = pi1010 & ~n12126;
  assign n12237 = pi2184 & n12126;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = pi1937 & ~n12238;
  assign po1061 = n12235 | n12239;
  assign n12241 = pi1011 & ~pi1937;
  assign n12242 = pi1011 & ~n12126;
  assign n12243 = pi2188 & n12126;
  assign n12244 = ~n12242 & ~n12243;
  assign n12245 = pi1937 & ~n12244;
  assign po1062 = n12241 | n12245;
  assign n12247 = ~pi1989 & pi2240;
  assign po1956 = n11504 & n12247;
  assign n12249 = pi1012 & ~po1956;
  assign n12250 = pi2176 & po1956;
  assign po1063 = n12249 | n12250;
  assign n12252 = pi1013 & ~pi1937;
  assign n12253 = pi1013 & ~n12126;
  assign n12254 = pi2193 & n12126;
  assign n12255 = ~n12253 & ~n12254;
  assign n12256 = pi1937 & ~n12255;
  assign po1064 = n12252 | n12256;
  assign n12258 = pi1014 & ~pi1941;
  assign n12259 = pi2189 & n11821;
  assign n12260 = pi1014 & ~n11821;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = pi1941 & ~n12261;
  assign po1065 = n12258 | n12262;
  assign n12264 = pi1015 & ~pi1940;
  assign n12265 = pi1015 & ~n12065;
  assign n12266 = pi2185 & n12065;
  assign n12267 = ~n12265 & ~n12266;
  assign n12268 = pi1940 & ~n12267;
  assign po1066 = n12264 | n12268;
  assign n12270 = pi1016 & ~pi1941;
  assign n12271 = pi2190 & n11821;
  assign n12272 = pi1016 & ~n11821;
  assign n12273 = ~n12271 & ~n12272;
  assign n12274 = pi1941 & ~n12273;
  assign po1067 = n12270 | n12274;
  assign n12276 = pi1017 & ~pi1941;
  assign n12277 = pi2182 & n11821;
  assign n12278 = pi1017 & ~n11821;
  assign n12279 = ~n12277 & ~n12278;
  assign n12280 = pi1941 & ~n12279;
  assign po1068 = n12276 | n12280;
  assign n12282 = pi1018 & ~pi1938;
  assign n12283 = pi2196 & n11837;
  assign n12284 = pi1018 & ~n11837;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = pi1938 & ~n12285;
  assign po1069 = n12282 | n12286;
  assign n12288 = pi1019 & ~pi1939;
  assign n12289 = pi2170 & n11745;
  assign n12290 = pi1019 & ~n11745;
  assign n12291 = ~n12289 & ~n12290;
  assign n12292 = pi1939 & ~n12291;
  assign po1070 = n12288 | n12292;
  assign n12294 = ~pi1989 & pi2238;
  assign n12295 = n5418 & n12294;
  assign n12296 = pi2172 & n12295;
  assign n12297 = pi1020 & ~n12295;
  assign po1071 = n12296 | n12297;
  assign n12299 = pi1021 & ~pi1939;
  assign n12300 = pi2176 & n11745;
  assign n12301 = pi1021 & ~n11745;
  assign n12302 = ~n12300 & ~n12301;
  assign n12303 = pi1939 & ~n12302;
  assign po1072 = n12299 | n12303;
  assign n12305 = pi1022 & ~pi1939;
  assign n12306 = pi2178 & n11745;
  assign n12307 = pi1022 & ~n11745;
  assign n12308 = ~n12306 & ~n12307;
  assign n12309 = pi1939 & ~n12308;
  assign po1073 = n12305 | n12309;
  assign n12311 = pi1023 & ~pi1939;
  assign n12312 = pi2179 & n11745;
  assign n12313 = pi1023 & ~n11745;
  assign n12314 = ~n12312 & ~n12313;
  assign n12315 = pi1939 & ~n12314;
  assign po1074 = n12311 | n12315;
  assign n12317 = pi1024 & ~pi1939;
  assign n12318 = pi2172 & n11745;
  assign n12319 = pi1024 & ~n11745;
  assign n12320 = ~n12318 & ~n12319;
  assign n12321 = pi1939 & ~n12320;
  assign po1075 = n12317 | n12321;
  assign n12323 = pi1025 & ~pi1937;
  assign n12324 = pi2176 & n11828;
  assign n12325 = pi1025 & ~n11828;
  assign n12326 = ~n12324 & ~n12325;
  assign n12327 = pi1937 & ~n12326;
  assign po1076 = n12323 | n12327;
  assign n12329 = pi1026 & ~pi1941;
  assign n12330 = pi2185 & n11821;
  assign n12331 = pi1026 & ~n11821;
  assign n12332 = ~n12330 & ~n12331;
  assign n12333 = pi1941 & ~n12332;
  assign po1077 = n12329 | n12333;
  assign n12335 = pi1027 & ~pi1938;
  assign n12336 = pi2192 & n11858;
  assign n12337 = pi1027 & ~n11858;
  assign n12338 = ~n12336 & ~n12337;
  assign n12339 = pi1938 & ~n12338;
  assign po1078 = n12335 | n12339;
  assign n12341 = pi1028 & ~pi1938;
  assign n12342 = pi2188 & n11858;
  assign n12343 = pi1028 & ~n11858;
  assign n12344 = ~n12342 & ~n12343;
  assign n12345 = pi1938 & ~n12344;
  assign po1079 = n12341 | n12345;
  assign n12347 = pi1029 & ~pi1938;
  assign n12348 = pi2177 & n11858;
  assign n12349 = pi1029 & ~n11858;
  assign n12350 = ~n12348 & ~n12349;
  assign n12351 = pi1938 & ~n12350;
  assign po1080 = n12347 | n12351;
  assign n12353 = pi1030 & ~pi1941;
  assign n12354 = pi1030 & ~n12145;
  assign n12355 = pi2178 & n12145;
  assign n12356 = ~n12354 & ~n12355;
  assign n12357 = pi1941 & ~n12356;
  assign po1081 = n12353 | n12357;
  assign n12359 = pi1031 & ~pi1937;
  assign n12360 = pi1031 & ~n12126;
  assign n12361 = pi2196 & n12126;
  assign n12362 = ~n12360 & ~n12361;
  assign n12363 = pi1937 & ~n12362;
  assign po1082 = n12359 | n12363;
  assign n12365 = pi1032 & ~pi1938;
  assign n12366 = pi2171 & n11858;
  assign n12367 = pi1032 & ~n11858;
  assign n12368 = ~n12366 & ~n12367;
  assign n12369 = pi1938 & ~n12368;
  assign po1083 = n12365 | n12369;
  assign n12371 = pi1033 & ~pi1938;
  assign n12372 = pi2181 & n11858;
  assign n12373 = pi1033 & ~n11858;
  assign n12374 = ~n12372 & ~n12373;
  assign n12375 = pi1938 & ~n12374;
  assign po1084 = n12371 | n12375;
  assign n12377 = pi1034 & ~pi1941;
  assign n12378 = pi2184 & n11820;
  assign n12379 = pi1034 & ~n11820;
  assign n12380 = ~n12378 & ~n12379;
  assign n12381 = pi1941 & ~n12380;
  assign po1085 = n12377 | n12381;
  assign n12383 = pi2195 & n12295;
  assign n12384 = pi1035 & ~n12295;
  assign po1086 = n12383 | n12384;
  assign n12386 = ~pi1989 & ~pi2240;
  assign n12387 = n11534 & n12386;
  assign n12388 = pi1036 & ~n12387;
  assign n12389 = pi2195 & n12387;
  assign po1087 = n12388 | n12389;
  assign n12391 = pi1037 & ~pi1941;
  assign n12392 = pi2174 & n11821;
  assign n12393 = pi1037 & ~n11821;
  assign n12394 = ~n12392 & ~n12393;
  assign n12395 = pi1941 & ~n12394;
  assign po1088 = n12391 | n12395;
  assign n12397 = pi1038 & ~pi1937;
  assign n12398 = pi2179 & n11828;
  assign n12399 = pi1038 & ~n11828;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = pi1937 & ~n12400;
  assign po1089 = n12397 | n12401;
  assign n12403 = pi1039 & ~pi1938;
  assign n12404 = pi2192 & n11837;
  assign n12405 = pi1039 & ~n11837;
  assign n12406 = ~n12404 & ~n12405;
  assign n12407 = pi1938 & ~n12406;
  assign po1090 = n12403 | n12407;
  assign n12409 = pi1040 & ~pi1938;
  assign n12410 = pi2196 & n11858;
  assign n12411 = pi1040 & ~n11858;
  assign n12412 = ~n12410 & ~n12411;
  assign n12413 = pi1938 & ~n12412;
  assign po1091 = n12409 | n12413;
  assign n12415 = pi1041 & ~pi1938;
  assign n12416 = pi2168 & n11858;
  assign n12417 = pi1041 & ~n11858;
  assign n12418 = ~n12416 & ~n12417;
  assign n12419 = pi1938 & ~n12418;
  assign po1092 = n12415 | n12419;
  assign n12421 = pi1042 & ~pi1938;
  assign n12422 = pi2188 & n11837;
  assign n12423 = pi1042 & ~n11837;
  assign n12424 = ~n12422 & ~n12423;
  assign n12425 = pi1938 & ~n12424;
  assign po1093 = n12421 | n12425;
  assign n12427 = pi1043 & ~pi1937;
  assign n12428 = pi2178 & n11828;
  assign n12429 = pi1043 & ~n11828;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = pi1937 & ~n12430;
  assign po1094 = n12427 | n12431;
  assign n12433 = pi1044 & ~pi1938;
  assign n12434 = pi2177 & n11837;
  assign n12435 = pi1044 & ~n11837;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = pi1938 & ~n12436;
  assign po1095 = n12433 | n12437;
  assign n12439 = pi1045 & ~pi1938;
  assign n12440 = pi2181 & n11837;
  assign n12441 = pi1045 & ~n11837;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = pi1938 & ~n12442;
  assign po1096 = n12439 | n12443;
  assign n12445 = pi1046 & ~pi1938;
  assign n12446 = pi2171 & n11837;
  assign n12447 = pi1046 & ~n11837;
  assign n12448 = ~n12446 & ~n12447;
  assign n12449 = pi1938 & ~n12448;
  assign po1097 = n12445 | n12449;
  assign n12451 = pi1047 & ~pi1940;
  assign n12452 = pi1047 & ~n12065;
  assign n12453 = pi2177 & n12065;
  assign n12454 = ~n12452 & ~n12453;
  assign n12455 = pi1940 & ~n12454;
  assign po1098 = n12451 | n12455;
  assign n12457 = pi1048 & ~pi1937;
  assign n12458 = pi2191 & n11829;
  assign n12459 = pi1048 & ~n11829;
  assign n12460 = ~n12458 & ~n12459;
  assign n12461 = pi1937 & ~n12460;
  assign po1099 = n12457 | n12461;
  assign n12463 = pi1049 & ~pi1941;
  assign n12464 = pi2187 & n11820;
  assign n12465 = pi1049 & ~n11820;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = pi1941 & ~n12466;
  assign po1100 = n12463 | n12467;
  assign n12469 = pi1050 & ~pi1937;
  assign n12470 = pi2172 & n11828;
  assign n12471 = pi1050 & ~n11828;
  assign n12472 = ~n12470 & ~n12471;
  assign n12473 = pi1937 & ~n12472;
  assign po1101 = n12469 | n12473;
  assign n12475 = pi1051 & ~pi1941;
  assign n12476 = pi2194 & n11820;
  assign n12477 = pi1051 & ~n11820;
  assign n12478 = ~n12476 & ~n12477;
  assign n12479 = pi1941 & ~n12478;
  assign po1102 = n12475 | n12479;
  assign n12481 = pi1052 & ~pi1938;
  assign n12482 = pi2168 & n11837;
  assign n12483 = pi1052 & ~n11837;
  assign n12484 = ~n12482 & ~n12483;
  assign n12485 = pi1938 & ~n12484;
  assign po1103 = n12481 | n12485;
  assign n12487 = pi1053 & ~pi1938;
  assign n12488 = pi2177 & n11836;
  assign n12489 = pi1053 & ~n11836;
  assign n12490 = ~n12488 & ~n12489;
  assign n12491 = pi1938 & ~n12490;
  assign po1104 = n12487 | n12491;
  assign n12493 = pi1054 & ~pi1938;
  assign n12494 = pi2192 & n11836;
  assign n12495 = pi1054 & ~n11836;
  assign n12496 = ~n12494 & ~n12495;
  assign n12497 = pi1938 & ~n12496;
  assign po1105 = n12493 | n12497;
  assign n12499 = pi1055 & ~pi1938;
  assign n12500 = pi2188 & n11836;
  assign n12501 = pi1055 & ~n11836;
  assign n12502 = ~n12500 & ~n12501;
  assign n12503 = pi1938 & ~n12502;
  assign po1106 = n12499 | n12503;
  assign n12505 = pi1056 & ~pi1938;
  assign n12506 = pi2181 & n11836;
  assign n12507 = pi1056 & ~n11836;
  assign n12508 = ~n12506 & ~n12507;
  assign n12509 = pi1938 & ~n12508;
  assign po1107 = n12505 | n12509;
  assign n12511 = pi1057 & ~pi1941;
  assign n12512 = pi2182 & n11820;
  assign n12513 = pi1057 & ~n11820;
  assign n12514 = ~n12512 & ~n12513;
  assign n12515 = pi1941 & ~n12514;
  assign po1108 = n12511 | n12515;
  assign n12517 = pi1058 & ~pi1937;
  assign n12518 = pi1058 & ~n12126;
  assign n12519 = pi2174 & n12126;
  assign n12520 = ~n12518 & ~n12519;
  assign n12521 = pi1937 & ~n12520;
  assign po1109 = n12517 | n12521;
  assign n12523 = pi1059 & ~pi1941;
  assign n12524 = pi2190 & n11820;
  assign n12525 = pi1059 & ~n11820;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = pi1941 & ~n12526;
  assign po1110 = n12523 | n12527;
  assign n12529 = pi1060 & ~pi1938;
  assign n12530 = pi2171 & n11836;
  assign n12531 = pi1060 & ~n11836;
  assign n12532 = ~n12530 & ~n12531;
  assign n12533 = pi1938 & ~n12532;
  assign po1111 = n12529 | n12533;
  assign n12535 = pi1061 & ~pi1938;
  assign n12536 = pi2196 & n11836;
  assign n12537 = pi1061 & ~n11836;
  assign n12538 = ~n12536 & ~n12537;
  assign n12539 = pi1938 & ~n12538;
  assign po1112 = n12535 | n12539;
  assign n12541 = pi1062 & ~pi1940;
  assign n12542 = pi1062 & ~n12065;
  assign n12543 = pi2184 & n12065;
  assign n12544 = ~n12542 & ~n12543;
  assign n12545 = pi1940 & ~n12544;
  assign po1113 = n12541 | n12545;
  assign n12547 = pi1063 & ~pi1940;
  assign n12548 = pi2190 & n11852;
  assign n12549 = pi1063 & ~n11852;
  assign n12550 = ~n12548 & ~n12549;
  assign n12551 = pi1940 & ~n12550;
  assign po1114 = n12547 | n12551;
  assign n12553 = pi1064 & ~pi1937;
  assign n12554 = pi2194 & n11778;
  assign n12555 = pi1064 & ~n11778;
  assign n12556 = ~n12554 & ~n12555;
  assign n12557 = pi1937 & ~n12556;
  assign po1115 = n12553 | n12557;
  assign n12559 = pi1065 & ~pi1938;
  assign n12560 = pi2168 & n11836;
  assign n12561 = pi1065 & ~n11836;
  assign n12562 = ~n12560 & ~n12561;
  assign n12563 = pi1938 & ~n12562;
  assign po1116 = n12559 | n12563;
  assign n12565 = pi1066 & ~pi1940;
  assign n12566 = pi2194 & n11794;
  assign n12567 = pi1066 & ~n11794;
  assign n12568 = ~n12566 & ~n12567;
  assign n12569 = pi1940 & ~n12568;
  assign po1117 = n12565 | n12569;
  assign n12571 = pi1067 & ~pi1941;
  assign n12572 = pi2197 & n11820;
  assign n12573 = pi1067 & ~n11820;
  assign n12574 = ~n12572 & ~n12573;
  assign n12575 = pi1941 & ~n12574;
  assign po1118 = n12571 | n12575;
  assign n12577 = pi1068 & ~pi1941;
  assign n12578 = pi2189 & n11820;
  assign n12579 = pi1068 & ~n11820;
  assign n12580 = ~n12578 & ~n12579;
  assign n12581 = pi1941 & ~n12580;
  assign po1119 = n12577 | n12581;
  assign n12583 = pi1069 & ~pi1937;
  assign n12584 = pi2184 & n11778;
  assign n12585 = pi1069 & ~n11778;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = pi1937 & ~n12586;
  assign po1120 = n12583 | n12587;
  assign n12589 = pi1070 & ~pi1937;
  assign n12590 = pi2176 & n11778;
  assign n12591 = pi1070 & ~n11778;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = pi1937 & ~n12592;
  assign po1121 = n12589 | n12593;
  assign n12595 = pi1071 & ~pi1937;
  assign n12596 = pi2177 & n11778;
  assign n12597 = pi1071 & ~n11778;
  assign n12598 = ~n12596 & ~n12597;
  assign n12599 = pi1937 & ~n12598;
  assign po1122 = n12595 | n12599;
  assign n12601 = pi1072 & ~pi1937;
  assign n12602 = pi2181 & n11778;
  assign n12603 = pi1072 & ~n11778;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = pi1937 & ~n12604;
  assign po1123 = n12601 | n12605;
  assign n12607 = pi1073 & ~pi1940;
  assign n12608 = pi1073 & ~n12065;
  assign n12609 = pi2171 & n12065;
  assign n12610 = ~n12608 & ~n12609;
  assign n12611 = pi1940 & ~n12610;
  assign po1124 = n12607 | n12611;
  assign n12613 = pi1074 & ~pi1937;
  assign n12614 = pi2179 & n11778;
  assign n12615 = pi1074 & ~n11778;
  assign n12616 = ~n12614 & ~n12615;
  assign n12617 = pi1937 & ~n12616;
  assign po1125 = n12613 | n12617;
  assign n12619 = pi1081 & ~pi1936;
  assign n12620 = pi1081 & ~n12004;
  assign n12621 = pi2168 & n12004;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = pi1936 & ~n12622;
  assign po1132 = n12619 | n12623;
  assign n12625 = pi1082 & ~pi1941;
  assign n12626 = pi2183 & n11820;
  assign n12627 = pi1082 & ~n11820;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = pi1941 & ~n12628;
  assign po1133 = n12625 | n12629;
  assign n12631 = pi1083 & ~pi1940;
  assign n12632 = pi2166 & n11794;
  assign n12633 = pi1083 & ~n11794;
  assign n12634 = ~n12632 & ~n12633;
  assign n12635 = pi1940 & ~n12634;
  assign po1134 = n12631 | n12635;
  assign n12637 = pi1084 & ~pi1937;
  assign n12638 = pi2178 & n11778;
  assign n12639 = pi1084 & ~n11778;
  assign n12640 = ~n12638 & ~n12639;
  assign n12641 = pi1937 & ~n12640;
  assign po1135 = n12637 | n12641;
  assign n12643 = pi1085 & ~pi1937;
  assign n12644 = pi2172 & n11778;
  assign n12645 = pi1085 & ~n11778;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = pi1937 & ~n12646;
  assign po1136 = n12643 | n12647;
  assign n12649 = pi1086 & ~pi1937;
  assign n12650 = pi2195 & n11829;
  assign n12651 = pi1086 & ~n11829;
  assign n12652 = ~n12650 & ~n12651;
  assign n12653 = pi1937 & ~n12652;
  assign po1137 = n12649 | n12653;
  assign n12655 = pi1087 & ~pi1940;
  assign n12656 = pi1087 & ~n12065;
  assign n12657 = pi2168 & n12065;
  assign n12658 = ~n12656 & ~n12657;
  assign n12659 = pi1940 & ~n12658;
  assign po1138 = n12655 | n12659;
  assign n12661 = pi1088 & ~pi1940;
  assign n12662 = pi2197 & n11794;
  assign n12663 = pi1088 & ~n11794;
  assign n12664 = ~n12662 & ~n12663;
  assign n12665 = pi1940 & ~n12664;
  assign po1139 = n12661 | n12665;
  assign n12667 = pi1089 & ~pi1940;
  assign n12668 = pi2190 & n11794;
  assign n12669 = pi1089 & ~n11794;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = pi1940 & ~n12670;
  assign po1140 = n12667 | n12671;
  assign n12673 = pi1090 & ~pi1940;
  assign n12674 = pi2175 & n11794;
  assign n12675 = pi1090 & ~n11794;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = pi1940 & ~n12676;
  assign po1141 = n12673 | n12677;
  assign n12679 = pi1091 & ~pi1937;
  assign n12680 = pi2170 & n11829;
  assign n12681 = pi1091 & ~n11829;
  assign n12682 = ~n12680 & ~n12681;
  assign n12683 = pi1937 & ~n12682;
  assign po1142 = n12679 | n12683;
  assign n12685 = pi1092 & ~pi1937;
  assign n12686 = pi2176 & n11829;
  assign n12687 = pi1092 & ~n11829;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = pi1937 & ~n12688;
  assign po1143 = n12685 | n12689;
  assign n12691 = pi1093 & ~pi1937;
  assign n12692 = pi2189 & n11829;
  assign n12693 = pi1093 & ~n11829;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = pi1937 & ~n12694;
  assign po1144 = n12691 | n12695;
  assign n12697 = pi1094 & ~pi1941;
  assign n12698 = pi2195 & n11770;
  assign n12699 = pi1094 & ~n11770;
  assign n12700 = ~n12698 & ~n12699;
  assign n12701 = pi1941 & ~n12700;
  assign po1145 = n12697 | n12701;
  assign n12703 = pi1095 & ~pi1941;
  assign n12704 = pi2184 & n11770;
  assign n12705 = pi1095 & ~n11770;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = pi1941 & ~n12706;
  assign po1146 = n12703 | n12707;
  assign n12709 = pi1096 & ~pi1940;
  assign n12710 = pi2187 & n11794;
  assign n12711 = pi1096 & ~n11794;
  assign n12712 = ~n12710 & ~n12711;
  assign n12713 = pi1940 & ~n12712;
  assign po1147 = n12709 | n12713;
  assign n12715 = pi1097 & ~pi1940;
  assign n12716 = pi2189 & n11794;
  assign n12717 = pi1097 & ~n11794;
  assign n12718 = ~n12716 & ~n12717;
  assign n12719 = pi1940 & ~n12718;
  assign po1148 = n12715 | n12719;
  assign n12721 = pi1098 & ~pi1941;
  assign n12722 = pi2194 & n11770;
  assign n12723 = pi1098 & ~n11770;
  assign n12724 = ~n12722 & ~n12723;
  assign n12725 = pi1941 & ~n12724;
  assign po1149 = n12721 | n12725;
  assign n12727 = pi1099 & ~pi1937;
  assign n12728 = pi2172 & n11829;
  assign n12729 = pi1099 & ~n11829;
  assign n12730 = ~n12728 & ~n12729;
  assign n12731 = pi1937 & ~n12730;
  assign po1150 = n12727 | n12731;
  assign n12733 = pi1100 & ~pi1941;
  assign n12734 = pi2182 & n11770;
  assign n12735 = pi1100 & ~n11770;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = pi1941 & ~n12736;
  assign po1151 = n12733 | n12737;
  assign n12739 = pi1101 & ~pi1940;
  assign n12740 = pi1101 & ~n12065;
  assign n12741 = pi2193 & n12065;
  assign n12742 = ~n12740 & ~n12741;
  assign n12743 = pi1940 & ~n12742;
  assign po1152 = n12739 | n12743;
  assign n12745 = pi1102 & ~pi1940;
  assign n12746 = pi1102 & ~n12065;
  assign n12747 = pi2186 & n12065;
  assign n12748 = ~n12746 & ~n12747;
  assign n12749 = pi1940 & ~n12748;
  assign po1153 = n12745 | n12749;
  assign n12751 = pi1103 & ~pi1941;
  assign n12752 = pi2176 & n11770;
  assign n12753 = pi1103 & ~n11770;
  assign n12754 = ~n12752 & ~n12753;
  assign n12755 = pi1941 & ~n12754;
  assign po1154 = n12751 | n12755;
  assign n12757 = pi1104 & ~pi1941;
  assign n12758 = pi2190 & n11770;
  assign n12759 = pi1104 & ~n11770;
  assign n12760 = ~n12758 & ~n12759;
  assign n12761 = pi1941 & ~n12760;
  assign po1155 = n12757 | n12761;
  assign n12763 = pi1105 & ~pi1940;
  assign n12764 = pi2190 & n11853;
  assign n12765 = pi1105 & ~n11853;
  assign n12766 = ~n12764 & ~n12765;
  assign n12767 = pi1940 & ~n12766;
  assign po1156 = n12763 | n12767;
  assign n12769 = pi1106 & ~pi1940;
  assign n12770 = pi2166 & n11853;
  assign n12771 = pi1106 & ~n11853;
  assign n12772 = ~n12770 & ~n12771;
  assign n12773 = pi1940 & ~n12772;
  assign po1157 = n12769 | n12773;
  assign n12775 = pi1107 & ~pi1940;
  assign n12776 = pi2183 & n11794;
  assign n12777 = pi1107 & ~n11794;
  assign n12778 = ~n12776 & ~n12777;
  assign n12779 = pi1940 & ~n12778;
  assign po1158 = n12775 | n12779;
  assign n12781 = pi1108 & ~pi1941;
  assign n12782 = pi2189 & n11770;
  assign n12783 = pi1108 & ~n11770;
  assign n12784 = ~n12782 & ~n12783;
  assign n12785 = pi1941 & ~n12784;
  assign po1159 = n12781 | n12785;
  assign n12787 = pi1109 & ~pi1937;
  assign n12788 = pi2194 & n11828;
  assign n12789 = pi1109 & ~n11828;
  assign n12790 = ~n12788 & ~n12789;
  assign n12791 = pi1937 & ~n12790;
  assign po1160 = n12787 | n12791;
  assign n12793 = pi1110 & ~pi1941;
  assign n12794 = pi2178 & n11770;
  assign n12795 = pi1110 & ~n11770;
  assign n12796 = ~n12794 & ~n12795;
  assign n12797 = pi1941 & ~n12796;
  assign po1161 = n12793 | n12797;
  assign n12799 = pi1111 & ~pi1941;
  assign n12800 = pi2183 & n11770;
  assign n12801 = pi1111 & ~n11770;
  assign n12802 = ~n12800 & ~n12801;
  assign n12803 = pi1941 & ~n12802;
  assign po1162 = n12799 | n12803;
  assign n12805 = pi1112 & ~pi1940;
  assign n12806 = pi2194 & n11853;
  assign n12807 = pi1112 & ~n11853;
  assign n12808 = ~n12806 & ~n12807;
  assign n12809 = pi1940 & ~n12808;
  assign po1163 = n12805 | n12809;
  assign n12811 = pi1113 & ~pi1940;
  assign n12812 = pi2175 & n11853;
  assign n12813 = pi1113 & ~n11853;
  assign n12814 = ~n12812 & ~n12813;
  assign n12815 = pi1940 & ~n12814;
  assign po1164 = n12811 | n12815;
  assign n12817 = pi1114 & ~pi1937;
  assign n12818 = pi2191 & n11828;
  assign n12819 = pi1114 & ~n11828;
  assign n12820 = ~n12818 & ~n12819;
  assign n12821 = pi1937 & ~n12820;
  assign po1165 = n12817 | n12821;
  assign n12823 = pi1115 & ~pi1940;
  assign n12824 = pi2187 & n11853;
  assign n12825 = pi1115 & ~n11853;
  assign n12826 = ~n12824 & ~n12825;
  assign n12827 = pi1940 & ~n12826;
  assign po1166 = n12823 | n12827;
  assign n12829 = pi1116 & ~pi1940;
  assign n12830 = pi2189 & n11853;
  assign n12831 = pi1116 & ~n11853;
  assign n12832 = ~n12830 & ~n12831;
  assign n12833 = pi1940 & ~n12832;
  assign po1167 = n12829 | n12833;
  assign n12835 = pi1117 & ~pi1936;
  assign n12836 = pi1117 & ~n12004;
  assign n12837 = pi2177 & n12004;
  assign n12838 = ~n12836 & ~n12837;
  assign n12839 = pi1936 & ~n12838;
  assign po1168 = n12835 | n12839;
  assign n12841 = pi1118 & ~pi1936;
  assign n12842 = pi1118 & ~n12004;
  assign n12843 = pi2184 & n12004;
  assign n12844 = ~n12842 & ~n12843;
  assign n12845 = pi1936 & ~n12844;
  assign po1169 = n12841 | n12845;
  assign n12847 = pi1119 & ~pi1940;
  assign n12848 = pi2197 & n11853;
  assign n12849 = pi1119 & ~n11853;
  assign n12850 = ~n12848 & ~n12849;
  assign n12851 = pi1940 & ~n12850;
  assign po1170 = n12847 | n12851;
  assign n12853 = pi1120 & ~pi1940;
  assign n12854 = pi2183 & n11853;
  assign n12855 = pi1120 & ~n11853;
  assign n12856 = ~n12854 & ~n12855;
  assign n12857 = pi1940 & ~n12856;
  assign po1171 = n12853 | n12857;
  assign n12859 = pi1121 & ~pi1941;
  assign n12860 = pi2184 & n11821;
  assign n12861 = pi1121 & ~n11821;
  assign n12862 = ~n12860 & ~n12861;
  assign n12863 = pi1941 & ~n12862;
  assign po1172 = n12859 | n12863;
  assign n12865 = pi1122 & ~pi1936;
  assign n12866 = pi1122 & ~n12004;
  assign n12867 = pi2182 & n12004;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = pi1936 & ~n12868;
  assign po1173 = n12865 | n12869;
  assign n12871 = pi1123 & ~pi1940;
  assign n12872 = pi2166 & n11852;
  assign n12873 = pi1123 & ~n11852;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = pi1940 & ~n12874;
  assign po1174 = n12871 | n12875;
  assign n12877 = pi1124 & ~pi1936;
  assign n12878 = pi2195 & n11751;
  assign n12879 = pi1124 & ~n11751;
  assign n12880 = ~n12878 & ~n12879;
  assign n12881 = pi1936 & ~n12880;
  assign po1175 = n12877 | n12881;
  assign n12883 = ~pi1125 & ~po1956;
  assign n12884 = pi2194 & po1956;
  assign po1176 = n12883 | n12884;
  assign n12886 = ~pi1126 & ~po1956;
  assign n12887 = pi2192 & po1956;
  assign po1177 = n12886 | n12887;
  assign n12889 = pi1127 & ~pi1940;
  assign n12890 = pi2194 & n11852;
  assign n12891 = pi1127 & ~n11852;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = pi1940 & ~n12892;
  assign po1178 = n12889 | n12893;
  assign n12895 = pi1128 & ~n12387;
  assign n12896 = pi2176 & n12387;
  assign po1179 = n12895 | n12896;
  assign n12898 = ~pi1129 & ~po1956;
  assign n12899 = pi2197 & po1956;
  assign po1180 = n12898 | n12899;
  assign n12901 = pi2191 & n12295;
  assign n12902 = pi1130 & ~n12295;
  assign po1181 = n12901 | n12902;
  assign n12904 = pi2167 & n12295;
  assign n12905 = pi1131 & ~n12295;
  assign po1182 = n12904 | n12905;
  assign n12907 = n11518 & n12247;
  assign n12908 = pi1132 & ~n12907;
  assign n12909 = pi2166 & n12907;
  assign po1183 = n12908 | n12909;
  assign n12911 = pi1133 & ~n12907;
  assign n12912 = pi2176 & n12907;
  assign po1184 = n12911 | n12912;
  assign n12914 = pi1134 & ~n12387;
  assign n12915 = pi2172 & n12387;
  assign po1185 = n12914 | n12915;
  assign n12917 = pi1135 & ~pi1940;
  assign n12918 = pi2175 & n11852;
  assign n12919 = pi1135 & ~n11852;
  assign n12920 = ~n12918 & ~n12919;
  assign n12921 = pi1940 & ~n12920;
  assign po1186 = n12917 | n12921;
  assign n12923 = pi1136 & ~pi1936;
  assign n12924 = pi1136 & ~n12004;
  assign n12925 = pi2171 & n12004;
  assign n12926 = ~n12924 & ~n12925;
  assign n12927 = pi1936 & ~n12926;
  assign po1187 = n12923 | n12927;
  assign n12929 = pi1137 & ~n12387;
  assign n12930 = pi2178 & n12387;
  assign po1188 = n12929 | n12930;
  assign n12932 = pi1138 & ~n12387;
  assign n12933 = pi2179 & n12387;
  assign po1189 = n12932 | n12933;
  assign n12935 = pi1139 & ~po1956;
  assign n12936 = pi2196 & po1956;
  assign po1190 = n12935 | n12936;
  assign n12938 = pi1140 & ~po1956;
  assign n12939 = pi2193 & po1956;
  assign po1191 = n12938 | n12939;
  assign n12941 = pi1141 & ~po1956;
  assign n12942 = pi2179 & po1956;
  assign po1192 = n12941 | n12942;
  assign n12944 = pi1142 & ~po1956;
  assign n12945 = pi2185 & po1956;
  assign po1193 = n12944 | n12945;
  assign n12947 = pi1143 & ~po1956;
  assign n12948 = pi2187 & po1956;
  assign po1194 = n12947 | n12948;
  assign n12950 = pi1144 & ~po1956;
  assign n12951 = pi2173 & po1956;
  assign po1195 = n12950 | n12951;
  assign n12953 = pi1145 & ~n12387;
  assign n12954 = pi2186 & n12387;
  assign po1196 = n12953 | n12954;
  assign n12956 = pi1146 & ~n12387;
  assign n12957 = pi2183 & n12387;
  assign po1197 = n12956 | n12957;
  assign n12959 = pi1147 & ~n12387;
  assign n12960 = pi2168 & n12387;
  assign po1198 = n12959 | n12960;
  assign n12962 = pi1148 & ~n12387;
  assign n12963 = pi2174 & n12387;
  assign po1199 = n12962 | n12963;
  assign n12965 = pi1149 & ~n12387;
  assign n12966 = pi2197 & n12387;
  assign po1200 = n12965 | n12966;
  assign n12968 = pi1150 & ~n12387;
  assign n12969 = pi2196 & n12387;
  assign po1201 = n12968 | n12969;
  assign n12971 = pi1151 & ~n12387;
  assign n12972 = pi2193 & n12387;
  assign po1202 = n12971 | n12972;
  assign n12974 = pi1152 & ~n12387;
  assign n12975 = pi2189 & n12387;
  assign po1203 = n12974 | n12975;
  assign n12977 = pi1153 & ~n12387;
  assign n12978 = pi2198 & n12387;
  assign po1204 = n12977 | n12978;
  assign n12980 = pi1154 & ~n12387;
  assign n12981 = pi2185 & n12387;
  assign po1205 = n12980 | n12981;
  assign n12983 = pi1155 & ~n12387;
  assign n12984 = pi2187 & n12387;
  assign po1206 = n12983 | n12984;
  assign n12986 = pi1156 & ~n12387;
  assign n12987 = pi2171 & n12387;
  assign po1207 = n12986 | n12987;
  assign n12989 = pi1157 & ~n12387;
  assign n12990 = pi2191 & n12387;
  assign po1208 = n12989 | n12990;
  assign n12992 = pi1158 & ~n12387;
  assign n12993 = pi2194 & n12387;
  assign po1209 = n12992 | n12993;
  assign n12995 = pi1159 & ~n12387;
  assign n12996 = pi2167 & n12387;
  assign po1210 = n12995 | n12996;
  assign n12998 = pi1160 & ~n12387;
  assign n12999 = pi2188 & n12387;
  assign po1211 = n12998 | n12999;
  assign n13001 = pi1161 & ~n12387;
  assign n13002 = pi2184 & n12387;
  assign po1212 = n13001 | n13002;
  assign n13004 = pi1162 & ~n12387;
  assign n13005 = pi2166 & n12387;
  assign po1213 = n13004 | n13005;
  assign n13007 = pi1163 & ~n12387;
  assign n13008 = pi2192 & n12387;
  assign po1214 = n13007 | n13008;
  assign n13010 = pi2186 & n12295;
  assign n13011 = pi1164 & ~n12295;
  assign po1215 = n13010 | n13011;
  assign n13013 = pi2183 & n12295;
  assign n13014 = pi1165 & ~n12295;
  assign po1216 = n13013 | n13014;
  assign n13016 = pi2168 & n12295;
  assign n13017 = pi1166 & ~n12295;
  assign po1217 = n13016 | n13017;
  assign n13019 = pi2174 & n12295;
  assign n13020 = pi1167 & ~n12295;
  assign po1218 = n13019 | n13020;
  assign n13022 = pi2197 & n12295;
  assign n13023 = pi1168 & ~n12295;
  assign po1219 = n13022 | n13023;
  assign n13025 = pi2196 & n12295;
  assign n13026 = pi1169 & ~n12295;
  assign po1220 = n13025 | n13026;
  assign n13028 = pi2193 & n12295;
  assign n13029 = pi1170 & ~n12295;
  assign po1221 = n13028 | n13029;
  assign n13031 = pi2189 & n12295;
  assign n13032 = pi1171 & ~n12295;
  assign po1222 = n13031 | n13032;
  assign n13034 = pi2198 & n12295;
  assign n13035 = pi1172 & ~n12295;
  assign po1223 = n13034 | n13035;
  assign n13037 = pi2185 & n12295;
  assign n13038 = pi1173 & ~n12295;
  assign po1224 = n13037 | n13038;
  assign n13040 = pi2187 & n12295;
  assign n13041 = pi1174 & ~n12295;
  assign po1225 = n13040 | n13041;
  assign n13043 = pi2171 & n12295;
  assign n13044 = pi1175 & ~n12295;
  assign po1226 = n13043 | n13044;
  assign n13046 = pi2169 & n12295;
  assign n13047 = pi1176 & ~n12295;
  assign po1227 = n13046 | n13047;
  assign n13049 = pi2190 & n12295;
  assign n13050 = pi1177 & ~n12295;
  assign po1228 = n13049 | n13050;
  assign n13052 = pi2181 & n12295;
  assign n13053 = pi1178 & ~n12295;
  assign po1229 = n13052 | n13053;
  assign n13055 = pi2182 & n12295;
  assign n13056 = pi1179 & ~n12295;
  assign po1230 = n13055 | n13056;
  assign n13058 = pi2175 & n12295;
  assign n13059 = pi1180 & ~n12295;
  assign po1231 = n13058 | n13059;
  assign n13061 = pi2177 & n12295;
  assign n13062 = pi1181 & ~n12295;
  assign po1232 = n13061 | n13062;
  assign n13064 = pi2173 & n12295;
  assign n13065 = pi1182 & ~n12295;
  assign po1233 = n13064 | n13065;
  assign n13067 = pi2194 & n12295;
  assign n13068 = pi1183 & ~n12295;
  assign po1234 = n13067 | n13068;
  assign n13070 = pi2188 & n12295;
  assign n13071 = pi1184 & ~n12295;
  assign po1235 = n13070 | n13071;
  assign n13073 = pi2184 & n12295;
  assign n13074 = pi1185 & ~n12295;
  assign po1236 = n13073 | n13074;
  assign n13076 = pi2166 & n12295;
  assign n13077 = pi1186 & ~n12295;
  assign po1237 = n13076 | n13077;
  assign n13079 = pi2192 & n12295;
  assign n13080 = pi1187 & ~n12295;
  assign po1238 = n13079 | n13080;
  assign n13082 = pi1188 & ~n12907;
  assign n13083 = pi2186 & n12907;
  assign po1239 = n13082 | n13083;
  assign n13085 = pi1189 & ~n12907;
  assign n13086 = pi2183 & n12907;
  assign po1240 = n13085 | n13086;
  assign n13088 = pi1190 & ~n12907;
  assign n13089 = pi2172 & n12907;
  assign po1241 = n13088 | n13089;
  assign n13091 = pi1191 & ~n12907;
  assign n13092 = pi2168 & n12907;
  assign po1242 = n13091 | n13092;
  assign n13094 = pi1192 & ~n12907;
  assign n13095 = pi2174 & n12907;
  assign po1243 = n13094 | n13095;
  assign n13097 = pi1193 & ~n12907;
  assign n13098 = pi2197 & n12907;
  assign po1244 = n13097 | n13098;
  assign n13100 = pi1194 & ~n12907;
  assign n13101 = pi2196 & n12907;
  assign po1245 = n13100 | n13101;
  assign n13103 = pi1195 & ~n12907;
  assign n13104 = pi2193 & n12907;
  assign po1246 = n13103 | n13104;
  assign n13106 = pi1196 & ~n12907;
  assign n13107 = pi2189 & n12907;
  assign po1247 = n13106 | n13107;
  assign n13109 = pi1197 & ~n12907;
  assign n13110 = pi2179 & n12907;
  assign po1248 = n13109 | n13110;
  assign n13112 = pi1198 & ~n12907;
  assign n13113 = pi2198 & n12907;
  assign po1249 = n13112 | n13113;
  assign n13115 = pi1199 & ~n12907;
  assign n13116 = pi2185 & n12907;
  assign po1250 = n13115 | n13116;
  assign n13118 = pi1200 & ~n12907;
  assign n13119 = pi2187 & n12907;
  assign po1251 = n13118 | n13119;
  assign n13121 = pi1201 & ~n12907;
  assign n13122 = pi2171 & n12907;
  assign po1252 = n13121 | n13122;
  assign n13124 = pi1202 & ~n12907;
  assign n13125 = pi2169 & n12907;
  assign po1253 = n13124 | n13125;
  assign n13127 = pi1203 & ~n12907;
  assign n13128 = pi2190 & n12907;
  assign po1254 = n13127 | n13128;
  assign n13130 = pi1204 & ~n12907;
  assign n13131 = pi2181 & n12907;
  assign po1255 = n13130 | n13131;
  assign n13133 = pi1205 & ~n12907;
  assign n13134 = pi2182 & n12907;
  assign po1256 = n13133 | n13134;
  assign n13136 = pi1206 & ~n12907;
  assign n13137 = pi2191 & n12907;
  assign po1257 = n13136 | n13137;
  assign n13139 = pi1207 & ~n12907;
  assign n13140 = pi2188 & n12907;
  assign po1258 = n13139 | n13140;
  assign n13142 = pi1208 & ~n12907;
  assign n13143 = pi2184 & n12907;
  assign po1259 = n13142 | n13143;
  assign n13145 = pi1209 & ~n12907;
  assign n13146 = pi2192 & n12907;
  assign po1260 = n13145 | n13146;
  assign n13148 = pi1210 & ~n12907;
  assign n13149 = pi2167 & n12907;
  assign po1261 = n13148 | n13149;
  assign n13151 = pi1211 & ~n12907;
  assign n13152 = pi2178 & n12907;
  assign po1262 = n13151 | n13152;
  assign n13154 = ~pi1212 & ~po1956;
  assign n13155 = pi2186 & po1956;
  assign po1263 = n13154 | n13155;
  assign n13157 = ~pi1213 & ~po1956;
  assign n13158 = pi2183 & po1956;
  assign po1264 = n13157 | n13158;
  assign n13160 = ~pi1214 & ~po1956;
  assign n13161 = pi2172 & po1956;
  assign po1265 = n13160 | n13161;
  assign n13163 = ~pi1215 & ~po1956;
  assign n13164 = pi2168 & po1956;
  assign po1266 = n13163 | n13164;
  assign n13166 = ~pi1216 & ~po1956;
  assign n13167 = pi2174 & po1956;
  assign po1267 = n13166 | n13167;
  assign n13169 = ~pi1217 & ~po1956;
  assign n13170 = pi2178 & po1956;
  assign po1268 = n13169 | n13170;
  assign n13172 = ~pi1218 & ~po1956;
  assign n13173 = pi2198 & po1956;
  assign po1269 = n13172 | n13173;
  assign n13175 = ~pi1219 & ~po1956;
  assign n13176 = pi2191 & po1956;
  assign po1270 = n13175 | n13176;
  assign n13178 = ~pi1220 & ~po1956;
  assign n13179 = pi2167 & po1956;
  assign po1271 = n13178 | n13179;
  assign n13181 = ~pi1221 & ~po1956;
  assign n13182 = pi2188 & po1956;
  assign po1272 = n13181 | n13182;
  assign n13184 = ~pi1222 & ~po1956;
  assign n13185 = pi2184 & po1956;
  assign po1273 = n13184 | n13185;
  assign n13187 = ~pi1223 & ~po1956;
  assign n13188 = pi2195 & po1956;
  assign po1274 = n13187 | n13188;
  assign n13190 = pi1224 & ~pi1941;
  assign n13191 = pi2167 & n11821;
  assign n13192 = pi1224 & ~n11821;
  assign n13193 = ~n13191 & ~n13192;
  assign n13194 = pi1941 & ~n13193;
  assign po1275 = n13190 | n13194;
  assign n13196 = pi1225 & ~pi1937;
  assign n13197 = pi2182 & n11828;
  assign n13198 = pi1225 & ~n11828;
  assign n13199 = ~n13197 & ~n13198;
  assign n13200 = pi1937 & ~n13199;
  assign po1276 = n13196 | n13200;
  assign n13202 = pi1226 & ~pi1941;
  assign n13203 = pi2188 & n11821;
  assign n13204 = pi1226 & ~n11821;
  assign n13205 = ~n13203 & ~n13204;
  assign n13206 = pi1941 & ~n13205;
  assign po1277 = n13202 | n13206;
  assign n13208 = pi1227 & ~pi1937;
  assign n13209 = pi2175 & n11828;
  assign n13210 = pi1227 & ~n11828;
  assign n13211 = ~n13209 & ~n13210;
  assign n13212 = pi1937 & ~n13211;
  assign po1278 = n13208 | n13212;
  assign n13214 = pi1228 & ~pi1941;
  assign n13215 = pi2166 & n11821;
  assign n13216 = pi1228 & ~n11821;
  assign n13217 = ~n13215 & ~n13216;
  assign n13218 = pi1941 & ~n13217;
  assign po1279 = n13214 | n13218;
  assign n13220 = pi1229 & ~pi1941;
  assign n13221 = pi2195 & n11821;
  assign n13222 = pi1229 & ~n11821;
  assign n13223 = ~n13221 & ~n13222;
  assign n13224 = pi1941 & ~n13223;
  assign po1280 = n13220 | n13224;
  assign n13226 = pi1230 & ~pi1941;
  assign n13227 = pi2192 & n11821;
  assign n13228 = pi1230 & ~n11821;
  assign n13229 = ~n13227 & ~n13228;
  assign n13230 = pi1941 & ~n13229;
  assign po1281 = n13226 | n13230;
  assign n13232 = pi1231 & ~pi1941;
  assign n13233 = pi2186 & n11770;
  assign n13234 = pi1231 & ~n11770;
  assign n13235 = ~n13233 & ~n13234;
  assign n13236 = pi1941 & ~n13235;
  assign po1282 = n13232 | n13236;
  assign n13238 = pi1232 & ~pi1937;
  assign n13239 = pi2177 & n11828;
  assign n13240 = pi1232 & ~n11828;
  assign n13241 = ~n13239 & ~n13240;
  assign n13242 = pi1937 & ~n13241;
  assign po1283 = n13238 | n13242;
  assign n13244 = pi1233 & ~pi1941;
  assign n13245 = pi2172 & n11770;
  assign n13246 = pi1233 & ~n11770;
  assign n13247 = ~n13245 & ~n13246;
  assign n13248 = pi1941 & ~n13247;
  assign po1284 = n13244 | n13248;
  assign n13250 = pi1234 & ~pi1937;
  assign n13251 = pi2173 & n11828;
  assign n13252 = pi1234 & ~n11828;
  assign n13253 = ~n13251 & ~n13252;
  assign n13254 = pi1937 & ~n13253;
  assign po1285 = n13250 | n13254;
  assign n13256 = pi1235 & ~pi1941;
  assign n13257 = pi2168 & n11770;
  assign n13258 = pi1235 & ~n11770;
  assign n13259 = ~n13257 & ~n13258;
  assign n13260 = pi1941 & ~n13259;
  assign po1286 = n13256 | n13260;
  assign n13262 = pi1236 & ~pi1941;
  assign n13263 = pi2174 & n11770;
  assign n13264 = pi1236 & ~n11770;
  assign n13265 = ~n13263 & ~n13264;
  assign n13266 = pi1941 & ~n13265;
  assign po1287 = n13262 | n13266;
  assign n13268 = pi1237 & ~pi1937;
  assign n13269 = pi2167 & n11828;
  assign n13270 = pi1237 & ~n11828;
  assign n13271 = ~n13269 & ~n13270;
  assign n13272 = pi1937 & ~n13271;
  assign po1288 = n13268 | n13272;
  assign n13274 = pi1238 & ~pi1941;
  assign n13275 = pi2197 & n11770;
  assign n13276 = pi1238 & ~n11770;
  assign n13277 = ~n13275 & ~n13276;
  assign n13278 = pi1941 & ~n13277;
  assign po1289 = n13274 | n13278;
  assign n13280 = pi1239 & ~pi1941;
  assign n13281 = pi2196 & n11770;
  assign n13282 = pi1239 & ~n11770;
  assign n13283 = ~n13281 & ~n13282;
  assign n13284 = pi1941 & ~n13283;
  assign po1290 = n13280 | n13284;
  assign n13286 = pi1240 & ~pi1941;
  assign n13287 = pi2193 & n11770;
  assign n13288 = pi1240 & ~n11770;
  assign n13289 = ~n13287 & ~n13288;
  assign n13290 = pi1941 & ~n13289;
  assign po1291 = n13286 | n13290;
  assign n13292 = pi1241 & ~pi1937;
  assign n13293 = pi2188 & n11828;
  assign n13294 = pi1241 & ~n11828;
  assign n13295 = ~n13293 & ~n13294;
  assign n13296 = pi1937 & ~n13295;
  assign po1292 = n13292 | n13296;
  assign n13298 = pi1242 & ~pi1941;
  assign n13299 = pi2179 & n11770;
  assign n13300 = pi1242 & ~n11770;
  assign n13301 = ~n13299 & ~n13300;
  assign n13302 = pi1941 & ~n13301;
  assign po1293 = n13298 | n13302;
  assign n13304 = pi1243 & ~pi1937;
  assign n13305 = pi2184 & n11828;
  assign n13306 = pi1243 & ~n11828;
  assign n13307 = ~n13305 & ~n13306;
  assign n13308 = pi1937 & ~n13307;
  assign po1294 = n13304 | n13308;
  assign n13310 = pi1244 & ~pi1941;
  assign n13311 = pi2198 & n11770;
  assign n13312 = pi1244 & ~n11770;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = pi1941 & ~n13313;
  assign po1295 = n13310 | n13314;
  assign n13316 = pi1245 & ~pi1937;
  assign n13317 = pi2166 & n11828;
  assign n13318 = pi1245 & ~n11828;
  assign n13319 = ~n13317 & ~n13318;
  assign n13320 = pi1937 & ~n13319;
  assign po1296 = n13316 | n13320;
  assign n13322 = pi1246 & ~pi1941;
  assign n13323 = pi2185 & n11770;
  assign n13324 = pi1246 & ~n11770;
  assign n13325 = ~n13323 & ~n13324;
  assign n13326 = pi1941 & ~n13325;
  assign po1297 = n13322 | n13326;
  assign n13328 = pi1247 & ~pi1941;
  assign n13329 = pi2187 & n11770;
  assign n13330 = pi1247 & ~n11770;
  assign n13331 = ~n13329 & ~n13330;
  assign n13332 = pi1941 & ~n13331;
  assign po1298 = n13328 | n13332;
  assign n13334 = pi1248 & ~pi1937;
  assign n13335 = pi2195 & n11828;
  assign n13336 = pi1248 & ~n11828;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = pi1937 & ~n13337;
  assign po1299 = n13334 | n13338;
  assign n13340 = pi1249 & ~pi1941;
  assign n13341 = pi2171 & n11770;
  assign n13342 = pi1249 & ~n11770;
  assign n13343 = ~n13341 & ~n13342;
  assign n13344 = pi1941 & ~n13343;
  assign po1300 = n13340 | n13344;
  assign n13346 = pi1250 & ~pi1941;
  assign n13347 = pi2169 & n11770;
  assign n13348 = pi1250 & ~n11770;
  assign n13349 = ~n13347 & ~n13348;
  assign n13350 = pi1941 & ~n13349;
  assign po1301 = n13346 | n13350;
  assign n13352 = pi1251 & ~pi1937;
  assign n13353 = pi2192 & n11828;
  assign n13354 = pi1251 & ~n11828;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = pi1937 & ~n13355;
  assign po1302 = n13352 | n13356;
  assign n13358 = pi1252 & ~pi1941;
  assign n13359 = pi2170 & n11770;
  assign n13360 = pi1252 & ~n11770;
  assign n13361 = ~n13359 & ~n13360;
  assign n13362 = pi1941 & ~n13361;
  assign po1303 = n13358 | n13362;
  assign n13364 = pi1253 & ~pi1937;
  assign n13365 = pi2186 & n11829;
  assign n13366 = pi1253 & ~n11829;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = pi1937 & ~n13367;
  assign po1304 = n13364 | n13368;
  assign n13370 = pi1254 & ~pi1941;
  assign n13371 = pi2181 & n11770;
  assign n13372 = pi1254 & ~n11770;
  assign n13373 = ~n13371 & ~n13372;
  assign n13374 = pi1941 & ~n13373;
  assign po1305 = n13370 | n13374;
  assign n13376 = pi1255 & ~pi1937;
  assign n13377 = pi2183 & n11829;
  assign n13378 = pi1255 & ~n11829;
  assign n13379 = ~n13377 & ~n13378;
  assign n13380 = pi1937 & ~n13379;
  assign po1306 = n13376 | n13380;
  assign n13382 = pi1256 & ~pi1941;
  assign n13383 = pi2175 & n11770;
  assign n13384 = pi1256 & ~n11770;
  assign n13385 = ~n13383 & ~n13384;
  assign n13386 = pi1941 & ~n13385;
  assign po1307 = n13382 | n13386;
  assign n13388 = pi1257 & ~pi1941;
  assign n13389 = pi2191 & n11770;
  assign n13390 = pi1257 & ~n11770;
  assign n13391 = ~n13389 & ~n13390;
  assign n13392 = pi1941 & ~n13391;
  assign po1308 = n13388 | n13392;
  assign n13394 = pi1258 & ~pi1941;
  assign n13395 = pi2177 & n11770;
  assign n13396 = pi1258 & ~n11770;
  assign n13397 = ~n13395 & ~n13396;
  assign n13398 = pi1941 & ~n13397;
  assign po1309 = n13394 | n13398;
  assign n13400 = pi1259 & ~pi1941;
  assign n13401 = pi2173 & n11770;
  assign n13402 = pi1259 & ~n11770;
  assign n13403 = ~n13401 & ~n13402;
  assign n13404 = pi1941 & ~n13403;
  assign po1310 = n13400 | n13404;
  assign n13406 = pi1260 & ~pi1937;
  assign n13407 = pi2168 & n11829;
  assign n13408 = pi1260 & ~n11829;
  assign n13409 = ~n13407 & ~n13408;
  assign n13410 = pi1937 & ~n13409;
  assign po1311 = n13406 | n13410;
  assign n13412 = pi1261 & ~pi1941;
  assign n13413 = pi2167 & n11770;
  assign n13414 = pi1261 & ~n11770;
  assign n13415 = ~n13413 & ~n13414;
  assign n13416 = pi1941 & ~n13415;
  assign po1312 = n13412 | n13416;
  assign n13418 = pi1262 & ~pi1937;
  assign n13419 = pi2174 & n11829;
  assign n13420 = pi1262 & ~n11829;
  assign n13421 = ~n13419 & ~n13420;
  assign n13422 = pi1937 & ~n13421;
  assign po1313 = n13418 | n13422;
  assign n13424 = pi1263 & ~pi1941;
  assign n13425 = pi2188 & n11770;
  assign n13426 = pi1263 & ~n11770;
  assign n13427 = ~n13425 & ~n13426;
  assign n13428 = pi1941 & ~n13427;
  assign po1314 = n13424 | n13428;
  assign n13430 = pi1264 & ~pi1937;
  assign n13431 = pi2197 & n11829;
  assign n13432 = pi1264 & ~n11829;
  assign n13433 = ~n13431 & ~n13432;
  assign n13434 = pi1937 & ~n13433;
  assign po1315 = n13430 | n13434;
  assign n13436 = pi1265 & ~pi1941;
  assign n13437 = pi2166 & n11770;
  assign n13438 = pi1265 & ~n11770;
  assign n13439 = ~n13437 & ~n13438;
  assign n13440 = pi1941 & ~n13439;
  assign po1316 = n13436 | n13440;
  assign n13442 = pi1266 & ~pi1937;
  assign n13443 = pi2178 & n11829;
  assign n13444 = pi1266 & ~n11829;
  assign n13445 = ~n13443 & ~n13444;
  assign n13446 = pi1937 & ~n13445;
  assign po1317 = n13442 | n13446;
  assign n13448 = pi1267 & ~pi1941;
  assign n13449 = pi2192 & n11770;
  assign n13450 = pi1267 & ~n11770;
  assign n13451 = ~n13449 & ~n13450;
  assign n13452 = pi1941 & ~n13451;
  assign po1318 = n13448 | n13452;
  assign n13454 = pi1268 & ~pi1937;
  assign n13455 = pi2196 & n11829;
  assign n13456 = pi1268 & ~n11829;
  assign n13457 = ~n13455 & ~n13456;
  assign n13458 = pi1937 & ~n13457;
  assign po1319 = n13454 | n13458;
  assign n13460 = pi1269 & ~pi1937;
  assign n13461 = pi2193 & n11829;
  assign n13462 = pi1269 & ~n11829;
  assign n13463 = ~n13461 & ~n13462;
  assign n13464 = pi1937 & ~n13463;
  assign po1320 = n13460 | n13464;
  assign n13466 = pi1270 & ~pi1937;
  assign n13467 = pi2179 & n11829;
  assign n13468 = pi1270 & ~n11829;
  assign n13469 = ~n13467 & ~n13468;
  assign n13470 = pi1937 & ~n13469;
  assign po1321 = n13466 | n13470;
  assign n13472 = pi1271 & ~pi1937;
  assign n13473 = pi2198 & n11829;
  assign n13474 = pi1271 & ~n11829;
  assign n13475 = ~n13473 & ~n13474;
  assign n13476 = pi1937 & ~n13475;
  assign po1322 = n13472 | n13476;
  assign n13478 = pi1272 & ~pi1937;
  assign n13479 = pi2187 & n11829;
  assign n13480 = pi1272 & ~n11829;
  assign n13481 = ~n13479 & ~n13480;
  assign n13482 = pi1937 & ~n13481;
  assign po1323 = n13478 | n13482;
  assign n13484 = pi1273 & ~pi1937;
  assign n13485 = pi2171 & n11829;
  assign n13486 = pi1273 & ~n11829;
  assign n13487 = ~n13485 & ~n13486;
  assign n13488 = pi1937 & ~n13487;
  assign po1324 = n13484 | n13488;
  assign n13490 = pi1274 & ~pi1937;
  assign n13491 = pi2169 & n11829;
  assign n13492 = pi1274 & ~n11829;
  assign n13493 = ~n13491 & ~n13492;
  assign n13494 = pi1937 & ~n13493;
  assign po1325 = n13490 | n13494;
  assign n13496 = pi1275 & ~pi1937;
  assign n13497 = pi2190 & n11829;
  assign n13498 = pi1275 & ~n11829;
  assign n13499 = ~n13497 & ~n13498;
  assign n13500 = pi1937 & ~n13499;
  assign po1326 = n13496 | n13500;
  assign n13502 = pi1276 & ~pi1937;
  assign n13503 = pi2181 & n11829;
  assign n13504 = pi1276 & ~n11829;
  assign n13505 = ~n13503 & ~n13504;
  assign n13506 = pi1937 & ~n13505;
  assign po1327 = n13502 | n13506;
  assign n13508 = pi1277 & ~pi1937;
  assign n13509 = pi2182 & n11829;
  assign n13510 = pi1277 & ~n11829;
  assign n13511 = ~n13509 & ~n13510;
  assign n13512 = pi1937 & ~n13511;
  assign po1328 = n13508 | n13512;
  assign n13514 = pi1278 & ~pi1937;
  assign n13515 = pi2175 & n11829;
  assign n13516 = pi1278 & ~n11829;
  assign n13517 = ~n13515 & ~n13516;
  assign n13518 = pi1937 & ~n13517;
  assign po1329 = n13514 | n13518;
  assign n13520 = pi1279 & ~pi1937;
  assign n13521 = pi2177 & n11829;
  assign n13522 = pi1279 & ~n11829;
  assign n13523 = ~n13521 & ~n13522;
  assign n13524 = pi1937 & ~n13523;
  assign po1330 = n13520 | n13524;
  assign n13526 = pi1280 & ~pi1937;
  assign n13527 = pi2173 & n11829;
  assign n13528 = pi1280 & ~n11829;
  assign n13529 = ~n13527 & ~n13528;
  assign n13530 = pi1937 & ~n13529;
  assign po1331 = n13526 | n13530;
  assign n13532 = pi1281 & ~pi1937;
  assign n13533 = pi2194 & n11829;
  assign n13534 = pi1281 & ~n11829;
  assign n13535 = ~n13533 & ~n13534;
  assign n13536 = pi1937 & ~n13535;
  assign po1332 = n13532 | n13536;
  assign n13538 = pi1282 & ~pi1937;
  assign n13539 = pi2167 & n11829;
  assign n13540 = pi1282 & ~n11829;
  assign n13541 = ~n13539 & ~n13540;
  assign n13542 = pi1937 & ~n13541;
  assign po1333 = n13538 | n13542;
  assign n13544 = pi1283 & ~pi1937;
  assign n13545 = pi2188 & n11829;
  assign n13546 = pi1283 & ~n11829;
  assign n13547 = ~n13545 & ~n13546;
  assign n13548 = pi1937 & ~n13547;
  assign po1334 = n13544 | n13548;
  assign n13550 = pi1284 & ~pi1937;
  assign n13551 = pi2184 & n11829;
  assign n13552 = pi1284 & ~n11829;
  assign n13553 = ~n13551 & ~n13552;
  assign n13554 = pi1937 & ~n13553;
  assign po1335 = n13550 | n13554;
  assign n13556 = pi1285 & ~pi1937;
  assign n13557 = pi2166 & n11829;
  assign n13558 = pi1285 & ~n11829;
  assign n13559 = ~n13557 & ~n13558;
  assign n13560 = pi1937 & ~n13559;
  assign po1336 = n13556 | n13560;
  assign n13562 = pi1286 & ~pi1937;
  assign n13563 = pi2192 & n11829;
  assign n13564 = pi1286 & ~n11829;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = pi1937 & ~n13565;
  assign po1337 = n13562 | n13566;
  assign n13568 = pi1287 & ~pi1937;
  assign n13569 = pi2186 & n11778;
  assign n13570 = pi1287 & ~n11778;
  assign n13571 = ~n13569 & ~n13570;
  assign n13572 = pi1937 & ~n13571;
  assign po1338 = n13568 | n13572;
  assign n13574 = pi1288 & ~pi1937;
  assign n13575 = pi2183 & n11778;
  assign n13576 = pi1288 & ~n11778;
  assign n13577 = ~n13575 & ~n13576;
  assign n13578 = pi1937 & ~n13577;
  assign po1339 = n13574 | n13578;
  assign n13580 = pi1289 & ~pi1937;
  assign n13581 = pi2168 & n11778;
  assign n13582 = pi1289 & ~n11778;
  assign n13583 = ~n13581 & ~n13582;
  assign n13584 = pi1937 & ~n13583;
  assign po1340 = n13580 | n13584;
  assign n13586 = pi1290 & ~pi1937;
  assign n13587 = pi2174 & n11778;
  assign n13588 = pi1290 & ~n11778;
  assign n13589 = ~n13587 & ~n13588;
  assign n13590 = pi1937 & ~n13589;
  assign po1341 = n13586 | n13590;
  assign n13592 = pi1291 & ~pi1937;
  assign n13593 = pi2197 & n11778;
  assign n13594 = pi1291 & ~n11778;
  assign n13595 = ~n13593 & ~n13594;
  assign n13596 = pi1937 & ~n13595;
  assign po1342 = n13592 | n13596;
  assign n13598 = pi1292 & ~pi1937;
  assign n13599 = pi2196 & n11778;
  assign n13600 = pi1292 & ~n11778;
  assign n13601 = ~n13599 & ~n13600;
  assign n13602 = pi1937 & ~n13601;
  assign po1343 = n13598 | n13602;
  assign n13604 = pi1293 & ~pi1937;
  assign n13605 = pi2193 & n11778;
  assign n13606 = pi1293 & ~n11778;
  assign n13607 = ~n13605 & ~n13606;
  assign n13608 = pi1937 & ~n13607;
  assign po1344 = n13604 | n13608;
  assign n13610 = pi1294 & ~pi1937;
  assign n13611 = pi2189 & n11778;
  assign n13612 = pi1294 & ~n11778;
  assign n13613 = ~n13611 & ~n13612;
  assign n13614 = pi1937 & ~n13613;
  assign po1345 = n13610 | n13614;
  assign n13616 = pi1295 & ~pi1937;
  assign n13617 = pi2198 & n11778;
  assign n13618 = pi1295 & ~n11778;
  assign n13619 = ~n13617 & ~n13618;
  assign n13620 = pi1937 & ~n13619;
  assign po1346 = n13616 | n13620;
  assign n13622 = pi1296 & ~pi1937;
  assign n13623 = pi2185 & n11778;
  assign n13624 = pi1296 & ~n11778;
  assign n13625 = ~n13623 & ~n13624;
  assign n13626 = pi1937 & ~n13625;
  assign po1347 = n13622 | n13626;
  assign n13628 = pi1297 & ~pi1937;
  assign n13629 = pi2187 & n11778;
  assign n13630 = pi1297 & ~n11778;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = pi1937 & ~n13631;
  assign po1348 = n13628 | n13632;
  assign n13634 = pi1298 & ~pi1937;
  assign n13635 = pi2171 & n11778;
  assign n13636 = pi1298 & ~n11778;
  assign n13637 = ~n13635 & ~n13636;
  assign n13638 = pi1937 & ~n13637;
  assign po1349 = n13634 | n13638;
  assign n13640 = pi1299 & ~pi1937;
  assign n13641 = pi2169 & n11778;
  assign n13642 = pi1299 & ~n11778;
  assign n13643 = ~n13641 & ~n13642;
  assign n13644 = pi1937 & ~n13643;
  assign po1350 = n13640 | n13644;
  assign n13646 = pi1300 & ~pi1937;
  assign n13647 = pi2170 & n11778;
  assign n13648 = pi1300 & ~n11778;
  assign n13649 = ~n13647 & ~n13648;
  assign n13650 = pi1937 & ~n13649;
  assign po1351 = n13646 | n13650;
  assign n13652 = pi1301 & ~pi1937;
  assign n13653 = pi2182 & n11778;
  assign n13654 = pi1301 & ~n11778;
  assign n13655 = ~n13653 & ~n13654;
  assign n13656 = pi1937 & ~n13655;
  assign po1352 = n13652 | n13656;
  assign n13658 = pi1302 & ~pi1937;
  assign n13659 = pi2175 & n11778;
  assign n13660 = pi1302 & ~n11778;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = pi1937 & ~n13661;
  assign po1353 = n13658 | n13662;
  assign n13664 = pi1303 & ~pi1937;
  assign n13665 = pi2191 & n11778;
  assign n13666 = pi1303 & ~n11778;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = pi1937 & ~n13667;
  assign po1354 = n13664 | n13668;
  assign n13670 = pi1304 & ~pi1937;
  assign n13671 = pi2173 & n11778;
  assign n13672 = pi1304 & ~n11778;
  assign n13673 = ~n13671 & ~n13672;
  assign n13674 = pi1937 & ~n13673;
  assign po1355 = n13670 | n13674;
  assign n13676 = pi1305 & ~pi1937;
  assign n13677 = pi2167 & n11778;
  assign n13678 = pi1305 & ~n11778;
  assign n13679 = ~n13677 & ~n13678;
  assign n13680 = pi1937 & ~n13679;
  assign po1356 = n13676 | n13680;
  assign n13682 = pi1306 & ~pi1937;
  assign n13683 = pi2188 & n11778;
  assign n13684 = pi1306 & ~n11778;
  assign n13685 = ~n13683 & ~n13684;
  assign n13686 = pi1937 & ~n13685;
  assign po1357 = n13682 | n13686;
  assign n13688 = pi1307 & ~pi1937;
  assign n13689 = pi2166 & n11778;
  assign n13690 = pi1307 & ~n11778;
  assign n13691 = ~n13689 & ~n13690;
  assign n13692 = pi1937 & ~n13691;
  assign po1358 = n13688 | n13692;
  assign n13694 = pi1308 & ~pi1937;
  assign n13695 = pi2192 & n11778;
  assign n13696 = pi1308 & ~n11778;
  assign n13697 = ~n13695 & ~n13696;
  assign n13698 = pi1937 & ~n13697;
  assign po1359 = n13694 | n13698;
  assign n13700 = pi1309 & ~pi1937;
  assign n13701 = pi2190 & n11778;
  assign n13702 = pi1309 & ~n11778;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = pi1937 & ~n13703;
  assign po1360 = n13700 | n13704;
  assign n13706 = pi1310 & ~pi1938;
  assign n13707 = pi2186 & n11836;
  assign n13708 = pi1310 & ~n11836;
  assign n13709 = ~n13707 & ~n13708;
  assign n13710 = pi1938 & ~n13709;
  assign po1361 = n13706 | n13710;
  assign n13712 = pi1311 & ~pi1938;
  assign n13713 = pi2183 & n11836;
  assign n13714 = pi1311 & ~n11836;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = pi1938 & ~n13715;
  assign po1362 = n13712 | n13716;
  assign n13718 = pi1312 & ~pi1938;
  assign n13719 = pi2172 & n11836;
  assign n13720 = pi1312 & ~n11836;
  assign n13721 = ~n13719 & ~n13720;
  assign n13722 = pi1938 & ~n13721;
  assign po1363 = n13718 | n13722;
  assign n13724 = pi1313 & ~pi1938;
  assign n13725 = pi2174 & n11836;
  assign n13726 = pi1313 & ~n11836;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = pi1938 & ~n13727;
  assign po1364 = n13724 | n13728;
  assign n13730 = pi1314 & ~pi1938;
  assign n13731 = pi2197 & n11836;
  assign n13732 = pi1314 & ~n11836;
  assign n13733 = ~n13731 & ~n13732;
  assign n13734 = pi1938 & ~n13733;
  assign po1365 = n13730 | n13734;
  assign n13736 = pi1315 & ~pi1938;
  assign n13737 = pi2178 & n11836;
  assign n13738 = pi1315 & ~n11836;
  assign n13739 = ~n13737 & ~n13738;
  assign n13740 = pi1938 & ~n13739;
  assign po1366 = n13736 | n13740;
  assign n13742 = pi1316 & ~pi1938;
  assign n13743 = pi2193 & n11836;
  assign n13744 = pi1316 & ~n11836;
  assign n13745 = ~n13743 & ~n13744;
  assign n13746 = pi1938 & ~n13745;
  assign po1367 = n13742 | n13746;
  assign n13748 = pi1317 & ~pi1938;
  assign n13749 = pi2189 & n11836;
  assign n13750 = pi1317 & ~n11836;
  assign n13751 = ~n13749 & ~n13750;
  assign n13752 = pi1938 & ~n13751;
  assign po1368 = n13748 | n13752;
  assign n13754 = pi1318 & ~pi1938;
  assign n13755 = pi2179 & n11836;
  assign n13756 = pi1318 & ~n11836;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = pi1938 & ~n13757;
  assign po1369 = n13754 | n13758;
  assign n13760 = pi1319 & ~pi1938;
  assign n13761 = pi2198 & n11836;
  assign n13762 = pi1319 & ~n11836;
  assign n13763 = ~n13761 & ~n13762;
  assign n13764 = pi1938 & ~n13763;
  assign po1370 = n13760 | n13764;
  assign n13766 = pi1320 & ~pi1938;
  assign n13767 = pi2185 & n11836;
  assign n13768 = pi1320 & ~n11836;
  assign n13769 = ~n13767 & ~n13768;
  assign n13770 = pi1938 & ~n13769;
  assign po1371 = n13766 | n13770;
  assign n13772 = pi1321 & ~pi1938;
  assign n13773 = pi2187 & n11836;
  assign n13774 = pi1321 & ~n11836;
  assign n13775 = ~n13773 & ~n13774;
  assign n13776 = pi1938 & ~n13775;
  assign po1372 = n13772 | n13776;
  assign n13778 = pi1322 & ~pi1938;
  assign n13779 = pi2176 & n11836;
  assign n13780 = pi1322 & ~n11836;
  assign n13781 = ~n13779 & ~n13780;
  assign n13782 = pi1938 & ~n13781;
  assign po1373 = n13778 | n13782;
  assign n13784 = pi1323 & ~pi1938;
  assign n13785 = pi2169 & n11836;
  assign n13786 = pi1323 & ~n11836;
  assign n13787 = ~n13785 & ~n13786;
  assign n13788 = pi1938 & ~n13787;
  assign po1374 = n13784 | n13788;
  assign n13790 = pi1324 & ~pi1938;
  assign n13791 = pi2190 & n11836;
  assign n13792 = pi1324 & ~n11836;
  assign n13793 = ~n13791 & ~n13792;
  assign n13794 = pi1938 & ~n13793;
  assign po1375 = n13790 | n13794;
  assign n13796 = pi1325 & ~pi1938;
  assign n13797 = pi2170 & n11836;
  assign n13798 = pi1325 & ~n11836;
  assign n13799 = ~n13797 & ~n13798;
  assign n13800 = pi1938 & ~n13799;
  assign po1376 = n13796 | n13800;
  assign n13802 = pi1326 & ~pi1938;
  assign n13803 = pi2182 & n11836;
  assign n13804 = pi1326 & ~n11836;
  assign n13805 = ~n13803 & ~n13804;
  assign n13806 = pi1938 & ~n13805;
  assign po1377 = n13802 | n13806;
  assign n13808 = pi1327 & ~pi1938;
  assign n13809 = pi2175 & n11836;
  assign n13810 = pi1327 & ~n11836;
  assign n13811 = ~n13809 & ~n13810;
  assign n13812 = pi1938 & ~n13811;
  assign po1378 = n13808 | n13812;
  assign n13814 = pi1328 & ~pi1938;
  assign n13815 = pi2191 & n11836;
  assign n13816 = pi1328 & ~n11836;
  assign n13817 = ~n13815 & ~n13816;
  assign n13818 = pi1938 & ~n13817;
  assign po1379 = n13814 | n13818;
  assign n13820 = pi1329 & ~pi1938;
  assign n13821 = pi2173 & n11836;
  assign n13822 = pi1329 & ~n11836;
  assign n13823 = ~n13821 & ~n13822;
  assign n13824 = pi1938 & ~n13823;
  assign po1380 = n13820 | n13824;
  assign n13826 = pi1330 & ~pi1938;
  assign n13827 = pi2194 & n11836;
  assign n13828 = pi1330 & ~n11836;
  assign n13829 = ~n13827 & ~n13828;
  assign n13830 = pi1938 & ~n13829;
  assign po1381 = n13826 | n13830;
  assign n13832 = pi1331 & ~pi1938;
  assign n13833 = pi2167 & n11836;
  assign n13834 = pi1331 & ~n11836;
  assign n13835 = ~n13833 & ~n13834;
  assign n13836 = pi1938 & ~n13835;
  assign po1382 = n13832 | n13836;
  assign n13838 = pi1332 & ~pi1938;
  assign n13839 = pi2184 & n11836;
  assign n13840 = pi1332 & ~n11836;
  assign n13841 = ~n13839 & ~n13840;
  assign n13842 = pi1938 & ~n13841;
  assign po1383 = n13838 | n13842;
  assign n13844 = pi1333 & ~pi1938;
  assign n13845 = pi2166 & n11836;
  assign n13846 = pi1333 & ~n11836;
  assign n13847 = ~n13845 & ~n13846;
  assign n13848 = pi1938 & ~n13847;
  assign po1384 = n13844 | n13848;
  assign n13850 = pi1334 & ~pi1938;
  assign n13851 = pi2195 & n11836;
  assign n13852 = pi1334 & ~n11836;
  assign n13853 = ~n13851 & ~n13852;
  assign n13854 = pi1938 & ~n13853;
  assign po1385 = n13850 | n13854;
  assign n13856 = pi1335 & ~pi1938;
  assign n13857 = pi2186 & n11837;
  assign n13858 = pi1335 & ~n11837;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = pi1938 & ~n13859;
  assign po1386 = n13856 | n13860;
  assign n13862 = pi1336 & ~pi1938;
  assign n13863 = pi2183 & n11837;
  assign n13864 = pi1336 & ~n11837;
  assign n13865 = ~n13863 & ~n13864;
  assign n13866 = pi1938 & ~n13865;
  assign po1387 = n13862 | n13866;
  assign n13868 = pi1337 & ~pi1938;
  assign n13869 = pi2172 & n11837;
  assign n13870 = pi1337 & ~n11837;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = pi1938 & ~n13871;
  assign po1388 = n13868 | n13872;
  assign n13874 = pi1338 & ~pi1938;
  assign n13875 = pi2174 & n11837;
  assign n13876 = pi1338 & ~n11837;
  assign n13877 = ~n13875 & ~n13876;
  assign n13878 = pi1938 & ~n13877;
  assign po1389 = n13874 | n13878;
  assign n13880 = pi1339 & ~pi1938;
  assign n13881 = pi2197 & n11837;
  assign n13882 = pi1339 & ~n11837;
  assign n13883 = ~n13881 & ~n13882;
  assign n13884 = pi1938 & ~n13883;
  assign po1390 = n13880 | n13884;
  assign n13886 = pi1340 & ~pi1938;
  assign n13887 = pi2178 & n11837;
  assign n13888 = pi1340 & ~n11837;
  assign n13889 = ~n13887 & ~n13888;
  assign n13890 = pi1938 & ~n13889;
  assign po1391 = n13886 | n13890;
  assign n13892 = pi1341 & ~pi1938;
  assign n13893 = pi2193 & n11837;
  assign n13894 = pi1341 & ~n11837;
  assign n13895 = ~n13893 & ~n13894;
  assign n13896 = pi1938 & ~n13895;
  assign po1392 = n13892 | n13896;
  assign n13898 = pi1342 & ~pi1938;
  assign n13899 = pi2189 & n11837;
  assign n13900 = pi1342 & ~n11837;
  assign n13901 = ~n13899 & ~n13900;
  assign n13902 = pi1938 & ~n13901;
  assign po1393 = n13898 | n13902;
  assign n13904 = pi1343 & ~pi1938;
  assign n13905 = pi2179 & n11837;
  assign n13906 = pi1343 & ~n11837;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = pi1938 & ~n13907;
  assign po1394 = n13904 | n13908;
  assign n13910 = pi1344 & ~pi1938;
  assign n13911 = pi2198 & n11837;
  assign n13912 = pi1344 & ~n11837;
  assign n13913 = ~n13911 & ~n13912;
  assign n13914 = pi1938 & ~n13913;
  assign po1395 = n13910 | n13914;
  assign n13916 = pi1345 & ~pi1938;
  assign n13917 = pi2185 & n11837;
  assign n13918 = pi1345 & ~n11837;
  assign n13919 = ~n13917 & ~n13918;
  assign n13920 = pi1938 & ~n13919;
  assign po1396 = n13916 | n13920;
  assign n13922 = pi1346 & ~pi1938;
  assign n13923 = pi2187 & n11837;
  assign n13924 = pi1346 & ~n11837;
  assign n13925 = ~n13923 & ~n13924;
  assign n13926 = pi1938 & ~n13925;
  assign po1397 = n13922 | n13926;
  assign n13928 = pi1347 & ~pi1938;
  assign n13929 = pi2176 & n11837;
  assign n13930 = pi1347 & ~n11837;
  assign n13931 = ~n13929 & ~n13930;
  assign n13932 = pi1938 & ~n13931;
  assign po1398 = n13928 | n13932;
  assign n13934 = pi1348 & ~pi1938;
  assign n13935 = pi2169 & n11837;
  assign n13936 = pi1348 & ~n11837;
  assign n13937 = ~n13935 & ~n13936;
  assign n13938 = pi1938 & ~n13937;
  assign po1399 = n13934 | n13938;
  assign n13940 = pi1349 & ~pi1938;
  assign n13941 = pi2190 & n11837;
  assign n13942 = pi1349 & ~n11837;
  assign n13943 = ~n13941 & ~n13942;
  assign n13944 = pi1938 & ~n13943;
  assign po1400 = n13940 | n13944;
  assign n13946 = pi1350 & ~pi1938;
  assign n13947 = pi2170 & n11837;
  assign n13948 = pi1350 & ~n11837;
  assign n13949 = ~n13947 & ~n13948;
  assign n13950 = pi1938 & ~n13949;
  assign po1401 = n13946 | n13950;
  assign n13952 = pi1351 & ~pi1938;
  assign n13953 = pi2182 & n11837;
  assign n13954 = pi1351 & ~n11837;
  assign n13955 = ~n13953 & ~n13954;
  assign n13956 = pi1938 & ~n13955;
  assign po1402 = n13952 | n13956;
  assign n13958 = pi1352 & ~pi1938;
  assign n13959 = pi2175 & n11837;
  assign n13960 = pi1352 & ~n11837;
  assign n13961 = ~n13959 & ~n13960;
  assign n13962 = pi1938 & ~n13961;
  assign po1403 = n13958 | n13962;
  assign n13964 = pi1353 & ~pi1938;
  assign n13965 = pi2191 & n11837;
  assign n13966 = pi1353 & ~n11837;
  assign n13967 = ~n13965 & ~n13966;
  assign n13968 = pi1938 & ~n13967;
  assign po1404 = n13964 | n13968;
  assign n13970 = pi1354 & ~pi1938;
  assign n13971 = pi2173 & n11837;
  assign n13972 = pi1354 & ~n11837;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = pi1938 & ~n13973;
  assign po1405 = n13970 | n13974;
  assign n13976 = pi1355 & ~pi1938;
  assign n13977 = pi2194 & n11837;
  assign n13978 = pi1355 & ~n11837;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = pi1938 & ~n13979;
  assign po1406 = n13976 | n13980;
  assign n13982 = pi1356 & ~pi1938;
  assign n13983 = pi2167 & n11837;
  assign n13984 = pi1356 & ~n11837;
  assign n13985 = ~n13983 & ~n13984;
  assign n13986 = pi1938 & ~n13985;
  assign po1407 = n13982 | n13986;
  assign n13988 = pi1357 & ~pi1938;
  assign n13989 = pi2184 & n11837;
  assign n13990 = pi1357 & ~n11837;
  assign n13991 = ~n13989 & ~n13990;
  assign n13992 = pi1938 & ~n13991;
  assign po1408 = n13988 | n13992;
  assign n13994 = pi1358 & ~pi1938;
  assign n13995 = pi2166 & n11837;
  assign n13996 = pi1358 & ~n11837;
  assign n13997 = ~n13995 & ~n13996;
  assign n13998 = pi1938 & ~n13997;
  assign po1409 = n13994 | n13998;
  assign n14000 = pi1359 & ~pi1938;
  assign n14001 = pi2195 & n11837;
  assign n14002 = pi1359 & ~n11837;
  assign n14003 = ~n14001 & ~n14002;
  assign n14004 = pi1938 & ~n14003;
  assign po1410 = n14000 | n14004;
  assign n14006 = pi1360 & ~pi1938;
  assign n14007 = pi2186 & n11858;
  assign n14008 = pi1360 & ~n11858;
  assign n14009 = ~n14007 & ~n14008;
  assign n14010 = pi1938 & ~n14009;
  assign po1411 = n14006 | n14010;
  assign n14012 = pi1361 & ~pi1938;
  assign n14013 = pi2183 & n11858;
  assign n14014 = pi1361 & ~n11858;
  assign n14015 = ~n14013 & ~n14014;
  assign n14016 = pi1938 & ~n14015;
  assign po1412 = n14012 | n14016;
  assign n14018 = pi1362 & ~pi1938;
  assign n14019 = pi2172 & n11858;
  assign n14020 = pi1362 & ~n11858;
  assign n14021 = ~n14019 & ~n14020;
  assign n14022 = pi1938 & ~n14021;
  assign po1413 = n14018 | n14022;
  assign n14024 = pi1363 & ~pi1938;
  assign n14025 = pi2174 & n11858;
  assign n14026 = pi1363 & ~n11858;
  assign n14027 = ~n14025 & ~n14026;
  assign n14028 = pi1938 & ~n14027;
  assign po1414 = n14024 | n14028;
  assign n14030 = pi1364 & ~pi1938;
  assign n14031 = pi2197 & n11858;
  assign n14032 = pi1364 & ~n11858;
  assign n14033 = ~n14031 & ~n14032;
  assign n14034 = pi1938 & ~n14033;
  assign po1415 = n14030 | n14034;
  assign n14036 = pi1365 & ~pi1938;
  assign n14037 = pi2178 & n11858;
  assign n14038 = pi1365 & ~n11858;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = pi1938 & ~n14039;
  assign po1416 = n14036 | n14040;
  assign n14042 = pi1366 & ~pi1938;
  assign n14043 = pi2193 & n11858;
  assign n14044 = pi1366 & ~n11858;
  assign n14045 = ~n14043 & ~n14044;
  assign n14046 = pi1938 & ~n14045;
  assign po1417 = n14042 | n14046;
  assign n14048 = pi1367 & ~pi1938;
  assign n14049 = pi2189 & n11858;
  assign n14050 = pi1367 & ~n11858;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = pi1938 & ~n14051;
  assign po1418 = n14048 | n14052;
  assign n14054 = pi1368 & ~pi1938;
  assign n14055 = pi2179 & n11858;
  assign n14056 = pi1368 & ~n11858;
  assign n14057 = ~n14055 & ~n14056;
  assign n14058 = pi1938 & ~n14057;
  assign po1419 = n14054 | n14058;
  assign n14060 = pi1369 & ~pi1938;
  assign n14061 = pi2198 & n11858;
  assign n14062 = pi1369 & ~n11858;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = pi1938 & ~n14063;
  assign po1420 = n14060 | n14064;
  assign n14066 = pi1370 & ~pi1938;
  assign n14067 = pi2185 & n11858;
  assign n14068 = pi1370 & ~n11858;
  assign n14069 = ~n14067 & ~n14068;
  assign n14070 = pi1938 & ~n14069;
  assign po1421 = n14066 | n14070;
  assign n14072 = pi1371 & ~pi1938;
  assign n14073 = pi2187 & n11858;
  assign n14074 = pi1371 & ~n11858;
  assign n14075 = ~n14073 & ~n14074;
  assign n14076 = pi1938 & ~n14075;
  assign po1422 = n14072 | n14076;
  assign n14078 = pi1372 & ~pi1938;
  assign n14079 = pi2176 & n11858;
  assign n14080 = pi1372 & ~n11858;
  assign n14081 = ~n14079 & ~n14080;
  assign n14082 = pi1938 & ~n14081;
  assign po1423 = n14078 | n14082;
  assign n14084 = pi1373 & ~pi1938;
  assign n14085 = pi2169 & n11858;
  assign n14086 = pi1373 & ~n11858;
  assign n14087 = ~n14085 & ~n14086;
  assign n14088 = pi1938 & ~n14087;
  assign po1424 = n14084 | n14088;
  assign n14090 = pi1374 & ~pi1938;
  assign n14091 = pi2190 & n11858;
  assign n14092 = pi1374 & ~n11858;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = pi1938 & ~n14093;
  assign po1425 = n14090 | n14094;
  assign n14096 = pi1375 & ~pi1938;
  assign n14097 = pi2170 & n11858;
  assign n14098 = pi1375 & ~n11858;
  assign n14099 = ~n14097 & ~n14098;
  assign n14100 = pi1938 & ~n14099;
  assign po1426 = n14096 | n14100;
  assign n14102 = pi1376 & ~pi1938;
  assign n14103 = pi2182 & n11858;
  assign n14104 = pi1376 & ~n11858;
  assign n14105 = ~n14103 & ~n14104;
  assign n14106 = pi1938 & ~n14105;
  assign po1427 = n14102 | n14106;
  assign n14108 = pi1377 & ~pi1938;
  assign n14109 = pi2175 & n11858;
  assign n14110 = pi1377 & ~n11858;
  assign n14111 = ~n14109 & ~n14110;
  assign n14112 = pi1938 & ~n14111;
  assign po1428 = n14108 | n14112;
  assign n14114 = pi1378 & ~pi1938;
  assign n14115 = pi2191 & n11858;
  assign n14116 = pi1378 & ~n11858;
  assign n14117 = ~n14115 & ~n14116;
  assign n14118 = pi1938 & ~n14117;
  assign po1429 = n14114 | n14118;
  assign n14120 = pi1379 & ~pi1938;
  assign n14121 = pi2173 & n11858;
  assign n14122 = pi1379 & ~n11858;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = pi1938 & ~n14123;
  assign po1430 = n14120 | n14124;
  assign n14126 = pi1380 & ~pi1938;
  assign n14127 = pi2194 & n11858;
  assign n14128 = pi1380 & ~n11858;
  assign n14129 = ~n14127 & ~n14128;
  assign n14130 = pi1938 & ~n14129;
  assign po1431 = n14126 | n14130;
  assign n14132 = pi1381 & ~pi1938;
  assign n14133 = pi2167 & n11858;
  assign n14134 = pi1381 & ~n11858;
  assign n14135 = ~n14133 & ~n14134;
  assign n14136 = pi1938 & ~n14135;
  assign po1432 = n14132 | n14136;
  assign n14138 = pi1382 & ~pi1938;
  assign n14139 = pi2184 & n11858;
  assign n14140 = pi1382 & ~n11858;
  assign n14141 = ~n14139 & ~n14140;
  assign n14142 = pi1938 & ~n14141;
  assign po1433 = n14138 | n14142;
  assign n14144 = pi1383 & ~pi1938;
  assign n14145 = pi2166 & n11858;
  assign n14146 = pi1383 & ~n11858;
  assign n14147 = ~n14145 & ~n14146;
  assign n14148 = pi1938 & ~n14147;
  assign po1434 = n14144 | n14148;
  assign n14150 = pi1384 & ~pi1938;
  assign n14151 = pi2195 & n11858;
  assign n14152 = pi1384 & ~n11858;
  assign n14153 = ~n14151 & ~n14152;
  assign n14154 = pi1938 & ~n14153;
  assign po1435 = n14150 | n14154;
  assign n14156 = pi1385 & ~pi1937;
  assign n14157 = pi2185 & n11829;
  assign n14158 = pi1385 & ~n11829;
  assign n14159 = ~n14157 & ~n14158;
  assign n14160 = pi1937 & ~n14159;
  assign po1436 = n14156 | n14160;
  assign n14162 = pi1386 & ~pi1939;
  assign n14163 = pi2186 & n11745;
  assign n14164 = pi1386 & ~n11745;
  assign n14165 = ~n14163 & ~n14164;
  assign n14166 = pi1939 & ~n14165;
  assign po1437 = n14162 | n14166;
  assign n14168 = pi1387 & ~pi1939;
  assign n14169 = pi2183 & n11745;
  assign n14170 = pi1387 & ~n11745;
  assign n14171 = ~n14169 & ~n14170;
  assign n14172 = pi1939 & ~n14171;
  assign po1438 = n14168 | n14172;
  assign n14174 = pi1388 & ~pi1939;
  assign n14175 = pi2168 & n11745;
  assign n14176 = pi1388 & ~n11745;
  assign n14177 = ~n14175 & ~n14176;
  assign n14178 = pi1939 & ~n14177;
  assign po1439 = n14174 | n14178;
  assign n14180 = pi1389 & ~pi1939;
  assign n14181 = pi2174 & n11745;
  assign n14182 = pi1389 & ~n11745;
  assign n14183 = ~n14181 & ~n14182;
  assign n14184 = pi1939 & ~n14183;
  assign po1440 = n14180 | n14184;
  assign n14186 = pi1390 & ~pi1939;
  assign n14187 = pi2197 & n11745;
  assign n14188 = pi1390 & ~n11745;
  assign n14189 = ~n14187 & ~n14188;
  assign n14190 = pi1939 & ~n14189;
  assign po1441 = n14186 | n14190;
  assign n14192 = pi1391 & ~pi1940;
  assign n14193 = pi2197 & n11852;
  assign n14194 = pi1391 & ~n11852;
  assign n14195 = ~n14193 & ~n14194;
  assign n14196 = pi1940 & ~n14195;
  assign po1442 = n14192 | n14196;
  assign n14198 = pi1392 & ~pi1939;
  assign n14199 = pi2196 & n11745;
  assign n14200 = pi1392 & ~n11745;
  assign n14201 = ~n14199 & ~n14200;
  assign n14202 = pi1939 & ~n14201;
  assign po1443 = n14198 | n14202;
  assign n14204 = pi1393 & ~pi1939;
  assign n14205 = pi2193 & n11745;
  assign n14206 = pi1393 & ~n11745;
  assign n14207 = ~n14205 & ~n14206;
  assign n14208 = pi1939 & ~n14207;
  assign po1444 = n14204 | n14208;
  assign n14210 = pi1394 & ~pi1939;
  assign n14211 = pi2189 & n11745;
  assign n14212 = pi1394 & ~n11745;
  assign n14213 = ~n14211 & ~n14212;
  assign n14214 = pi1939 & ~n14213;
  assign po1445 = n14210 | n14214;
  assign n14216 = pi1395 & ~pi1939;
  assign n14217 = pi2198 & n11745;
  assign n14218 = pi1395 & ~n11745;
  assign n14219 = ~n14217 & ~n14218;
  assign n14220 = pi1939 & ~n14219;
  assign po1446 = n14216 | n14220;
  assign n14222 = pi1396 & ~pi1939;
  assign n14223 = pi2185 & n11745;
  assign n14224 = pi1396 & ~n11745;
  assign n14225 = ~n14223 & ~n14224;
  assign n14226 = pi1939 & ~n14225;
  assign po1447 = n14222 | n14226;
  assign n14228 = pi1397 & ~pi1939;
  assign n14229 = pi2187 & n11745;
  assign n14230 = pi1397 & ~n11745;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = pi1939 & ~n14231;
  assign po1448 = n14228 | n14232;
  assign n14234 = pi1398 & ~pi1939;
  assign n14235 = pi2171 & n11745;
  assign n14236 = pi1398 & ~n11745;
  assign n14237 = ~n14235 & ~n14236;
  assign n14238 = pi1939 & ~n14237;
  assign po1449 = n14234 | n14238;
  assign n14240 = pi1399 & ~pi1939;
  assign n14241 = pi2169 & n11745;
  assign n14242 = pi1399 & ~n11745;
  assign n14243 = ~n14241 & ~n14242;
  assign n14244 = pi1939 & ~n14243;
  assign po1450 = n14240 | n14244;
  assign n14246 = pi1400 & ~pi1939;
  assign n14247 = pi2190 & n11745;
  assign n14248 = pi1400 & ~n11745;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = pi1939 & ~n14249;
  assign po1451 = n14246 | n14250;
  assign n14252 = pi1401 & ~pi1939;
  assign n14253 = pi2181 & n11745;
  assign n14254 = pi1401 & ~n11745;
  assign n14255 = ~n14253 & ~n14254;
  assign n14256 = pi1939 & ~n14255;
  assign po1452 = n14252 | n14256;
  assign n14258 = pi1402 & ~pi1939;
  assign n14259 = pi2182 & n11745;
  assign n14260 = pi1402 & ~n11745;
  assign n14261 = ~n14259 & ~n14260;
  assign n14262 = pi1939 & ~n14261;
  assign po1453 = n14258 | n14262;
  assign n14264 = pi1403 & ~pi1939;
  assign n14265 = pi2175 & n11745;
  assign n14266 = pi1403 & ~n11745;
  assign n14267 = ~n14265 & ~n14266;
  assign n14268 = pi1939 & ~n14267;
  assign po1454 = n14264 | n14268;
  assign n14270 = pi1404 & ~pi1939;
  assign n14271 = pi2177 & n11745;
  assign n14272 = pi1404 & ~n11745;
  assign n14273 = ~n14271 & ~n14272;
  assign n14274 = pi1939 & ~n14273;
  assign po1455 = n14270 | n14274;
  assign n14276 = pi1405 & ~pi1939;
  assign n14277 = pi2173 & n11745;
  assign n14278 = pi1405 & ~n11745;
  assign n14279 = ~n14277 & ~n14278;
  assign n14280 = pi1939 & ~n14279;
  assign po1456 = n14276 | n14280;
  assign n14282 = pi1406 & ~pi1939;
  assign n14283 = pi2194 & n11745;
  assign n14284 = pi1406 & ~n11745;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = pi1939 & ~n14285;
  assign po1457 = n14282 | n14286;
  assign n14288 = pi1407 & ~pi1939;
  assign n14289 = pi2188 & n11745;
  assign n14290 = pi1407 & ~n11745;
  assign n14291 = ~n14289 & ~n14290;
  assign n14292 = pi1939 & ~n14291;
  assign po1458 = n14288 | n14292;
  assign n14294 = pi1408 & ~pi1939;
  assign n14295 = pi2184 & n11745;
  assign n14296 = pi1408 & ~n11745;
  assign n14297 = ~n14295 & ~n14296;
  assign n14298 = pi1939 & ~n14297;
  assign po1459 = n14294 | n14298;
  assign n14300 = pi1409 & ~pi1939;
  assign n14301 = pi2166 & n11745;
  assign n14302 = pi1409 & ~n11745;
  assign n14303 = ~n14301 & ~n14302;
  assign n14304 = pi1939 & ~n14303;
  assign po1460 = n14300 | n14304;
  assign n14306 = pi1410 & ~pi1939;
  assign n14307 = pi2192 & n11745;
  assign n14308 = pi1410 & ~n11745;
  assign n14309 = ~n14307 & ~n14308;
  assign n14310 = pi1939 & ~n14309;
  assign po1461 = n14306 | n14310;
  assign n14312 = pi1411 & ~pi1939;
  assign n14313 = pi2186 & n11746;
  assign n14314 = pi1411 & ~n11746;
  assign n14315 = ~n14313 & ~n14314;
  assign n14316 = pi1939 & ~n14315;
  assign po1462 = n14312 | n14316;
  assign n14318 = pi1412 & ~pi1939;
  assign n14319 = pi2183 & n11746;
  assign n14320 = pi1412 & ~n11746;
  assign n14321 = ~n14319 & ~n14320;
  assign n14322 = pi1939 & ~n14321;
  assign po1463 = n14318 | n14322;
  assign n14324 = pi1413 & ~pi1939;
  assign n14325 = pi2168 & n11746;
  assign n14326 = pi1413 & ~n11746;
  assign n14327 = ~n14325 & ~n14326;
  assign n14328 = pi1939 & ~n14327;
  assign po1464 = n14324 | n14328;
  assign n14330 = pi1414 & ~pi1939;
  assign n14331 = pi2174 & n11746;
  assign n14332 = pi1414 & ~n11746;
  assign n14333 = ~n14331 & ~n14332;
  assign n14334 = pi1939 & ~n14333;
  assign po1465 = n14330 | n14334;
  assign n14336 = pi1415 & ~pi1939;
  assign n14337 = pi2197 & n11746;
  assign n14338 = pi1415 & ~n11746;
  assign n14339 = ~n14337 & ~n14338;
  assign n14340 = pi1939 & ~n14339;
  assign po1466 = n14336 | n14340;
  assign n14342 = pi1416 & ~pi1939;
  assign n14343 = pi2196 & n11746;
  assign n14344 = pi1416 & ~n11746;
  assign n14345 = ~n14343 & ~n14344;
  assign n14346 = pi1939 & ~n14345;
  assign po1467 = n14342 | n14346;
  assign n14348 = pi1417 & ~pi1939;
  assign n14349 = pi2193 & n11746;
  assign n14350 = pi1417 & ~n11746;
  assign n14351 = ~n14349 & ~n14350;
  assign n14352 = pi1939 & ~n14351;
  assign po1468 = n14348 | n14352;
  assign n14354 = pi1418 & ~pi1939;
  assign n14355 = pi2189 & n11746;
  assign n14356 = pi1418 & ~n11746;
  assign n14357 = ~n14355 & ~n14356;
  assign n14358 = pi1939 & ~n14357;
  assign po1469 = n14354 | n14358;
  assign n14360 = pi1419 & ~pi1939;
  assign n14361 = pi2198 & n11746;
  assign n14362 = pi1419 & ~n11746;
  assign n14363 = ~n14361 & ~n14362;
  assign n14364 = pi1939 & ~n14363;
  assign po1470 = n14360 | n14364;
  assign n14366 = pi1420 & ~pi1939;
  assign n14367 = pi2185 & n11746;
  assign n14368 = pi1420 & ~n11746;
  assign n14369 = ~n14367 & ~n14368;
  assign n14370 = pi1939 & ~n14369;
  assign po1471 = n14366 | n14370;
  assign n14372 = pi1421 & ~pi1939;
  assign n14373 = pi2187 & n11746;
  assign n14374 = pi1421 & ~n11746;
  assign n14375 = ~n14373 & ~n14374;
  assign n14376 = pi1939 & ~n14375;
  assign po1472 = n14372 | n14376;
  assign n14378 = pi1422 & ~pi1939;
  assign n14379 = pi2171 & n11746;
  assign n14380 = pi1422 & ~n11746;
  assign n14381 = ~n14379 & ~n14380;
  assign n14382 = pi1939 & ~n14381;
  assign po1473 = n14378 | n14382;
  assign n14384 = pi1423 & ~pi1939;
  assign n14385 = pi2169 & n11746;
  assign n14386 = pi1423 & ~n11746;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = pi1939 & ~n14387;
  assign po1474 = n14384 | n14388;
  assign n14390 = pi1424 & ~pi1939;
  assign n14391 = pi2190 & n11746;
  assign n14392 = pi1424 & ~n11746;
  assign n14393 = ~n14391 & ~n14392;
  assign n14394 = pi1939 & ~n14393;
  assign po1475 = n14390 | n14394;
  assign n14396 = pi1425 & ~pi1939;
  assign n14397 = pi2181 & n11746;
  assign n14398 = pi1425 & ~n11746;
  assign n14399 = ~n14397 & ~n14398;
  assign n14400 = pi1939 & ~n14399;
  assign po1476 = n14396 | n14400;
  assign n14402 = pi1426 & ~pi1939;
  assign n14403 = pi2182 & n11746;
  assign n14404 = pi1426 & ~n11746;
  assign n14405 = ~n14403 & ~n14404;
  assign n14406 = pi1939 & ~n14405;
  assign po1477 = n14402 | n14406;
  assign n14408 = pi1427 & ~pi1939;
  assign n14409 = pi2175 & n11746;
  assign n14410 = pi1427 & ~n11746;
  assign n14411 = ~n14409 & ~n14410;
  assign n14412 = pi1939 & ~n14411;
  assign po1478 = n14408 | n14412;
  assign n14414 = pi1428 & ~pi1939;
  assign n14415 = pi2177 & n11746;
  assign n14416 = pi1428 & ~n11746;
  assign n14417 = ~n14415 & ~n14416;
  assign n14418 = pi1939 & ~n14417;
  assign po1479 = n14414 | n14418;
  assign n14420 = pi1429 & ~pi1939;
  assign n14421 = pi2173 & n11746;
  assign n14422 = pi1429 & ~n11746;
  assign n14423 = ~n14421 & ~n14422;
  assign n14424 = pi1939 & ~n14423;
  assign po1480 = n14420 | n14424;
  assign n14426 = pi1430 & ~pi1939;
  assign n14427 = pi2194 & n11746;
  assign n14428 = pi1430 & ~n11746;
  assign n14429 = ~n14427 & ~n14428;
  assign n14430 = pi1939 & ~n14429;
  assign po1481 = n14426 | n14430;
  assign n14432 = pi1431 & ~pi1939;
  assign n14433 = pi2167 & n11746;
  assign n14434 = pi1431 & ~n11746;
  assign n14435 = ~n14433 & ~n14434;
  assign n14436 = pi1939 & ~n14435;
  assign po1482 = n14432 | n14436;
  assign n14438 = pi1432 & ~pi1939;
  assign n14439 = pi2188 & n11746;
  assign n14440 = pi1432 & ~n11746;
  assign n14441 = ~n14439 & ~n14440;
  assign n14442 = pi1939 & ~n14441;
  assign po1483 = n14438 | n14442;
  assign n14444 = pi1433 & ~pi1939;
  assign n14445 = pi2184 & n11746;
  assign n14446 = pi1433 & ~n11746;
  assign n14447 = ~n14445 & ~n14446;
  assign n14448 = pi1939 & ~n14447;
  assign po1484 = n14444 | n14448;
  assign n14450 = pi1434 & ~pi1939;
  assign n14451 = pi2166 & n11746;
  assign n14452 = pi1434 & ~n11746;
  assign n14453 = ~n14451 & ~n14452;
  assign n14454 = pi1939 & ~n14453;
  assign po1485 = n14450 | n14454;
  assign n14456 = pi1435 & ~pi1939;
  assign n14457 = pi2192 & n11746;
  assign n14458 = pi1435 & ~n11746;
  assign n14459 = ~n14457 & ~n14458;
  assign n14460 = pi1939 & ~n14459;
  assign po1486 = n14456 | n14460;
  assign n14462 = pi1436 & ~pi1939;
  assign n14463 = pi2186 & n11786;
  assign n14464 = pi1436 & ~n11786;
  assign n14465 = ~n14463 & ~n14464;
  assign n14466 = pi1939 & ~n14465;
  assign po1487 = n14462 | n14466;
  assign n14468 = pi1437 & ~pi1939;
  assign n14469 = pi2183 & n11786;
  assign n14470 = pi1437 & ~n11786;
  assign n14471 = ~n14469 & ~n14470;
  assign n14472 = pi1939 & ~n14471;
  assign po1488 = n14468 | n14472;
  assign n14474 = pi1438 & ~pi1939;
  assign n14475 = pi2168 & n11786;
  assign n14476 = pi1438 & ~n11786;
  assign n14477 = ~n14475 & ~n14476;
  assign n14478 = pi1939 & ~n14477;
  assign po1489 = n14474 | n14478;
  assign n14480 = pi1439 & ~pi1939;
  assign n14481 = pi2174 & n11786;
  assign n14482 = pi1439 & ~n11786;
  assign n14483 = ~n14481 & ~n14482;
  assign n14484 = pi1939 & ~n14483;
  assign po1490 = n14480 | n14484;
  assign n14486 = pi1440 & ~pi1939;
  assign n14487 = pi2197 & n11786;
  assign n14488 = pi1440 & ~n11786;
  assign n14489 = ~n14487 & ~n14488;
  assign n14490 = pi1939 & ~n14489;
  assign po1491 = n14486 | n14490;
  assign n14492 = pi1441 & ~pi1939;
  assign n14493 = pi2196 & n11786;
  assign n14494 = pi1441 & ~n11786;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = pi1939 & ~n14495;
  assign po1492 = n14492 | n14496;
  assign n14498 = pi1442 & ~pi1939;
  assign n14499 = pi2193 & n11786;
  assign n14500 = pi1442 & ~n11786;
  assign n14501 = ~n14499 & ~n14500;
  assign n14502 = pi1939 & ~n14501;
  assign po1493 = n14498 | n14502;
  assign n14504 = pi1443 & ~pi1939;
  assign n14505 = pi2189 & n11786;
  assign n14506 = pi1443 & ~n11786;
  assign n14507 = ~n14505 & ~n14506;
  assign n14508 = pi1939 & ~n14507;
  assign po1494 = n14504 | n14508;
  assign n14510 = pi1444 & ~pi1939;
  assign n14511 = pi2198 & n11786;
  assign n14512 = pi1444 & ~n11786;
  assign n14513 = ~n14511 & ~n14512;
  assign n14514 = pi1939 & ~n14513;
  assign po1495 = n14510 | n14514;
  assign n14516 = pi1445 & ~pi1939;
  assign n14517 = pi2185 & n11786;
  assign n14518 = pi1445 & ~n11786;
  assign n14519 = ~n14517 & ~n14518;
  assign n14520 = pi1939 & ~n14519;
  assign po1496 = n14516 | n14520;
  assign n14522 = pi1446 & ~pi1939;
  assign n14523 = pi2187 & n11786;
  assign n14524 = pi1446 & ~n11786;
  assign n14525 = ~n14523 & ~n14524;
  assign n14526 = pi1939 & ~n14525;
  assign po1497 = n14522 | n14526;
  assign n14528 = pi1447 & ~pi1936;
  assign n14529 = pi1447 & ~n12004;
  assign n14530 = pi2193 & n12004;
  assign n14531 = ~n14529 & ~n14530;
  assign n14532 = pi1936 & ~n14531;
  assign po1498 = n14528 | n14532;
  assign n14534 = pi1448 & ~pi1939;
  assign n14535 = pi2171 & n11786;
  assign n14536 = pi1448 & ~n11786;
  assign n14537 = ~n14535 & ~n14536;
  assign n14538 = pi1939 & ~n14537;
  assign po1499 = n14534 | n14538;
  assign n14540 = pi1449 & ~pi1939;
  assign n14541 = pi2169 & n11786;
  assign n14542 = pi1449 & ~n11786;
  assign n14543 = ~n14541 & ~n14542;
  assign n14544 = pi1939 & ~n14543;
  assign po1500 = n14540 | n14544;
  assign n14546 = pi1450 & ~pi1939;
  assign n14547 = pi2190 & n11786;
  assign n14548 = pi1450 & ~n11786;
  assign n14549 = ~n14547 & ~n14548;
  assign n14550 = pi1939 & ~n14549;
  assign po1501 = n14546 | n14550;
  assign n14552 = pi1451 & ~pi1939;
  assign n14553 = pi2181 & n11786;
  assign n14554 = pi1451 & ~n11786;
  assign n14555 = ~n14553 & ~n14554;
  assign n14556 = pi1939 & ~n14555;
  assign po1502 = n14552 | n14556;
  assign n14558 = pi1452 & ~pi1939;
  assign n14559 = pi2182 & n11786;
  assign n14560 = pi1452 & ~n11786;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = pi1939 & ~n14561;
  assign po1503 = n14558 | n14562;
  assign n14564 = pi1453 & ~pi1939;
  assign n14565 = pi2175 & n11786;
  assign n14566 = pi1453 & ~n11786;
  assign n14567 = ~n14565 & ~n14566;
  assign n14568 = pi1939 & ~n14567;
  assign po1504 = n14564 | n14568;
  assign n14570 = pi1454 & ~pi1939;
  assign n14571 = pi2177 & n11786;
  assign n14572 = pi1454 & ~n11786;
  assign n14573 = ~n14571 & ~n14572;
  assign n14574 = pi1939 & ~n14573;
  assign po1505 = n14570 | n14574;
  assign n14576 = pi1455 & ~pi1939;
  assign n14577 = pi2173 & n11786;
  assign n14578 = pi1455 & ~n11786;
  assign n14579 = ~n14577 & ~n14578;
  assign n14580 = pi1939 & ~n14579;
  assign po1506 = n14576 | n14580;
  assign n14582 = pi1456 & ~pi1939;
  assign n14583 = pi2194 & n11786;
  assign n14584 = pi1456 & ~n11786;
  assign n14585 = ~n14583 & ~n14584;
  assign n14586 = pi1939 & ~n14585;
  assign po1507 = n14582 | n14586;
  assign n14588 = pi1457 & ~pi1939;
  assign n14589 = pi2188 & n11786;
  assign n14590 = pi1457 & ~n11786;
  assign n14591 = ~n14589 & ~n14590;
  assign n14592 = pi1939 & ~n14591;
  assign po1508 = n14588 | n14592;
  assign n14594 = pi1458 & ~pi1939;
  assign n14595 = pi2184 & n11786;
  assign n14596 = pi1458 & ~n11786;
  assign n14597 = ~n14595 & ~n14596;
  assign n14598 = pi1939 & ~n14597;
  assign po1509 = n14594 | n14598;
  assign n14600 = pi1459 & ~pi1939;
  assign n14601 = pi2166 & n11786;
  assign n14602 = pi1459 & ~n11786;
  assign n14603 = ~n14601 & ~n14602;
  assign n14604 = pi1939 & ~n14603;
  assign po1510 = n14600 | n14604;
  assign n14606 = pi1460 & ~pi1939;
  assign n14607 = pi2192 & n11786;
  assign n14608 = pi1460 & ~n11786;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = pi1939 & ~n14609;
  assign po1511 = n14606 | n14610;
  assign n14612 = pi1461 & ~pi1936;
  assign n14613 = pi2186 & n11844;
  assign n14614 = pi1461 & ~n11844;
  assign n14615 = ~n14613 & ~n14614;
  assign n14616 = pi1936 & ~n14615;
  assign po1512 = n14612 | n14616;
  assign n14618 = pi1462 & ~pi1936;
  assign n14619 = pi2183 & n11844;
  assign n14620 = pi1462 & ~n11844;
  assign n14621 = ~n14619 & ~n14620;
  assign n14622 = pi1936 & ~n14621;
  assign po1513 = n14618 | n14622;
  assign n14624 = pi1463 & ~pi1936;
  assign n14625 = pi2168 & n11844;
  assign n14626 = pi1463 & ~n11844;
  assign n14627 = ~n14625 & ~n14626;
  assign n14628 = pi1936 & ~n14627;
  assign po1514 = n14624 | n14628;
  assign n14630 = pi1464 & ~pi1936;
  assign n14631 = pi2174 & n11844;
  assign n14632 = pi1464 & ~n11844;
  assign n14633 = ~n14631 & ~n14632;
  assign n14634 = pi1936 & ~n14633;
  assign po1515 = n14630 | n14634;
  assign n14636 = pi1465 & ~pi1936;
  assign n14637 = pi2197 & n11844;
  assign n14638 = pi1465 & ~n11844;
  assign n14639 = ~n14637 & ~n14638;
  assign n14640 = pi1936 & ~n14639;
  assign po1516 = n14636 | n14640;
  assign n14642 = pi1466 & ~pi1936;
  assign n14643 = pi2196 & n11844;
  assign n14644 = pi1466 & ~n11844;
  assign n14645 = ~n14643 & ~n14644;
  assign n14646 = pi1936 & ~n14645;
  assign po1517 = n14642 | n14646;
  assign n14648 = pi1467 & ~pi1936;
  assign n14649 = pi2193 & n11844;
  assign n14650 = pi1467 & ~n11844;
  assign n14651 = ~n14649 & ~n14650;
  assign n14652 = pi1936 & ~n14651;
  assign po1518 = n14648 | n14652;
  assign n14654 = pi1468 & ~pi1936;
  assign n14655 = pi2189 & n11844;
  assign n14656 = pi1468 & ~n11844;
  assign n14657 = ~n14655 & ~n14656;
  assign n14658 = pi1936 & ~n14657;
  assign po1519 = n14654 | n14658;
  assign n14660 = pi1469 & ~pi1936;
  assign n14661 = pi2179 & n11844;
  assign n14662 = pi1469 & ~n11844;
  assign n14663 = ~n14661 & ~n14662;
  assign n14664 = pi1936 & ~n14663;
  assign po1520 = n14660 | n14664;
  assign n14666 = pi1470 & ~pi1936;
  assign n14667 = pi2198 & n11844;
  assign n14668 = pi1470 & ~n11844;
  assign n14669 = ~n14667 & ~n14668;
  assign n14670 = pi1936 & ~n14669;
  assign po1521 = n14666 | n14670;
  assign n14672 = pi1471 & ~pi1936;
  assign n14673 = pi2185 & n11844;
  assign n14674 = pi1471 & ~n11844;
  assign n14675 = ~n14673 & ~n14674;
  assign n14676 = pi1936 & ~n14675;
  assign po1522 = n14672 | n14676;
  assign n14678 = pi1472 & ~pi1936;
  assign n14679 = pi2187 & n11844;
  assign n14680 = pi1472 & ~n11844;
  assign n14681 = ~n14679 & ~n14680;
  assign n14682 = pi1936 & ~n14681;
  assign po1523 = n14678 | n14682;
  assign n14684 = pi1473 & ~pi1936;
  assign n14685 = pi2171 & n11844;
  assign n14686 = pi1473 & ~n11844;
  assign n14687 = ~n14685 & ~n14686;
  assign n14688 = pi1936 & ~n14687;
  assign po1524 = n14684 | n14688;
  assign n14690 = pi1474 & ~pi1936;
  assign n14691 = pi2169 & n11844;
  assign n14692 = pi1474 & ~n11844;
  assign n14693 = ~n14691 & ~n14692;
  assign n14694 = pi1936 & ~n14693;
  assign po1525 = n14690 | n14694;
  assign n14696 = pi1475 & ~pi1936;
  assign n14697 = pi2190 & n11844;
  assign n14698 = pi1475 & ~n11844;
  assign n14699 = ~n14697 & ~n14698;
  assign n14700 = pi1936 & ~n14699;
  assign po1526 = n14696 | n14700;
  assign n14702 = pi1476 & ~pi1936;
  assign n14703 = pi2181 & n11844;
  assign n14704 = pi1476 & ~n11844;
  assign n14705 = ~n14703 & ~n14704;
  assign n14706 = pi1936 & ~n14705;
  assign po1527 = n14702 | n14706;
  assign n14708 = pi1477 & ~pi1936;
  assign n14709 = pi2182 & n11844;
  assign n14710 = pi1477 & ~n11844;
  assign n14711 = ~n14709 & ~n14710;
  assign n14712 = pi1936 & ~n14711;
  assign po1528 = n14708 | n14712;
  assign n14714 = pi1478 & ~pi1936;
  assign n14715 = pi2175 & n11844;
  assign n14716 = pi1478 & ~n11844;
  assign n14717 = ~n14715 & ~n14716;
  assign n14718 = pi1936 & ~n14717;
  assign po1529 = n14714 | n14718;
  assign n14720 = pi1479 & ~pi1936;
  assign n14721 = pi2177 & n11844;
  assign n14722 = pi1479 & ~n11844;
  assign n14723 = ~n14721 & ~n14722;
  assign n14724 = pi1936 & ~n14723;
  assign po1530 = n14720 | n14724;
  assign n14726 = pi1480 & ~pi1936;
  assign n14727 = pi2173 & n11844;
  assign n14728 = pi1480 & ~n11844;
  assign n14729 = ~n14727 & ~n14728;
  assign n14730 = pi1936 & ~n14729;
  assign po1531 = n14726 | n14730;
  assign n14732 = pi1481 & ~pi1936;
  assign n14733 = pi2194 & n11844;
  assign n14734 = pi1481 & ~n11844;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = pi1936 & ~n14735;
  assign po1532 = n14732 | n14736;
  assign n14738 = pi1482 & ~pi1936;
  assign n14739 = pi2188 & n11844;
  assign n14740 = pi1482 & ~n11844;
  assign n14741 = ~n14739 & ~n14740;
  assign n14742 = pi1936 & ~n14741;
  assign po1533 = n14738 | n14742;
  assign n14744 = pi1483 & ~pi1936;
  assign n14745 = pi2184 & n11844;
  assign n14746 = pi1483 & ~n11844;
  assign n14747 = ~n14745 & ~n14746;
  assign n14748 = pi1936 & ~n14747;
  assign po1534 = n14744 | n14748;
  assign n14750 = pi1484 & ~pi1936;
  assign n14751 = pi2166 & n11844;
  assign n14752 = pi1484 & ~n11844;
  assign n14753 = ~n14751 & ~n14752;
  assign n14754 = pi1936 & ~n14753;
  assign po1535 = n14750 | n14754;
  assign n14756 = pi1485 & ~pi1936;
  assign n14757 = pi2192 & n11844;
  assign n14758 = pi1485 & ~n11844;
  assign n14759 = ~n14757 & ~n14758;
  assign n14760 = pi1936 & ~n14759;
  assign po1536 = n14756 | n14760;
  assign n14762 = pi1486 & ~pi1936;
  assign n14763 = pi2186 & n11845;
  assign n14764 = pi1486 & ~n11845;
  assign n14765 = ~n14763 & ~n14764;
  assign n14766 = pi1936 & ~n14765;
  assign po1537 = n14762 | n14766;
  assign n14768 = pi1487 & ~pi1936;
  assign n14769 = pi2183 & n11845;
  assign n14770 = pi1487 & ~n11845;
  assign n14771 = ~n14769 & ~n14770;
  assign n14772 = pi1936 & ~n14771;
  assign po1538 = n14768 | n14772;
  assign n14774 = pi1488 & ~pi1936;
  assign n14775 = pi2168 & n11845;
  assign n14776 = pi1488 & ~n11845;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = pi1936 & ~n14777;
  assign po1539 = n14774 | n14778;
  assign n14780 = pi1489 & ~pi1936;
  assign n14781 = pi2174 & n11845;
  assign n14782 = pi1489 & ~n11845;
  assign n14783 = ~n14781 & ~n14782;
  assign n14784 = pi1936 & ~n14783;
  assign po1540 = n14780 | n14784;
  assign n14786 = pi1490 & ~pi1936;
  assign n14787 = pi2197 & n11845;
  assign n14788 = pi1490 & ~n11845;
  assign n14789 = ~n14787 & ~n14788;
  assign n14790 = pi1936 & ~n14789;
  assign po1541 = n14786 | n14790;
  assign n14792 = pi1491 & ~pi1936;
  assign n14793 = pi2196 & n11845;
  assign n14794 = pi1491 & ~n11845;
  assign n14795 = ~n14793 & ~n14794;
  assign n14796 = pi1936 & ~n14795;
  assign po1542 = n14792 | n14796;
  assign n14798 = pi1492 & ~pi1936;
  assign n14799 = pi2193 & n11845;
  assign n14800 = pi1492 & ~n11845;
  assign n14801 = ~n14799 & ~n14800;
  assign n14802 = pi1936 & ~n14801;
  assign po1543 = n14798 | n14802;
  assign n14804 = pi1493 & ~pi1936;
  assign n14805 = pi2189 & n11845;
  assign n14806 = pi1493 & ~n11845;
  assign n14807 = ~n14805 & ~n14806;
  assign n14808 = pi1936 & ~n14807;
  assign po1544 = n14804 | n14808;
  assign n14810 = pi1494 & ~pi1936;
  assign n14811 = pi2198 & n11845;
  assign n14812 = pi1494 & ~n11845;
  assign n14813 = ~n14811 & ~n14812;
  assign n14814 = pi1936 & ~n14813;
  assign po1545 = n14810 | n14814;
  assign n14816 = pi1495 & ~pi1936;
  assign n14817 = pi2185 & n11845;
  assign n14818 = pi1495 & ~n11845;
  assign n14819 = ~n14817 & ~n14818;
  assign n14820 = pi1936 & ~n14819;
  assign po1546 = n14816 | n14820;
  assign n14822 = pi1496 & ~pi1936;
  assign n14823 = pi2187 & n11845;
  assign n14824 = pi1496 & ~n11845;
  assign n14825 = ~n14823 & ~n14824;
  assign n14826 = pi1936 & ~n14825;
  assign po1547 = n14822 | n14826;
  assign n14828 = pi1497 & ~pi1936;
  assign n14829 = pi2171 & n11845;
  assign n14830 = pi1497 & ~n11845;
  assign n14831 = ~n14829 & ~n14830;
  assign n14832 = pi1936 & ~n14831;
  assign po1548 = n14828 | n14832;
  assign n14834 = pi1498 & ~pi1936;
  assign n14835 = pi2169 & n11845;
  assign n14836 = pi1498 & ~n11845;
  assign n14837 = ~n14835 & ~n14836;
  assign n14838 = pi1936 & ~n14837;
  assign po1549 = n14834 | n14838;
  assign n14840 = pi1499 & ~pi1936;
  assign n14841 = pi2190 & n11845;
  assign n14842 = pi1499 & ~n11845;
  assign n14843 = ~n14841 & ~n14842;
  assign n14844 = pi1936 & ~n14843;
  assign po1550 = n14840 | n14844;
  assign n14846 = pi1500 & ~pi1936;
  assign n14847 = pi2181 & n11845;
  assign n14848 = pi1500 & ~n11845;
  assign n14849 = ~n14847 & ~n14848;
  assign n14850 = pi1936 & ~n14849;
  assign po1551 = n14846 | n14850;
  assign n14852 = pi1501 & ~pi1936;
  assign n14853 = pi2182 & n11845;
  assign n14854 = pi1501 & ~n11845;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = pi1936 & ~n14855;
  assign po1552 = n14852 | n14856;
  assign n14858 = pi1502 & ~pi1936;
  assign n14859 = pi2175 & n11845;
  assign n14860 = pi1502 & ~n11845;
  assign n14861 = ~n14859 & ~n14860;
  assign n14862 = pi1936 & ~n14861;
  assign po1553 = n14858 | n14862;
  assign n14864 = pi1503 & ~pi1936;
  assign n14865 = pi2177 & n11845;
  assign n14866 = pi1503 & ~n11845;
  assign n14867 = ~n14865 & ~n14866;
  assign n14868 = pi1936 & ~n14867;
  assign po1554 = n14864 | n14868;
  assign n14870 = pi1504 & ~pi1936;
  assign n14871 = pi2173 & n11845;
  assign n14872 = pi1504 & ~n11845;
  assign n14873 = ~n14871 & ~n14872;
  assign n14874 = pi1936 & ~n14873;
  assign po1555 = n14870 | n14874;
  assign n14876 = pi1505 & ~pi1936;
  assign n14877 = pi2194 & n11845;
  assign n14878 = pi1505 & ~n11845;
  assign n14879 = ~n14877 & ~n14878;
  assign n14880 = pi1936 & ~n14879;
  assign po1556 = n14876 | n14880;
  assign n14882 = pi1506 & ~pi1936;
  assign n14883 = pi2188 & n11845;
  assign n14884 = pi1506 & ~n11845;
  assign n14885 = ~n14883 & ~n14884;
  assign n14886 = pi1936 & ~n14885;
  assign po1557 = n14882 | n14886;
  assign n14888 = pi1507 & ~pi1936;
  assign n14889 = pi2184 & n11845;
  assign n14890 = pi1507 & ~n11845;
  assign n14891 = ~n14889 & ~n14890;
  assign n14892 = pi1936 & ~n14891;
  assign po1558 = n14888 | n14892;
  assign n14894 = pi1508 & ~pi1936;
  assign n14895 = pi2166 & n11845;
  assign n14896 = pi1508 & ~n11845;
  assign n14897 = ~n14895 & ~n14896;
  assign n14898 = pi1936 & ~n14897;
  assign po1559 = n14894 | n14898;
  assign n14900 = pi1509 & ~pi1936;
  assign n14901 = pi2192 & n11845;
  assign n14902 = pi1509 & ~n11845;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = pi1936 & ~n14903;
  assign po1560 = n14900 | n14904;
  assign n14906 = pi1510 & ~pi1936;
  assign n14907 = pi2186 & n11751;
  assign n14908 = pi1510 & ~n11751;
  assign n14909 = ~n14907 & ~n14908;
  assign n14910 = pi1936 & ~n14909;
  assign po1561 = n14906 | n14910;
  assign n14912 = pi1511 & ~pi1936;
  assign n14913 = pi2183 & n11751;
  assign n14914 = pi1511 & ~n11751;
  assign n14915 = ~n14913 & ~n14914;
  assign n14916 = pi1936 & ~n14915;
  assign po1562 = n14912 | n14916;
  assign n14918 = pi1512 & ~pi1936;
  assign n14919 = pi2168 & n11751;
  assign n14920 = pi1512 & ~n11751;
  assign n14921 = ~n14919 & ~n14920;
  assign n14922 = pi1936 & ~n14921;
  assign po1563 = n14918 | n14922;
  assign n14924 = pi1513 & ~pi1936;
  assign n14925 = pi2174 & n11751;
  assign n14926 = pi1513 & ~n11751;
  assign n14927 = ~n14925 & ~n14926;
  assign n14928 = pi1936 & ~n14927;
  assign po1564 = n14924 | n14928;
  assign n14930 = pi1514 & ~pi1936;
  assign n14931 = pi2197 & n11751;
  assign n14932 = pi1514 & ~n11751;
  assign n14933 = ~n14931 & ~n14932;
  assign n14934 = pi1936 & ~n14933;
  assign po1565 = n14930 | n14934;
  assign n14936 = pi1515 & ~pi1936;
  assign n14937 = pi2196 & n11751;
  assign n14938 = pi1515 & ~n11751;
  assign n14939 = ~n14937 & ~n14938;
  assign n14940 = pi1936 & ~n14939;
  assign po1566 = n14936 | n14940;
  assign n14942 = pi1516 & ~pi1936;
  assign n14943 = pi2193 & n11751;
  assign n14944 = pi1516 & ~n11751;
  assign n14945 = ~n14943 & ~n14944;
  assign n14946 = pi1936 & ~n14945;
  assign po1567 = n14942 | n14946;
  assign n14948 = pi1517 & ~pi1936;
  assign n14949 = pi2189 & n11751;
  assign n14950 = pi1517 & ~n11751;
  assign n14951 = ~n14949 & ~n14950;
  assign n14952 = pi1936 & ~n14951;
  assign po1568 = n14948 | n14952;
  assign n14954 = pi1518 & ~pi1936;
  assign n14955 = pi2198 & n11751;
  assign n14956 = pi1518 & ~n11751;
  assign n14957 = ~n14955 & ~n14956;
  assign n14958 = pi1936 & ~n14957;
  assign po1569 = n14954 | n14958;
  assign n14960 = pi1519 & ~pi1936;
  assign n14961 = pi2185 & n11751;
  assign n14962 = pi1519 & ~n11751;
  assign n14963 = ~n14961 & ~n14962;
  assign n14964 = pi1936 & ~n14963;
  assign po1570 = n14960 | n14964;
  assign n14966 = pi1520 & ~pi1936;
  assign n14967 = pi2187 & n11751;
  assign n14968 = pi1520 & ~n11751;
  assign n14969 = ~n14967 & ~n14968;
  assign n14970 = pi1936 & ~n14969;
  assign po1571 = n14966 | n14970;
  assign n14972 = pi1521 & ~pi1936;
  assign n14973 = pi2171 & n11751;
  assign n14974 = pi1521 & ~n11751;
  assign n14975 = ~n14973 & ~n14974;
  assign n14976 = pi1936 & ~n14975;
  assign po1572 = n14972 | n14976;
  assign n14978 = pi1522 & ~pi1936;
  assign n14979 = pi2169 & n11751;
  assign n14980 = pi1522 & ~n11751;
  assign n14981 = ~n14979 & ~n14980;
  assign n14982 = pi1936 & ~n14981;
  assign po1573 = n14978 | n14982;
  assign n14984 = pi1523 & ~pi1936;
  assign n14985 = pi2190 & n11751;
  assign n14986 = pi1523 & ~n11751;
  assign n14987 = ~n14985 & ~n14986;
  assign n14988 = pi1936 & ~n14987;
  assign po1574 = n14984 | n14988;
  assign n14990 = pi1524 & ~pi1936;
  assign n14991 = pi2181 & n11751;
  assign n14992 = pi1524 & ~n11751;
  assign n14993 = ~n14991 & ~n14992;
  assign n14994 = pi1936 & ~n14993;
  assign po1575 = n14990 | n14994;
  assign n14996 = pi1525 & ~pi1936;
  assign n14997 = pi2182 & n11751;
  assign n14998 = pi1525 & ~n11751;
  assign n14999 = ~n14997 & ~n14998;
  assign n15000 = pi1936 & ~n14999;
  assign po1576 = n14996 | n15000;
  assign n15002 = pi1526 & ~pi1936;
  assign n15003 = pi2175 & n11751;
  assign n15004 = pi1526 & ~n11751;
  assign n15005 = ~n15003 & ~n15004;
  assign n15006 = pi1936 & ~n15005;
  assign po1577 = n15002 | n15006;
  assign n15008 = pi1527 & ~pi1936;
  assign n15009 = pi2177 & n11751;
  assign n15010 = pi1527 & ~n11751;
  assign n15011 = ~n15009 & ~n15010;
  assign n15012 = pi1936 & ~n15011;
  assign po1578 = n15008 | n15012;
  assign n15014 = pi1528 & ~pi1936;
  assign n15015 = pi2173 & n11751;
  assign n15016 = pi1528 & ~n11751;
  assign n15017 = ~n15015 & ~n15016;
  assign n15018 = pi1936 & ~n15017;
  assign po1579 = n15014 | n15018;
  assign n15020 = pi1529 & ~pi1936;
  assign n15021 = pi2194 & n11751;
  assign n15022 = pi1529 & ~n11751;
  assign n15023 = ~n15021 & ~n15022;
  assign n15024 = pi1936 & ~n15023;
  assign po1580 = n15020 | n15024;
  assign n15026 = pi1530 & ~pi1936;
  assign n15027 = pi2188 & n11751;
  assign n15028 = pi1530 & ~n11751;
  assign n15029 = ~n15027 & ~n15028;
  assign n15030 = pi1936 & ~n15029;
  assign po1581 = n15026 | n15030;
  assign n15032 = pi1531 & ~pi1936;
  assign n15033 = pi2184 & n11751;
  assign n15034 = pi1531 & ~n11751;
  assign n15035 = ~n15033 & ~n15034;
  assign n15036 = pi1936 & ~n15035;
  assign po1582 = n15032 | n15036;
  assign n15038 = pi1532 & ~pi1936;
  assign n15039 = pi2166 & n11751;
  assign n15040 = pi1532 & ~n11751;
  assign n15041 = ~n15039 & ~n15040;
  assign n15042 = pi1936 & ~n15041;
  assign po1583 = n15038 | n15042;
  assign n15044 = pi1533 & ~pi1936;
  assign n15045 = pi2192 & n11751;
  assign n15046 = pi1533 & ~n11751;
  assign n15047 = ~n15045 & ~n15046;
  assign n15048 = pi1936 & ~n15047;
  assign po1584 = n15044 | n15048;
  assign n15050 = pi1534 & ~pi1937;
  assign n15051 = pi2195 & n11778;
  assign n15052 = pi1534 & ~n11778;
  assign n15053 = ~n15051 & ~n15052;
  assign n15054 = pi1937 & ~n15053;
  assign po1585 = n15050 | n15054;
  assign n15056 = pi1535 & ~pi1940;
  assign n15057 = pi2186 & n11852;
  assign n15058 = pi1535 & ~n11852;
  assign n15059 = ~n15057 & ~n15058;
  assign n15060 = pi1940 & ~n15059;
  assign po1586 = n15056 | n15060;
  assign n15062 = pi1536 & ~pi1940;
  assign n15063 = pi2172 & n11852;
  assign n15064 = pi1536 & ~n11852;
  assign n15065 = ~n15063 & ~n15064;
  assign n15066 = pi1940 & ~n15065;
  assign po1587 = n15062 | n15066;
  assign n15068 = pi1537 & ~pi1940;
  assign n15069 = pi2168 & n11852;
  assign n15070 = pi1537 & ~n11852;
  assign n15071 = ~n15069 & ~n15070;
  assign n15072 = pi1940 & ~n15071;
  assign po1588 = n15068 | n15072;
  assign n15074 = pi1538 & ~pi1940;
  assign n15075 = pi2174 & n11852;
  assign n15076 = pi1538 & ~n11852;
  assign n15077 = ~n15075 & ~n15076;
  assign n15078 = pi1940 & ~n15077;
  assign po1589 = n15074 | n15078;
  assign n15080 = pi1539 & ~pi1940;
  assign n15081 = pi2178 & n11852;
  assign n15082 = pi1539 & ~n11852;
  assign n15083 = ~n15081 & ~n15082;
  assign n15084 = pi1940 & ~n15083;
  assign po1590 = n15080 | n15084;
  assign n15086 = pi1540 & ~pi1940;
  assign n15087 = pi2196 & n11852;
  assign n15088 = pi1540 & ~n11852;
  assign n15089 = ~n15087 & ~n15088;
  assign n15090 = pi1940 & ~n15089;
  assign po1591 = n15086 | n15090;
  assign n15092 = pi1541 & ~pi1940;
  assign n15093 = pi2193 & n11852;
  assign n15094 = pi1541 & ~n11852;
  assign n15095 = ~n15093 & ~n15094;
  assign n15096 = pi1940 & ~n15095;
  assign po1592 = n15092 | n15096;
  assign n15098 = pi1542 & ~pi1940;
  assign n15099 = pi2189 & n11852;
  assign n15100 = pi1542 & ~n11852;
  assign n15101 = ~n15099 & ~n15100;
  assign n15102 = pi1940 & ~n15101;
  assign po1593 = n15098 | n15102;
  assign n15104 = pi1543 & ~pi1940;
  assign n15105 = pi2179 & n11852;
  assign n15106 = pi1543 & ~n11852;
  assign n15107 = ~n15105 & ~n15106;
  assign n15108 = pi1940 & ~n15107;
  assign po1594 = n15104 | n15108;
  assign n15110 = pi1544 & ~pi1940;
  assign n15111 = pi2198 & n11852;
  assign n15112 = pi1544 & ~n11852;
  assign n15113 = ~n15111 & ~n15112;
  assign n15114 = pi1940 & ~n15113;
  assign po1595 = n15110 | n15114;
  assign n15116 = pi1545 & ~pi1940;
  assign n15117 = pi2185 & n11852;
  assign n15118 = pi1545 & ~n11852;
  assign n15119 = ~n15117 & ~n15118;
  assign n15120 = pi1940 & ~n15119;
  assign po1596 = n15116 | n15120;
  assign n15122 = pi1546 & ~pi1940;
  assign n15123 = pi2176 & n11852;
  assign n15124 = pi1546 & ~n11852;
  assign n15125 = ~n15123 & ~n15124;
  assign n15126 = pi1940 & ~n15125;
  assign po1597 = n15122 | n15126;
  assign n15128 = pi1547 & ~pi1940;
  assign n15129 = pi2171 & n11852;
  assign n15130 = pi1547 & ~n11852;
  assign n15131 = ~n15129 & ~n15130;
  assign n15132 = pi1940 & ~n15131;
  assign po1598 = n15128 | n15132;
  assign n15134 = pi1548 & ~pi1940;
  assign n15135 = pi2169 & n11852;
  assign n15136 = pi1548 & ~n11852;
  assign n15137 = ~n15135 & ~n15136;
  assign n15138 = pi1940 & ~n15137;
  assign po1599 = n15134 | n15138;
  assign n15140 = pi1549 & ~pi1940;
  assign n15141 = pi2170 & n11852;
  assign n15142 = pi1549 & ~n11852;
  assign n15143 = ~n15141 & ~n15142;
  assign n15144 = pi1940 & ~n15143;
  assign po1600 = n15140 | n15144;
  assign n15146 = pi1550 & ~pi1940;
  assign n15147 = pi2181 & n11852;
  assign n15148 = pi1550 & ~n11852;
  assign n15149 = ~n15147 & ~n15148;
  assign n15150 = pi1940 & ~n15149;
  assign po1601 = n15146 | n15150;
  assign n15152 = pi1551 & ~pi1940;
  assign n15153 = pi2182 & n11852;
  assign n15154 = pi1551 & ~n11852;
  assign n15155 = ~n15153 & ~n15154;
  assign n15156 = pi1940 & ~n15155;
  assign po1602 = n15152 | n15156;
  assign n15158 = pi1552 & ~pi1940;
  assign n15159 = pi2191 & n11852;
  assign n15160 = pi1552 & ~n11852;
  assign n15161 = ~n15159 & ~n15160;
  assign n15162 = pi1940 & ~n15161;
  assign po1603 = n15158 | n15162;
  assign n15164 = pi1553 & ~pi1940;
  assign n15165 = pi2177 & n11852;
  assign n15166 = pi1553 & ~n11852;
  assign n15167 = ~n15165 & ~n15166;
  assign n15168 = pi1940 & ~n15167;
  assign po1604 = n15164 | n15168;
  assign n15170 = pi1554 & ~pi1940;
  assign n15171 = pi2173 & n11852;
  assign n15172 = pi1554 & ~n11852;
  assign n15173 = ~n15171 & ~n15172;
  assign n15174 = pi1940 & ~n15173;
  assign po1605 = n15170 | n15174;
  assign n15176 = pi1555 & ~pi1940;
  assign n15177 = pi2167 & n11852;
  assign n15178 = pi1555 & ~n11852;
  assign n15179 = ~n15177 & ~n15178;
  assign n15180 = pi1940 & ~n15179;
  assign po1606 = n15176 | n15180;
  assign n15182 = pi1556 & ~pi1940;
  assign n15183 = pi2188 & n11852;
  assign n15184 = pi1556 & ~n11852;
  assign n15185 = ~n15183 & ~n15184;
  assign n15186 = pi1940 & ~n15185;
  assign po1607 = n15182 | n15186;
  assign n15188 = pi1557 & ~pi1940;
  assign n15189 = pi2184 & n11852;
  assign n15190 = pi1557 & ~n11852;
  assign n15191 = ~n15189 & ~n15190;
  assign n15192 = pi1940 & ~n15191;
  assign po1608 = n15188 | n15192;
  assign n15194 = pi1558 & ~pi1940;
  assign n15195 = pi2195 & n11852;
  assign n15196 = pi1558 & ~n11852;
  assign n15197 = ~n15195 & ~n15196;
  assign n15198 = pi1940 & ~n15197;
  assign po1609 = n15194 | n15198;
  assign n15200 = pi1559 & ~pi1940;
  assign n15201 = pi2192 & n11852;
  assign n15202 = pi1559 & ~n11852;
  assign n15203 = ~n15201 & ~n15202;
  assign n15204 = pi1940 & ~n15203;
  assign po1610 = n15200 | n15204;
  assign n15206 = pi1560 & ~pi1940;
  assign n15207 = pi2186 & n11853;
  assign n15208 = pi1560 & ~n11853;
  assign n15209 = ~n15207 & ~n15208;
  assign n15210 = pi1940 & ~n15209;
  assign po1611 = n15206 | n15210;
  assign n15212 = pi1561 & ~pi1940;
  assign n15213 = pi2172 & n11853;
  assign n15214 = pi1561 & ~n11853;
  assign n15215 = ~n15213 & ~n15214;
  assign n15216 = pi1940 & ~n15215;
  assign po1612 = n15212 | n15216;
  assign n15218 = pi1562 & ~pi1940;
  assign n15219 = pi2168 & n11853;
  assign n15220 = pi1562 & ~n11853;
  assign n15221 = ~n15219 & ~n15220;
  assign n15222 = pi1940 & ~n15221;
  assign po1613 = n15218 | n15222;
  assign n15224 = pi1563 & ~pi1940;
  assign n15225 = pi2174 & n11853;
  assign n15226 = pi1563 & ~n11853;
  assign n15227 = ~n15225 & ~n15226;
  assign n15228 = pi1940 & ~n15227;
  assign po1614 = n15224 | n15228;
  assign n15230 = pi1564 & ~pi1940;
  assign n15231 = pi2178 & n11853;
  assign n15232 = pi1564 & ~n11853;
  assign n15233 = ~n15231 & ~n15232;
  assign n15234 = pi1940 & ~n15233;
  assign po1615 = n15230 | n15234;
  assign n15236 = pi1565 & ~pi1940;
  assign n15237 = pi2196 & n11853;
  assign n15238 = pi1565 & ~n11853;
  assign n15239 = ~n15237 & ~n15238;
  assign n15240 = pi1940 & ~n15239;
  assign po1616 = n15236 | n15240;
  assign n15242 = pi1566 & ~pi1940;
  assign n15243 = pi2193 & n11853;
  assign n15244 = pi1566 & ~n11853;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = pi1940 & ~n15245;
  assign po1617 = n15242 | n15246;
  assign n15248 = pi1567 & ~pi1940;
  assign n15249 = pi2179 & n11853;
  assign n15250 = pi1567 & ~n11853;
  assign n15251 = ~n15249 & ~n15250;
  assign n15252 = pi1940 & ~n15251;
  assign po1618 = n15248 | n15252;
  assign n15254 = pi1568 & ~pi1940;
  assign n15255 = pi2198 & n11853;
  assign n15256 = pi1568 & ~n11853;
  assign n15257 = ~n15255 & ~n15256;
  assign n15258 = pi1940 & ~n15257;
  assign po1619 = n15254 | n15258;
  assign n15260 = pi1569 & ~pi1940;
  assign n15261 = pi2185 & n11853;
  assign n15262 = pi1569 & ~n11853;
  assign n15263 = ~n15261 & ~n15262;
  assign n15264 = pi1940 & ~n15263;
  assign po1620 = n15260 | n15264;
  assign n15266 = pi1570 & ~pi1940;
  assign n15267 = pi2176 & n11853;
  assign n15268 = pi1570 & ~n11853;
  assign n15269 = ~n15267 & ~n15268;
  assign n15270 = pi1940 & ~n15269;
  assign po1621 = n15266 | n15270;
  assign n15272 = pi1571 & ~pi1940;
  assign n15273 = pi2171 & n11853;
  assign n15274 = pi1571 & ~n11853;
  assign n15275 = ~n15273 & ~n15274;
  assign n15276 = pi1940 & ~n15275;
  assign po1622 = n15272 | n15276;
  assign n15278 = pi1572 & ~pi1940;
  assign n15279 = pi2169 & n11853;
  assign n15280 = pi1572 & ~n11853;
  assign n15281 = ~n15279 & ~n15280;
  assign n15282 = pi1940 & ~n15281;
  assign po1623 = n15278 | n15282;
  assign n15284 = pi1573 & ~pi1940;
  assign n15285 = pi2170 & n11853;
  assign n15286 = pi1573 & ~n11853;
  assign n15287 = ~n15285 & ~n15286;
  assign n15288 = pi1940 & ~n15287;
  assign po1624 = n15284 | n15288;
  assign n15290 = pi1574 & ~pi1940;
  assign n15291 = pi2181 & n11853;
  assign n15292 = pi1574 & ~n11853;
  assign n15293 = ~n15291 & ~n15292;
  assign n15294 = pi1940 & ~n15293;
  assign po1625 = n15290 | n15294;
  assign n15296 = pi1575 & ~pi1940;
  assign n15297 = pi2182 & n11853;
  assign n15298 = pi1575 & ~n11853;
  assign n15299 = ~n15297 & ~n15298;
  assign n15300 = pi1940 & ~n15299;
  assign po1626 = n15296 | n15300;
  assign n15302 = pi1576 & ~pi1940;
  assign n15303 = pi2191 & n11853;
  assign n15304 = pi1576 & ~n11853;
  assign n15305 = ~n15303 & ~n15304;
  assign n15306 = pi1940 & ~n15305;
  assign po1627 = n15302 | n15306;
  assign n15308 = pi1577 & ~pi1940;
  assign n15309 = pi2177 & n11853;
  assign n15310 = pi1577 & ~n11853;
  assign n15311 = ~n15309 & ~n15310;
  assign n15312 = pi1940 & ~n15311;
  assign po1628 = n15308 | n15312;
  assign n15314 = pi1578 & ~pi1940;
  assign n15315 = pi2173 & n11853;
  assign n15316 = pi1578 & ~n11853;
  assign n15317 = ~n15315 & ~n15316;
  assign n15318 = pi1940 & ~n15317;
  assign po1629 = n15314 | n15318;
  assign n15320 = pi1579 & ~pi1940;
  assign n15321 = pi2167 & n11853;
  assign n15322 = pi1579 & ~n11853;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = pi1940 & ~n15323;
  assign po1630 = n15320 | n15324;
  assign n15326 = pi1580 & ~pi1940;
  assign n15327 = pi2188 & n11853;
  assign n15328 = pi1580 & ~n11853;
  assign n15329 = ~n15327 & ~n15328;
  assign n15330 = pi1940 & ~n15329;
  assign po1631 = n15326 | n15330;
  assign n15332 = pi1581 & ~pi1940;
  assign n15333 = pi2184 & n11853;
  assign n15334 = pi1581 & ~n11853;
  assign n15335 = ~n15333 & ~n15334;
  assign n15336 = pi1940 & ~n15335;
  assign po1632 = n15332 | n15336;
  assign n15338 = pi1582 & ~pi1940;
  assign n15339 = pi2195 & n11853;
  assign n15340 = pi1582 & ~n11853;
  assign n15341 = ~n15339 & ~n15340;
  assign n15342 = pi1940 & ~n15341;
  assign po1633 = n15338 | n15342;
  assign n15344 = pi1583 & ~pi1940;
  assign n15345 = pi2192 & n11853;
  assign n15346 = pi1583 & ~n11853;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = pi1940 & ~n15347;
  assign po1634 = n15344 | n15348;
  assign n15350 = pi1584 & ~pi1940;
  assign n15351 = pi2186 & n11794;
  assign n15352 = pi1584 & ~n11794;
  assign n15353 = ~n15351 & ~n15352;
  assign n15354 = pi1940 & ~n15353;
  assign po1635 = n15350 | n15354;
  assign n15356 = pi1585 & ~pi1940;
  assign n15357 = pi2172 & n11794;
  assign n15358 = pi1585 & ~n11794;
  assign n15359 = ~n15357 & ~n15358;
  assign n15360 = pi1940 & ~n15359;
  assign po1636 = n15356 | n15360;
  assign n15362 = pi1586 & ~pi1940;
  assign n15363 = pi2168 & n11794;
  assign n15364 = pi1586 & ~n11794;
  assign n15365 = ~n15363 & ~n15364;
  assign n15366 = pi1940 & ~n15365;
  assign po1637 = n15362 | n15366;
  assign n15368 = pi1587 & ~pi1940;
  assign n15369 = pi2174 & n11794;
  assign n15370 = pi1587 & ~n11794;
  assign n15371 = ~n15369 & ~n15370;
  assign n15372 = pi1940 & ~n15371;
  assign po1638 = n15368 | n15372;
  assign n15374 = pi1588 & ~pi1940;
  assign n15375 = pi2178 & n11794;
  assign n15376 = pi1588 & ~n11794;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = pi1940 & ~n15377;
  assign po1639 = n15374 | n15378;
  assign n15380 = pi1589 & ~pi1940;
  assign n15381 = pi2196 & n11794;
  assign n15382 = pi1589 & ~n11794;
  assign n15383 = ~n15381 & ~n15382;
  assign n15384 = pi1940 & ~n15383;
  assign po1640 = n15380 | n15384;
  assign n15386 = pi1590 & ~pi1940;
  assign n15387 = pi2193 & n11794;
  assign n15388 = pi1590 & ~n11794;
  assign n15389 = ~n15387 & ~n15388;
  assign n15390 = pi1940 & ~n15389;
  assign po1641 = n15386 | n15390;
  assign n15392 = pi1591 & ~pi1940;
  assign n15393 = pi2179 & n11794;
  assign n15394 = pi1591 & ~n11794;
  assign n15395 = ~n15393 & ~n15394;
  assign n15396 = pi1940 & ~n15395;
  assign po1642 = n15392 | n15396;
  assign n15398 = pi1592 & ~pi1940;
  assign n15399 = pi2198 & n11794;
  assign n15400 = pi1592 & ~n11794;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = pi1940 & ~n15401;
  assign po1643 = n15398 | n15402;
  assign n15404 = pi1593 & ~pi1940;
  assign n15405 = pi2185 & n11794;
  assign n15406 = pi1593 & ~n11794;
  assign n15407 = ~n15405 & ~n15406;
  assign n15408 = pi1940 & ~n15407;
  assign po1644 = n15404 | n15408;
  assign n15410 = pi1594 & ~pi1936;
  assign n15411 = pi1594 & ~n12004;
  assign n15412 = pi2185 & n12004;
  assign n15413 = ~n15411 & ~n15412;
  assign n15414 = pi1936 & ~n15413;
  assign po1645 = n15410 | n15414;
  assign n15416 = pi1595 & ~pi1940;
  assign n15417 = pi2176 & n11794;
  assign n15418 = pi1595 & ~n11794;
  assign n15419 = ~n15417 & ~n15418;
  assign n15420 = pi1940 & ~n15419;
  assign po1646 = n15416 | n15420;
  assign n15422 = pi1596 & ~pi1940;
  assign n15423 = pi2171 & n11794;
  assign n15424 = pi1596 & ~n11794;
  assign n15425 = ~n15423 & ~n15424;
  assign n15426 = pi1940 & ~n15425;
  assign po1647 = n15422 | n15426;
  assign n15428 = pi1597 & ~pi1940;
  assign n15429 = pi2169 & n11794;
  assign n15430 = pi1597 & ~n11794;
  assign n15431 = ~n15429 & ~n15430;
  assign n15432 = pi1940 & ~n15431;
  assign po1648 = n15428 | n15432;
  assign n15434 = pi1598 & ~pi1940;
  assign n15435 = pi2170 & n11794;
  assign n15436 = pi1598 & ~n11794;
  assign n15437 = ~n15435 & ~n15436;
  assign n15438 = pi1940 & ~n15437;
  assign po1649 = n15434 | n15438;
  assign n15440 = pi1599 & ~pi1940;
  assign n15441 = pi2181 & n11794;
  assign n15442 = pi1599 & ~n11794;
  assign n15443 = ~n15441 & ~n15442;
  assign n15444 = pi1940 & ~n15443;
  assign po1650 = n15440 | n15444;
  assign n15446 = pi1600 & ~pi1940;
  assign n15447 = pi2182 & n11794;
  assign n15448 = pi1600 & ~n11794;
  assign n15449 = ~n15447 & ~n15448;
  assign n15450 = pi1940 & ~n15449;
  assign po1651 = n15446 | n15450;
  assign n15452 = pi1601 & ~pi1940;
  assign n15453 = pi2191 & n11794;
  assign n15454 = pi1601 & ~n11794;
  assign n15455 = ~n15453 & ~n15454;
  assign n15456 = pi1940 & ~n15455;
  assign po1652 = n15452 | n15456;
  assign n15458 = pi1602 & ~pi1940;
  assign n15459 = pi2177 & n11794;
  assign n15460 = pi1602 & ~n11794;
  assign n15461 = ~n15459 & ~n15460;
  assign n15462 = pi1940 & ~n15461;
  assign po1653 = n15458 | n15462;
  assign n15464 = pi1603 & ~pi1940;
  assign n15465 = pi2173 & n11794;
  assign n15466 = pi1603 & ~n11794;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = pi1940 & ~n15467;
  assign po1654 = n15464 | n15468;
  assign n15470 = pi1604 & ~pi1940;
  assign n15471 = pi2167 & n11794;
  assign n15472 = pi1604 & ~n11794;
  assign n15473 = ~n15471 & ~n15472;
  assign n15474 = pi1940 & ~n15473;
  assign po1655 = n15470 | n15474;
  assign n15476 = pi1605 & ~pi1940;
  assign n15477 = pi2188 & n11794;
  assign n15478 = pi1605 & ~n11794;
  assign n15479 = ~n15477 & ~n15478;
  assign n15480 = pi1940 & ~n15479;
  assign po1656 = n15476 | n15480;
  assign n15482 = pi1606 & ~pi1940;
  assign n15483 = pi2184 & n11794;
  assign n15484 = pi1606 & ~n11794;
  assign n15485 = ~n15483 & ~n15484;
  assign n15486 = pi1940 & ~n15485;
  assign po1657 = n15482 | n15486;
  assign n15488 = pi1607 & ~pi1940;
  assign n15489 = pi2195 & n11794;
  assign n15490 = pi1607 & ~n11794;
  assign n15491 = ~n15489 & ~n15490;
  assign n15492 = pi1940 & ~n15491;
  assign po1658 = n15488 | n15492;
  assign n15494 = pi1608 & ~pi1940;
  assign n15495 = pi2192 & n11794;
  assign n15496 = pi1608 & ~n11794;
  assign n15497 = ~n15495 & ~n15496;
  assign n15498 = pi1940 & ~n15497;
  assign po1659 = n15494 | n15498;
  assign n15500 = pi1609 & ~pi1941;
  assign n15501 = pi2186 & n11820;
  assign n15502 = pi1609 & ~n11820;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = pi1941 & ~n15503;
  assign po1660 = n15500 | n15504;
  assign n15506 = pi1610 & ~pi1941;
  assign n15507 = pi2172 & n11820;
  assign n15508 = pi1610 & ~n11820;
  assign n15509 = ~n15507 & ~n15508;
  assign n15510 = pi1941 & ~n15509;
  assign po1661 = n15506 | n15510;
  assign n15512 = pi1611 & ~pi1941;
  assign n15513 = pi2168 & n11820;
  assign n15514 = pi1611 & ~n11820;
  assign n15515 = ~n15513 & ~n15514;
  assign n15516 = pi1941 & ~n15515;
  assign po1662 = n15512 | n15516;
  assign n15518 = pi1612 & ~pi1941;
  assign n15519 = pi2174 & n11820;
  assign n15520 = pi1612 & ~n11820;
  assign n15521 = ~n15519 & ~n15520;
  assign n15522 = pi1941 & ~n15521;
  assign po1663 = n15518 | n15522;
  assign n15524 = pi1613 & ~pi1941;
  assign n15525 = pi2178 & n11820;
  assign n15526 = pi1613 & ~n11820;
  assign n15527 = ~n15525 & ~n15526;
  assign n15528 = pi1941 & ~n15527;
  assign po1664 = n15524 | n15528;
  assign n15530 = pi1614 & ~pi1941;
  assign n15531 = pi2196 & n11820;
  assign n15532 = pi1614 & ~n11820;
  assign n15533 = ~n15531 & ~n15532;
  assign n15534 = pi1941 & ~n15533;
  assign po1665 = n15530 | n15534;
  assign n15536 = pi1615 & ~pi1941;
  assign n15537 = pi2193 & n11820;
  assign n15538 = pi1615 & ~n11820;
  assign n15539 = ~n15537 & ~n15538;
  assign n15540 = pi1941 & ~n15539;
  assign po1666 = n15536 | n15540;
  assign n15542 = pi1616 & ~pi1941;
  assign n15543 = pi2179 & n11820;
  assign n15544 = pi1616 & ~n11820;
  assign n15545 = ~n15543 & ~n15544;
  assign n15546 = pi1941 & ~n15545;
  assign po1667 = n15542 | n15546;
  assign n15548 = pi1617 & ~pi1941;
  assign n15549 = pi2198 & n11820;
  assign n15550 = pi1617 & ~n11820;
  assign n15551 = ~n15549 & ~n15550;
  assign n15552 = pi1941 & ~n15551;
  assign po1668 = n15548 | n15552;
  assign n15554 = pi1618 & ~pi1941;
  assign n15555 = pi2185 & n11820;
  assign n15556 = pi1618 & ~n11820;
  assign n15557 = ~n15555 & ~n15556;
  assign n15558 = pi1941 & ~n15557;
  assign po1669 = n15554 | n15558;
  assign n15560 = pi1619 & ~pi1941;
  assign n15561 = pi2176 & n11820;
  assign n15562 = pi1619 & ~n11820;
  assign n15563 = ~n15561 & ~n15562;
  assign n15564 = pi1941 & ~n15563;
  assign po1670 = n15560 | n15564;
  assign n15566 = pi1620 & ~pi1941;
  assign n15567 = pi2171 & n11820;
  assign n15568 = pi1620 & ~n11820;
  assign n15569 = ~n15567 & ~n15568;
  assign n15570 = pi1941 & ~n15569;
  assign po1671 = n15566 | n15570;
  assign n15572 = pi1621 & ~pi1941;
  assign n15573 = pi2169 & n11820;
  assign n15574 = pi1621 & ~n11820;
  assign n15575 = ~n15573 & ~n15574;
  assign n15576 = pi1941 & ~n15575;
  assign po1672 = n15572 | n15576;
  assign n15578 = pi1622 & ~pi1941;
  assign n15579 = pi2170 & n11820;
  assign n15580 = pi1622 & ~n11820;
  assign n15581 = ~n15579 & ~n15580;
  assign n15582 = pi1941 & ~n15581;
  assign po1673 = n15578 | n15582;
  assign n15584 = pi1623 & ~pi1937;
  assign n15585 = pi2186 & n11828;
  assign n15586 = pi1623 & ~n11828;
  assign n15587 = ~n15585 & ~n15586;
  assign n15588 = pi1937 & ~n15587;
  assign po1674 = n15584 | n15588;
  assign n15590 = pi1624 & ~pi1941;
  assign n15591 = pi2181 & n11820;
  assign n15592 = pi1624 & ~n11820;
  assign n15593 = ~n15591 & ~n15592;
  assign n15594 = pi1941 & ~n15593;
  assign po1675 = n15590 | n15594;
  assign n15596 = pi1625 & ~pi1937;
  assign n15597 = pi2183 & n11828;
  assign n15598 = pi1625 & ~n11828;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = pi1937 & ~n15599;
  assign po1676 = n15596 | n15600;
  assign n15602 = pi1626 & ~pi1941;
  assign n15603 = pi2175 & n11820;
  assign n15604 = pi1626 & ~n11820;
  assign n15605 = ~n15603 & ~n15604;
  assign n15606 = pi1941 & ~n15605;
  assign po1677 = n15602 | n15606;
  assign n15608 = pi1627 & ~pi1941;
  assign n15609 = pi2191 & n11820;
  assign n15610 = pi1627 & ~n11820;
  assign n15611 = ~n15609 & ~n15610;
  assign n15612 = pi1941 & ~n15611;
  assign po1678 = n15608 | n15612;
  assign n15614 = pi1628 & ~pi1941;
  assign n15615 = pi2177 & n11820;
  assign n15616 = pi1628 & ~n11820;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = pi1941 & ~n15617;
  assign po1679 = n15614 | n15618;
  assign n15620 = pi1629 & ~pi1941;
  assign n15621 = pi2173 & n11820;
  assign n15622 = pi1629 & ~n11820;
  assign n15623 = ~n15621 & ~n15622;
  assign n15624 = pi1941 & ~n15623;
  assign po1680 = n15620 | n15624;
  assign n15626 = pi1630 & ~pi1937;
  assign n15627 = pi2168 & n11828;
  assign n15628 = pi1630 & ~n11828;
  assign n15629 = ~n15627 & ~n15628;
  assign n15630 = pi1937 & ~n15629;
  assign po1681 = n15626 | n15630;
  assign n15632 = pi1631 & ~pi1941;
  assign n15633 = pi2167 & n11820;
  assign n15634 = pi1631 & ~n11820;
  assign n15635 = ~n15633 & ~n15634;
  assign n15636 = pi1941 & ~n15635;
  assign po1682 = n15632 | n15636;
  assign n15638 = pi1632 & ~pi1937;
  assign n15639 = pi2174 & n11828;
  assign n15640 = pi1632 & ~n11828;
  assign n15641 = ~n15639 & ~n15640;
  assign n15642 = pi1937 & ~n15641;
  assign po1683 = n15638 | n15642;
  assign n15644 = pi1633 & ~pi1941;
  assign n15645 = pi2188 & n11820;
  assign n15646 = pi1633 & ~n11820;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = pi1941 & ~n15647;
  assign po1684 = n15644 | n15648;
  assign n15650 = pi1634 & ~pi1937;
  assign n15651 = pi2197 & n11828;
  assign n15652 = pi1634 & ~n11828;
  assign n15653 = ~n15651 & ~n15652;
  assign n15654 = pi1937 & ~n15653;
  assign po1685 = n15650 | n15654;
  assign n15656 = pi1635 & ~pi1941;
  assign n15657 = pi2166 & n11820;
  assign n15658 = pi1635 & ~n11820;
  assign n15659 = ~n15657 & ~n15658;
  assign n15660 = pi1941 & ~n15659;
  assign po1686 = n15656 | n15660;
  assign n15662 = pi1636 & ~pi1941;
  assign n15663 = pi2195 & n11820;
  assign n15664 = pi1636 & ~n11820;
  assign n15665 = ~n15663 & ~n15664;
  assign n15666 = pi1941 & ~n15665;
  assign po1687 = n15662 | n15666;
  assign n15668 = pi1637 & ~pi1941;
  assign n15669 = pi2192 & n11820;
  assign n15670 = pi1637 & ~n11820;
  assign n15671 = ~n15669 & ~n15670;
  assign n15672 = pi1941 & ~n15671;
  assign po1688 = n15668 | n15672;
  assign n15674 = pi1638 & ~pi1941;
  assign n15675 = pi2186 & n11821;
  assign n15676 = pi1638 & ~n11821;
  assign n15677 = ~n15675 & ~n15676;
  assign n15678 = pi1941 & ~n15677;
  assign po1689 = n15674 | n15678;
  assign n15680 = pi1639 & ~pi1937;
  assign n15681 = pi2196 & n11828;
  assign n15682 = pi1639 & ~n11828;
  assign n15683 = ~n15681 & ~n15682;
  assign n15684 = pi1937 & ~n15683;
  assign po1690 = n15680 | n15684;
  assign n15686 = pi1640 & ~pi1941;
  assign n15687 = pi2183 & n11821;
  assign n15688 = pi1640 & ~n11821;
  assign n15689 = ~n15687 & ~n15688;
  assign n15690 = pi1941 & ~n15689;
  assign po1691 = n15686 | n15690;
  assign n15692 = pi1641 & ~pi1941;
  assign n15693 = pi2172 & n11821;
  assign n15694 = pi1641 & ~n11821;
  assign n15695 = ~n15693 & ~n15694;
  assign n15696 = pi1941 & ~n15695;
  assign po1692 = n15692 | n15696;
  assign n15698 = pi1642 & ~pi1937;
  assign n15699 = pi2193 & n11828;
  assign n15700 = pi1642 & ~n11828;
  assign n15701 = ~n15699 & ~n15700;
  assign n15702 = pi1937 & ~n15701;
  assign po1693 = n15698 | n15702;
  assign n15704 = pi1643 & ~pi1941;
  assign n15705 = pi2168 & n11821;
  assign n15706 = pi1643 & ~n11821;
  assign n15707 = ~n15705 & ~n15706;
  assign n15708 = pi1941 & ~n15707;
  assign po1694 = n15704 | n15708;
  assign n15710 = pi1644 & ~pi1937;
  assign n15711 = pi2189 & n11828;
  assign n15712 = pi1644 & ~n11828;
  assign n15713 = ~n15711 & ~n15712;
  assign n15714 = pi1937 & ~n15713;
  assign po1695 = n15710 | n15714;
  assign n15716 = pi1645 & ~pi1941;
  assign n15717 = pi2197 & n11821;
  assign n15718 = pi1645 & ~n11821;
  assign n15719 = ~n15717 & ~n15718;
  assign n15720 = pi1941 & ~n15719;
  assign po1696 = n15716 | n15720;
  assign n15722 = pi1646 & ~pi1941;
  assign n15723 = pi2178 & n11821;
  assign n15724 = pi1646 & ~n11821;
  assign n15725 = ~n15723 & ~n15724;
  assign n15726 = pi1941 & ~n15725;
  assign po1697 = n15722 | n15726;
  assign n15728 = pi1647 & ~pi1941;
  assign n15729 = pi2196 & n11821;
  assign n15730 = pi1647 & ~n11821;
  assign n15731 = ~n15729 & ~n15730;
  assign n15732 = pi1941 & ~n15731;
  assign po1698 = n15728 | n15732;
  assign n15734 = pi1648 & ~pi1941;
  assign n15735 = pi2193 & n11821;
  assign n15736 = pi1648 & ~n11821;
  assign n15737 = ~n15735 & ~n15736;
  assign n15738 = pi1941 & ~n15737;
  assign po1699 = n15734 | n15738;
  assign n15740 = pi1649 & ~pi1937;
  assign n15741 = pi2198 & n11828;
  assign n15742 = pi1649 & ~n11828;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = pi1937 & ~n15743;
  assign po1700 = n15740 | n15744;
  assign n15746 = pi1650 & ~pi1941;
  assign n15747 = pi2179 & n11821;
  assign n15748 = pi1650 & ~n11821;
  assign n15749 = ~n15747 & ~n15748;
  assign n15750 = pi1941 & ~n15749;
  assign po1701 = n15746 | n15750;
  assign n15752 = pi1651 & ~pi1937;
  assign n15753 = pi2185 & n11828;
  assign n15754 = pi1651 & ~n11828;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = pi1937 & ~n15755;
  assign po1702 = n15752 | n15756;
  assign n15758 = pi1652 & ~pi1941;
  assign n15759 = pi2198 & n11821;
  assign n15760 = pi1652 & ~n11821;
  assign n15761 = ~n15759 & ~n15760;
  assign n15762 = pi1941 & ~n15761;
  assign po1703 = n15758 | n15762;
  assign n15764 = pi1653 & ~pi1937;
  assign n15765 = pi2187 & n11828;
  assign n15766 = pi1653 & ~n11828;
  assign n15767 = ~n15765 & ~n15766;
  assign n15768 = pi1937 & ~n15767;
  assign po1704 = n15764 | n15768;
  assign n15770 = pi1654 & ~pi1941;
  assign n15771 = pi2187 & n11821;
  assign n15772 = pi1654 & ~n11821;
  assign n15773 = ~n15771 & ~n15772;
  assign n15774 = pi1941 & ~n15773;
  assign po1705 = n15770 | n15774;
  assign n15776 = pi1655 & ~pi1941;
  assign n15777 = pi2176 & n11821;
  assign n15778 = pi1655 & ~n11821;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = pi1941 & ~n15779;
  assign po1706 = n15776 | n15780;
  assign n15782 = pi1656 & ~pi1941;
  assign n15783 = pi2171 & n11821;
  assign n15784 = pi1656 & ~n11821;
  assign n15785 = ~n15783 & ~n15784;
  assign n15786 = pi1941 & ~n15785;
  assign po1707 = n15782 | n15786;
  assign n15788 = pi1657 & ~pi1941;
  assign n15789 = pi2169 & n11821;
  assign n15790 = pi1657 & ~n11821;
  assign n15791 = ~n15789 & ~n15790;
  assign n15792 = pi1941 & ~n15791;
  assign po1708 = n15788 | n15792;
  assign n15794 = pi1658 & ~pi1937;
  assign n15795 = pi2171 & n11828;
  assign n15796 = pi1658 & ~n11828;
  assign n15797 = ~n15795 & ~n15796;
  assign n15798 = pi1937 & ~n15797;
  assign po1709 = n15794 | n15798;
  assign n15800 = pi1659 & ~pi1941;
  assign n15801 = pi2170 & n11821;
  assign n15802 = pi1659 & ~n11821;
  assign n15803 = ~n15801 & ~n15802;
  assign n15804 = pi1941 & ~n15803;
  assign po1710 = n15800 | n15804;
  assign n15806 = pi1660 & ~pi1937;
  assign n15807 = pi2169 & n11828;
  assign n15808 = pi1660 & ~n11828;
  assign n15809 = ~n15807 & ~n15808;
  assign n15810 = pi1937 & ~n15809;
  assign po1711 = n15806 | n15810;
  assign n15812 = pi1661 & ~pi1941;
  assign n15813 = pi2181 & n11821;
  assign n15814 = pi1661 & ~n11821;
  assign n15815 = ~n15813 & ~n15814;
  assign n15816 = pi1941 & ~n15815;
  assign po1712 = n15812 | n15816;
  assign n15818 = pi1662 & ~pi1937;
  assign n15819 = pi2190 & n11828;
  assign n15820 = pi1662 & ~n11828;
  assign n15821 = ~n15819 & ~n15820;
  assign n15822 = pi1937 & ~n15821;
  assign po1713 = n15818 | n15822;
  assign n15824 = pi1663 & ~pi1941;
  assign n15825 = pi2175 & n11821;
  assign n15826 = pi1663 & ~n11821;
  assign n15827 = ~n15825 & ~n15826;
  assign n15828 = pi1941 & ~n15827;
  assign po1714 = n15824 | n15828;
  assign n15830 = pi1664 & ~pi1941;
  assign n15831 = pi2191 & n11821;
  assign n15832 = pi1664 & ~n11821;
  assign n15833 = ~n15831 & ~n15832;
  assign n15834 = pi1941 & ~n15833;
  assign po1715 = n15830 | n15834;
  assign n15836 = pi1665 & ~pi1941;
  assign n15837 = pi2177 & n11821;
  assign n15838 = pi1665 & ~n11821;
  assign n15839 = ~n15837 & ~n15838;
  assign n15840 = pi1941 & ~n15839;
  assign po1716 = n15836 | n15840;
  assign n15842 = pi1666 & ~pi1941;
  assign n15843 = pi2173 & n11821;
  assign n15844 = pi1666 & ~n11821;
  assign n15845 = ~n15843 & ~n15844;
  assign n15846 = pi1941 & ~n15845;
  assign po1717 = n15842 | n15846;
  assign n15848 = pi1667 & ~pi1937;
  assign n15849 = pi2181 & n11828;
  assign n15850 = pi1667 & ~n11828;
  assign n15851 = ~n15849 & ~n15850;
  assign n15852 = pi1937 & ~n15851;
  assign po1718 = n15848 | n15852;
  assign n15854 = pi1668 & ~pi1938;
  assign n15855 = pi1668 & ~n11882;
  assign n15856 = pi2186 & n11882;
  assign n15857 = ~n15855 & ~n15856;
  assign n15858 = pi1938 & ~n15857;
  assign po1719 = n15854 | n15858;
  assign n15860 = pi1669 & ~pi1938;
  assign n15861 = pi1669 & ~n11882;
  assign n15862 = pi2183 & n11882;
  assign n15863 = ~n15861 & ~n15862;
  assign n15864 = pi1938 & ~n15863;
  assign po1720 = n15860 | n15864;
  assign n15866 = pi1670 & ~pi1938;
  assign n15867 = pi1670 & ~n11882;
  assign n15868 = pi2172 & n11882;
  assign n15869 = ~n15867 & ~n15868;
  assign n15870 = pi1938 & ~n15869;
  assign po1721 = n15866 | n15870;
  assign n15872 = pi1671 & ~pi1938;
  assign n15873 = pi1671 & ~n11882;
  assign n15874 = pi2178 & n11882;
  assign n15875 = ~n15873 & ~n15874;
  assign n15876 = pi1938 & ~n15875;
  assign po1722 = n15872 | n15876;
  assign n15878 = pi1672 & ~pi1938;
  assign n15879 = pi1672 & ~n11882;
  assign n15880 = pi2189 & n11882;
  assign n15881 = ~n15879 & ~n15880;
  assign n15882 = pi1938 & ~n15881;
  assign po1723 = n15878 | n15882;
  assign n15884 = pi1673 & ~pi1938;
  assign n15885 = pi1673 & ~n11882;
  assign n15886 = pi2198 & n11882;
  assign n15887 = ~n15885 & ~n15886;
  assign n15888 = pi1938 & ~n15887;
  assign po1724 = n15884 | n15888;
  assign n15890 = pi1674 & ~pi1938;
  assign n15891 = pi1674 & ~n11882;
  assign n15892 = pi2187 & n11882;
  assign n15893 = ~n15891 & ~n15892;
  assign n15894 = pi1938 & ~n15893;
  assign po1725 = n15890 | n15894;
  assign n15896 = pi1675 & ~pi1938;
  assign n15897 = pi1675 & ~n11882;
  assign n15898 = pi2190 & n11882;
  assign n15899 = ~n15897 & ~n15898;
  assign n15900 = pi1938 & ~n15899;
  assign po1726 = n15896 | n15900;
  assign n15902 = pi1676 & ~pi1938;
  assign n15903 = pi1676 & ~n11882;
  assign n15904 = pi2181 & n11882;
  assign n15905 = ~n15903 & ~n15904;
  assign n15906 = pi1938 & ~n15905;
  assign po1727 = n15902 | n15906;
  assign n15908 = pi1677 & ~pi1938;
  assign n15909 = pi1677 & ~n11882;
  assign n15910 = pi2182 & n11882;
  assign n15911 = ~n15909 & ~n15910;
  assign n15912 = pi1938 & ~n15911;
  assign po1728 = n15908 | n15912;
  assign n15914 = pi1678 & ~pi1938;
  assign n15915 = pi1678 & ~n11882;
  assign n15916 = pi2170 & n11882;
  assign n15917 = ~n15915 & ~n15916;
  assign n15918 = pi1938 & ~n15917;
  assign po1729 = n15914 | n15918;
  assign n15920 = pi1679 & ~pi1938;
  assign n15921 = pi1679 & ~n11882;
  assign n15922 = pi2191 & n11882;
  assign n15923 = ~n15921 & ~n15922;
  assign n15924 = pi1938 & ~n15923;
  assign po1730 = n15920 | n15924;
  assign n15926 = pi1680 & ~pi1938;
  assign n15927 = pi1680 & ~n11882;
  assign n15928 = pi2175 & n11882;
  assign n15929 = ~n15927 & ~n15928;
  assign n15930 = pi1938 & ~n15929;
  assign po1731 = n15926 | n15930;
  assign n15932 = pi1681 & ~pi1938;
  assign n15933 = pi1681 & ~n11882;
  assign n15934 = pi2194 & n11882;
  assign n15935 = ~n15933 & ~n15934;
  assign n15936 = pi1938 & ~n15935;
  assign po1732 = n15932 | n15936;
  assign n15938 = pi1682 & ~pi1938;
  assign n15939 = pi1682 & ~n11882;
  assign n15940 = pi2188 & n11882;
  assign n15941 = ~n15939 & ~n15940;
  assign n15942 = pi1938 & ~n15941;
  assign po1733 = n15938 | n15942;
  assign n15944 = pi1683 & ~pi1938;
  assign n15945 = pi1683 & ~n11882;
  assign n15946 = pi2195 & n11882;
  assign n15947 = ~n15945 & ~n15946;
  assign n15948 = pi1938 & ~n15947;
  assign po1734 = n15944 | n15948;
  assign n15950 = pi1684 & ~pi1939;
  assign n15951 = pi1684 & ~n11943;
  assign n15952 = pi2183 & n11943;
  assign n15953 = ~n15951 & ~n15952;
  assign n15954 = pi1939 & ~n15953;
  assign po1735 = n15950 | n15954;
  assign n15956 = pi1685 & ~pi1939;
  assign n15957 = pi1685 & ~n11943;
  assign n15958 = pi2172 & n11943;
  assign n15959 = ~n15957 & ~n15958;
  assign n15960 = pi1939 & ~n15959;
  assign po1736 = n15956 | n15960;
  assign n15962 = pi1686 & ~pi1939;
  assign n15963 = pi1686 & ~n11943;
  assign n15964 = pi2178 & n11943;
  assign n15965 = ~n15963 & ~n15964;
  assign n15966 = pi1939 & ~n15965;
  assign po1737 = n15962 | n15966;
  assign n15968 = pi1687 & ~pi1939;
  assign n15969 = pi1687 & ~n11943;
  assign n15970 = pi2189 & n11943;
  assign n15971 = ~n15969 & ~n15970;
  assign n15972 = pi1939 & ~n15971;
  assign po1738 = n15968 | n15972;
  assign n15974 = pi1688 & ~pi1939;
  assign n15975 = pi1688 & ~n11943;
  assign n15976 = pi2198 & n11943;
  assign n15977 = ~n15975 & ~n15976;
  assign n15978 = pi1939 & ~n15977;
  assign po1739 = n15974 | n15978;
  assign n15980 = pi1689 & ~pi1939;
  assign n15981 = pi1689 & ~n11943;
  assign n15982 = pi2187 & n11943;
  assign n15983 = ~n15981 & ~n15982;
  assign n15984 = pi1939 & ~n15983;
  assign po1740 = n15980 | n15984;
  assign n15986 = pi1690 & ~n12907;
  assign n15987 = pi2195 & n12907;
  assign po1741 = n15986 | n15987;
  assign n15989 = pi1691 & ~pi1939;
  assign n15990 = pi1691 & ~n11943;
  assign n15991 = pi2170 & n11943;
  assign n15992 = ~n15990 & ~n15991;
  assign n15993 = pi1939 & ~n15992;
  assign po1742 = n15989 | n15993;
  assign n15995 = pi1692 & ~pi1939;
  assign n15996 = pi1692 & ~n11943;
  assign n15997 = pi2181 & n11943;
  assign n15998 = ~n15996 & ~n15997;
  assign n15999 = pi1939 & ~n15998;
  assign po1743 = n15995 | n15999;
  assign n16001 = pi1693 & ~pi1939;
  assign n16002 = pi1693 & ~n11943;
  assign n16003 = pi2190 & n11943;
  assign n16004 = ~n16002 & ~n16003;
  assign n16005 = pi1939 & ~n16004;
  assign po1744 = n16001 | n16005;
  assign n16007 = pi1694 & ~pi1939;
  assign n16008 = pi1694 & ~n11943;
  assign n16009 = pi2191 & n11943;
  assign n16010 = ~n16008 & ~n16009;
  assign n16011 = pi1939 & ~n16010;
  assign po1745 = n16007 | n16011;
  assign n16013 = pi1695 & ~pi1939;
  assign n16014 = pi1695 & ~n11943;
  assign n16015 = pi2175 & n11943;
  assign n16016 = ~n16014 & ~n16015;
  assign n16017 = pi1939 & ~n16016;
  assign po1746 = n16013 | n16017;
  assign n16019 = pi1696 & ~pi1939;
  assign n16020 = pi1696 & ~n11943;
  assign n16021 = pi2194 & n11943;
  assign n16022 = ~n16020 & ~n16021;
  assign n16023 = pi1939 & ~n16022;
  assign po1747 = n16019 | n16023;
  assign n16025 = pi1697 & ~pi1939;
  assign n16026 = pi1697 & ~n11943;
  assign n16027 = pi2188 & n11943;
  assign n16028 = ~n16026 & ~n16027;
  assign n16029 = pi1939 & ~n16028;
  assign po1748 = n16025 | n16029;
  assign n16031 = pi1698 & ~pi1939;
  assign n16032 = pi1698 & ~n11943;
  assign n16033 = pi2195 & n11943;
  assign n16034 = ~n16032 & ~n16033;
  assign n16035 = pi1939 & ~n16034;
  assign po1749 = n16031 | n16035;
  assign n16037 = pi1699 & ~pi1936;
  assign n16038 = pi1699 & ~n12004;
  assign n16039 = pi2183 & n12004;
  assign n16040 = ~n16038 & ~n16039;
  assign n16041 = pi1936 & ~n16040;
  assign po1750 = n16037 | n16041;
  assign n16043 = pi1700 & ~pi1936;
  assign n16044 = pi1700 & ~n12004;
  assign n16045 = pi2172 & n12004;
  assign n16046 = ~n16044 & ~n16045;
  assign n16047 = pi1936 & ~n16046;
  assign po1751 = n16043 | n16047;
  assign n16049 = pi1701 & ~pi1936;
  assign n16050 = pi1701 & ~n12004;
  assign n16051 = pi2178 & n12004;
  assign n16052 = ~n16050 & ~n16051;
  assign n16053 = pi1936 & ~n16052;
  assign po1752 = n16049 | n16053;
  assign n16055 = pi1702 & ~pi1940;
  assign n16056 = pi2187 & n11852;
  assign n16057 = pi1702 & ~n11852;
  assign n16058 = ~n16056 & ~n16057;
  assign n16059 = pi1940 & ~n16058;
  assign po1753 = n16055 | n16059;
  assign n16061 = pi1703 & ~pi1936;
  assign n16062 = pi1703 & ~n12004;
  assign n16063 = pi2189 & n12004;
  assign n16064 = ~n16062 & ~n16063;
  assign n16065 = pi1936 & ~n16064;
  assign po1754 = n16061 | n16065;
  assign n16067 = pi1704 & ~pi1936;
  assign n16068 = pi1704 & ~n12004;
  assign n16069 = pi2198 & n12004;
  assign n16070 = ~n16068 & ~n16069;
  assign n16071 = pi1936 & ~n16070;
  assign po1755 = n16067 | n16071;
  assign n16073 = pi1705 & ~pi1936;
  assign n16074 = pi1705 & ~n12004;
  assign n16075 = pi2187 & n12004;
  assign n16076 = ~n16074 & ~n16075;
  assign n16077 = pi1936 & ~n16076;
  assign po1756 = n16073 | n16077;
  assign n16079 = pi1706 & ~pi1936;
  assign n16080 = pi1706 & ~n12004;
  assign n16081 = pi2170 & n12004;
  assign n16082 = ~n16080 & ~n16081;
  assign n16083 = pi1936 & ~n16082;
  assign po1757 = n16079 | n16083;
  assign n16085 = pi1707 & ~pi1936;
  assign n16086 = pi1707 & ~n12004;
  assign n16087 = pi2181 & n12004;
  assign n16088 = ~n16086 & ~n16087;
  assign n16089 = pi1936 & ~n16088;
  assign po1758 = n16085 | n16089;
  assign n16091 = pi1708 & ~pi1936;
  assign n16092 = pi1708 & ~n12004;
  assign n16093 = pi2190 & n12004;
  assign n16094 = ~n16092 & ~n16093;
  assign n16095 = pi1936 & ~n16094;
  assign po1759 = n16091 | n16095;
  assign n16097 = pi1709 & ~pi1936;
  assign n16098 = pi1709 & ~n12004;
  assign n16099 = pi2191 & n12004;
  assign n16100 = ~n16098 & ~n16099;
  assign n16101 = pi1936 & ~n16100;
  assign po1760 = n16097 | n16101;
  assign n16103 = pi1710 & ~pi1936;
  assign n16104 = pi1710 & ~n12004;
  assign n16105 = pi2175 & n12004;
  assign n16106 = ~n16104 & ~n16105;
  assign n16107 = pi1936 & ~n16106;
  assign po1761 = n16103 | n16107;
  assign n16109 = pi1711 & ~pi1936;
  assign n16110 = pi1711 & ~n12004;
  assign n16111 = pi2194 & n12004;
  assign n16112 = ~n16110 & ~n16111;
  assign n16113 = pi1936 & ~n16112;
  assign po1762 = n16109 | n16113;
  assign n16115 = pi1712 & ~pi1936;
  assign n16116 = pi1712 & ~n12004;
  assign n16117 = pi2188 & n12004;
  assign n16118 = ~n16116 & ~n16117;
  assign n16119 = pi1936 & ~n16118;
  assign po1763 = n16115 | n16119;
  assign n16121 = pi1713 & ~pi1936;
  assign n16122 = pi1713 & ~n12004;
  assign n16123 = pi2195 & n12004;
  assign n16124 = ~n16122 & ~n16123;
  assign n16125 = pi1936 & ~n16124;
  assign po1764 = n16121 | n16125;
  assign n16127 = pi1714 & ~pi1940;
  assign n16128 = pi1714 & ~n12065;
  assign n16129 = pi2183 & n12065;
  assign n16130 = ~n16128 & ~n16129;
  assign n16131 = pi1940 & ~n16130;
  assign po1765 = n16127 | n16131;
  assign n16133 = pi1715 & ~pi1940;
  assign n16134 = pi1715 & ~n12065;
  assign n16135 = pi2172 & n12065;
  assign n16136 = ~n16134 & ~n16135;
  assign n16137 = pi1940 & ~n16136;
  assign po1766 = n16133 | n16137;
  assign n16139 = pi1716 & ~pi1940;
  assign n16140 = pi1716 & ~n12065;
  assign n16141 = pi2178 & n12065;
  assign n16142 = ~n16140 & ~n16141;
  assign n16143 = pi1940 & ~n16142;
  assign po1767 = n16139 | n16143;
  assign n16145 = pi1717 & ~pi1940;
  assign n16146 = pi1717 & ~n12065;
  assign n16147 = pi2189 & n12065;
  assign n16148 = ~n16146 & ~n16147;
  assign n16149 = pi1940 & ~n16148;
  assign po1768 = n16145 | n16149;
  assign n16151 = pi1718 & ~pi1940;
  assign n16152 = pi1718 & ~n12065;
  assign n16153 = pi2198 & n12065;
  assign n16154 = ~n16152 & ~n16153;
  assign n16155 = pi1940 & ~n16154;
  assign po1769 = n16151 | n16155;
  assign n16157 = pi1719 & ~pi1940;
  assign n16158 = pi1719 & ~n12065;
  assign n16159 = pi2187 & n12065;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = pi1940 & ~n16160;
  assign po1770 = n16157 | n16161;
  assign n16163 = pi1720 & ~pi1940;
  assign n16164 = pi1720 & ~n12065;
  assign n16165 = pi2190 & n12065;
  assign n16166 = ~n16164 & ~n16165;
  assign n16167 = pi1940 & ~n16166;
  assign po1771 = n16163 | n16167;
  assign n16169 = pi1721 & ~pi1940;
  assign n16170 = pi1721 & ~n12065;
  assign n16171 = pi2181 & n12065;
  assign n16172 = ~n16170 & ~n16171;
  assign n16173 = pi1940 & ~n16172;
  assign po1772 = n16169 | n16173;
  assign n16175 = pi1722 & ~pi1940;
  assign n16176 = pi1722 & ~n12065;
  assign n16177 = pi2182 & n12065;
  assign n16178 = ~n16176 & ~n16177;
  assign n16179 = pi1940 & ~n16178;
  assign po1773 = n16175 | n16179;
  assign n16181 = pi1723 & ~pi1940;
  assign n16182 = pi1723 & ~n12065;
  assign n16183 = pi2170 & n12065;
  assign n16184 = ~n16182 & ~n16183;
  assign n16185 = pi1940 & ~n16184;
  assign po1774 = n16181 | n16185;
  assign n16187 = pi1724 & ~pi1940;
  assign n16188 = pi1724 & ~n12065;
  assign n16189 = pi2191 & n12065;
  assign n16190 = ~n16188 & ~n16189;
  assign n16191 = pi1940 & ~n16190;
  assign po1775 = n16187 | n16191;
  assign n16193 = pi1725 & ~pi1940;
  assign n16194 = pi1725 & ~n12065;
  assign n16195 = pi2175 & n12065;
  assign n16196 = ~n16194 & ~n16195;
  assign n16197 = pi1940 & ~n16196;
  assign po1776 = n16193 | n16197;
  assign n16199 = pi1726 & ~pi1940;
  assign n16200 = pi1726 & ~n12065;
  assign n16201 = pi2194 & n12065;
  assign n16202 = ~n16200 & ~n16201;
  assign n16203 = pi1940 & ~n16202;
  assign po1777 = n16199 | n16203;
  assign n16205 = pi1727 & ~pi1940;
  assign n16206 = pi1727 & ~n12065;
  assign n16207 = pi2188 & n12065;
  assign n16208 = ~n16206 & ~n16207;
  assign n16209 = pi1940 & ~n16208;
  assign po1778 = n16205 | n16209;
  assign n16211 = pi1728 & ~pi1940;
  assign n16212 = pi1728 & ~n12065;
  assign n16213 = pi2195 & n12065;
  assign n16214 = ~n16212 & ~n16213;
  assign n16215 = pi1940 & ~n16214;
  assign po1779 = n16211 | n16215;
  assign n16217 = pi1729 & ~pi1937;
  assign n16218 = pi1729 & ~n12126;
  assign n16219 = pi2183 & n12126;
  assign n16220 = ~n16218 & ~n16219;
  assign n16221 = pi1937 & ~n16220;
  assign po1780 = n16217 | n16221;
  assign n16223 = pi1730 & ~pi1941;
  assign n16224 = pi1730 & ~n12145;
  assign n16225 = pi2183 & n12145;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = pi1941 & ~n16226;
  assign po1781 = n16223 | n16227;
  assign n16229 = pi1731 & ~pi1941;
  assign n16230 = pi1731 & ~n12145;
  assign n16231 = pi2174 & n12145;
  assign n16232 = ~n16230 & ~n16231;
  assign n16233 = pi1941 & ~n16232;
  assign po1782 = n16229 | n16233;
  assign n16235 = pi1732 & ~pi1937;
  assign n16236 = pi1732 & ~n12126;
  assign n16237 = pi2189 & n12126;
  assign n16238 = ~n16236 & ~n16237;
  assign n16239 = pi1937 & ~n16238;
  assign po1783 = n16235 | n16239;
  assign n16241 = pi1733 & ~pi1941;
  assign n16242 = pi1733 & ~n12145;
  assign n16243 = pi2197 & n12145;
  assign n16244 = ~n16242 & ~n16243;
  assign n16245 = pi1941 & ~n16244;
  assign po1784 = n16241 | n16245;
  assign n16247 = pi1734 & ~pi1937;
  assign n16248 = pi1734 & ~n12126;
  assign n16249 = pi2179 & n12126;
  assign n16250 = ~n16248 & ~n16249;
  assign n16251 = pi1937 & ~n16250;
  assign po1785 = n16247 | n16251;
  assign n16253 = pi1735 & ~pi1941;
  assign n16254 = pi1735 & ~n12145;
  assign n16255 = pi2189 & n12145;
  assign n16256 = ~n16254 & ~n16255;
  assign n16257 = pi1941 & ~n16256;
  assign po1786 = n16253 | n16257;
  assign n16259 = pi1736 & ~pi1941;
  assign n16260 = pi1736 & ~n12145;
  assign n16261 = pi2179 & n12145;
  assign n16262 = ~n16260 & ~n16261;
  assign n16263 = pi1941 & ~n16262;
  assign po1787 = n16259 | n16263;
  assign n16265 = pi1737 & ~pi1937;
  assign n16266 = pi1737 & ~n12126;
  assign n16267 = pi2185 & n12126;
  assign n16268 = ~n16266 & ~n16267;
  assign n16269 = pi1937 & ~n16268;
  assign po1788 = n16265 | n16269;
  assign n16271 = pi1738 & ~pi1941;
  assign n16272 = pi1738 & ~n12145;
  assign n16273 = pi2185 & n12145;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = pi1941 & ~n16274;
  assign po1789 = n16271 | n16275;
  assign n16277 = pi1739 & ~pi1941;
  assign n16278 = pi1739 & ~n12145;
  assign n16279 = pi2187 & n12145;
  assign n16280 = ~n16278 & ~n16279;
  assign n16281 = pi1941 & ~n16280;
  assign po1790 = n16277 | n16281;
  assign n16283 = pi1740 & ~pi1937;
  assign n16284 = pi1740 & ~n12126;
  assign n16285 = pi2176 & n12126;
  assign n16286 = ~n16284 & ~n16285;
  assign n16287 = pi1937 & ~n16286;
  assign po1791 = n16283 | n16287;
  assign n16289 = pi1741 & ~pi1941;
  assign n16290 = pi1741 & ~n12145;
  assign n16291 = pi2171 & n12145;
  assign n16292 = ~n16290 & ~n16291;
  assign n16293 = pi1941 & ~n16292;
  assign po1792 = n16289 | n16293;
  assign n16295 = pi1742 & ~pi1941;
  assign n16296 = pi1742 & ~n12145;
  assign n16297 = pi2169 & n12145;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = pi1941 & ~n16298;
  assign po1793 = n16295 | n16299;
  assign n16301 = pi1743 & ~pi1941;
  assign n16302 = pi1743 & ~n12145;
  assign n16303 = pi2190 & n12145;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = pi1941 & ~n16304;
  assign po1794 = n16301 | n16305;
  assign n16307 = pi1744 & ~pi1937;
  assign n16308 = pi1744 & ~n12126;
  assign n16309 = pi2169 & n12126;
  assign n16310 = ~n16308 & ~n16309;
  assign n16311 = pi1937 & ~n16310;
  assign po1795 = n16307 | n16311;
  assign n16313 = pi1745 & ~pi1937;
  assign n16314 = pi1745 & ~n12126;
  assign n16315 = pi2190 & n12126;
  assign n16316 = ~n16314 & ~n16315;
  assign n16317 = pi1937 & ~n16316;
  assign po1796 = n16313 | n16317;
  assign n16319 = pi1746 & ~pi1937;
  assign n16320 = pi1746 & ~n12126;
  assign n16321 = pi2170 & n12126;
  assign n16322 = ~n16320 & ~n16321;
  assign n16323 = pi1937 & ~n16322;
  assign po1797 = n16319 | n16323;
  assign n16325 = pi1747 & ~pi1937;
  assign n16326 = pi1747 & ~n12126;
  assign n16327 = pi2182 & n12126;
  assign n16328 = ~n16326 & ~n16327;
  assign n16329 = pi1937 & ~n16328;
  assign po1798 = n16325 | n16329;
  assign n16331 = pi1748 & ~pi1941;
  assign n16332 = pi1748 & ~n12145;
  assign n16333 = pi2166 & n12145;
  assign n16334 = ~n16332 & ~n16333;
  assign n16335 = pi1941 & ~n16334;
  assign po1799 = n16331 | n16335;
  assign n16337 = pi1749 & ~pi1941;
  assign n16338 = pi1749 & ~n12145;
  assign n16339 = pi2195 & n12145;
  assign n16340 = ~n16338 & ~n16339;
  assign n16341 = pi1941 & ~n16340;
  assign po1800 = n16337 | n16341;
  assign n16343 = pi1750 & ~pi1941;
  assign n16344 = pi1750 & ~n12145;
  assign n16345 = pi2184 & n12145;
  assign n16346 = ~n16344 & ~n16345;
  assign n16347 = pi1941 & ~n16346;
  assign po1801 = n16343 | n16347;
  assign n16349 = pi1751 & ~pi1941;
  assign n16350 = pi1751 & ~n12145;
  assign n16351 = pi2192 & n12145;
  assign n16352 = ~n16350 & ~n16351;
  assign n16353 = pi1941 & ~n16352;
  assign po1802 = n16349 | n16353;
  assign n16355 = pi1752 & ~pi1937;
  assign n16356 = pi1752 & ~n12126;
  assign n16357 = pi2177 & n12126;
  assign n16358 = ~n16356 & ~n16357;
  assign n16359 = pi1937 & ~n16358;
  assign po1803 = n16355 | n16359;
  assign n16361 = pi1753 & ~pi1937;
  assign n16362 = pi1753 & ~n12126;
  assign n16363 = pi2194 & n12126;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = pi1937 & ~n16364;
  assign po1804 = n16361 | n16365;
  assign n16367 = pi1754 & ~pi1937;
  assign n16368 = pi1754 & ~n12126;
  assign n16369 = pi2195 & n12126;
  assign n16370 = ~n16368 & ~n16369;
  assign n16371 = pi1937 & ~n16370;
  assign po1805 = n16367 | n16371;
  assign n16373 = pi1755 & ~pi1940;
  assign n16374 = pi2183 & n11852;
  assign n16375 = pi1755 & ~n11852;
  assign n16376 = ~n16374 & ~n16375;
  assign n16377 = pi1940 & ~n16376;
  assign po1806 = n16373 | n16377;
  assign n16379 = ~pi1756 & ~po1956;
  assign n16380 = pi2166 & po1956;
  assign po1807 = n16379 | n16380;
  assign n16382 = pi1757 & ~pi1936;
  assign n16383 = pi2176 & n11845;
  assign n16384 = pi1757 & ~n11845;
  assign n16385 = ~n16383 & ~n16384;
  assign n16386 = pi1936 & ~n16385;
  assign po1808 = n16382 | n16386;
  assign n16388 = pi1758 & ~pi1936;
  assign n16389 = pi1758 & ~n12004;
  assign n16390 = pi2186 & n12004;
  assign n16391 = ~n16389 & ~n16390;
  assign n16392 = pi1936 & ~n16391;
  assign po1809 = n16388 | n16392;
  assign n16394 = pi1759 & ~pi1936;
  assign n16395 = pi2167 & n11751;
  assign n16396 = pi1759 & ~n11751;
  assign n16397 = ~n16395 & ~n16396;
  assign n16398 = pi1936 & ~n16397;
  assign po1810 = n16394 | n16398;
  assign n16400 = pi1760 & ~n12907;
  assign n16401 = pi2170 & n12907;
  assign po1811 = n16400 | n16401;
  assign n16403 = pi1761 & ~pi1936;
  assign n16404 = pi2191 & n11751;
  assign n16405 = pi1761 & ~n11751;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = pi1936 & ~n16406;
  assign po1812 = n16403 | n16407;
  assign n16409 = pi2176 & n12295;
  assign n16410 = pi1762 & ~n12295;
  assign po1813 = n16409 | n16410;
  assign n16412 = pi1763 & ~pi1936;
  assign n16413 = pi2170 & n11751;
  assign n16414 = pi1763 & ~n11751;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = pi1936 & ~n16415;
  assign po1814 = n16412 | n16416;
  assign n16418 = pi1764 & ~pi1936;
  assign n16419 = pi2176 & n11751;
  assign n16420 = pi1764 & ~n11751;
  assign n16421 = ~n16419 & ~n16420;
  assign n16422 = pi1936 & ~n16421;
  assign po1815 = n16418 | n16422;
  assign n16424 = pi1765 & ~pi1936;
  assign n16425 = pi2178 & n11751;
  assign n16426 = pi1765 & ~n11751;
  assign n16427 = ~n16425 & ~n16426;
  assign n16428 = pi1936 & ~n16427;
  assign po1816 = n16424 | n16428;
  assign n16430 = pi1766 & ~pi1939;
  assign n16431 = pi1766 & ~n11943;
  assign n16432 = pi2184 & n11943;
  assign n16433 = ~n16431 & ~n16432;
  assign n16434 = pi1939 & ~n16433;
  assign po1817 = n16430 | n16434;
  assign n16436 = pi1767 & ~pi1936;
  assign n16437 = pi2179 & n11751;
  assign n16438 = pi1767 & ~n11751;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = pi1936 & ~n16439;
  assign po1818 = n16436 | n16440;
  assign n16442 = pi1769 & ~pi1939;
  assign n16443 = pi1769 & ~n11943;
  assign n16444 = pi2177 & n11943;
  assign n16445 = ~n16443 & ~n16444;
  assign n16446 = pi1939 & ~n16445;
  assign po1820 = n16442 | n16446;
  assign n16448 = pi1770 & ~pi1939;
  assign n16449 = pi1770 & ~n11943;
  assign n16450 = pi2171 & n11943;
  assign n16451 = ~n16449 & ~n16450;
  assign n16452 = pi1939 & ~n16451;
  assign po1821 = n16448 | n16452;
  assign n16454 = pi1771 & ~po1956;
  assign n16455 = pi2189 & po1956;
  assign po1822 = n16454 | n16455;
  assign n16457 = pi1772 & ~pi1936;
  assign n16458 = pi2167 & n11845;
  assign n16459 = pi1772 & ~n11845;
  assign n16460 = ~n16458 & ~n16459;
  assign n16461 = pi1936 & ~n16460;
  assign po1823 = n16457 | n16461;
  assign n16463 = pi1773 & ~pi1936;
  assign n16464 = pi2172 & n11751;
  assign n16465 = pi1773 & ~n11751;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = pi1936 & ~n16466;
  assign po1824 = n16463 | n16467;
  assign n16469 = pi1774 & ~pi1936;
  assign n16470 = pi2195 & n11845;
  assign n16471 = pi1774 & ~n11845;
  assign n16472 = ~n16470 & ~n16471;
  assign n16473 = pi1936 & ~n16472;
  assign po1825 = n16469 | n16473;
  assign n16475 = pi1775 & ~pi1936;
  assign n16476 = pi2191 & n11845;
  assign n16477 = pi1775 & ~n11845;
  assign n16478 = ~n16476 & ~n16477;
  assign n16479 = pi1936 & ~n16478;
  assign po1826 = n16475 | n16479;
  assign n16481 = pi1776 & ~pi1937;
  assign n16482 = pi1776 & ~n12126;
  assign n16483 = pi2192 & n12126;
  assign n16484 = ~n16482 & ~n16483;
  assign n16485 = pi1937 & ~n16484;
  assign po1827 = n16481 | n16485;
  assign n16487 = pi2170 & n12295;
  assign n16488 = pi1777 & ~n12295;
  assign po1828 = n16487 | n16488;
  assign n16490 = pi1778 & ~pi1939;
  assign n16491 = pi1778 & ~n11943;
  assign n16492 = pi2182 & n11943;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = pi1939 & ~n16493;
  assign po1829 = n16490 | n16494;
  assign n16496 = pi1779 & ~n12907;
  assign n16497 = pi2194 & n12907;
  assign po1830 = n16496 | n16497;
  assign n16499 = pi1780 & ~pi1936;
  assign n16500 = pi2170 & n11845;
  assign n16501 = pi1780 & ~n11845;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = pi1936 & ~n16502;
  assign po1831 = n16499 | n16503;
  assign n16505 = pi1781 & ~pi1937;
  assign n16506 = pi1781 & ~n12126;
  assign n16507 = pi2167 & n12126;
  assign n16508 = ~n16506 & ~n16507;
  assign n16509 = pi1937 & ~n16508;
  assign po1832 = n16505 | n16509;
  assign n16511 = pi1782 & ~pi1939;
  assign n16512 = pi1782 & ~n11943;
  assign n16513 = pi2185 & n11943;
  assign n16514 = ~n16512 & ~n16513;
  assign n16515 = pi1939 & ~n16514;
  assign po1833 = n16511 | n16515;
  assign n16517 = pi1783 & ~pi1941;
  assign n16518 = pi1783 & ~n12145;
  assign n16519 = pi2173 & n12145;
  assign n16520 = ~n16518 & ~n16519;
  assign n16521 = pi1941 & ~n16520;
  assign po1834 = n16517 | n16521;
  assign n16523 = pi1784 & ~pi1936;
  assign n16524 = pi2178 & n11845;
  assign n16525 = pi1784 & ~n11845;
  assign n16526 = ~n16524 & ~n16525;
  assign n16527 = pi1936 & ~n16526;
  assign po1835 = n16523 | n16527;
  assign n16529 = pi1785 & ~pi1936;
  assign n16530 = pi2178 & n11844;
  assign n16531 = pi1785 & ~n11844;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = pi1936 & ~n16532;
  assign po1836 = n16529 | n16533;
  assign n16535 = pi1786 & ~pi1936;
  assign n16536 = pi2179 & n11845;
  assign n16537 = pi1786 & ~n11845;
  assign n16538 = ~n16536 & ~n16537;
  assign n16539 = pi1936 & ~n16538;
  assign po1837 = n16535 | n16539;
  assign n16541 = pi1787 & ~pi1936;
  assign n16542 = pi2172 & n11845;
  assign n16543 = pi1787 & ~n11845;
  assign n16544 = ~n16542 & ~n16543;
  assign n16545 = pi1936 & ~n16544;
  assign po1838 = n16541 | n16545;
  assign n16547 = pi1788 & ~pi1939;
  assign n16548 = pi1788 & ~n11943;
  assign n16549 = pi2193 & n11943;
  assign n16550 = ~n16548 & ~n16549;
  assign n16551 = pi1939 & ~n16550;
  assign po1839 = n16547 | n16551;
  assign n16553 = pi2179 & n12295;
  assign n16554 = pi1789 & ~n12295;
  assign po1840 = n16553 | n16554;
  assign n16556 = pi1790 & ~pi1939;
  assign n16557 = pi1790 & ~n11943;
  assign n16558 = pi2168 & n11943;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = pi1939 & ~n16559;
  assign po1841 = n16556 | n16560;
  assign n16562 = pi1791 & ~pi1936;
  assign n16563 = pi2170 & n11844;
  assign n16564 = pi1791 & ~n11844;
  assign n16565 = ~n16563 & ~n16564;
  assign n16566 = pi1936 & ~n16565;
  assign po1842 = n16562 | n16566;
  assign n16568 = pi1792 & ~pi1938;
  assign n16569 = pi1792 & ~n11882;
  assign n16570 = pi2184 & n11882;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = pi1938 & ~n16571;
  assign po1843 = n16568 | n16572;
  assign n16574 = pi1793 & ~pi1936;
  assign n16575 = pi2167 & n11844;
  assign n16576 = pi1793 & ~n11844;
  assign n16577 = ~n16575 & ~n16576;
  assign n16578 = pi1936 & ~n16577;
  assign po1844 = n16574 | n16578;
  assign n16580 = pi1794 & ~pi1936;
  assign n16581 = pi2195 & n11844;
  assign n16582 = pi1794 & ~n11844;
  assign n16583 = ~n16581 & ~n16582;
  assign n16584 = pi1936 & ~n16583;
  assign po1845 = n16580 | n16584;
  assign n16586 = pi1795 & ~pi1936;
  assign n16587 = pi2191 & n11844;
  assign n16588 = pi1795 & ~n11844;
  assign n16589 = ~n16587 & ~n16588;
  assign n16590 = pi1936 & ~n16589;
  assign po1846 = n16586 | n16590;
  assign n16592 = pi1796 & ~pi1939;
  assign n16593 = pi1796 & ~n11943;
  assign n16594 = pi2186 & n11943;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = pi1939 & ~n16595;
  assign po1847 = n16592 | n16596;
  assign n16598 = pi1797 & ~pi1936;
  assign n16599 = pi2176 & n11844;
  assign n16600 = pi1797 & ~n11844;
  assign n16601 = ~n16599 & ~n16600;
  assign n16602 = pi1936 & ~n16601;
  assign po1848 = n16598 | n16602;
  assign n16604 = pi1798 & ~pi1941;
  assign n16605 = pi1798 & ~n12145;
  assign n16606 = pi2194 & n12145;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = pi1941 & ~n16607;
  assign po1849 = n16604 | n16608;
  assign n16610 = pi1799 & ~pi1938;
  assign n16611 = pi1799 & ~n11882;
  assign n16612 = pi2177 & n11882;
  assign n16613 = ~n16611 & ~n16612;
  assign n16614 = pi1938 & ~n16613;
  assign po1850 = n16610 | n16614;
  assign n16616 = pi1800 & ~pi1941;
  assign n16617 = pi1800 & ~n12145;
  assign n16618 = pi2196 & n12145;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = pi1941 & ~n16619;
  assign po1851 = n16616 | n16620;
  assign n16622 = pi1801 & ~pi1939;
  assign n16623 = pi2195 & n11786;
  assign n16624 = pi1801 & ~n11786;
  assign n16625 = ~n16623 & ~n16624;
  assign n16626 = pi1939 & ~n16625;
  assign po1852 = n16622 | n16626;
  assign n16628 = pi1802 & ~pi1936;
  assign n16629 = pi2172 & n11844;
  assign n16630 = pi1802 & ~n11844;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = pi1936 & ~n16631;
  assign po1853 = n16628 | n16632;
  assign n16634 = pi1803 & ~pi1939;
  assign n16635 = pi2167 & n11786;
  assign n16636 = pi1803 & ~n11786;
  assign n16637 = ~n16635 & ~n16636;
  assign n16638 = pi1939 & ~n16637;
  assign po1854 = n16634 | n16638;
  assign n16640 = pi1804 & ~pi1941;
  assign n16641 = pi1804 & ~n12145;
  assign n16642 = pi2191 & n12145;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = pi1941 & ~n16643;
  assign po1855 = n16640 | n16644;
  assign n16646 = pi1805 & ~pi1939;
  assign n16647 = pi2195 & n11746;
  assign n16648 = pi1805 & ~n11746;
  assign n16649 = ~n16647 & ~n16648;
  assign n16650 = pi1939 & ~n16649;
  assign po1856 = n16646 | n16650;
  assign n16652 = pi1806 & ~pi1938;
  assign n16653 = pi1806 & ~n11882;
  assign n16654 = pi2171 & n11882;
  assign n16655 = ~n16653 & ~n16654;
  assign n16656 = pi1938 & ~n16655;
  assign po1857 = n16652 | n16656;
  assign n16658 = pi1807 & ~pi1937;
  assign n16659 = pi1807 & ~n12126;
  assign n16660 = pi2171 & n12126;
  assign n16661 = ~n16659 & ~n16660;
  assign n16662 = pi1937 & ~n16661;
  assign po1858 = n16658 | n16662;
  assign n16664 = pi1808 & ~pi1938;
  assign n16665 = pi1808 & ~n11882;
  assign n16666 = pi2193 & n11882;
  assign n16667 = ~n16665 & ~n16666;
  assign n16668 = pi1938 & ~n16667;
  assign po1859 = n16664 | n16668;
  assign n16670 = pi1809 & ~pi1939;
  assign n16671 = pi2179 & n11786;
  assign n16672 = pi1809 & ~n11786;
  assign n16673 = ~n16671 & ~n16672;
  assign n16674 = pi1939 & ~n16673;
  assign po1860 = n16670 | n16674;
  assign n16676 = pi1810 & ~pi1939;
  assign n16677 = pi2170 & n11786;
  assign n16678 = pi1810 & ~n11786;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = pi1939 & ~n16679;
  assign po1861 = n16676 | n16680;
  assign n16682 = pi1811 & ~pi1939;
  assign n16683 = pi2191 & n11786;
  assign n16684 = pi1811 & ~n11786;
  assign n16685 = ~n16683 & ~n16684;
  assign n16686 = pi1939 & ~n16685;
  assign po1862 = n16682 | n16686;
  assign n16688 = pi1812 & ~pi1939;
  assign n16689 = pi2176 & n11786;
  assign n16690 = pi1812 & ~n11786;
  assign n16691 = ~n16689 & ~n16690;
  assign n16692 = pi1939 & ~n16691;
  assign po1863 = n16688 | n16692;
  assign n16694 = pi1813 & ~pi1939;
  assign n16695 = pi2178 & n11786;
  assign n16696 = pi1813 & ~n11786;
  assign n16697 = ~n16695 & ~n16696;
  assign n16698 = pi1939 & ~n16697;
  assign po1864 = n16694 | n16698;
  assign n16700 = pi1814 & ~pi1941;
  assign n16701 = pi1814 & ~n12145;
  assign n16702 = pi2181 & n12145;
  assign n16703 = ~n16701 & ~n16702;
  assign n16704 = pi1941 & ~n16703;
  assign po1865 = n16700 | n16704;
  assign n16706 = pi1815 & ~pi1938;
  assign n16707 = pi1815 & ~n11882;
  assign n16708 = pi2185 & n11882;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = pi1938 & ~n16709;
  assign po1866 = n16706 | n16710;
  assign n16712 = pi1816 & ~pi1939;
  assign n16713 = pi2172 & n11786;
  assign n16714 = pi1816 & ~n11786;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 = pi1939 & ~n16715;
  assign po1867 = n16712 | n16716;
  assign n16718 = pi1817 & ~pi1939;
  assign n16719 = pi2191 & n11746;
  assign n16720 = pi1817 & ~n11746;
  assign n16721 = ~n16719 & ~n16720;
  assign n16722 = pi1939 & ~n16721;
  assign po1868 = n16718 | n16722;
  assign n16724 = pi1818 & ~pi1938;
  assign n16725 = pi1818 & ~n11882;
  assign n16726 = pi2168 & n11882;
  assign n16727 = ~n16725 & ~n16726;
  assign n16728 = pi1938 & ~n16727;
  assign po1869 = n16724 | n16728;
  assign n16730 = pi1819 & ~pi1939;
  assign n16731 = pi2170 & n11746;
  assign n16732 = pi1819 & ~n11746;
  assign n16733 = ~n16731 & ~n16732;
  assign n16734 = pi1939 & ~n16733;
  assign po1870 = n16730 | n16734;
  assign n16736 = pi1820 & ~pi1941;
  assign n16737 = pi1820 & ~n12145;
  assign n16738 = pi2176 & n12145;
  assign n16739 = ~n16737 & ~n16738;
  assign n16740 = pi1941 & ~n16739;
  assign po1871 = n16736 | n16740;
  assign n16742 = pi2178 & n12295;
  assign n16743 = pi1821 & ~n12295;
  assign po1872 = n16742 | n16743;
  assign n16745 = pi1822 & ~pi1939;
  assign n16746 = pi2191 & n11745;
  assign n16747 = pi1822 & ~n11745;
  assign n16748 = ~n16746 & ~n16747;
  assign n16749 = pi1939 & ~n16748;
  assign po1873 = n16745 | n16749;
  assign n16751 = pi1823 & ~pi1939;
  assign n16752 = pi2172 & n11746;
  assign n16753 = pi1823 & ~n11746;
  assign n16754 = ~n16752 & ~n16753;
  assign n16755 = pi1939 & ~n16754;
  assign po1874 = n16751 | n16755;
  assign n16757 = pi1824 & ~pi1937;
  assign n16758 = pi2170 & n11828;
  assign n16759 = pi1824 & ~n11828;
  assign n16760 = ~n16758 & ~n16759;
  assign n16761 = pi1937 & ~n16760;
  assign po1875 = n16757 | n16761;
  assign n16763 = pi1825 & ~pi1939;
  assign n16764 = pi2179 & n11746;
  assign n16765 = pi1825 & ~n11746;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = pi1939 & ~n16766;
  assign po1876 = n16763 | n16767;
  assign n16769 = pi1826 & ~pi1939;
  assign n16770 = pi2176 & n11746;
  assign n16771 = pi1826 & ~n11746;
  assign n16772 = ~n16770 & ~n16771;
  assign n16773 = pi1939 & ~n16772;
  assign po1877 = n16769 | n16773;
  assign n16775 = pi1827 & ~pi1939;
  assign n16776 = pi2178 & n11746;
  assign n16777 = pi1827 & ~n11746;
  assign n16778 = ~n16776 & ~n16777;
  assign n16779 = pi1939 & ~n16778;
  assign po1878 = n16775 | n16779;
  assign n16781 = pi1828 & ~pi1941;
  assign n16782 = pi2194 & n11821;
  assign n16783 = pi1828 & ~n11821;
  assign n16784 = ~n16782 & ~n16783;
  assign n16785 = pi1941 & ~n16784;
  assign po1879 = n16781 | n16785;
  assign n16787 = pi1829 & ~pi1939;
  assign n16788 = pi2195 & n11745;
  assign n16789 = pi1829 & ~n11745;
  assign n16790 = ~n16788 & ~n16789;
  assign n16791 = pi1939 & ~n16790;
  assign po1880 = n16787 | n16791;
  assign n16793 = pi1830 & ~pi1939;
  assign n16794 = pi2167 & n11745;
  assign n16795 = pi1830 & ~n11745;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = pi1939 & ~n16796;
  assign po1881 = n16793 | n16797;
  assign n16799 = pi1831 & ~pi1941;
  assign n16800 = pi1831 & ~n12145;
  assign n16801 = pi2198 & n12145;
  assign n16802 = ~n16800 & ~n16801;
  assign n16803 = pi1941 & ~n16802;
  assign po1882 = n16799 | n16803;
  assign n16805 = n5422 & n12386;
  assign n16806 = pi2172 & n16805;
  assign n16807 = pi1832 & ~n16805;
  assign po1883 = n16806 | n16807;
  assign n16809 = pi1833 & ~pi1937;
  assign n16810 = pi1833 & ~n12126;
  assign n16811 = pi2186 & n12126;
  assign n16812 = ~n16810 & ~n16811;
  assign n16813 = pi1937 & ~n16812;
  assign po1884 = n16809 | n16813;
  assign n16815 = pi2119 & n11507;
  assign n16816 = pi2082 & n11512;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = pi1210 & n11519;
  assign n16819 = pi2151 & n11521;
  assign n16820 = ~n16818 & ~n16819;
  assign n16821 = pi1975 & n5423;
  assign n16822 = n16820 & ~n16821;
  assign n16823 = pi1131 & n11529;
  assign n16824 = n16822 & ~n16823;
  assign n16825 = pi1873 & n11532;
  assign n16826 = pi1159 & n11535;
  assign n16827 = ~n16825 & ~n16826;
  assign n16828 = n16824 & n16827;
  assign n16829 = n11517 & ~n16828;
  assign n16830 = pi2050 & n11515;
  assign n16831 = ~n16829 & ~n16830;
  assign po1886 = ~n16817 | ~n16831;
  assign n16833 = pi2121 & n11507;
  assign n16834 = pi2084 & n11512;
  assign n16835 = ~n16833 & ~n16834;
  assign n16836 = pi1208 & n11519;
  assign n16837 = pi2143 & n11521;
  assign n16838 = ~n16836 & ~n16837;
  assign n16839 = pi1977 & n5423;
  assign n16840 = n16838 & ~n16839;
  assign n16841 = pi1185 & n11529;
  assign n16842 = n16840 & ~n16841;
  assign n16843 = pi1848 & n11532;
  assign n16844 = pi1161 & n11535;
  assign n16845 = ~n16843 & ~n16844;
  assign n16846 = n16842 & n16845;
  assign n16847 = n11517 & ~n16846;
  assign n16848 = pi2051 & n11515;
  assign n16849 = ~n16847 & ~n16848;
  assign po1887 = ~n16835 | ~n16849;
  assign n16851 = pi2092 & n11507;
  assign n16852 = pi2129 & n11512;
  assign n16853 = ~n16851 & ~n16852;
  assign n16854 = pi1189 & n11519;
  assign n16855 = pi2149 & n11521;
  assign n16856 = ~n16854 & ~n16855;
  assign n16857 = pi1964 & n5423;
  assign n16858 = n16856 & ~n16857;
  assign n16859 = pi1165 & n11529;
  assign n16860 = n16858 & ~n16859;
  assign n16861 = pi1840 & n11532;
  assign n16862 = pi1146 & n11535;
  assign n16863 = ~n16861 & ~n16862;
  assign n16864 = n16860 & n16863;
  assign n16865 = n11517 & ~n16864;
  assign n16866 = pi2040 & n11515;
  assign n16867 = ~n16865 & ~n16866;
  assign po1888 = ~n16853 | ~n16867;
  assign n16869 = pi2195 & n16805;
  assign n16870 = pi1838 & ~n16805;
  assign po1889 = n16869 | n16870;
  assign n16872 = pi2186 & n16805;
  assign n16873 = pi1839 & ~n16805;
  assign po1890 = n16872 | n16873;
  assign n16875 = pi2183 & n16805;
  assign n16876 = pi1840 & ~n16805;
  assign po1891 = n16875 | n16876;
  assign n16878 = pi2168 & n16805;
  assign n16879 = pi1841 & ~n16805;
  assign po1892 = n16878 | n16879;
  assign n16881 = pi2174 & n16805;
  assign n16882 = pi1842 & ~n16805;
  assign po1893 = n16881 | n16882;
  assign n16884 = pi2197 & n16805;
  assign n16885 = pi1843 & ~n16805;
  assign po1894 = n16884 | n16885;
  assign n16887 = pi2198 & n16805;
  assign n16888 = pi1844 & ~n16805;
  assign po1895 = n16887 | n16888;
  assign n16890 = pi2191 & n16805;
  assign n16891 = pi1845 & ~n16805;
  assign po1896 = n16890 | n16891;
  assign n16893 = pi2194 & n16805;
  assign n16894 = pi1846 & ~n16805;
  assign po1897 = n16893 | n16894;
  assign n16896 = pi2188 & n16805;
  assign n16897 = pi1847 & ~n16805;
  assign po1898 = n16896 | n16897;
  assign n16899 = pi2184 & n16805;
  assign n16900 = pi1848 & ~n16805;
  assign po1899 = n16899 | n16900;
  assign n16902 = pi2166 & n16805;
  assign n16903 = pi1849 & ~n16805;
  assign po1900 = n16902 | n16903;
  assign n16905 = pi1928 & ~pi2035;
  assign n16906 = pi1850 & pi2035;
  assign po1901 = n16905 | n16906;
  assign n16908 = pi1928 & ~pi2056;
  assign n16909 = pi1851 & pi2056;
  assign po1902 = n16908 | n16909;
  assign n16911 = pi1928 & ~pi2057;
  assign n16912 = pi1852 & pi2057;
  assign po1903 = n16911 | n16912;
  assign n16914 = pi1928 & ~pi2059;
  assign n16915 = pi1853 & pi2059;
  assign po1904 = n16914 | n16915;
  assign n16917 = pi1854 & ~pi1937;
  assign n16918 = pi1854 & ~n12126;
  assign n16919 = pi2197 & n12126;
  assign n16920 = ~n16918 & ~n16919;
  assign n16921 = pi1937 & ~n16920;
  assign po1905 = n16917 | n16921;
  assign n16923 = pi1855 & ~pi1937;
  assign n16924 = pi1855 & ~n12126;
  assign n16925 = pi2166 & n12126;
  assign n16926 = ~n16924 & ~n16925;
  assign n16927 = pi1937 & ~n16926;
  assign po1906 = n16923 | n16927;
  assign n16929 = pi1931 & pi2033;
  assign n16930 = pi1856 & ~pi1931;
  assign po1907 = n16929 | n16930;
  assign n16932 = ~pi1943 & pi2020;
  assign n16933 = pi1857 & pi1943;
  assign po1908 = n16932 | n16933;
  assign n16935 = pi2091 & n11507;
  assign n16936 = pi2127 & n11512;
  assign n16937 = ~n16935 & ~n16936;
  assign n16938 = pi1188 & n11519;
  assign n16939 = pi2156 & n11521;
  assign n16940 = ~n16938 & ~n16939;
  assign n16941 = pi1948 & n5423;
  assign n16942 = n16940 & ~n16941;
  assign n16943 = pi1164 & n11529;
  assign n16944 = n16942 & ~n16943;
  assign n16945 = pi1839 & n11532;
  assign n16946 = pi1145 & n11535;
  assign n16947 = ~n16945 & ~n16946;
  assign n16948 = n16944 & n16947;
  assign n16949 = n11517 & ~n16948;
  assign n16950 = pi2039 & n11515;
  assign n16951 = ~n16949 & ~n16950;
  assign po1909 = ~n16937 | ~n16951;
  assign n16953 = pi2097 & n11507;
  assign n16954 = pi2062 & n11512;
  assign n16955 = ~n16953 & ~n16954;
  assign n16956 = pi1193 & n11519;
  assign n16957 = pi2148 & n11521;
  assign n16958 = ~n16956 & ~n16957;
  assign n16959 = pi0248 & n5423;
  assign n16960 = n16958 & ~n16959;
  assign n16961 = pi1168 & n11529;
  assign n16962 = n16960 & ~n16961;
  assign n16963 = pi1843 & n11532;
  assign n16964 = pi1149 & n11535;
  assign n16965 = ~n16963 & ~n16964;
  assign n16966 = n16962 & n16965;
  assign n16967 = n11517 & ~n16966;
  assign n16968 = pi2021 & n11515;
  assign n16969 = ~n16967 & ~n16968;
  assign po1910 = ~n16955 | ~n16969;
  assign n16971 = pi2095 & n11507;
  assign n16972 = pi2090 & n11512;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = pi1192 & n11519;
  assign n16975 = pi2154 & n11521;
  assign n16976 = ~n16974 & ~n16975;
  assign n16977 = pi1966 & n5423;
  assign n16978 = n16976 & ~n16977;
  assign n16979 = pi1167 & n11529;
  assign n16980 = n16978 & ~n16979;
  assign n16981 = pi1842 & n11532;
  assign n16982 = pi1148 & n11535;
  assign n16983 = ~n16981 & ~n16982;
  assign n16984 = n16980 & n16983;
  assign n16985 = n11517 & ~n16984;
  assign n16986 = pi2042 & n11515;
  assign n16987 = ~n16985 & ~n16986;
  assign po1911 = ~n16973 | ~n16987;
  assign n16989 = pi2094 & n11507;
  assign n16990 = pi2128 & n11512;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = pi1191 & n11519;
  assign n16993 = pi2145 & n11521;
  assign n16994 = ~n16992 & ~n16993;
  assign n16995 = pi1965 & n5423;
  assign n16996 = n16994 & ~n16995;
  assign n16997 = pi1166 & n11529;
  assign n16998 = n16996 & ~n16997;
  assign n16999 = pi1841 & n11532;
  assign n17000 = pi1147 & n11535;
  assign n17001 = ~n16999 & ~n17000;
  assign n17002 = n16998 & n17001;
  assign n17003 = n11517 & ~n17002;
  assign n17004 = pi2041 & n11515;
  assign n17005 = ~n17003 & ~n17004;
  assign po1912 = ~n16991 | ~n17005;
  assign n17007 = pi2093 & n11507;
  assign n17008 = pi2061 & n11512;
  assign n17009 = ~n17007 & ~n17008;
  assign n17010 = pi1190 & n11519;
  assign n17011 = pi2153 & n11521;
  assign n17012 = ~n17010 & ~n17011;
  assign n17013 = pi0229 & n5423;
  assign n17014 = n17012 & ~n17013;
  assign n17015 = pi1020 & n11529;
  assign n17016 = n17014 & ~n17015;
  assign n17017 = pi1832 & n11532;
  assign n17018 = pi1134 & n11535;
  assign n17019 = ~n17017 & ~n17018;
  assign n17020 = n17016 & n17019;
  assign n17021 = n11517 & ~n17020;
  assign n17022 = pi2038 & n11515;
  assign n17023 = ~n17021 & ~n17022;
  assign po1913 = ~n17009 | ~n17023;
  assign n17025 = pi2124 & n11507;
  assign n17026 = pi2087 & n11512;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = pi1209 & n11519;
  assign n17029 = pi2144 & n11521;
  assign n17030 = ~n17028 & ~n17029;
  assign n17031 = pi1982 & n5423;
  assign n17032 = n17030 & ~n17031;
  assign n17033 = pi1187 & n11529;
  assign n17034 = n17032 & ~n17033;
  assign n17035 = pi1870 & n11532;
  assign n17036 = pi1163 & n11535;
  assign n17037 = ~n17035 & ~n17036;
  assign n17038 = n17034 & n17037;
  assign n17039 = n11517 & ~n17038;
  assign n17040 = pi2054 & n11515;
  assign n17041 = ~n17039 & ~n17040;
  assign po1914 = ~n17027 | ~n17041;
  assign n17043 = pi2122 & n11507;
  assign n17044 = pi2085 & n11512;
  assign n17045 = ~n17043 & ~n17044;
  assign n17046 = pi1132 & n11519;
  assign n17047 = pi2147 & n11521;
  assign n17048 = ~n17046 & ~n17047;
  assign n17049 = pi1976 & n5423;
  assign n17050 = n17048 & ~n17049;
  assign n17051 = pi1186 & n11529;
  assign n17052 = n17050 & ~n17051;
  assign n17053 = pi1849 & n11532;
  assign n17054 = pi1162 & n11535;
  assign n17055 = ~n17053 & ~n17054;
  assign n17056 = n17052 & n17055;
  assign n17057 = n11517 & ~n17056;
  assign n17058 = pi2052 & n11515;
  assign n17059 = ~n17057 & ~n17058;
  assign po1915 = ~n17045 | ~n17059;
  assign n17061 = pi2098 & n11507;
  assign n17062 = pi2125 & n11512;
  assign n17063 = ~n17061 & ~n17062;
  assign n17064 = pi1211 & n11519;
  assign n17065 = pi2150 & n11521;
  assign n17066 = ~n17064 & ~n17065;
  assign n17067 = pi1950 & n5423;
  assign n17068 = n17066 & ~n17067;
  assign n17069 = pi1821 & n11529;
  assign n17070 = n17068 & ~n17069;
  assign n17071 = pi1871 & n11532;
  assign n17072 = pi1137 & n11535;
  assign n17073 = ~n17071 & ~n17072;
  assign n17074 = n17070 & n17073;
  assign n17075 = n11517 & ~n17074;
  assign n17076 = pi2022 & n11515;
  assign n17077 = ~n17075 & ~n17076;
  assign po1916 = ~n17063 | ~n17077;
  assign n17079 = pi2120 & n11507;
  assign n17080 = pi2083 & n11512;
  assign n17081 = ~n17079 & ~n17080;
  assign n17082 = pi1207 & n11519;
  assign n17083 = pi2157 & n11521;
  assign n17084 = ~n17082 & ~n17083;
  assign n17085 = pi0230 & n5423;
  assign n17086 = n17084 & ~n17085;
  assign n17087 = pi1184 & n11529;
  assign n17088 = n17086 & ~n17087;
  assign n17089 = pi1847 & n11532;
  assign n17090 = pi1160 & n11535;
  assign n17091 = ~n17089 & ~n17090;
  assign n17092 = n17088 & n17091;
  assign n17093 = n11517 & ~n17092;
  assign n17094 = pi2103 & n11515;
  assign n17095 = ~n17093 & ~n17094;
  assign po1917 = ~n17081 | ~n17095;
  assign n17097 = pi2118 & n11507;
  assign n17098 = pi2080 & n11512;
  assign n17099 = ~n17097 & ~n17098;
  assign n17100 = pi1779 & n11519;
  assign n17101 = pi2160 & n11521;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = pi1974 & n5423;
  assign n17104 = n17102 & ~n17103;
  assign n17105 = pi1183 & n11529;
  assign n17106 = n17104 & ~n17105;
  assign n17107 = pi1846 & n11532;
  assign n17108 = pi1158 & n11535;
  assign n17109 = ~n17107 & ~n17108;
  assign n17110 = n17106 & n17109;
  assign n17111 = n11517 & ~n17110;
  assign n17112 = pi2049 & n11515;
  assign n17113 = ~n17111 & ~n17112;
  assign po1918 = ~n17099 | ~n17113;
  assign n17115 = pi2123 & n11507;
  assign n17116 = pi2086 & n11512;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = pi1690 & n11519;
  assign n17119 = pi2152 & n11521;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = pi0251 & n5423;
  assign n17122 = n17120 & ~n17121;
  assign n17123 = pi1035 & n11529;
  assign n17124 = n17122 & ~n17123;
  assign n17125 = pi1838 & n11532;
  assign n17126 = pi1036 & n11535;
  assign n17127 = ~n17125 & ~n17126;
  assign n17128 = n17124 & n17127;
  assign n17129 = n11517 & ~n17128;
  assign n17130 = pi2053 & n11515;
  assign n17131 = ~n17129 & ~n17130;
  assign po1919 = ~n17117 | ~n17131;
  assign n17133 = pi2115 & n11507;
  assign n17134 = pi2077 & n11512;
  assign n17135 = ~n17133 & ~n17134;
  assign n17136 = pi1206 & n11519;
  assign n17137 = pi2155 & n11521;
  assign n17138 = ~n17136 & ~n17137;
  assign n17139 = pi0250 & n5423;
  assign n17140 = n17138 & ~n17139;
  assign n17141 = pi1130 & n11529;
  assign n17142 = n17140 & ~n17141;
  assign n17143 = pi1845 & n11532;
  assign n17144 = pi1157 & n11535;
  assign n17145 = ~n17143 & ~n17144;
  assign n17146 = n17142 & n17145;
  assign n17147 = n11517 & ~n17146;
  assign n17148 = pi2047 & n11515;
  assign n17149 = ~n17147 & ~n17148;
  assign po1920 = ~n17135 | ~n17149;
  assign n17151 = pi2192 & n16805;
  assign n17152 = pi1870 & ~n16805;
  assign po1921 = n17151 | n17152;
  assign n17154 = pi2178 & n16805;
  assign n17155 = pi1871 & ~n16805;
  assign po1922 = n17154 | n17155;
  assign n17157 = pi1872 & ~pi1937;
  assign n17158 = pi1872 & ~n12126;
  assign n17159 = pi2173 & n12126;
  assign n17160 = ~n17158 & ~n17159;
  assign n17161 = pi1937 & ~n17160;
  assign po1923 = n17157 | n17161;
  assign n17163 = pi2167 & n16805;
  assign n17164 = pi1873 & ~n16805;
  assign po1924 = n17163 | n17164;
  assign n17166 = ~pi0259 & ~pi2032;
  assign n17167 = pi1929 & pi2032;
  assign po1925 = n17166 | n17167;
  assign n17169 = pi1928 & ~pi2058;
  assign n17170 = pi1875 & pi2058;
  assign po1926 = n17169 | n17170;
  assign n17172 = ~pi1952 & pi2055;
  assign n17173 = pi1877 & pi1952;
  assign po1928 = n17172 | n17173;
  assign n17175 = ~pi1989 & ~pi2238;
  assign n17176 = n5418 & n17175;
  assign po1929 = pi2186 & n17176;
  assign po1930 = pi2198 & n17176;
  assign n17179 = pi2117 & n11507;
  assign n17180 = pi2079 & n11512;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = pi1144 & n11521;
  assign n17183 = pi1182 & n11529;
  assign n17184 = ~n17182 & ~n17183;
  assign n17185 = n11517 & ~n17184;
  assign n17186 = pi2096 & n11515;
  assign n17187 = ~n17185 & ~n17186;
  assign po1933 = ~n17181 | ~n17187;
  assign n17189 = pi1942 & ~pi2059;
  assign n17190 = pi1883 & pi2059;
  assign po1934 = n17189 | n17190;
  assign n17192 = pi1942 & ~pi2035;
  assign n17193 = pi1884 & pi2035;
  assign po1935 = n17192 | n17193;
  assign n17195 = pi1942 & ~pi2056;
  assign n17196 = pi1885 & pi2056;
  assign po1936 = n17195 | n17196;
  assign n17198 = pi1942 & ~pi2057;
  assign n17199 = pi1886 & pi2057;
  assign po1937 = n17198 | n17199;
  assign n17201 = pi1175 & n11529;
  assign n17202 = pi0841 & n5423;
  assign n17203 = ~n17201 & ~n17202;
  assign n17204 = pi1156 & n11535;
  assign n17205 = n17203 & ~n17204;
  assign n17206 = pi1201 & n11519;
  assign n17207 = n17205 & ~n17206;
  assign n17208 = n11517 & ~n17207;
  assign n17209 = pi2030 & n11515;
  assign n17210 = ~n17208 & ~n17209;
  assign n17211 = pi2108 & n11507;
  assign n17212 = pi2068 & n11512;
  assign n17213 = ~n17211 & ~n17212;
  assign po1938 = ~n17210 | ~n17213;
  assign n17215 = pi2107 & n11507;
  assign n17216 = pi2067 & n11512;
  assign n17217 = ~n17215 & ~n17216;
  assign n17218 = pi1012 & n11521;
  assign n17219 = pi1762 & n11529;
  assign n17220 = ~n17218 & ~n17219;
  assign n17221 = pi1128 & n11535;
  assign n17222 = n17220 & ~n17221;
  assign n17223 = pi1133 & n11519;
  assign n17224 = pi1970 & n5423;
  assign n17225 = ~n17223 & ~n17224;
  assign n17226 = n17222 & n17225;
  assign n17227 = n11517 & ~n17226;
  assign n17228 = pi2029 & n11515;
  assign n17229 = ~n17227 & ~n17228;
  assign po1939 = ~n17217 | ~n17229;
  assign n17231 = pi2106 & n11507;
  assign n17232 = pi2066 & n11512;
  assign n17233 = ~n17231 & ~n17232;
  assign n17234 = pi1143 & n11521;
  assign n17235 = pi1174 & n11529;
  assign n17236 = ~n17234 & ~n17235;
  assign n17237 = pi1155 & n11535;
  assign n17238 = n17236 & ~n17237;
  assign n17239 = pi1200 & n11519;
  assign n17240 = pi1946 & n5423;
  assign n17241 = ~n17239 & ~n17240;
  assign n17242 = n17238 & n17241;
  assign n17243 = n11517 & ~n17242;
  assign n17244 = pi2028 & n11515;
  assign n17245 = ~n17243 & ~n17244;
  assign po1940 = ~n17233 | ~n17245;
  assign n17247 = pi2099 & n11507;
  assign n17248 = pi2072 & n11515;
  assign n17249 = ~n17247 & ~n17248;
  assign n17250 = pi1139 & n11521;
  assign n17251 = pi1150 & n11535;
  assign n17252 = pi1169 & n11529;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = ~n17250 & n17253;
  assign n17255 = pi1194 & n11519;
  assign n17256 = pi1967 & n5423;
  assign n17257 = ~n17255 & ~n17256;
  assign n17258 = n17254 & n17257;
  assign n17259 = n11517 & ~n17258;
  assign n17260 = pi2071 & n11512;
  assign n17261 = ~n17259 & ~n17260;
  assign po1941 = ~n17249 | ~n17261;
  assign n17263 = pi2105 & n11507;
  assign n17264 = pi2027 & n11515;
  assign n17265 = ~n17263 & ~n17264;
  assign n17266 = pi1142 & n11521;
  assign n17267 = pi1173 & n11529;
  assign n17268 = ~n17266 & ~n17267;
  assign n17269 = pi1154 & n11535;
  assign n17270 = n17268 & ~n17269;
  assign n17271 = pi1199 & n11519;
  assign n17272 = pi0842 & n5423;
  assign n17273 = ~n17271 & ~n17272;
  assign n17274 = n17270 & n17273;
  assign n17275 = n11517 & ~n17274;
  assign n17276 = pi2065 & n11512;
  assign n17277 = ~n17275 & ~n17276;
  assign po1942 = ~n17265 | ~n17277;
  assign n17279 = pi2102 & n11507;
  assign n17280 = pi2064 & n11512;
  assign n17281 = ~n17279 & ~n17280;
  assign n17282 = pi1141 & n11521;
  assign n17283 = pi1138 & n11535;
  assign n17284 = pi1789 & n11529;
  assign n17285 = ~n17283 & ~n17284;
  assign n17286 = ~n17282 & n17285;
  assign n17287 = pi1197 & n11519;
  assign n17288 = pi1969 & n5423;
  assign n17289 = ~n17287 & ~n17288;
  assign n17290 = n17286 & n17289;
  assign n17291 = n11517 & ~n17290;
  assign n17292 = pi2025 & n11515;
  assign n17293 = ~n17291 & ~n17292;
  assign po1943 = ~n17281 | ~n17293;
  assign n17295 = pi2100 & n11507;
  assign n17296 = pi2126 & n11512;
  assign n17297 = ~n17295 & ~n17296;
  assign n17298 = pi1140 & n11521;
  assign n17299 = pi1170 & n11529;
  assign n17300 = ~n17298 & ~n17299;
  assign n17301 = pi1151 & n11535;
  assign n17302 = n17300 & ~n17301;
  assign n17303 = pi1195 & n11519;
  assign n17304 = pi0249 & n5423;
  assign n17305 = ~n17303 & ~n17304;
  assign n17306 = n17302 & n17305;
  assign n17307 = n11517 & ~n17306;
  assign n17308 = pi2023 & n11515;
  assign n17309 = ~n17307 & ~n17308;
  assign po1944 = ~n17297 | ~n17309;
  assign n17311 = pi1971 & n5423;
  assign n17312 = pi1202 & n11519;
  assign n17313 = pi1176 & n11529;
  assign n17314 = ~n17312 & ~n17313;
  assign n17315 = ~n17311 & n17314;
  assign n17316 = n11517 & ~n17315;
  assign n17317 = pi2069 & n11512;
  assign n17318 = ~n17316 & ~n17317;
  assign n17319 = pi2109 & n11507;
  assign n17320 = pi2088 & n11515;
  assign n17321 = ~n17319 & ~n17320;
  assign po1945 = ~n17318 | ~n17321;
  assign n17323 = pi1181 & n11529;
  assign n17324 = n11517 & n17323;
  assign n17325 = pi2048 & n11515;
  assign n17326 = ~n17324 & ~n17325;
  assign n17327 = pi2116 & n11507;
  assign n17328 = pi2078 & n11512;
  assign n17329 = ~n17327 & ~n17328;
  assign po1946 = ~n17326 | ~n17329;
  assign n17331 = pi1973 & n5423;
  assign n17332 = pi1205 & n11519;
  assign n17333 = pi1179 & n11529;
  assign n17334 = ~n17332 & ~n17333;
  assign n17335 = ~n17331 & n17334;
  assign n17336 = n11517 & ~n17335;
  assign n17337 = pi2045 & n11515;
  assign n17338 = ~n17336 & ~n17337;
  assign n17339 = pi2113 & n11507;
  assign n17340 = pi2075 & n11512;
  assign n17341 = ~n17339 & ~n17340;
  assign po1947 = ~n17338 | ~n17341;
  assign n17343 = pi1949 & n5423;
  assign n17344 = pi1204 & n11519;
  assign n17345 = pi1178 & n11529;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = ~n17343 & n17346;
  assign n17348 = n11517 & ~n17347;
  assign n17349 = pi2044 & n11515;
  assign n17350 = ~n17348 & ~n17349;
  assign n17351 = pi2112 & n11507;
  assign n17352 = pi2074 & n11512;
  assign n17353 = ~n17351 & ~n17352;
  assign po1948 = ~n17350 | ~n17353;
  assign n17355 = pi0815 & n5423;
  assign n17356 = pi1760 & n11519;
  assign n17357 = pi1777 & n11529;
  assign n17358 = ~n17356 & ~n17357;
  assign n17359 = ~n17355 & n17358;
  assign n17360 = n11517 & ~n17359;
  assign n17361 = pi2089 & n11515;
  assign n17362 = ~n17360 & ~n17361;
  assign n17363 = pi2111 & n11507;
  assign n17364 = pi2073 & n11512;
  assign n17365 = ~n17363 & ~n17364;
  assign po1949 = ~n17362 | ~n17365;
  assign n17367 = pi1180 & n11529;
  assign n17368 = n11517 & n17367;
  assign n17369 = pi2046 & n11515;
  assign n17370 = ~n17368 & ~n17369;
  assign n17371 = pi2114 & n11507;
  assign n17372 = pi2076 & n11512;
  assign n17373 = ~n17371 & ~n17372;
  assign po1950 = ~n17370 | ~n17373;
  assign n17375 = pi1972 & n5423;
  assign n17376 = pi1203 & n11519;
  assign n17377 = pi1177 & n11529;
  assign n17378 = ~n17376 & ~n17377;
  assign n17379 = ~n17375 & n17378;
  assign n17380 = n11517 & ~n17379;
  assign n17381 = pi2070 & n11512;
  assign n17382 = ~n17380 & ~n17381;
  assign n17383 = pi2110 & n11507;
  assign n17384 = pi2043 & n11515;
  assign n17385 = ~n17383 & ~n17384;
  assign po1951 = ~n17382 | ~n17385;
  assign n17387 = pi1942 & ~pi2058;
  assign n17388 = pi1901 & pi2058;
  assign po1952 = n17387 | n17388;
  assign n17390 = pi2101 & n11507;
  assign n17391 = pi2063 & n11512;
  assign n17392 = ~n17390 & ~n17391;
  assign n17393 = pi1771 & n11521;
  assign n17394 = pi1152 & n11535;
  assign n17395 = pi1171 & n11529;
  assign n17396 = ~n17394 & ~n17395;
  assign n17397 = ~n17393 & n17396;
  assign n17398 = pi1196 & n11519;
  assign n17399 = pi1968 & n5423;
  assign n17400 = ~n17398 & ~n17399;
  assign n17401 = n17397 & n17400;
  assign n17402 = n11517 & ~n17401;
  assign n17403 = pi2024 & n11515;
  assign n17404 = ~n17402 & ~n17403;
  assign po1953 = ~n17392 | ~n17404;
  assign n17406 = pi0353 & n5197;
  assign n17407 = pi0942 & ~n5210;
  assign n17408 = ~pi0942 & n5210;
  assign n17409 = ~n17407 & ~n17408;
  assign n17410 = ~pi0945 & n5460;
  assign n17411 = pi0945 & ~n5460;
  assign n17412 = ~n17410 & ~n17411;
  assign n17413 = ~n17409 & ~n17412;
  assign n17414 = ~n17406 & n17413;
  assign n17415 = pi0919 & n5446;
  assign n17416 = ~pi0919 & ~n5446;
  assign n17417 = ~n17415 & ~n17416;
  assign po1954 = n17414 & n17417;
  assign n17419 = pi0262 & n5273;
  assign n17420 = pi0943 & ~n5286;
  assign n17421 = ~pi0943 & n5286;
  assign n17422 = ~n17420 & ~n17421;
  assign n17423 = ~pi0931 & n5353;
  assign n17424 = pi0931 & ~n5353;
  assign n17425 = ~n17423 & ~n17424;
  assign n17426 = ~n17422 & ~n17425;
  assign n17427 = ~n17419 & n17426;
  assign n17428 = pi0921 & n5409;
  assign n17429 = ~pi0921 & ~n5409;
  assign n17430 = ~n17428 & ~n17429;
  assign po1955 = n17427 & n17430;
  assign n17432 = pi0941 & ~n5267;
  assign n17433 = ~pi0941 & n5267;
  assign n17434 = ~n17432 & ~n17433;
  assign n17435 = ~pi0935 & n5337;
  assign n17436 = pi0935 & ~n5337;
  assign n17437 = ~n17435 & ~n17436;
  assign n17438 = ~n17434 & ~n17437;
  assign n17439 = ~n6573 & n17438;
  assign n17440 = pi0918 & n5385;
  assign n17441 = ~pi0918 & ~n5385;
  assign n17442 = ~n17440 & ~n17441;
  assign po1958 = n17439 & n17442;
  assign n17444 = pi0354 & n5216;
  assign n17445 = pi0930 & ~n5229;
  assign n17446 = ~pi0930 & n5229;
  assign n17447 = ~n17445 & ~n17446;
  assign n17448 = ~pi0936 & n5486;
  assign n17449 = pi0936 & ~n5486;
  assign n17450 = ~n17448 & ~n17449;
  assign n17451 = ~n17447 & ~n17450;
  assign n17452 = ~n17444 & n17451;
  assign n17453 = pi0920 & n5472;
  assign n17454 = ~pi0920 & ~n5472;
  assign n17455 = ~n17453 & ~n17454;
  assign po1959 = n17452 & n17455;
  assign n17457 = pi0922 & n5399;
  assign n17458 = ~pi0922 & ~n5399;
  assign n17459 = ~n17457 & ~n17458;
  assign n17460 = pi0944 & ~n5305;
  assign n17461 = ~pi0944 & n5305;
  assign n17462 = ~n17460 & ~n17461;
  assign n17463 = ~pi0937 & n5369;
  assign n17464 = pi0937 & ~n5369;
  assign n17465 = ~n17463 & ~n17464;
  assign n17466 = ~n17462 & ~n17465;
  assign n17467 = ~n6320 & n17466;
  assign po1960 = n17459 & n17467;
  assign n17469 = pi0260 & n5235;
  assign n17470 = pi0940 & ~n5248;
  assign n17471 = ~pi0940 & n5248;
  assign n17472 = ~n17470 & ~n17471;
  assign n17473 = ~pi0934 & n5321;
  assign n17474 = pi0934 & ~n5321;
  assign n17475 = ~n17473 & ~n17474;
  assign n17476 = ~n17472 & ~n17475;
  assign n17477 = ~n17469 & n17476;
  assign n17478 = pi0917 & n5379;
  assign n17479 = ~pi0917 & ~n5379;
  assign n17480 = ~n17478 & ~n17479;
  assign po1961 = n17477 & n17480;
  assign n17482 = pi1917 & pi1921;
  assign n17483 = pi1911 & n17482;
  assign n17484 = ~pi1911 & ~n17482;
  assign n17485 = ~n17483 & ~n17484;
  assign n17486 = ~pi2031 & n17485;
  assign n17487 = pi1911 & pi2031;
  assign n17488 = ~n17486 & ~n17487;
  assign po1962 = pi1036 & ~n17488;
  assign n17490 = pi1915 & pi1918;
  assign n17491 = pi1912 & n17490;
  assign n17492 = ~pi1912 & ~n17490;
  assign n17493 = ~n17491 & ~n17492;
  assign n17494 = ~pi2034 & n17493;
  assign n17495 = pi1912 & pi2034;
  assign n17496 = ~n17494 & ~n17495;
  assign po1963 = pi1150 & ~n17496;
  assign n17498 = ~pi2010 & ~pi2036;
  assign po1964 = pi1913 | n17498;
  assign n17500 = ~pi2009 & ~pi2031;
  assign po1965 = pi1914 | n17500;
  assign n17502 = ~pi1915 & pi1918;
  assign n17503 = pi1915 & ~pi1918;
  assign n17504 = ~n17502 & ~n17503;
  assign n17505 = ~pi2034 & ~n17504;
  assign n17506 = pi1915 & pi2034;
  assign n17507 = ~n17505 & ~n17506;
  assign po1966 = pi1150 & ~n17507;
  assign n17509 = ~pi1916 & pi1919;
  assign n17510 = pi1916 & ~pi1919;
  assign n17511 = ~n17509 & ~n17510;
  assign n17512 = ~pi2036 & ~n17511;
  assign n17513 = pi1916 & pi2036;
  assign n17514 = ~n17512 & ~n17513;
  assign po1967 = pi1145 & ~n17514;
  assign n17516 = pi1917 & ~pi1921;
  assign n17517 = ~pi1917 & pi1921;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = ~pi2031 & ~n17518;
  assign n17520 = pi1917 & pi2031;
  assign n17521 = ~n17519 & ~n17520;
  assign po1968 = pi1036 & ~n17521;
  assign n17523 = ~pi1918 & ~pi2034;
  assign n17524 = pi1918 & pi2034;
  assign n17525 = ~n17523 & ~n17524;
  assign po1969 = pi1150 & ~n17525;
  assign n17527 = ~pi1919 & ~pi2036;
  assign n17528 = pi1919 & pi2036;
  assign n17529 = ~n17527 & ~n17528;
  assign po1970 = pi1145 & ~n17529;
  assign n17531 = pi1916 & pi1919;
  assign n17532 = pi1920 & n17531;
  assign n17533 = ~pi1920 & ~n17531;
  assign n17534 = ~n17532 & ~n17533;
  assign n17535 = ~pi2036 & n17534;
  assign n17536 = pi1920 & pi2036;
  assign n17537 = ~n17535 & ~n17536;
  assign po1971 = pi1145 & ~n17537;
  assign n17539 = ~pi1921 & ~pi2031;
  assign n17540 = pi1921 & pi2031;
  assign n17541 = ~n17539 & ~n17540;
  assign po1972 = pi1036 & ~n17541;
  assign n17543 = pi1992 & ~pi2035;
  assign n17544 = pi1922 & pi2035;
  assign po1973 = n17543 | n17544;
  assign n17546 = pi1992 & ~pi2056;
  assign n17547 = pi1923 & pi2056;
  assign po1974 = n17546 | n17547;
  assign n17549 = pi1992 & ~pi2057;
  assign n17550 = pi1924 & pi2057;
  assign po1975 = n17549 | n17550;
  assign n17552 = pi1992 & ~pi2059;
  assign n17553 = pi1925 & pi2059;
  assign po1976 = n17552 | n17553;
  assign n17555 = pi1992 & ~pi2058;
  assign n17556 = pi1926 & pi2058;
  assign po1977 = n17555 | n17556;
  assign n17558 = ~pi2018 & ~pi2034;
  assign po1978 = pi1927 | n17558;
  assign po1980 = ~pi0257 & ~pi2032;
  assign n17561 = pi2014 & ~pi2056;
  assign n17562 = pi1932 & pi2056;
  assign po1983 = n17561 | n17562;
  assign n17564 = pi2014 & ~pi2059;
  assign n17565 = pi1933 & pi2059;
  assign po1984 = n17564 | n17565;
  assign n17567 = pi2014 & ~pi2057;
  assign n17568 = pi1934 & pi2057;
  assign po1985 = n17567 | n17568;
  assign n17570 = pi2014 & ~pi2058;
  assign n17571 = pi1935 & pi2058;
  assign po1986 = n17570 | n17571;
  assign n17573 = pi2201 & pi2203;
  assign n17574 = pi2202 & n17573;
  assign n17575 = pi2162 & n17574;
  assign n17576 = pi2013 & n17575;
  assign n17577 = ~pi2242 & n17576;
  assign n17578 = n11534 & n17577;
  assign n17579 = ~pi2240 & pi2241;
  assign po1987 = n17578 & n17579;
  assign n17581 = pi2241 & n17577;
  assign po1988 = n11505 & n17581;
  assign n17583 = n11518 & n17577;
  assign po1989 = n17579 & n17583;
  assign po1990 = n11532 & n17581;
  assign po1991 = n11521 & n17581;
  assign n17587 = pi2240 & pi2241;
  assign po1992 = n17583 & n17587;
  assign n17589 = pi1944 & ~pi1955;
  assign n17590 = ~pi1996 & n17589;
  assign n17591 = ~pi1957 & n17590;
  assign n17592 = ~pi1986 & n17591;
  assign po2185 = pi1995 & n17592;
  assign n17594 = pi1944 & po2185;
  assign n17595 = pi1995 & pi1996;
  assign n17596 = pi1955 & pi1986;
  assign n17597 = n17595 & n17596;
  assign n17598 = pi1957 & n17597;
  assign n17599 = pi1944 & ~n17598;
  assign n17600 = ~pi1944 & n17598;
  assign n17601 = ~n17599 & ~n17600;
  assign n17602 = ~po2185 & ~n17601;
  assign n17603 = ~n17594 & ~n17602;
  assign po1995 = ~pi2133 & ~n17603;
  assign n17605 = pi1200 & pi1946;
  assign n17606 = pi1133 & pi1970;
  assign n17607 = ~n17605 & ~n17606;
  assign n17608 = pi1203 & pi1972;
  assign n17609 = pi0815 & pi1760;
  assign n17610 = ~n17608 & ~n17609;
  assign n17611 = pi1132 & pi1976;
  assign n17612 = pi0251 & pi1690;
  assign n17613 = ~n17611 & ~n17612;
  assign n17614 = pi0230 & pi1207;
  assign n17615 = pi1208 & pi1977;
  assign n17616 = ~n17614 & ~n17615;
  assign n17617 = pi0810 & pi1198;
  assign n17618 = pi1779 & pi1974;
  assign n17619 = ~n17617 & ~n17618;
  assign n17620 = pi0250 & pi1206;
  assign n17621 = pi1210 & pi1975;
  assign n17622 = ~n17620 & ~n17621;
  assign n17623 = n17619 & n17622;
  assign n17624 = n17616 & n17623;
  assign n17625 = n17613 & n17624;
  assign n17626 = pi0229 & pi1190;
  assign n17627 = pi1191 & pi1965;
  assign n17628 = ~n17626 & ~n17627;
  assign n17629 = pi1189 & pi1964;
  assign n17630 = pi1209 & pi1982;
  assign n17631 = ~n17629 & ~n17630;
  assign n17632 = pi0248 & pi1193;
  assign n17633 = pi1194 & pi1967;
  assign n17634 = ~n17632 & ~n17633;
  assign n17635 = pi1192 & pi1966;
  assign n17636 = pi1211 & pi1950;
  assign n17637 = ~n17635 & ~n17636;
  assign n17638 = n17634 & n17637;
  assign n17639 = n17631 & n17638;
  assign n17640 = n17628 & n17639;
  assign n17641 = n17625 & n17640;
  assign n17642 = pi1204 & pi1949;
  assign n17643 = pi1205 & pi1973;
  assign n17644 = ~n17642 & ~n17643;
  assign n17645 = n17641 & n17644;
  assign n17646 = n17610 & n17645;
  assign n17647 = pi1197 & pi1969;
  assign n17648 = pi0842 & pi1199;
  assign n17649 = ~n17647 & ~n17648;
  assign n17650 = pi0249 & pi1195;
  assign n17651 = pi1196 & pi1968;
  assign n17652 = ~n17650 & ~n17651;
  assign n17653 = pi1188 & pi1948;
  assign n17654 = n17652 & ~n17653;
  assign n17655 = n17649 & n17654;
  assign n17656 = n17646 & n17655;
  assign n17657 = pi0841 & pi1201;
  assign n17658 = pi1202 & pi1971;
  assign n17659 = ~n17657 & ~n17658;
  assign n17660 = n17656 & n17659;
  assign po1996 = ~n17607 | ~n17660;
  assign n17662 = ~pi1913 & ~pi1946;
  assign po1997 = ~n5425 & ~n17662;
  assign n17664 = ~pi2059 & pi2164;
  assign n17665 = pi1947 & pi2059;
  assign po1998 = n17664 | n17665;
  assign n17667 = ~pi0873 & ~pi1948;
  assign po1999 = ~n5425 & ~n17667;
  assign n17669 = ~pi1927 & ~pi1949;
  assign po2000 = ~n5425 & ~n17669;
  assign n17671 = pi0452 & ~pi1950;
  assign po2001 = ~n5425 & ~n17671;
  assign n17673 = pi1985 & pi1999;
  assign n17674 = pi2000 & n17673;
  assign n17675 = pi1994 & n17674;
  assign n17676 = pi1997 & n17675;
  assign n17677 = pi1998 & n17676;
  assign n17678 = pi1993 & n17677;
  assign n17679 = pi1951 & n17678;
  assign n17680 = ~pi1951 & ~n17678;
  assign n17681 = ~n17679 & ~n17680;
  assign po2002 = pi2134 | n17681;
  assign n17683 = pi1955 & po2185;
  assign n17684 = pi1986 & n17595;
  assign n17685 = pi1955 & ~n17684;
  assign n17686 = ~pi1955 & n17684;
  assign n17687 = ~n17685 & ~n17686;
  assign n17688 = ~po2185 & ~n17687;
  assign n17689 = ~n17683 & ~n17688;
  assign po2006 = ~pi2133 & ~n17689;
  assign n17691 = pi1990 & pi2003;
  assign n17692 = pi2001 & n17691;
  assign n17693 = pi1956 & ~n17692;
  assign n17694 = ~pi1956 & n17692;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = n11481 & ~n17695;
  assign n17697 = pi1956 & ~n11481;
  assign n17698 = ~n17696 & ~n17697;
  assign po2007 = pi0880 & ~n17698;
  assign n17700 = pi1957 & po2185;
  assign n17701 = pi1957 & ~n17597;
  assign n17702 = ~pi1957 & n17597;
  assign n17703 = ~n17701 & ~n17702;
  assign n17704 = ~po2185 & ~n17703;
  assign n17705 = ~n17700 & ~n17704;
  assign po2008 = ~pi2133 & ~n17705;
  assign n17707 = ~pi2059 & pi2142;
  assign n17708 = pi1958 & pi2059;
  assign po2009 = n17707 | n17708;
  assign n17710 = ~pi2059 & pi2161;
  assign n17711 = pi1959 & pi2059;
  assign po2010 = n17710 | n17711;
  assign n17713 = ~pi2057 & pi2161;
  assign n17714 = pi1960 & pi2057;
  assign po2011 = n17713 | n17714;
  assign n17716 = ~pi2058 & pi2161;
  assign n17717 = pi1961 & pi2058;
  assign po2012 = n17716 | n17717;
  assign n17719 = ~pi2058 & pi2142;
  assign n17720 = pi1962 & pi2058;
  assign po2013 = n17719 | n17720;
  assign n17722 = ~n5417 & ~n17576;
  assign n17723 = pi2202 & ~n17722;
  assign n17724 = ~pi1963 & n17723;
  assign po2014 = pi2203 & n17724;
  assign n17726 = pi0905 & ~pi1964;
  assign po2015 = ~n5425 & ~n17726;
  assign n17728 = pi0451 & ~pi1965;
  assign po2016 = ~n5425 & ~n17728;
  assign n17730 = pi0902 & ~pi1966;
  assign po2017 = ~n5425 & ~n17730;
  assign n17732 = pi0901 & ~pi1967;
  assign po2018 = ~n5425 & ~n17732;
  assign n17734 = pi0453 & ~pi1968;
  assign po2019 = ~n5425 & ~n17734;
  assign n17736 = pi0904 & ~pi1969;
  assign po2020 = ~n5425 & ~n17736;
  assign n17738 = pi0872 & ~pi1970;
  assign po2021 = ~n5425 & ~n17738;
  assign n17740 = ~pi1914 & ~pi1971;
  assign po2022 = ~n5425 & ~n17740;
  assign n17742 = pi0808 & ~pi1972;
  assign po2023 = ~n5425 & ~n17742;
  assign n17744 = pi0636 & ~pi1973;
  assign po2024 = ~n5425 & ~n17744;
  assign n17746 = pi0450 & ~pi1974;
  assign po2025 = ~n5425 & ~n17746;
  assign n17748 = pi0899 & ~pi1975;
  assign po2026 = ~n5425 & ~n17748;
  assign n17750 = pi0900 & ~pi1976;
  assign po2027 = ~n5425 & ~n17750;
  assign n17752 = pi0806 & ~pi1977;
  assign po2028 = ~n5425 & ~n17752;
  assign n17754 = ~pi2058 & pi2081;
  assign n17755 = pi1978 & pi2058;
  assign po2029 = n17754 | n17755;
  assign n17757 = ~pi2058 & pi2164;
  assign n17758 = pi1979 & pi2058;
  assign po2030 = n17757 | n17758;
  assign n17760 = ~pi2057 & pi2081;
  assign n17761 = pi1980 & pi2057;
  assign po2031 = n17760 | n17761;
  assign n17763 = ~pi2059 & pi2081;
  assign n17764 = pi1981 & pi2059;
  assign po2032 = n17763 | n17764;
  assign n17766 = pi0807 & ~pi1982;
  assign po2033 = ~n5425 & ~n17766;
  assign n17768 = ~pi2057 & pi2142;
  assign n17769 = pi1983 & pi2057;
  assign po2034 = n17768 | n17769;
  assign n17771 = ~pi2057 & pi2164;
  assign n17772 = pi1984 & pi2057;
  assign po2035 = n17771 | n17772;
  assign n17774 = ~pi1985 & pi1999;
  assign n17775 = pi1985 & ~pi1999;
  assign n17776 = ~n17774 & ~n17775;
  assign po2036 = pi2134 | ~n17776;
  assign n17778 = pi1986 & po2185;
  assign n17779 = pi1986 & ~n17595;
  assign n17780 = ~pi1986 & n17595;
  assign n17781 = ~n17779 & ~n17780;
  assign n17782 = ~po2185 & ~n17781;
  assign n17783 = ~n17778 & ~n17782;
  assign po2037 = ~pi2133 & ~n17783;
  assign n17785 = pi0236 & ~pi0919;
  assign n17786 = ~pi0214 & pi0942;
  assign n17787 = pi0214 & ~pi0942;
  assign n17788 = ~n17786 & ~n17787;
  assign n17789 = n17785 & n17788;
  assign n17790 = ~n17785 & ~n17788;
  assign n17791 = ~n17789 & ~n17790;
  assign n17792 = po2191 & n17791;
  assign n17793 = ~po2191 & ~n17791;
  assign po2038 = n17792 | n17793;
  assign n17795 = pi0238 & ~pi0920;
  assign n17796 = ~pi0215 & pi0930;
  assign n17797 = pi0215 & ~pi0930;
  assign n17798 = ~n17796 & ~n17797;
  assign n17799 = n17795 & n17798;
  assign n17800 = ~n17795 & ~n17798;
  assign n17801 = ~n17799 & ~n17800;
  assign n17802 = po2209 & n17801;
  assign n17803 = ~po2209 & ~n17801;
  assign po2039 = n17802 | n17803;
  assign n17805 = ~pi2241 & n17576;
  assign po2040 = n5420 & n17805;
  assign n17807 = pi1990 & ~n11481;
  assign n17808 = ~pi1990 & n11481;
  assign n17809 = ~n17807 & ~n17808;
  assign po2041 = pi0880 & ~n17809;
  assign n17811 = pi1993 & n17675;
  assign n17812 = ~pi1993 & ~n17675;
  assign n17813 = ~n17811 & ~n17812;
  assign po2044 = pi2134 | n17813;
  assign n17815 = ~pi1994 & ~n17674;
  assign n17816 = ~n17675 & ~n17815;
  assign po2045 = pi2134 | n17816;
  assign n17818 = pi1995 & ~po2185;
  assign n17819 = ~pi1995 & po2185;
  assign n17820 = ~n17818 & ~n17819;
  assign po2046 = ~pi2133 & n17820;
  assign n17822 = pi1996 & po2185;
  assign n17823 = pi1995 & ~pi1996;
  assign n17824 = ~pi1995 & pi1996;
  assign n17825 = ~n17823 & ~n17824;
  assign n17826 = ~po2185 & ~n17825;
  assign n17827 = ~n17822 & ~n17826;
  assign po2047 = ~pi2133 & ~n17827;
  assign n17829 = pi1994 & pi2000;
  assign n17830 = pi1985 & n17829;
  assign n17831 = pi1999 & n17830;
  assign n17832 = pi1993 & n17831;
  assign n17833 = pi1997 & n17832;
  assign n17834 = ~pi1997 & ~n17832;
  assign n17835 = ~n17833 & ~n17834;
  assign po2048 = pi2134 | n17835;
  assign n17837 = n17673 & n17829;
  assign n17838 = pi1993 & n17837;
  assign n17839 = pi1997 & n17838;
  assign n17840 = ~pi1998 & n17839;
  assign n17841 = pi1998 & ~n17839;
  assign n17842 = ~n17840 & ~n17841;
  assign po2049 = pi2134 | ~n17842;
  assign po2050 = ~pi1999 | pi2134;
  assign n17845 = ~pi2000 & ~n17673;
  assign n17846 = ~n17674 & ~n17845;
  assign po2051 = pi2134 | n17846;
  assign n17848 = pi2001 & ~n17691;
  assign n17849 = ~pi2001 & n17691;
  assign n17850 = ~n17848 & ~n17849;
  assign n17851 = n11481 & ~n17850;
  assign n17852 = pi2001 & ~n11481;
  assign n17853 = ~n17851 & ~n17852;
  assign po2052 = pi0880 & ~n17853;
  assign n17855 = ~pi1951 & ~pi1998;
  assign n17856 = ~pi1997 & n17855;
  assign n17857 = ~pi1985 & ~pi2000;
  assign n17858 = pi1994 & ~n17857;
  assign n17859 = pi1993 & n17858;
  assign n17860 = n17855 & ~n17859;
  assign po2053 = ~n17856 & ~n17860;
  assign n17862 = ~pi1990 & pi2003;
  assign n17863 = pi1990 & ~pi2003;
  assign n17864 = ~n17862 & ~n17863;
  assign n17865 = n11481 & ~n17864;
  assign n17866 = pi2003 & ~n11481;
  assign n17867 = ~n17865 & ~n17866;
  assign po2054 = pi0880 & ~n17867;
  assign n17869 = pi0225 & ~pi0918;
  assign n17870 = ~pi0217 & pi0941;
  assign n17871 = pi0217 & ~pi0941;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = n17869 & n17872;
  assign n17874 = ~n17869 & ~n17872;
  assign n17875 = ~n17873 & ~n17874;
  assign n17876 = po2190 & n17875;
  assign n17877 = ~po2190 & ~n17875;
  assign po2055 = n17876 | n17877;
  assign n17879 = pi0227 & ~pi0921;
  assign n17880 = ~pi0218 & pi0943;
  assign n17881 = pi0218 & ~pi0943;
  assign n17882 = ~n17880 & ~n17881;
  assign n17883 = n17879 & n17882;
  assign n17884 = ~n17879 & ~n17882;
  assign n17885 = ~n17883 & ~n17884;
  assign n17886 = po2189 & n17885;
  assign n17887 = ~po2189 & ~n17885;
  assign po2056 = n17886 | n17887;
  assign n17889 = pi0226 & ~pi0922;
  assign n17890 = ~pi0219 & pi0944;
  assign n17891 = pi0219 & ~pi0944;
  assign n17892 = ~n17890 & ~n17891;
  assign n17893 = n17889 & n17892;
  assign n17894 = ~n17889 & ~n17892;
  assign n17895 = ~n17893 & ~n17894;
  assign n17896 = po2192 & n17895;
  assign n17897 = ~po2192 & ~n17895;
  assign po2057 = n17896 | n17897;
  assign n17899 = pi0224 & ~pi0917;
  assign n17900 = ~pi0216 & pi0940;
  assign n17901 = pi0216 & ~pi0940;
  assign n17902 = ~n17900 & ~n17901;
  assign n17903 = n17899 & n17902;
  assign n17904 = ~n17899 & ~n17902;
  assign n17905 = ~n17903 & ~n17904;
  assign n17906 = po2210 & n17905;
  assign n17907 = ~po2210 & ~n17905;
  assign po2058 = n17906 | n17907;
  assign n17909 = ~pi0411 & ~pi1918;
  assign n17910 = pi0411 & pi1918;
  assign po2188 = n17909 | n17910;
  assign n17912 = pi0411 & ~pi1918;
  assign n17913 = ~pi0412 & pi1915;
  assign n17914 = pi0412 & ~pi1915;
  assign n17915 = ~n17913 & ~n17914;
  assign n17916 = ~n17912 & n17915;
  assign n17917 = n17912 & ~n17915;
  assign n17918 = ~n17916 & ~n17917;
  assign n17919 = ~po2188 & n17918;
  assign n17920 = po2188 & ~n17918;
  assign po2059 = n17919 | n17920;
  assign n17922 = ~pi0601 & ~pi1921;
  assign n17923 = pi0601 & pi1921;
  assign po2186 = n17922 | n17923;
  assign n17925 = pi0602 & pi1917;
  assign n17926 = ~pi0602 & ~pi1917;
  assign n17927 = ~n17925 & ~n17926;
  assign n17928 = po2186 & ~n17927;
  assign n17929 = ~pi0463 & ~pi1911;
  assign n17930 = pi0463 & pi1911;
  assign n17931 = ~n17929 & ~n17930;
  assign n17932 = n8807 & ~n17931;
  assign po2060 = n17928 & n17932;
  assign n17934 = ~pi0843 & ~pi1919;
  assign n17935 = pi0843 & pi1919;
  assign po2187 = n17934 | n17935;
  assign n17937 = pi0746 & pi1916;
  assign n17938 = ~pi0746 & ~pi1916;
  assign n17939 = ~n17937 & ~n17938;
  assign n17940 = po2187 & ~n17939;
  assign n17941 = ~pi0643 & ~pi1920;
  assign n17942 = pi0643 & pi1920;
  assign n17943 = ~n17941 & ~n17942;
  assign n17944 = n8838 & ~n17943;
  assign po2061 = n17940 & n17944;
  assign n17946 = ~pi1993 & ~pi1997;
  assign n17947 = ~n17830 & n17946;
  assign n17948 = pi1998 & ~n17947;
  assign po2063 = pi1951 | n17948;
  assign n17950 = ~pi2243 & ~pi2245;
  assign n17951 = ~pi2244 & n17950;
  assign n17952 = n17574 & n17951;
  assign po2064 = ~n17576 & n17952;
  assign n17954 = ~pi1997 & ~n17858;
  assign n17955 = ~pi1998 & n17954;
  assign n17956 = ~pi1993 & n17955;
  assign po2066 = pi1951 & ~n17956;
  assign n17958 = ~pi0602 & pi1917;
  assign n17959 = pi0602 & ~pi1917;
  assign n17960 = ~n17958 & ~n17959;
  assign n17961 = pi0601 & ~pi1921;
  assign n17962 = ~n17960 & n17961;
  assign n17963 = n17960 & ~n17961;
  assign n17964 = ~n17962 & ~n17963;
  assign n17965 = po2186 & ~n17964;
  assign n17966 = ~po2186 & n17964;
  assign po2067 = n17965 | n17966;
  assign n17968 = ~pi0746 & pi1916;
  assign n17969 = pi0746 & ~pi1916;
  assign n17970 = ~n17968 & ~n17969;
  assign n17971 = pi0843 & ~pi1919;
  assign n17972 = ~n17970 & n17971;
  assign n17973 = n17970 & ~n17971;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = ~po2187 & n17974;
  assign n17976 = po2187 & ~n17974;
  assign po2068 = n17975 | n17976;
  assign n17978 = pi0412 & pi1915;
  assign n17979 = ~pi0412 & ~pi1915;
  assign n17980 = ~n17978 & ~n17979;
  assign n17981 = po2188 & ~n17980;
  assign n17982 = ~pi0346 & ~pi1912;
  assign n17983 = pi0346 & pi1912;
  assign n17984 = ~n17982 & ~n17983;
  assign n17985 = n7543 & ~n17984;
  assign po2069 = n17981 & n17985;
  assign n17987 = ~pi1985 & ~pi1994;
  assign n17988 = ~pi2000 & n17987;
  assign n17989 = ~pi1999 & n17988;
  assign n17990 = n17946 & ~n17989;
  assign n17991 = n17855 & n17990;
  assign n17992 = ~pi1999 & n17857;
  assign n17993 = ~pi1994 & n17992;
  assign n17994 = ~pi1993 & n17993;
  assign po2083 = n17856 & n17994;
  assign po2070 = n17991 | po2083;
  assign n17997 = ~n17980 & n17984;
  assign po2071 = po2188 & n17997;
  assign n17999 = ~pi0671 & n17516;
  assign n18000 = ~pi0726 & n17482;
  assign n18001 = ~n17999 & ~n18000;
  assign n18002 = ~pi0736 & n17517;
  assign n18003 = ~pi1917 & ~pi1921;
  assign n18004 = ~pi0780 & n18003;
  assign n18005 = ~n18002 & ~n18004;
  assign po2072 = ~n18001 | ~n18005;
  assign n18007 = ~pi0781 & n18003;
  assign n18008 = ~pi0672 & n17516;
  assign n18009 = ~n18007 & ~n18008;
  assign n18010 = ~pi0652 & n17517;
  assign n18011 = ~pi0727 & n17482;
  assign n18012 = ~n18010 & ~n18011;
  assign po2073 = ~n18009 | ~n18012;
  assign n18014 = ~pi0737 & n17517;
  assign n18015 = ~pi0749 & n17516;
  assign n18016 = ~n18014 & ~n18015;
  assign n18017 = ~pi0783 & n18003;
  assign n18018 = ~pi0639 & n17482;
  assign n18019 = ~n18017 & ~n18018;
  assign po2074 = ~n18016 | ~n18019;
  assign n18021 = ~pi0458 & n18003;
  assign n18022 = ~pi0482 & n17516;
  assign n18023 = ~n18021 & ~n18022;
  assign n18024 = ~pi0543 & n17517;
  assign n18025 = ~pi0530 & n17482;
  assign n18026 = ~n18024 & ~n18025;
  assign po2075 = ~n18023 | ~n18026;
  assign n18028 = ~pi0544 & n17517;
  assign n18029 = ~pi0483 & n17516;
  assign n18030 = ~n18028 & ~n18029;
  assign n18031 = ~pi0542 & n18003;
  assign n18032 = ~pi0531 & n17482;
  assign n18033 = ~n18031 & ~n18032;
  assign po2076 = ~n18030 | ~n18033;
  assign n18035 = ~pi0637 & n18003;
  assign n18036 = ~pi0559 & n17516;
  assign n18037 = ~n18035 & ~n18036;
  assign n18038 = ~pi0651 & n17517;
  assign n18039 = ~pi0729 & n17482;
  assign n18040 = ~n18038 & ~n18039;
  assign po2077 = ~n18037 | ~n18040;
  assign n18042 = ~pi0554 & n17517;
  assign n18043 = ~pi0484 & n17516;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = ~pi0811 & n18003;
  assign n18046 = ~pi0532 & n17482;
  assign n18047 = ~n18045 & ~n18046;
  assign po2078 = ~n18044 | ~n18047;
  assign n18049 = ~pi0545 & n17517;
  assign n18050 = ~pi0485 & n17516;
  assign n18051 = ~n18049 & ~n18050;
  assign n18052 = ~pi0614 & n18003;
  assign n18053 = ~pi0533 & n17482;
  assign n18054 = ~n18052 & ~n18053;
  assign po2079 = ~n18051 | ~n18054;
  assign n18056 = ~pi0617 & n18003;
  assign n18057 = ~pi0486 & n17516;
  assign n18058 = ~n18056 & ~n18057;
  assign n18059 = ~pi0546 & n17517;
  assign n18060 = ~pi0534 & n17482;
  assign n18061 = ~n18059 & ~n18060;
  assign po2080 = ~n18058 | ~n18061;
  assign n18063 = ~pi0547 & n17517;
  assign n18064 = ~pi0489 & n17516;
  assign n18065 = ~n18063 & ~n18064;
  assign n18066 = ~pi0656 & n18003;
  assign n18067 = ~pi0535 & n17482;
  assign n18068 = ~n18066 & ~n18067;
  assign po2081 = ~n18065 | ~n18068;
  assign n18070 = n11534 & n17587;
  assign n18071 = ~pi2242 & n5417;
  assign po2082 = n18070 & n18071;
  assign n18073 = ~n17939 & n17943;
  assign po2084 = po2187 & n18073;
  assign n18075 = pi2242 & n5417;
  assign n18076 = ~pi2241 & n5418;
  assign n18077 = ~pi2238 & n18076;
  assign po2085 = n18075 & n18077;
  assign n18079 = pi1997 & pi1999;
  assign n18080 = pi2000 & n18079;
  assign n18081 = n17855 & n18080;
  assign n18082 = ~pi1993 & n18081;
  assign po2086 = n17987 & n18082;
  assign n18084 = pi2241 & n5423;
  assign po2087 = n18071 & n18084;
  assign n18086 = pi1997 & pi1998;
  assign n18087 = ~pi1993 & n17988;
  assign n18088 = n18086 & ~n18087;
  assign po2088 = pi1951 | n18088;
  assign n18090 = ~pi0641 & n18003;
  assign n18091 = ~pi0734 & n17517;
  assign n18092 = ~n18090 & ~n18091;
  assign n18093 = ~pi0668 & n17516;
  assign n18094 = ~pi0724 & n17482;
  assign n18095 = ~n18093 & ~n18094;
  assign po2089 = ~n18092 | ~n18095;
  assign n18097 = ~pi0778 & n18003;
  assign n18098 = ~pi0667 & n17516;
  assign n18099 = ~n18097 & ~n18098;
  assign n18100 = ~pi0475 & n17517;
  assign n18101 = ~pi0660 & n17482;
  assign n18102 = ~n18100 & ~n18101;
  assign po2090 = ~n18099 | ~n18102;
  assign n18104 = ~pi0779 & n18003;
  assign n18105 = ~pi0674 & n17516;
  assign n18106 = ~n18104 & ~n18105;
  assign n18107 = ~pi0654 & n17517;
  assign n18108 = ~pi0723 & n17482;
  assign n18109 = ~n18107 & ~n18108;
  assign po2091 = ~n18106 | ~n18109;
  assign n18111 = ~pi0606 & n18003;
  assign n18112 = ~pi0735 & n17517;
  assign n18113 = ~n18111 & ~n18112;
  assign n18114 = ~pi0669 & n17516;
  assign n18115 = ~pi0725 & n17482;
  assign n18116 = ~n18114 & ~n18115;
  assign po2092 = ~n18113 | ~n18116;
  assign n18118 = ~pi0605 & n18003;
  assign n18119 = ~pi0670 & n17516;
  assign n18120 = ~n18118 & ~n18119;
  assign n18121 = ~pi0653 & n17517;
  assign n18122 = ~pi0659 & n17482;
  assign n18123 = ~n18121 & ~n18122;
  assign po2093 = ~n18120 | ~n18123;
  assign n18125 = ~pi0624 & n18003;
  assign n18126 = ~pi0490 & n17516;
  assign n18127 = ~n18125 & ~n18126;
  assign n18128 = ~pi0549 & n17517;
  assign n18129 = ~pi0536 & n17482;
  assign n18130 = ~n18128 & ~n18129;
  assign po2094 = ~n18127 | ~n18130;
  assign n18132 = ~pi0551 & n17517;
  assign n18133 = ~pi0492 & n17516;
  assign n18134 = ~n18132 & ~n18133;
  assign n18135 = ~pi0627 & n18003;
  assign n18136 = ~pi0538 & n17482;
  assign n18137 = ~n18135 & ~n18136;
  assign po2095 = ~n18134 | ~n18137;
  assign n18139 = ~pi0552 & n17517;
  assign n18140 = ~pi0497 & n17516;
  assign n18141 = ~n18139 & ~n18140;
  assign n18142 = ~pi0629 & n18003;
  assign n18143 = ~pi0459 & n17482;
  assign n18144 = ~n18142 & ~n18143;
  assign po2096 = ~n18141 | ~n18144;
  assign n18146 = ~pi0632 & n18003;
  assign n18147 = ~pi0553 & n17517;
  assign n18148 = ~n18146 & ~n18147;
  assign n18149 = ~pi0501 & n17516;
  assign n18150 = ~pi0539 & n17482;
  assign n18151 = ~n18149 & ~n18150;
  assign po2097 = ~n18148 | ~n18151;
  assign n18153 = ~pi0743 & n17517;
  assign n18154 = ~pi0744 & n17516;
  assign n18155 = ~n18153 & ~n18154;
  assign n18156 = ~pi0603 & n18003;
  assign n18157 = ~pi0567 & n17482;
  assign n18158 = ~n18156 & ~n18157;
  assign po2098 = ~n18155 | ~n18158;
  assign n18160 = ~pi0555 & n17517;
  assign n18161 = ~pi0506 & n17516;
  assign n18162 = ~n18160 & ~n18161;
  assign n18163 = ~pi0786 & n18003;
  assign n18164 = ~pi0540 & n17482;
  assign n18165 = ~n18163 & ~n18164;
  assign po2099 = ~n18162 | ~n18165;
  assign n18167 = ~pi0740 & n17517;
  assign n18168 = ~pi0698 & n17516;
  assign n18169 = ~n18167 & ~n18168;
  assign n18170 = ~pi0785 & n18003;
  assign n18171 = ~pi0562 & n17482;
  assign n18172 = ~n18170 & ~n18171;
  assign po2100 = ~n18169 | ~n18172;
  assign n18174 = ~pi0741 & n17517;
  assign n18175 = ~pi0700 & n17516;
  assign n18176 = ~n18174 & ~n18175;
  assign n18177 = ~pi0753 & n18003;
  assign n18178 = ~pi0730 & n17482;
  assign n18179 = ~n18177 & ~n18178;
  assign po2101 = ~n18176 | ~n18179;
  assign n18181 = ~pi0648 & n17517;
  assign n18182 = ~pi0561 & n17516;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = ~pi0787 & n18003;
  assign n18185 = ~pi0732 & n17482;
  assign n18186 = ~n18184 & ~n18185;
  assign po2102 = ~n18183 | ~n18186;
  assign n18188 = ~pi0745 & n17517;
  assign n18189 = ~pi0714 & n17516;
  assign n18190 = ~n18188 & ~n18189;
  assign n18191 = ~pi0788 & n18003;
  assign n18192 = ~pi0733 & n17482;
  assign n18193 = ~n18191 & ~n18192;
  assign po2103 = ~n18190 | ~n18193;
  assign n18195 = ~pi0752 & n18003;
  assign n18196 = ~pi0720 & n17516;
  assign n18197 = ~n18195 & ~n18196;
  assign n18198 = ~pi0645 & n17517;
  assign n18199 = ~pi0655 & n17482;
  assign n18200 = ~n18198 & ~n18199;
  assign po2104 = ~n18197 | ~n18200;
  assign n18202 = ~pi0789 & n18003;
  assign n18203 = ~pi0666 & n17517;
  assign n18204 = ~n18202 & ~n18203;
  assign n18205 = ~pi0563 & n17516;
  assign n18206 = ~pi0568 & n17482;
  assign n18207 = ~n18205 & ~n18206;
  assign po2105 = ~n18204 | ~n18207;
  assign n18209 = ~n17927 & n17931;
  assign po2106 = po2186 & n18209;
  assign n18211 = pi1993 & n17855;
  assign n18212 = pi1997 & n18211;
  assign n18213 = ~pi2000 & n17774;
  assign n18214 = pi1994 & n18213;
  assign po2107 = n18212 & n18214;
  assign n18216 = ~pi1993 & pi1998;
  assign n18217 = n17774 & n18216;
  assign n18218 = ~pi2000 & n18217;
  assign n18219 = ~pi1994 & pi1997;
  assign n18220 = ~pi1951 & n18219;
  assign po2108 = n18218 & n18220;
  assign n18222 = pi1951 & ~pi1993;
  assign n18223 = ~pi1998 & n18222;
  assign n18224 = n18214 & n18223;
  assign po2109 = ~pi1997 & n18224;
  assign n18226 = pi2000 & n18217;
  assign n18227 = pi1994 & ~pi1997;
  assign n18228 = ~pi1951 & n18227;
  assign po2110 = n18226 & n18228;
  assign n18230 = n17988 & n18211;
  assign n18231 = ~pi1997 & n18230;
  assign po2111 = pi1999 & n18231;
  assign n18233 = ~pi1916 & ~pi1919;
  assign n18234 = ~pi0756 & n18233;
  assign n18235 = ~pi0748 & n17509;
  assign n18236 = ~n18234 & ~n18235;
  assign n18237 = ~pi0692 & n17510;
  assign n18238 = ~pi0707 & n17531;
  assign n18239 = ~n18237 & ~n18238;
  assign po2112 = ~n18236 | ~n18239;
  assign n18241 = ~pi0758 & n18233;
  assign n18242 = ~pi0679 & n17509;
  assign n18243 = ~n18241 & ~n18242;
  assign n18244 = ~pi0693 & n17510;
  assign n18245 = ~pi0710 & n17531;
  assign n18246 = ~n18244 & ~n18245;
  assign po2113 = ~n18243 | ~n18246;
  assign n18248 = ~pi0487 & n18233;
  assign n18249 = ~pi0507 & n17510;
  assign n18250 = ~n18248 & ~n18249;
  assign n18251 = ~pi0493 & n17509;
  assign n18252 = ~pi0519 & n17531;
  assign n18253 = ~n18251 & ~n18252;
  assign po2114 = ~n18250 | ~n18253;
  assign n18255 = ~pi0488 & n18233;
  assign n18256 = ~pi0494 & n17509;
  assign n18257 = ~n18255 & ~n18256;
  assign n18258 = ~pi0508 & n17510;
  assign n18259 = ~pi0520 & n17531;
  assign n18260 = ~n18258 & ~n18259;
  assign po2115 = ~n18257 | ~n18260;
  assign n18262 = ~pi0495 & n17509;
  assign n18263 = ~pi0467 & n17510;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = ~pi0762 & n18233;
  assign n18266 = ~pi0521 & n17531;
  assign n18267 = ~n18265 & ~n18266;
  assign po2116 = ~n18264 | ~n18267;
  assign n18269 = ~pi0763 & n18233;
  assign n18270 = ~pi0496 & n17509;
  assign n18271 = ~n18269 & ~n18270;
  assign n18272 = ~pi0510 & n17510;
  assign n18273 = ~pi0522 & n17531;
  assign n18274 = ~n18272 & ~n18273;
  assign po2117 = ~n18271 | ~n18274;
  assign n18276 = ~pi0764 & n18233;
  assign n18277 = ~pi0470 & n17509;
  assign n18278 = ~n18276 & ~n18277;
  assign n18279 = ~pi0511 & n17510;
  assign n18280 = ~pi0464 & n17531;
  assign n18281 = ~n18279 & ~n18280;
  assign po2118 = ~n18278 | ~n18281;
  assign n18283 = ~pi0765 & n18233;
  assign n18284 = ~pi0512 & n17510;
  assign n18285 = ~n18283 & ~n18284;
  assign n18286 = ~pi0498 & n17509;
  assign n18287 = ~pi0523 & n17531;
  assign n18288 = ~n18286 & ~n18287;
  assign po2119 = ~n18285 | ~n18288;
  assign n18290 = ~pi0766 & n18233;
  assign n18291 = ~pi0499 & n17509;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = ~pi0466 & n17510;
  assign n18294 = ~pi0524 & n17531;
  assign n18295 = ~n18293 & ~n18294;
  assign po2120 = ~n18292 | ~n18295;
  assign n18297 = ~pi0767 & n18233;
  assign n18298 = ~pi0513 & n17510;
  assign n18299 = ~n18297 & ~n18298;
  assign n18300 = ~pi0469 & n17509;
  assign n18301 = ~pi0525 & n17531;
  assign n18302 = ~n18300 & ~n18301;
  assign po2121 = ~n18299 | ~n18302;
  assign n18304 = ~pi0680 & n17509;
  assign n18305 = ~pi0695 & n17510;
  assign n18306 = ~n18304 & ~n18305;
  assign n18307 = ~pi0760 & n18233;
  assign n18308 = ~pi0712 & n17531;
  assign n18309 = ~n18307 & ~n18308;
  assign po2122 = ~n18306 | ~n18309;
  assign n18311 = ~pi0782 & n18003;
  assign n18312 = ~pi0738 & n17517;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = ~pi0673 & n17516;
  assign n18315 = ~pi0728 & n17482;
  assign n18316 = ~n18314 & ~n18315;
  assign po2123 = ~n18313 | ~n18316;
  assign n18318 = ~pi0647 & n18233;
  assign n18319 = ~pi0500 & n17509;
  assign n18320 = ~n18318 & ~n18319;
  assign n18321 = ~pi0514 & n17510;
  assign n18322 = ~pi0462 & n17531;
  assign n18323 = ~n18321 & ~n18322;
  assign po2124 = ~n18320 | ~n18323;
  assign n18325 = ~pi0768 & n18233;
  assign n18326 = ~pi0502 & n17509;
  assign n18327 = ~n18325 & ~n18326;
  assign n18328 = ~pi0515 & n17510;
  assign n18329 = ~pi0526 & n17531;
  assign n18330 = ~n18328 & ~n18329;
  assign po2125 = ~n18327 | ~n18330;
  assign n18332 = ~pi0769 & n18233;
  assign n18333 = ~pi0468 & n17509;
  assign n18334 = ~n18332 & ~n18333;
  assign n18335 = ~pi0465 & n17510;
  assign n18336 = ~pi0527 & n17531;
  assign n18337 = ~n18335 & ~n18336;
  assign po2126 = ~n18334 | ~n18337;
  assign n18339 = ~pi0770 & n18233;
  assign n18340 = ~pi0516 & n17510;
  assign n18341 = ~n18339 & ~n18340;
  assign n18342 = ~pi0503 & n17509;
  assign n18343 = ~pi0528 & n17531;
  assign n18344 = ~n18342 & ~n18343;
  assign po2127 = ~n18341 | ~n18344;
  assign n18346 = ~pi0646 & n18233;
  assign n18347 = ~pi0683 & n17509;
  assign n18348 = ~n18346 & ~n18347;
  assign n18349 = ~pi0665 & n17510;
  assign n18350 = ~pi0715 & n17531;
  assign n18351 = ~n18349 & ~n18350;
  assign po2128 = ~n18348 | ~n18351;
  assign n18353 = ~pi0771 & n18233;
  assign n18354 = ~pi0504 & n17509;
  assign n18355 = ~n18353 & ~n18354;
  assign n18356 = ~pi0517 & n17510;
  assign n18357 = ~pi0461 & n17531;
  assign n18358 = ~n18356 & ~n18357;
  assign po2129 = ~n18355 | ~n18358;
  assign n18360 = ~pi0772 & n18233;
  assign n18361 = ~pi0505 & n17509;
  assign n18362 = ~n18360 & ~n18361;
  assign n18363 = ~pi0518 & n17510;
  assign n18364 = ~pi0529 & n17531;
  assign n18365 = ~n18363 & ~n18364;
  assign po2130 = ~n18362 | ~n18365;
  assign n18367 = ~pi0773 & n18233;
  assign n18368 = ~pi0684 & n17509;
  assign n18369 = ~n18367 & ~n18368;
  assign n18370 = ~pi0699 & n17510;
  assign n18371 = ~pi0716 & n17531;
  assign n18372 = ~n18370 & ~n18371;
  assign po2131 = ~n18369 | ~n18372;
  assign n18374 = ~pi0642 & n18233;
  assign n18375 = ~pi0685 & n17509;
  assign n18376 = ~n18374 & ~n18375;
  assign n18377 = ~pi0701 & n17510;
  assign n18378 = ~pi0661 & n17531;
  assign n18379 = ~n18377 & ~n18378;
  assign po2133 = ~n18376 | ~n18379;
  assign n18381 = ~pi0774 & n18233;
  assign n18382 = ~pi0686 & n17509;
  assign n18383 = ~n18381 & ~n18382;
  assign n18384 = ~pi0664 & n17510;
  assign n18385 = ~pi0717 & n17531;
  assign n18386 = ~n18384 & ~n18385;
  assign po2134 = ~n18383 | ~n18386;
  assign n18388 = ~pi0687 & n17509;
  assign n18389 = ~pi0702 & n17510;
  assign n18390 = ~n18388 & ~n18389;
  assign n18391 = ~pi0775 & n18233;
  assign n18392 = ~pi0718 & n17531;
  assign n18393 = ~n18391 & ~n18392;
  assign po2135 = ~n18390 | ~n18393;
  assign n18395 = ~pi0776 & n18233;
  assign n18396 = ~pi0703 & n17510;
  assign n18397 = ~n18395 & ~n18396;
  assign n18398 = ~pi0688 & n17509;
  assign n18399 = ~pi0719 & n17531;
  assign n18400 = ~n18398 & ~n18399;
  assign po2136 = ~n18397 | ~n18400;
  assign n18402 = ~pi0644 & n18233;
  assign n18403 = ~pi0689 & n17509;
  assign n18404 = ~n18402 & ~n18403;
  assign n18405 = ~pi0704 & n17510;
  assign n18406 = ~pi0722 & n17531;
  assign n18407 = ~n18405 & ~n18406;
  assign po2137 = ~n18404 | ~n18407;
  assign n18409 = ~pi0777 & n18233;
  assign n18410 = ~pi0739 & n17509;
  assign n18411 = ~n18409 & ~n18410;
  assign n18412 = ~pi0805 & n17510;
  assign n18413 = ~pi0721 & n17531;
  assign n18414 = ~n18412 & ~n18413;
  assign po2138 = ~n18411 | ~n18414;
  assign n18416 = ~pi0750 & n18003;
  assign n18417 = ~pi0548 & n17517;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = ~pi0471 & n17516;
  assign n18420 = ~pi0460 & n17482;
  assign n18421 = ~n18419 & ~n18420;
  assign po2139 = ~n18418 | ~n18421;
  assign n18423 = ~pi0626 & n18003;
  assign n18424 = ~pi0550 & n17517;
  assign n18425 = ~n18423 & ~n18424;
  assign n18426 = ~pi0491 & n17516;
  assign n18427 = ~pi0537 & n17482;
  assign n18428 = ~n18426 & ~n18427;
  assign po2140 = ~n18425 | ~n18428;
  assign n18430 = ~pi0650 & n18233;
  assign n18431 = ~pi0678 & n17509;
  assign n18432 = ~n18430 & ~n18431;
  assign n18433 = ~pi0711 & n17510;
  assign n18434 = ~pi0709 & n17531;
  assign n18435 = ~n18433 & ~n18434;
  assign po2141 = ~n18432 | ~n18435;
  assign n18437 = ~pi1915 & ~pi1918;
  assign n18438 = ~pi0441 & n18437;
  assign n18439 = ~pi0564 & n17502;
  assign n18440 = ~n18438 & ~n18439;
  assign n18441 = ~pi0578 & n17503;
  assign n18442 = ~pi0473 & n17490;
  assign n18443 = ~n18441 & ~n18442;
  assign po2142 = ~n18440 | ~n18443;
  assign n18445 = ~pi0442 & n18437;
  assign n18446 = ~pi0565 & n17502;
  assign n18447 = ~n18445 & ~n18446;
  assign n18448 = ~pi0579 & n17503;
  assign n18449 = ~pi0596 & n17490;
  assign n18450 = ~n18448 & ~n18449;
  assign po2143 = ~n18447 | ~n18450;
  assign n18452 = ~pi0443 & n18437;
  assign n18453 = ~pi0566 & n17502;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = ~pi0580 & n17503;
  assign n18456 = ~pi0593 & n17490;
  assign n18457 = ~n18455 & ~n18456;
  assign po2144 = ~n18454 | ~n18457;
  assign n18459 = ~pi0444 & n18437;
  assign n18460 = ~pi0400 & n17502;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = ~pi0586 & n17503;
  assign n18463 = ~pi0594 & n17490;
  assign n18464 = ~n18462 & ~n18463;
  assign po2145 = ~n18461 | ~n18464;
  assign n18466 = ~pi0445 & n18437;
  assign n18467 = ~pi0401 & n17502;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = ~pi0581 & n17503;
  assign n18470 = ~pi0474 & n17490;
  assign n18471 = ~n18469 & ~n18470;
  assign po2146 = ~n18468 | ~n18471;
  assign n18473 = ~pi0784 & n18003;
  assign n18474 = ~pi0509 & n17516;
  assign n18475 = ~n18473 & ~n18474;
  assign n18476 = ~pi0556 & n17517;
  assign n18477 = ~pi0541 & n17482;
  assign n18478 = ~n18476 & ~n18477;
  assign po2147 = ~n18475 | ~n18478;
  assign n18480 = ~pi0446 & n18437;
  assign n18481 = ~pi0582 & n17503;
  assign n18482 = ~n18480 & ~n18481;
  assign n18483 = ~pi0569 & n17502;
  assign n18484 = ~pi0472 & n17490;
  assign n18485 = ~n18483 & ~n18484;
  assign po2148 = ~n18482 | ~n18485;
  assign n18487 = ~pi0447 & n18437;
  assign n18488 = ~pi0476 & n17502;
  assign n18489 = ~n18487 & ~n18488;
  assign n18490 = ~pi0583 & n17503;
  assign n18491 = ~pi0595 & n17490;
  assign n18492 = ~n18490 & ~n18491;
  assign po2149 = ~n18489 | ~n18492;
  assign n18494 = ~pi0607 & n18437;
  assign n18495 = ~pi0402 & n17502;
  assign n18496 = ~n18494 & ~n18495;
  assign n18497 = ~pi0584 & n17503;
  assign n18498 = ~pi0407 & n17490;
  assign n18499 = ~n18497 & ~n18498;
  assign po2150 = ~n18496 | ~n18499;
  assign n18501 = ~pi0638 & n18437;
  assign n18502 = ~pi0585 & n17502;
  assign n18503 = ~n18501 & ~n18502;
  assign n18504 = ~pi0403 & n17503;
  assign n18505 = ~pi0408 & n17490;
  assign n18506 = ~n18504 & ~n18505;
  assign po2151 = ~n18503 | ~n18506;
  assign n18508 = ~pi0355 & n18437;
  assign n18509 = ~pi0357 & n17502;
  assign n18510 = ~n18508 & ~n18509;
  assign n18511 = ~pi0371 & n17503;
  assign n18512 = ~pi0385 & n17490;
  assign n18513 = ~n18511 & ~n18512;
  assign po2152 = ~n18510 | ~n18513;
  assign n18515 = ~pi0356 & n18437;
  assign n18516 = ~pi0358 & n17502;
  assign n18517 = ~n18515 & ~n18516;
  assign n18518 = ~pi0372 & n17503;
  assign n18519 = ~pi0386 & n17490;
  assign n18520 = ~n18518 & ~n18519;
  assign po2153 = ~n18517 | ~n18520;
  assign n18522 = ~pi0634 & n18003;
  assign n18523 = ~pi0560 & n17516;
  assign n18524 = ~n18522 & ~n18523;
  assign n18525 = ~pi0742 & n17517;
  assign n18526 = ~pi0731 & n17482;
  assign n18527 = ~n18525 & ~n18526;
  assign po2154 = ~n18524 | ~n18527;
  assign n18529 = ~pi0448 & n18437;
  assign n18530 = ~pi0570 & n17502;
  assign n18531 = ~n18529 & ~n18530;
  assign n18532 = ~pi0404 & n17503;
  assign n18533 = ~pi0600 & n17490;
  assign n18534 = ~n18532 & ~n18533;
  assign po2155 = ~n18531 | ~n18534;
  assign n18536 = ~pi0608 & n18437;
  assign n18537 = ~pi0359 & n17502;
  assign n18538 = ~n18536 & ~n18537;
  assign n18539 = ~pi0373 & n17503;
  assign n18540 = ~pi0387 & n17490;
  assign n18541 = ~n18539 & ~n18540;
  assign po2156 = ~n18538 | ~n18541;
  assign n18543 = ~pi0609 & n18437;
  assign n18544 = ~pi0374 & n17503;
  assign n18545 = ~n18543 & ~n18544;
  assign n18546 = ~pi0360 & n17502;
  assign n18547 = ~pi0388 & n17490;
  assign n18548 = ~n18546 & ~n18547;
  assign po2157 = ~n18545 | ~n18548;
  assign n18550 = ~pi0610 & n18437;
  assign n18551 = ~pi0361 & n17502;
  assign n18552 = ~n18550 & ~n18551;
  assign n18553 = ~pi0375 & n17503;
  assign n18554 = ~pi0389 & n17490;
  assign n18555 = ~n18553 & ~n18554;
  assign po2158 = ~n18552 | ~n18555;
  assign n18557 = ~pi0611 & n18437;
  assign n18558 = ~pi0362 & n17502;
  assign n18559 = ~n18557 & ~n18558;
  assign n18560 = ~pi0376 & n17503;
  assign n18561 = ~pi0390 & n17490;
  assign n18562 = ~n18560 & ~n18561;
  assign po2159 = ~n18559 | ~n18562;
  assign n18564 = ~pi0612 & n18437;
  assign n18565 = ~pi0363 & n17502;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = ~pi0377 & n17503;
  assign n18568 = ~pi0391 & n17490;
  assign n18569 = ~n18567 & ~n18568;
  assign po2160 = ~n18566 | ~n18569;
  assign n18571 = ~pi0613 & n18437;
  assign n18572 = ~pi0364 & n17502;
  assign n18573 = ~n18571 & ~n18572;
  assign n18574 = ~pi0378 & n17503;
  assign n18575 = ~pi0392 & n17490;
  assign n18576 = ~n18574 & ~n18575;
  assign po2161 = ~n18573 | ~n18576;
  assign n18578 = ~pi0615 & n18437;
  assign n18579 = ~pi0365 & n17502;
  assign n18580 = ~n18578 & ~n18579;
  assign n18581 = ~pi0379 & n17503;
  assign n18582 = ~pi0393 & n17490;
  assign n18583 = ~n18581 & ~n18582;
  assign po2162 = ~n18580 | ~n18583;
  assign n18585 = ~pi0616 & n18437;
  assign n18586 = ~pi0366 & n17502;
  assign n18587 = ~n18585 & ~n18586;
  assign n18588 = ~pi0380 & n17503;
  assign n18589 = ~pi0394 & n17490;
  assign n18590 = ~n18588 & ~n18589;
  assign po2163 = ~n18587 | ~n18590;
  assign n18592 = ~pi0618 & n18437;
  assign n18593 = ~pi0367 & n17502;
  assign n18594 = ~n18592 & ~n18593;
  assign n18595 = ~pi0381 & n17503;
  assign n18596 = ~pi0395 & n17490;
  assign n18597 = ~n18595 & ~n18596;
  assign po2164 = ~n18594 | ~n18597;
  assign n18599 = ~pi0619 & n18437;
  assign n18600 = ~pi0368 & n17502;
  assign n18601 = ~n18599 & ~n18600;
  assign n18602 = ~pi0382 & n17503;
  assign n18603 = ~pi0396 & n17490;
  assign n18604 = ~n18602 & ~n18603;
  assign po2165 = ~n18601 | ~n18604;
  assign n18606 = ~pi0620 & n18437;
  assign n18607 = ~pi0571 & n17502;
  assign n18608 = ~n18606 & ~n18607;
  assign n18609 = ~pi0587 & n17503;
  assign n18610 = ~pi0597 & n17490;
  assign n18611 = ~n18609 & ~n18610;
  assign po2166 = ~n18608 | ~n18611;
  assign n18613 = ~pi0621 & n18437;
  assign n18614 = ~pi0369 & n17502;
  assign n18615 = ~n18613 & ~n18614;
  assign n18616 = ~pi0383 & n17503;
  assign n18617 = ~pi0397 & n17490;
  assign n18618 = ~n18616 & ~n18617;
  assign po2167 = ~n18615 | ~n18618;
  assign n18620 = ~pi0622 & n18437;
  assign n18621 = ~pi0370 & n17502;
  assign n18622 = ~n18620 & ~n18621;
  assign n18623 = ~pi0384 & n17503;
  assign n18624 = ~pi0398 & n17490;
  assign n18625 = ~n18623 & ~n18624;
  assign po2168 = ~n18622 | ~n18625;
  assign n18627 = ~pi0623 & n18437;
  assign n18628 = ~pi0572 & n17502;
  assign n18629 = ~n18627 & ~n18628;
  assign n18630 = ~pi0588 & n17503;
  assign n18631 = ~pi0598 & n17490;
  assign n18632 = ~n18630 & ~n18631;
  assign po2169 = ~n18629 | ~n18632;
  assign n18634 = ~pi0625 & n18437;
  assign n18635 = ~pi0573 & n17502;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = ~pi0590 & n17503;
  assign n18638 = ~pi0599 & n17490;
  assign n18639 = ~n18637 & ~n18638;
  assign po2170 = ~n18636 | ~n18639;
  assign n18641 = ~pi0604 & n18437;
  assign n18642 = ~pi0574 & n17502;
  assign n18643 = ~n18641 & ~n18642;
  assign n18644 = ~pi0591 & n17503;
  assign n18645 = ~pi0409 & n17490;
  assign n18646 = ~n18644 & ~n18645;
  assign po2171 = ~n18643 | ~n18646;
  assign n18648 = ~pi0628 & n18437;
  assign n18649 = ~pi0477 & n17502;
  assign n18650 = ~n18648 & ~n18649;
  assign n18651 = ~pi0589 & n17503;
  assign n18652 = ~pi0410 & n17490;
  assign n18653 = ~n18651 & ~n18652;
  assign po2172 = ~n18650 | ~n18653;
  assign n18655 = ~pi0630 & n18437;
  assign n18656 = ~pi0405 & n17503;
  assign n18657 = ~n18655 & ~n18656;
  assign n18658 = ~pi0575 & n17502;
  assign n18659 = ~pi0399 & n17490;
  assign n18660 = ~n18658 & ~n18659;
  assign po2173 = ~n18657 | ~n18660;
  assign n18662 = ~pi0631 & n18437;
  assign n18663 = ~pi0576 & n17502;
  assign n18664 = ~n18662 & ~n18663;
  assign n18665 = ~pi0406 & n17503;
  assign n18666 = ~pi0557 & n17490;
  assign n18667 = ~n18665 & ~n18666;
  assign po2174 = ~n18664 | ~n18667;
  assign n18669 = ~pi0633 & n18437;
  assign n18670 = ~pi0577 & n17502;
  assign n18671 = ~n18669 & ~n18670;
  assign n18672 = ~pi0592 & n17503;
  assign n18673 = ~pi0558 & n17490;
  assign n18674 = ~n18672 & ~n18673;
  assign po2175 = ~n18671 | ~n18674;
  assign n18676 = ~pi0759 & n18233;
  assign n18677 = ~pi0747 & n17509;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 = ~pi0694 & n17510;
  assign n18680 = ~pi0663 & n17531;
  assign n18681 = ~n18679 & ~n18680;
  assign po2176 = ~n18678 | ~n18681;
  assign n18683 = ~pi0649 & n18233;
  assign n18684 = ~pi0681 & n17509;
  assign n18685 = ~n18683 & ~n18684;
  assign n18686 = ~pi0696 & n17510;
  assign n18687 = ~pi0713 & n17531;
  assign n18688 = ~n18686 & ~n18687;
  assign po2177 = ~n18685 | ~n18688;
  assign n18690 = ~pi0754 & n18233;
  assign n18691 = ~pi0675 & n17509;
  assign n18692 = ~n18690 & ~n18691;
  assign n18693 = ~pi0690 & n17510;
  assign n18694 = ~pi0705 & n17531;
  assign n18695 = ~n18693 & ~n18694;
  assign po2178 = ~n18692 | ~n18695;
  assign n18697 = ~pi0757 & n18233;
  assign n18698 = ~pi0677 & n17509;
  assign n18699 = ~n18697 & ~n18698;
  assign n18700 = ~pi0658 & n17510;
  assign n18701 = ~pi0708 & n17531;
  assign n18702 = ~n18700 & ~n18701;
  assign po2179 = ~n18699 | ~n18702;
  assign n18704 = ~pi0755 & n18233;
  assign n18705 = ~pi0691 & n17510;
  assign n18706 = ~n18704 & ~n18705;
  assign n18707 = ~pi0676 & n17509;
  assign n18708 = ~pi0706 & n17531;
  assign n18709 = ~n18707 & ~n18708;
  assign po2180 = ~n18706 | ~n18709;
  assign n18711 = ~pi0761 & n18233;
  assign n18712 = ~pi0682 & n17509;
  assign n18713 = ~n18711 & ~n18712;
  assign n18714 = ~pi0697 & n17510;
  assign n18715 = ~pi0662 & n17531;
  assign n18716 = ~n18714 & ~n18715;
  assign po2181 = ~n18713 | ~n18716;
  assign n18718 = ~pi2201 & n5417;
  assign po2182 = n5414 & n18718;
  assign n18720 = n5415 & n17951;
  assign po2183 = n5414 & n18720;
  assign n18722 = pi2163 & ~pi2180;
  assign n18723 = ~pi2163 & pi2180;
  assign po2184 = n18722 | n18723;
  assign n18725 = ~pi0873 & pi2143;
  assign n18726 = pi0873 & pi0878;
  assign po2194 = n18725 | n18726;
  assign n18728 = ~pi0873 & pi2144;
  assign n18729 = pi0478 & pi0873;
  assign po2195 = n18728 | n18729;
  assign n18731 = ~pi0873 & pi2145;
  assign n18732 = pi0210 & pi0873;
  assign po2196 = n18731 | n18732;
  assign n18734 = ~pi0873 & pi2146;
  assign n18735 = pi0873 & pi1923;
  assign po2197 = n18734 | n18735;
  assign n18737 = ~pi0873 & pi2147;
  assign n18738 = pi0869 & pi0873;
  assign po2198 = n18737 | n18738;
  assign n18740 = ~pi0873 & pi2148;
  assign n18741 = pi0194 & pi0873;
  assign po2199 = n18740 | n18741;
  assign n18743 = ~pi0873 & pi2149;
  assign n18744 = pi0336 & pi0873;
  assign po2200 = n18743 | n18744;
  assign n18746 = ~pi0873 & pi2150;
  assign n18747 = pi0190 & pi0873;
  assign po2201 = n18746 | n18747;
  assign n18749 = ~pi0873 & pi2151;
  assign n18750 = pi0873 & pi0948;
  assign po2202 = n18749 | n18750;
  assign n18752 = ~pi0873 & pi2152;
  assign n18753 = pi0817 & pi0873;
  assign po2203 = n18752 | n18753;
  assign n18755 = ~pi0873 & pi2153;
  assign n18756 = pi0234 & pi0873;
  assign po2204 = n18755 | n18756;
  assign n18758 = ~pi0873 & pi2154;
  assign n18759 = pi0205 & pi0873;
  assign po2205 = n18758 | n18759;
  assign n18761 = ~pi0873 & pi2155;
  assign n18762 = pi0873 & pi1885;
  assign po2206 = n18761 | n18762;
  assign n18764 = ~pi0873 & pi2156;
  assign n18765 = pi0873 & pi1932;
  assign po2207 = n18764 | n18765;
  assign n18767 = ~pi0873 & pi2157;
  assign n18768 = pi0873 & pi0906;
  assign po2208 = n18767 | n18768;
  assign n18770 = ~pi0873 & pi2160;
  assign n18771 = pi0873 & pi1851;
  assign po2211 = n18770 | n18771;
  assign n18773 = pi2013 & pi2202;
  assign po2213 = n17573 & n18773;
  assign po0247 = 1'b1;
  assign po2214 = ~pi2180;
  assign po2216 = ~pi2204;
  assign po0000 = pi1858;
  assign po0001 = pi0898;
  assign po0002 = pi1869;
  assign po0003 = pi1867;
  assign po0004 = pi1835;
  assign po0005 = pi1866;
  assign po0006 = pi1836;
  assign po0007 = pi1864;
  assign po0008 = pi1868;
  assign po0009 = pi1863;
  assign po0010 = pi1837;
  assign po0011 = pi1862;
  assign po0012 = pi1861;
  assign po0013 = pi1860;
  assign po0014 = pi1859;
  assign po0015 = pi1865;
  assign po0016 = pi1890;
  assign po0017 = pi1893;
  assign po0018 = pi1902;
  assign po0019 = pi1892;
  assign po0020 = pi1891;
  assign po0021 = pi1889;
  assign po0022 = pi1888;
  assign po0023 = pi1887;
  assign po0024 = pi1894;
  assign po0025 = pi1900;
  assign po0026 = pi1898;
  assign po0027 = pi1897;
  assign po0028 = pi1896;
  assign po0029 = pi1899;
  assign po0030 = pi1895;
  assign po0031 = pi1882;
  assign po0032 = pi1963;
  assign po0033 = pi1945;
  assign po0034 = pi2134;
  assign po0036 = pi0000;
  assign po0037 = pi0924;
  assign po0038 = pi0201;
  assign po0039 = pi0198;
  assign po0040 = pi0202;
  assign po0041 = pi0199;
  assign po0042 = pi0203;
  assign po0043 = pi0204;
  assign po0044 = pi0347;
  assign po0045 = pi0348;
  assign po0046 = pi0332;
  assign po0047 = pi2204;
  assign po0246 = pi2200;
  assign po0248 = pi2199;
  assign po0260 = pi0228;
  assign po0279 = pi0331;
  assign po0382 = pi0456;
  assign po0507 = pi0640;
  assign po0691 = pi0840;
  assign po0891 = pi0876;
  assign po0927 = pi0891;
  assign po0942 = pi0925;
  assign po0976 = pi1768;
  assign po0997 = pi1930;
  assign po1819 = pi1880;
  assign po1931 = pi1906;
  assign po1957 = pi1928;
  assign po1979 = pi1942;
  assign po1981 = pi1953;
  assign po1982 = pi1954;
  assign po1993 = pi1992;
  assign po1994 = pi1991;
  assign po2003 = pi2011;
  assign po2004 = pi2002;
  assign po2005 = pi2012;
  assign po2042 = pi2015;
  assign po2043 = pi2014;
  assign po2062 = pi2037;
  assign po2065 = pi2081;
  assign po2132 = pi2142;
  assign po2193 = pi2161;
  assign po2212 = pi2164;
  assign po2215 = pi2165;
  assign po2217 = pi2205;
  assign po2218 = pi2213;
  assign po2219 = pi2210;
  assign po2220 = pi2218;
  assign po2221 = pi2230;
  assign po2222 = pi2232;
  assign po2223 = pi2229;
  assign po2224 = pi2217;
  assign po2225 = pi2237;
  assign po2226 = pi2219;
  assign po2227 = pi2235;
  assign po2228 = pi2228;
  assign po2229 = pi2236;
  assign po2230 = pi2221;
  assign po2231 = pi2225;
  assign po2232 = pi2233;
  assign po2233 = pi2234;
  assign po2234 = pi2216;
  assign po2235 = pi2212;
  assign po2236 = pi2226;
  assign po2237 = pi2206;
  assign po2238 = pi2227;
  assign po2239 = pi2211;
  assign po2240 = pi2224;
  assign po2241 = pi2231;
  assign po2242 = pi2208;
  assign po2243 = pi2215;
  assign po2244 = pi2223;
  assign po2245 = pi2209;
  assign po2246 = pi2214;
  assign po2247 = pi2222;
  assign po2248 = pi2220;
  assign po2249 = pi2207;
endmodule


