// Benchmark "C17.iscas" written by ABC on Fri Mar  3 17:59:48 2017

module \C17.iscas  ( 
    pi0, pi1, pi2, pi3, pi4,
    po0, po1  );
  input  pi0, pi1, pi2, pi3, pi4;
  output po0, po1;
  wire n9, n10,n11 ,n12;
  assign n9 = pi2 & pi3;
  assign n10 = pi0 & pi2;
  assign n11 = ~n9 & pi1;
  assign n12 = pi1 | pi4;
  assign po0 = n10 | n11;
  assign po1 = ~n9 & n12;
endmodule


